netcdf ecmwf_r24_2018062300_f096 {
dimensions: 
 lat = 601; 
 lon = 701; 
variables:  
float lat(lat) ; 
   lat:long_name = "latitude" ;
   lat:units = "degrees_north" ;
   lat:standard_name = "latitude" ;
float lon(lon) ;
   lon:long_name = "longitude" ;
   lon:units = "degrees_east" ;
   lon:standard_name = "longitude" ;
float APCP_24(lat, lon) ;
   APCP_24:name = "APCP_24" ;
   APCP_24:long_name = "Total Precipitation" ;
   APCP_24:level = "A24" ;
   APCP_24:units = "kg/m^2" ;
   APCP_24:_FillValue = -9999.f ;
   APCP_24:init_time = "20180623_000000" ;
   APCP_24:init_time_ut = "1529712000.0" ;
   APCP_24:valid_time = "20180627_000000" ;
   APCP_24:valid_time_ut = "1530057600.0" ;
   APCP_24:accum_time = "240000" ;
   APCP_24:_FillValue = 65535 ;
   APCP_24:accum_time_sec = 86400 ;
 // global attributes: 
 :_NCProperties = "version=1|netcdflibversion=4.4.1.1" ;
	:FileOrigins = "ECMWF_HR_APCP24" ; 
	:MET_version = "V7.0" ;
	:Projection = "LatLon" ;
	:lat_ll = "0.0 degrees_north" ; 
	:lon_ll = "70.0 degrees_east" ; 
	:delta_lat = "0.10 degrees" ;
	:delta_lon = "0.10 degrees" ;
	:Nlat = "601 grid_points" ; 
	:Nlon = "701 grid_points" ; 
data:
lat = 0.0,0.1,0.2,0.3,0.4,0.5,0.6,0.7,0.8,0.90000004,1.0,1.1,1.2,1.3000001,1.4,1.5,1.6,1.7,1.8000001,1.9,2.0,2.1000001,2.2,2.3,2.4,2.5,2.6000001,2.7,2.8,2.9,3.0,3.1000001,3.2,3.3,3.4,3.5,3.6000001,3.7,3.8,3.9,4.0,4.1,4.2000003,4.3,4.4,4.5,4.6,4.7000003,4.8,4.9,5.0,5.1,5.2000003,5.3,5.4,5.5,5.6,5.7000003,5.8,5.9,6.0,6.1,6.2000003,6.3,6.4,6.5,6.6,6.7000003,6.8,6.9,7.0,7.1,7.2000003,7.3,7.4,7.5,7.6,7.7000003,7.8,7.9,8.0,8.1,8.2,8.3,8.400001,8.5,8.6,8.7,8.8,8.900001,9.0,9.1,9.2,9.3,9.400001,9.5,9.6,9.7,9.8,9.900001,10.0,10.1,10.2,10.3,10.400001,10.5,10.6,10.7,10.8,10.900001,11.0,11.1,11.2,11.3,11.400001,11.5,11.6,11.7,11.8,11.900001,12.0,12.1,12.2,12.3,12.400001,12.5,12.6,12.7,12.8,12.900001,13.0,13.1,13.2,13.3,13.400001,13.5,13.6,13.7,13.8,13.900001,14.0,14.1,14.2,14.3,14.400001,14.5,14.6,14.7,14.8,14.900001,15.0,15.1,15.2,15.3,15.400001,15.5,15.6,15.7,15.8,15.900001,16.0,16.1,16.2,16.300001,16.4,16.5,16.6,16.7,16.800001,16.9,17.0,17.1,17.2,17.300001,17.4,17.5,17.6,17.7,17.800001,17.9,18.0,18.1,18.2,18.300001,18.4,18.5,18.6,18.7,18.800001,18.9,19.0,19.1,19.2,19.300001,19.4,19.5,19.6,19.7,19.800001,19.9,20.0,20.1,20.2,20.300001,20.4,20.5,20.6,20.7,20.800001,20.9,21.0,21.1,21.2,21.300001,21.4,21.5,21.6,21.7,21.800001,21.9,22.0,22.1,22.2,22.300001,22.4,22.5,22.6,22.7,22.800001,22.9,23.0,23.1,23.2,23.300001,23.4,23.5,23.6,23.7,23.800001,23.9,24.0,24.1,24.2,24.300001,24.4,24.5,24.6,24.7,24.800001,24.9,25.0,25.1,25.2,25.300001,25.4,25.5,25.6,25.7,25.800001,25.9,26.0,26.1,26.2,26.300001,26.4,26.5,26.6,26.7,26.800001,26.9,27.0,27.1,27.2,27.300001,27.4,27.5,27.6,27.7,27.800001,27.9,28.0,28.1,28.2,28.300001,28.4,28.5,28.6,28.7,28.800001,28.9,29.0,29.1,29.2,29.300001,29.4,29.5,29.6,29.7,29.800001,29.9,30.0,30.1,30.2,30.300001,30.4,30.5,30.6,30.7,30.800001,30.9,31.0,31.1,31.2,31.300001,31.4,31.5,31.6,31.7,31.800001,31.9,32.0,32.100002,32.2,32.3,32.4,32.5,32.600002,32.7,32.8,32.9,33.0,33.100002,33.2,33.3,33.4,33.5,33.600002,33.7,33.8,33.9,34.0,34.100002,34.2,34.3,34.4,34.5,34.600002,34.7,34.8,34.9,35.0,35.100002,35.2,35.3,35.4,35.5,35.600002,35.7,35.8,35.9,36.0,36.100002,36.2,36.3,36.4,36.5,36.600002,36.7,36.8,36.9,37.0,37.100002,37.2,37.3,37.4,37.5,37.600002,37.7,37.8,37.9,38.0,38.100002,38.2,38.3,38.4,38.5,38.600002,38.7,38.8,38.9,39.0,39.100002,39.2,39.3,39.4,39.5,39.600002,39.7,39.8,39.9,40.0,40.100002,40.2,40.3,40.4,40.5,40.600002,40.7,40.8,40.9,41.0,41.100002,41.2,41.3,41.4,41.5,41.600002,41.7,41.8,41.9,42.0,42.100002,42.2,42.3,42.4,42.5,42.600002,42.7,42.8,42.9,43.0,43.100002,43.2,43.3,43.4,43.5,43.600002,43.7,43.8,43.9,44.0,44.100002,44.2,44.3,44.4,44.5,44.600002,44.7,44.8,44.9,45.0,45.100002,45.2,45.3,45.4,45.5,45.600002,45.7,45.8,45.9,46.0,46.100002,46.2,46.3,46.4,46.5,46.600002,46.7,46.8,46.9,47.0,47.100002,47.2,47.3,47.4,47.5,47.600002,47.7,47.8,47.9,48.0,48.100002,48.2,48.3,48.4,48.5,48.600002,48.7,48.8,48.9,49.0,49.100002,49.2,49.3,49.4,49.5,49.600002,49.7,49.8,49.9,50.0,50.100002,50.2,50.3,50.4,50.5,50.600002,50.7,50.8,50.9,51.0,51.100002,51.2,51.3,51.4,51.5,51.600002,51.7,51.8,51.9,52.0,52.100002,52.2,52.3,52.4,52.5,52.600002,52.7,52.8,52.9,53.0,53.100002,53.2,53.3,53.4,53.5,53.600002,53.7,53.8,53.9,54.0,54.100002,54.2,54.3,54.4,54.5,54.600002,54.7,54.8,54.9,55.0,55.100002,55.2,55.3,55.4,55.5,55.600002,55.7,55.8,55.9,56.0,56.100002,56.2,56.3,56.4,56.5,56.600002,56.7,56.8,56.9,57.0,57.100002,57.2,57.3,57.4,57.5,57.600002,57.7,57.8,57.9,58.0,58.100002,58.2,58.3,58.4,58.5,58.600002,58.7,58.8,58.9,59.0,59.100002,59.2,59.3,59.4,59.5,59.600002,59.7,59.8,59.9,60.0;
lon = 70.0,70.1,70.2,70.3,70.4,70.5,70.6,70.7,70.8,70.9,71.0,71.1,71.2,71.3,71.4,71.5,71.6,71.7,71.8,71.9,72.0,72.1,72.2,72.3,72.4,72.5,72.6,72.7,72.8,72.9,73.0,73.1,73.2,73.3,73.4,73.5,73.6,73.7,73.8,73.9,74.0,74.1,74.2,74.3,74.4,74.5,74.6,74.7,74.8,74.9,75.0,75.1,75.2,75.3,75.4,75.5,75.6,75.7,75.8,75.9,76.0,76.1,76.2,76.3,76.4,76.5,76.6,76.7,76.8,76.9,77.0,77.1,77.2,77.3,77.4,77.5,77.6,77.7,77.8,77.9,78.0,78.1,78.2,78.3,78.4,78.5,78.6,78.7,78.8,78.9,79.0,79.1,79.2,79.3,79.4,79.5,79.6,79.7,79.8,79.9,80.0,80.1,80.2,80.3,80.4,80.5,80.6,80.7,80.8,80.9,81.0,81.1,81.2,81.3,81.4,81.5,81.6,81.7,81.8,81.9,82.0,82.1,82.2,82.3,82.4,82.5,82.6,82.7,82.8,82.9,83.0,83.1,83.2,83.3,83.4,83.5,83.6,83.7,83.8,83.9,84.0,84.1,84.2,84.3,84.4,84.5,84.6,84.7,84.8,84.9,85.0,85.1,85.2,85.3,85.4,85.5,85.6,85.7,85.8,85.9,86.0,86.1,86.2,86.3,86.4,86.5,86.6,86.7,86.8,86.9,87.0,87.1,87.2,87.3,87.4,87.5,87.6,87.7,87.8,87.9,88.0,88.1,88.2,88.3,88.4,88.5,88.6,88.7,88.8,88.9,89.0,89.1,89.2,89.3,89.4,89.5,89.6,89.7,89.8,89.9,90.0,90.1,90.2,90.3,90.4,90.5,90.6,90.7,90.8,90.9,91.0,91.1,91.2,91.3,91.4,91.5,91.6,91.7,91.8,91.9,92.0,92.1,92.2,92.3,92.4,92.5,92.6,92.7,92.8,92.9,93.0,93.1,93.2,93.3,93.4,93.5,93.6,93.7,93.8,93.9,94.0,94.1,94.2,94.3,94.4,94.5,94.6,94.7,94.8,94.9,95.0,95.1,95.2,95.3,95.4,95.5,95.6,95.7,95.8,95.9,96.0,96.1,96.2,96.3,96.4,96.5,96.6,96.7,96.8,96.9,97.0,97.1,97.2,97.3,97.4,97.5,97.6,97.7,97.8,97.9,98.0,98.1,98.2,98.3,98.4,98.5,98.6,98.7,98.8,98.9,99.0,99.1,99.2,99.3,99.4,99.5,99.6,99.7,99.8,99.9,100.0,100.1,100.2,100.3,100.4,100.5,100.6,100.7,100.8,100.9,101.0,101.1,101.2,101.3,101.4,101.5,101.6,101.7,101.8,101.9,102.0,102.100006,102.2,102.3,102.4,102.5,102.600006,102.7,102.8,102.9,103.0,103.100006,103.2,103.3,103.4,103.5,103.600006,103.7,103.8,103.9,104.0,104.100006,104.2,104.3,104.4,104.5,104.600006,104.7,104.8,104.9,105.0,105.100006,105.2,105.3,105.4,105.5,105.600006,105.7,105.8,105.9,106.0,106.100006,106.2,106.3,106.4,106.5,106.600006,106.7,106.8,106.9,107.0,107.100006,107.2,107.3,107.4,107.5,107.600006,107.7,107.8,107.9,108.0,108.100006,108.2,108.3,108.4,108.5,108.600006,108.7,108.8,108.9,109.0,109.100006,109.2,109.3,109.4,109.5,109.600006,109.7,109.8,109.9,110.0,110.100006,110.2,110.3,110.4,110.5,110.600006,110.7,110.8,110.9,111.0,111.100006,111.2,111.3,111.4,111.5,111.600006,111.7,111.8,111.9,112.0,112.100006,112.2,112.3,112.4,112.5,112.600006,112.7,112.8,112.9,113.0,113.100006,113.2,113.3,113.4,113.5,113.600006,113.7,113.8,113.9,114.0,114.100006,114.2,114.3,114.4,114.5,114.600006,114.7,114.8,114.9,115.0,115.100006,115.2,115.3,115.4,115.5,115.600006,115.7,115.8,115.9,116.0,116.100006,116.2,116.3,116.4,116.5,116.600006,116.7,116.8,116.9,117.0,117.100006,117.2,117.3,117.4,117.5,117.600006,117.7,117.8,117.9,118.0,118.100006,118.2,118.3,118.4,118.5,118.600006,118.7,118.8,118.9,119.0,119.100006,119.2,119.3,119.4,119.5,119.600006,119.7,119.8,119.9,120.0,120.100006,120.2,120.3,120.4,120.5,120.600006,120.7,120.8,120.9,121.0,121.100006,121.2,121.3,121.4,121.5,121.600006,121.7,121.8,121.9,122.0,122.100006,122.2,122.3,122.4,122.5,122.600006,122.7,122.8,122.9,123.0,123.100006,123.2,123.3,123.4,123.5,123.600006,123.7,123.8,123.9,124.0,124.100006,124.2,124.3,124.4,124.5,124.600006,124.7,124.8,124.9,125.0,125.100006,125.2,125.3,125.4,125.5,125.600006,125.7,125.8,125.9,126.0,126.100006,126.2,126.3,126.4,126.5,126.600006,126.7,126.8,126.9,127.0,127.100006,127.2,127.3,127.4,127.5,127.600006,127.7,127.8,127.9,128.0,128.1,128.2,128.3,128.4,128.5,128.6,128.7,128.8,128.9,129.0,129.1,129.2,129.3,129.4,129.5,129.6,129.7,129.8,129.9,130.0,130.1,130.2,130.3,130.4,130.5,130.6,130.7,130.8,130.9,131.0,131.1,131.2,131.3,131.4,131.5,131.6,131.7,131.8,131.9,132.0,132.1,132.2,132.3,132.4,132.5,132.6,132.7,132.8,132.9,133.0,133.1,133.2,133.3,133.4,133.5,133.6,133.7,133.8,133.9,134.0,134.1,134.20001,134.3,134.4,134.5,134.6,134.70001,134.8,134.9,135.0,135.1,135.20001,135.3,135.4,135.5,135.6,135.70001,135.8,135.9,136.0,136.1,136.20001,136.3,136.4,136.5,136.6,136.70001,136.8,136.9,137.0,137.1,137.20001,137.3,137.4,137.5,137.6,137.70001,137.8,137.9,138.0,138.1,138.20001,138.3,138.4,138.5,138.6,138.70001,138.8,138.9,139.0,139.1,139.20001,139.3,139.4,139.5,139.6,139.70001,139.8,139.9,140.0;
APCP_24 = 10.725573,11.080199,12.15917,13.505998,14.509516,14.388792,12.898605,12.445889,12.774108,13.309821,13.13628,12.049765,11.955449,12.098808,12.366665,13.245687,13.36641,14.011529,15.230087,16.920223,18.814081,18.580177,18.040693,18.006739,18.342503,17.912424,17.644567,17.338985,16.358103,15.015047,14.588741,14.234114,13.679539,13.36641,13.151371,12.283667,11.076427,10.891568,11.076427,11.155652,10.86516,9.740918,9.480607,8.880759,7.6697464,6.485142,6.387054,5.915476,5.304311,4.678055,4.044254,4.5912848,5.342037,6.368191,7.3415284,7.537705,6.587003,5.8626595,5.5985756,5.670255,5.583485,4.9987283,4.402653,4.304565,4.5724216,4.425289,4.6554193,4.979865,5.27413,5.485397,5.643847,5.413717,5.1534057,5.1232247,5.4250345,6.013564,5.7419353,5.4212623,5.194905,5.243949,5.7683434,5.7683434,5.3910813,5.2099953,5.5683947,6.6058664,7.6207023,7.8923316,7.673519,7.2094865,6.760544,6.307829,6.2323766,6.2361493,6.0701537,5.5080323,5.119452,5.413717,5.926794,6.387054,6.730363,6.6813188,6.6134114,6.741681,7.1076255,7.5829763,7.865923,7.8508325,7.7112455,7.699928,8.16396,7.748972,7.0849895,7.4471617,8.820397,9.918231,10.076681,9.9257765,9.733373,9.703192,9.933322,10.982111,11.970539,12.830698,13.321139,13.015556,12.038446,11.136789,10.419991,9.895596,9.446653,9.175024,8.514814,7.598067,6.828451,6.851087,6.779407,6.8435416,6.6662283,6.2436943,5.9494295,5.4250345,5.4703064,5.613666,5.6061206,5.3873086,5.4703064,5.3194013,5.081726,4.9157305,4.991183,4.9534564,4.447925,4.002755,3.7914882,3.6330378,3.5689032,3.5387223,3.6669915,3.9008942,3.9989824,3.85185,3.7952607,3.6669915,3.3727267,2.8822856,2.2598023,1.8297231,1.5882751,1.4713237,1.3732355,1.1544232,1.0978339,1.0789708,1.0450171,1.0072908,0.8224323,0.8224323,0.87902164,0.8941121,0.80734175,0.79602385,0.694163,0.47912338,0.2565385,0.24522063,0.2565385,0.29426476,0.27917424,0.19994913,0.1358145,0.1358145,0.10940613,0.071679875,0.0452715,0.0452715,0.0452715,0.0452715,0.0452715,0.049044125,0.060362,0.060362,0.060362,0.060362,0.06790725,0.090543,0.12826926,0.120724,0.094315626,0.0754525,0.0754525,0.11317875,0.13204187,0.14335975,0.150905,0.150905,0.18863125,0.181086,0.1659955,0.16222288,0.1358145,0.11317875,0.124496624,0.13204187,0.13204187,0.1659955,0.13204187,0.11317875,0.10186087,0.08677038,0.060362,0.060362,0.07922512,0.08677038,0.071679875,0.060362,0.071679875,0.1056335,0.08677038,0.033953626,0.0452715,0.1056335,0.1659955,0.20372175,0.21881226,0.24522063,0.29426476,0.452715,0.5319401,0.5772116,0.87147635,1.0035182,0.7809334,0.6149379,0.63002837,0.6413463,0.8601585,1.0148361,0.90543,0.80734175,1.4637785,1.6109109,1.750498,1.5279131,1.0487897,0.8526133,0.965792,0.73566186,0.80356914,1.2411937,1.5731846,0.9016574,0.8224323,0.86770374,0.8563859,0.9318384,0.9922004,1.2713746,2.1013522,3.663219,5.994701,4.2517486,2.305074,2.8106055,4.3800178,1.5731846,2.7313805,3.4783602,4.61392,5.666483,4.8968673,4.9723196,6.590776,6.571913,4.4630156,2.5314314,2.9464202,4.112161,7.3377557,11.6875925,14.007756,8.345046,10.442626,14.777372,17.795471,17.927513,14.1926155,11.200924,8.394091,6.1078796,5.5683947,3.591539,1.7165444,0.90920264,1.0676528,1.0072908,0.45648763,0.422534,0.9016574,1.3204187,0.5055317,0.49044126,0.41498876,0.3169005,0.29049212,0.47157812,0.30181,0.41498876,0.67152727,0.8563859,0.68661773,0.7582976,0.6790725,0.7582976,1.2336484,2.2598023,3.187868,4.8100967,5.462761,5.342037,6.515323,5.8211603,7.2472124,7.0812173,4.938366,3.7537618,2.4974778,3.0709167,3.682082,4.425289,7.2924843,7.3415284,8.224322,8.786444,8.707218,8.499724,10.231359,10.510533,9.978593,9.688101,11.091517,10.823661,11.306557,10.7218,9.0957985,8.314865,8.548768,8.854351,9.378746,9.786189,9.261794,8.89585,8.8769865,8.137552,7.145352,7.888559,8.3525915,9.842778,10.989656,11.068882,9.993684,9.590013,9.967276,10.106862,10.197406,11.61214,12.245941,10.985884,8.258276,5.0666356,2.9916916,2.0372176,5.3080835,7.2358947,6.270103,4.8666863,3.6481283,6.7944975,8.654402,7.707473,6.5455046,5.300538,6.205968,5.8173876,4.274384,5.3269467,7.54525,7.020855,5.617439,4.0970707,2.1051247,3.1312788,2.161714,2.263575,4.1310244,6.0739264,3.0218725,1.3807807,1.9579924,3.9688015,5.0213637,3.3463185,3.3764994,5.0251365,8.13378,12.464753,10.367173,8.533678,7.5188417,6.9869013,5.692891,2.969056,3.0860074,4.715781,6.6624556,7.858378,6.6247296,8.367682,8.2507305,6.255012,7.1566696,4.678055,2.4861598,3.6179473,8.537451,15.0905,16.433554,12.804289,7.6395655,5.032682,9.718282,9.439108,10.220041,11.642321,11.830952,7.462252,9.597558,10.423763,10.469034,9.88805,8.484633,9.337247,9.87296,9.854096,9.57115,9.827688,10.167224,10.144588,10.627484,11.136789,9.842778,8.718536,11.714001,12.155397,10.080454,12.253486,16.780636,23.058285,23.292187,16.38451,7.9489207,8.29223,9.58624,9.782416,8.375228,6.40969,6.432326,9.578695,13.343775,14.992412,11.551778,11.136789,9.556059,7.7942433,6.1720147,4.3649273,4.889322,3.7386713,3.9159849,6.587003,11.091517,11.947904,12.664702,12.242168,10.93684,10.253995,9.020347,9.235386,9.623966,9.971047,11.091517,12.521342,12.117672,12.479843,14.02662,15.015047,13.29473,11.876224,9.390063,8.00551,13.411682,18.87067,18.704676,18.900852,20.013775,17.180534,12.932558,10.770844,12.083718,15.656394,17.686066,23.824127,26.540417,25.204908,21.798227,20.919205,18.844261,17.052265,16.791954,16.603323,12.344029,10.367173,11.00852,11.502733,10.895341,10.038955,6.571913,8.058327,9.378746,9.242931,10.208723,10.770844,11.038701,10.47658,9.891823,11.427281,12.196897,11.959221,11.208468,10.023865,8.073418,7.6923823,8.552541,9.265567,9.148616,8.209232,7.281166,6.1795597,5.704209,5.9984736,6.5455046,6.741681,6.9567204,8.047009,8.933576,6.590776,5.8211603,9.393836,12.310076,13.456953,15.580941,14.626467,13.226823,12.909923,13.754991,14.388792,14.241659,15.845025,17.13149,17.557796,18.082191,17.912424,18.02183,17.72002,16.923996,16.203424,14.875461,13.389046,11.555551,9.446653,7.3868,7.567886,7.6508837,7.115171,6.270103,6.255012,3.5462675,4.644101,7.220804,9.22784,8.91094,7.8017883,6.205968,5.270357,5.13077,4.8968673,5.4476705,5.402399,5.6476197,6.379509,7.1264887,8.039464,8.13378,7.6697464,7.375482,8.439363,9.329701,9.442881,9.258021,9.431562,10.770844,12.004493,12.917468,13.162688,13.155144,14.083209,15.120681,15.811071,15.701665,14.920732,14.173752,14.713238,14.332202,14.071891,13.909668,12.785426,12.67602,12.540206,12.868423,13.992666,16.06761,15.739391,15.4074,15.860115,16.935314,17.53139,19.960958,19.662922,18.587723,17.731337,17.120173,16.776863,16.361876,17.139036,19.032892,20.643805,19.31584,18.599041,18.293459,18.082191,17.53139,17.84829,19.017803,19.7761,19.670467,19.074392,19.806282,20.621168,20.594759,19.466745,17.625704,15.961976,15.675257,15.041456,13.81158,13.215506,13.494679,14.177525,14.856597,15.241405,15.165953,14.1926155,13.864397,14.456699,15.773345,17.165443,17.546478,18.116146,18.648085,19.021576,19.240387,11.751727,11.59705,11.808316,12.468526,13.298503,13.656902,13.230596,13.890805,14.634012,14.954685,14.871688,14.743419,14.626467,14.2944765,13.72481,13.109872,13.86817,15.335721,17.45971,19.557287,20.326904,18.395319,16.535416,15.158407,14.50197,14.641558,15.124454,15.82239,15.890297,15.067864,13.6833105,13.057055,12.842015,12.50248,11.808316,10.842525,9.820143,9.80128,10.174769,10.27663,9.4013815,8.412953,7.5037513,6.651138,5.994701,5.824933,5.9418845,5.9909286,5.7909794,5.462761,5.4363527,6.0739264,6.4134626,6.25124,5.7117543,5.243949,4.9157305,4.5761943,4.4516973,4.67051,5.2665844,5.2099953,5.0515447,4.991183,5.0553174,5.1345425,5.093044,5.3986263,5.617439,5.5268955,5.119452,5.221313,4.870459,4.5761943,4.5422406,4.67051,4.6629643,4.436607,4.4139714,4.768598,5.3910813,5.613666,5.7117543,5.8211603,6.217286,7.3151197,7.3113475,6.802043,6.3455553,6.19465,6.307829,6.217286,5.938112,5.613666,5.379763,5.3759904,5.304311,5.462761,5.5495315,5.587258,5.9003854,6.4474163,6.5945487,6.960493,7.541477,7.6923823,7.466025,7.303802,7.032173,6.8397694,7.284939,7.816879,8.6732645,9.971047,11.314102,11.796998,11.947904,11.740409,11.3820095,11.114153,11.23865,11.830952,11.148107,10.355856,9.929549,9.684328,8.571404,7.7942433,7.6508837,7.8810134,7.6622014,8.126234,7.99042,7.6093845,7.24344,7.069899,7.0963078,6.620957,6.228604,6.1041074,6.0248823,6.085244,6.273875,6.477597,6.515323,6.119198,5.9003854,5.7909794,5.73439,5.6476197,5.4288073,5.458988,4.9459114,4.515832,4.323428,4.0593443,3.8707132,3.783943,3.9499383,4.274384,4.4139714,4.1989317,4.236658,4.1762958,3.8858037,3.4557245,2.795515,2.1881225,1.7731338,1.5656394,1.4600059,1.237421,1.1695137,1.1619685,1.1544232,1.116697,1.0110635,0.9280658,0.875249,0.8299775,0.724344,0.6526641,0.7394345,0.69793564,0.5319401,0.55080324,0.55080324,0.49421388,0.392353,0.29049212,0.26031113,0.19994913,0.181086,0.14713238,0.09808825,0.056589376,0.049044125,0.05281675,0.056589376,0.060362,0.071679875,0.05281675,0.071679875,0.0754525,0.06790725,0.090543,0.12826926,0.120724,0.094315626,0.07922512,0.08677038,0.094315626,0.1056335,0.120724,0.1358145,0.1659955,0.211267,0.211267,0.18863125,0.16222288,0.1358145,0.11317875,0.10940613,0.124496624,0.14713238,0.15467763,0.120724,0.116951376,0.09808825,0.06790725,0.071679875,0.08299775,0.0754525,0.071679875,0.06790725,0.03772625,0.049044125,0.049044125,0.0452715,0.049044125,0.08299775,0.15467763,0.181086,0.19240387,0.1961765,0.18485862,0.241448,0.3734899,0.43385187,0.5470306,1.1129243,1.0223814,0.8111144,0.694163,0.68661773,0.58098423,0.6451189,0.995973,1.2223305,1.3505998,1.8448136,1.9693103,1.8448136,1.327964,0.80734175,1.20724,0.995973,1.146878,1.1355602,0.8941121,0.80356914,0.66775465,0.73188925,0.90920264,1.0487897,0.95447415,1.3204187,1.931584,3.4444065,5.5004873,6.730363,6.458734,4.666737,2.8445592,1.8674494,1.9994912,3.3161373,5.304311,5.87775,5.1534057,5.4476705,6.379509,6.85486,5.794752,4.4177437,6.221059,9.348565,7.8244243,8.3525915,12.653384,17.474798,15.588487,16.58446,15.856343,11.921495,6.3832817,4.8138695,6.436098,7.835742,7.8696957,7.6584287,4.323428,3.1840954,2.463524,1.7957695,2.203213,1.2034674,0.7130261,0.84129536,1.1242423,0.5017591,0.6375736,0.38480774,0.2263575,0.26408374,0.25276586,0.2678564,0.56589377,0.72811663,0.66775465,0.6149379,0.7469798,0.86770374,1.146878,1.6071383,2.1353056,2.867195,4.2027044,5.2250857,5.753253,6.319147,5.1571784,6.7152724,7.1378064,5.413717,3.399135,5.3269467,6.089017,5.926794,5.6476197,6.620957,7.1679873,8.190369,8.782671,8.714764,8.439363,9.0957985,10.133271,10.336992,9.986138,10.812344,10.34831,10.834979,10.710483,9.650374,8.537451,8.797762,8.771353,8.692128,8.499724,7.858378,7.111398,7.752744,7.77538,7.043491,7.2924843,6.8850408,8.084735,9.710737,10.533169,9.261794,9.163706,9.567377,10.329447,11.249968,12.098808,11.3971,10.608622,8.461998,5.462761,3.904667,2.0070364,4.304565,5.1081343,4.6327834,9.016574,6.3908267,7.8319697,7.6886096,5.6476197,6.7039547,6.006019,7.201941,6.779407,4.515832,3.4934506,5.383536,5.032682,4.2064767,3.5538127,2.6182017,1.9429018,1.9542197,2.8785129,4.085753,4.08198,2.3013012,1.056335,1.026154,1.841041,2.0900342,2.957738,4.961002,7.5905213,10.510533,13.5663595,7.069899,5.828706,6.1644692,6.3719635,6.7152724,6.730363,6.1229706,6.085244,6.609639,6.466279,5.243949,9.49947,9.944639,6.126743,6.4247804,6.688864,4.353609,5.6589375,10.872705,14.27184,9.276885,7.303802,7.8621507,9.635284,10.465261,7.54525,7.7338815,11.604594,15.150862,9.793735,8.122461,8.062099,9.110889,10.4049,10.729345,10.79348,9.1976595,10.114408,12.657157,10.86516,11.46878,11.891314,11.449917,10.917976,12.50248,9.397609,9.439108,9.5032425,9.21275,10.948157,15.8676605,20.19109,19.908142,14.656648,7.707473,9.367428,10.291721,10.880251,10.850069,9.265567,8.975075,9.635284,13.58145,17.101309,10.416218,9.989911,8.167733,6.862405,6.48137,5.915476,4.8553686,3.832987,3.591539,5.5306683,11.664956,10.831206,12.728837,13.65313,13.241914,14.50197,11.891314,11.498961,12.268577,13.249459,13.570132,13.788944,13.200415,12.287439,11.5857315,11.695138,13.245687,13.962485,14.158662,14.713238,17.074902,19.678013,20.53817,20.889025,20.168453,15.99593,12.442118,12.196897,14.132254,17.757746,23.250689,25.514263,23.337458,19.478064,15.999702,14.241659,14.317112,14.70192,15.056546,14.547242,11.879996,10.480352,9.295748,8.499724,8.480861,9.831461,8.405409,8.484633,8.650629,8.771353,10.001229,10.970794,11.751727,11.242422,10.201178,11.268831,11.6875925,11.506506,10.646348,9.329701,8.107371,8.160188,8.582722,9.092027,9.216523,8.307321,7.7225633,7.020855,6.802043,7.111398,7.424526,7.1038527,7.1340337,7.914967,8.541223,6.8246784,6.983129,9.495697,12.577931,14.962231,15.882751,15.041456,14.777372,14.600059,14.162435,13.302276,13.830443,15.218769,16.746683,17.765291,17.70493,17.112627,17.437073,17.365393,16.618414,15.946886,14.490653,12.491161,10.38981,8.499724,6.983129,7.7225633,7.877241,7.1340337,5.855114,5.05909,4.52715,5.3571277,5.907931,5.7192993,5.5193505,5.9418845,5.553304,5.3684454,5.323174,4.3007927,4.8968673,5.070408,5.160951,5.300538,5.3910813,5.945657,6.907676,7.3717093,7.273621,7.3868,8.590267,9.076936,9.582467,10.465261,11.69891,11.879996,12.242168,12.672247,13.298503,14.498198,15.762027,16.029884,15.848798,15.799753,16.531643,16.463736,15.558306,14.93205,14.856597,14.78869,14.600059,14.2077055,14.211478,14.856597,16.044973,15.252723,14.958458,15.667711,17.014538,17.738882,19.134754,19.081938,18.723537,18.75372,19.40261,18.79899,17.731337,17.25976,17.640795,18.327412,18.704676,18.795218,18.666948,18.421728,18.214233,18.221779,19.312067,20.225042,20.387266,19.915688,19.817598,19.383747,18.983849,18.621677,17.927513,17.022083,16.248695,15.188588,13.909668,12.970284,13.43809,14.252977,14.811326,14.886778,14.667966,13.962485,13.837989,14.27184,15.150862,16.237377,17.074902,17.53516,17.904879,18.41041,19.217752,13.336229,13.011784,12.423254,11.823407,11.589504,12.2119875,12.0724,11.981857,12.491161,13.358865,13.536179,14.124708,14.48688,14.151116,13.400364,13.2607765,13.913441,14.347293,15.460217,17.033401,17.712475,15.912932,14.558559,13.943622,14.094527,14.777372,15.490398,16.373192,16.403374,15.290449,13.449409,12.261031,11.917723,11.604594,11.027383,10.427535,9.891823,10.091772,10.18986,9.578695,7.914967,7.7037,7.277394,6.8699503,6.5945487,6.477597,6.858632,7.1906233,7.484888,7.7602897,8.043237,7.413208,6.417235,5.5759397,5.0666356,4.7233267,4.5761943,4.3913355,4.183841,4.1800685,4.8327327,5.1081343,5.2628117,5.0741806,4.617693,4.285702,4.425289,4.745962,5.1760416,5.4740787,5.2175403,5.3194013,4.859141,4.425289,4.221567,4.0593443,4.29702,4.5196047,4.7006907,4.9044123,5.292993,5.3194013,5.6023483,5.9984736,6.458734,7.0359454,6.72659,6.3719635,6.515323,7.032173,7.1302614,6.828451,6.6813188,6.462507,6.1606965,5.9720654,5.594803,5.323174,5.270357,5.492942,6.013564,7.152897,7.6584287,7.967784,8.239413,8.371455,8.179051,7.986647,7.911195,8.07719,8.601585,8.835487,9.435335,10.631257,12.038446,12.623203,12.559069,12.098808,11.981857,12.396846,12.992921,12.709973,11.283921,9.789962,8.869441,8.703445,8.024373,7.7716074,7.8244243,8.013056,8.096053,8.495952,8.439363,8.031919,7.356619,6.485142,6.3229194,6.115425,5.9230213,5.8626595,6.089017,6.2436943,6.2663302,6.0324273,5.692891,5.670255,5.832478,5.9532022,6.017337,5.9607477,5.666483,5.2779026,4.8365054,4.636556,4.708236,4.7874613,4.678055,4.610148,4.666737,4.8629136,5.1571784,4.8968673,4.7648253,4.6856003,4.52715,4.06689,3.361409,2.7087448,2.1994405,1.8749946,1.7354075,1.5165952,1.3732355,1.2940104,1.2449663,1.1732863,1.0336993,0.8639311,0.7582976,0.73188925,0.70170826,0.7130261,0.8601585,0.9280658,0.88279426,0.8526133,0.7582976,0.66775465,0.6413463,0.60362,0.33576363,0.211267,0.18485862,0.17731337,0.14713238,0.09808825,0.071679875,0.071679875,0.0754525,0.071679875,0.08677038,0.0754525,0.06790725,0.06413463,0.06790725,0.090543,0.120724,0.116951376,0.10940613,0.10940613,0.090543,0.090543,0.13204187,0.14335975,0.116951376,0.13958712,0.15845025,0.18863125,0.17731337,0.14335975,0.14713238,0.12826926,0.124496624,0.124496624,0.13204187,0.150905,0.124496624,0.10940613,0.08299775,0.056589376,0.06790725,0.07922512,0.07922512,0.071679875,0.05281675,0.041498873,0.094315626,0.06790725,0.0452715,0.06413463,0.10940613,0.16976812,0.23767537,0.26408374,0.24522063,0.241448,0.271629,0.38480774,0.41498876,0.4376245,0.77338815,0.69793564,0.66775465,0.6413463,0.63002837,0.65643674,0.7922512,1.0902886,1.4713237,1.7467253,1.6373192,1.6637276,1.358145,1.1129243,1.116697,1.3430545,1.086516,1.2751472,1.2449663,0.86770374,0.5470306,0.59607476,0.814887,1.1619685,1.3505998,0.8526133,1.2487389,2.5804756,4.5761943,6.5002327,7.1679873,7.492433,5.59103,3.048281,1.4071891,2.1315331,3.5387223,5.2250857,5.764571,5.3948536,6.0248823,5.5382137,6.56814,8.379,9.318384,6.8397694,11.649866,13.65313,11.69891,8.677037,11.521597,17.40689,17.003222,12.408164,6.470052,2.7728794,6.40969,8.039464,8.050782,7.394345,7.5829763,3.9386206,3.2670932,3.0935526,2.6182017,2.704972,1.8485862,1.6976813,1.3958713,0.8337501,0.6488915,0.6526641,0.4678055,0.33576363,0.32821837,0.362172,0.58475685,0.935611,0.8526133,0.422534,0.3772625,0.5357128,1.0148361,1.7240896,2.3993895,2.6182017,2.3993895,3.5424948,5.13077,6.3644185,6.537959,5.138315,6.436098,6.790725,5.383536,4.255521,7.854605,7.967784,6.9869013,6.5341864,7.443389,8.326183,8.707218,9.239159,9.748463,9.220296,8.854351,9.669238,9.812597,9.325929,10.148361,9.986138,10.26154,10.782163,10.86516,9.333474,9.235386,8.892077,8.469543,7.986647,7.3151197,6.5530496,7.3075747,7.5037513,6.8473144,6.828451,6.221059,6.6586833,7.7602897,8.714764,8.29223,8.514814,8.899622,9.982366,11.578186,12.800517,11.514051,10.899114,9.291975,6.3153744,2.8822856,2.444661,3.4972234,5.613666,7.4735703,6.8774953,6.9680386,5.926794,5.7419353,7.5301595,11.521597,7.122716,4.9723196,4.146115,4.406426,6.221059,4.014073,2.9615107,2.584248,2.4182527,2.033445,1.8334957,3.240685,3.9725742,3.5500402,3.2670932,4.3121104,3.7198083,3.097325,2.686109,1.3656902,3.0746894,3.4481792,5.142088,9.012801,14.132254,8.16396,9.26934,12.1101265,14.34352,16.622187,17.836971,18.002966,17.527617,14.50197,4.719554,4.4139714,8.507269,9.26934,5.8664317,4.3724723,6.8774953,4.9647746,4.9534564,8.771353,13.977575,7.726336,5.6325293,7.654656,10.853842,9.386291,6.2436943,5.7494807,7.888559,10.155907,7.5565677,7.0774446,7.7716074,9.348565,11.174516,12.298758,11.631002,9.488152,9.303293,11.189606,11.921495,12.494934,12.996693,12.393073,11.370691,12.31762,9.967276,8.458225,8.14887,9.092027,11.02361,15.07541,19.496925,18.440592,12.958967,11.02361,12.777881,11.144334,10.265312,10.555805,8.714764,10.401127,9.695646,11.706455,14.898096,11.091517,8.499724,7.3868,8.152642,9.005256,5.9720654,4.168751,3.6254926,4.38379,6.990674,12.479843,8.790216,8.748717,8.967529,8.726082,9.989911,9.107117,9.159933,9.65792,10.016319,9.567377,9.914458,10.657665,11.378237,11.691365,11.219787,10.989656,11.227332,12.67602,15.01882,16.882498,19.719511,20.65135,19.900597,17.727566,14.445381,13.585222,13.7700815,14.400109,15.705438,18.757492,17.282394,16.158154,15.701665,15.214996,13.004238,13.004238,12.366665,11.00852,9.276885,7.964011,10.891568,11.827179,10.827434,8.8618965,7.8319697,9.631512,9.258021,8.458225,8.59404,10.63503,10.514306,11.351829,11.521597,10.884023,10.782163,10.680302,11.389555,10.876478,9.186342,8.465771,8.544995,8.446907,8.89585,9.465516,8.605357,8.16396,8.16396,7.964011,7.598067,7.7829256,7.2358947,6.79827,7.6697464,9.012801,7.9715567,7.7829256,8.552541,11.691365,15.294222,14.139798,13.72481,14.498198,14.524607,13.532406,12.921241,14.460471,14.611377,15.520579,16.976812,16.41092,15.433809,15.577168,15.848798,15.577168,14.381247,13.419228,11.566868,9.567377,7.745199,5.994701,6.1531515,6.319147,6.0701537,5.5193505,5.300538,5.2099953,5.3609,5.43258,5.342037,5.247721,4.930821,4.5950575,4.8365054,5.270357,4.515832,4.3422914,4.5120597,4.7912335,5.0515447,5.243949,5.451443,6.2021956,7.2585306,8.428044,9.552286,10.63503,10.846297,11.09529,11.631002,12.042219,12.404391,12.921241,13.615403,14.7321005,16.77309,17.312576,16.467508,16.376965,17.437073,18.263277,17.003222,16.056292,15.645076,15.803526,16.376965,16.565596,15.645076,14.905642,14.984866,15.852571,15.924251,15.218769,14.962231,15.652621,17.067356,17.4333,17.976559,18.489635,19.240387,20.979568,21.145563,20.33822,18.817854,17.497435,17.957695,18.153872,18.059555,18.176508,18.531134,18.678267,18.19537,18.715992,19.364883,19.56106,18.991394,18.384,18.16519,18.059555,17.91997,17.72002,17.04472,16.705183,15.912932,14.649103,13.6682205,13.370183,13.758763,14.060574,13.920986,13.407909,13.204187,13.340002,13.43809,13.65313,14.698147,16.16947,17.003222,17.587978,18.0671,18.368912,14.037937,14.034165,13.815352,12.728837,11.329193,11.385782,11.000975,10.423763,10.47658,11.1631975,11.68382,12.687338,13.513543,13.479589,12.883514,13.008011,13.072145,12.902377,13.268322,14.109617,14.57365,13.849306,13.788944,14.211478,14.93205,15.739391,16.293968,16.754227,16.403374,15.260268,14.079436,12.860879,12.370438,12.147853,11.902632,11.52537,11.129244,10.9594755,10.56335,9.623966,7.9413757,8.073418,8.390318,8.627994,8.582722,8.130007,8.118689,8.058327,7.911195,7.748972,7.7338815,6.7341356,5.564622,4.821415,4.5724216,4.353609,4.357382,4.293247,4.1310244,4.0103,4.2630663,4.504514,4.689373,4.5837393,4.247976,4.032936,4.191386,4.3649273,4.6629643,4.961002,4.8968673,4.9534564,4.689373,4.3649273,4.1083884,3.9386206,4.2064767,4.5799665,4.8365054,4.9685473,5.172269,5.5193505,5.8588867,6.2436943,6.6020937,6.7341356,6.719045,6.900131,7.4509344,8.07719,7.9941926,7.8017883,7.7640624,7.605612,7.1868505,6.485142,6.2851934,5.87775,5.726845,6.047518,6.7944975,8.031919,8.733627,9.084481,9.250477,9.397609,9.537196,9.4127,9.435335,9.695646,9.989911,9.933322,10.1294985,10.872705,11.940358,12.593022,12.3289385,11.680047,11.465008,11.962994,12.909923,12.626976,11.823407,10.9594755,10.325675,10.035183,9.529651,9.348565,9.175024,8.89585,8.620448,8.605357,8.439363,7.9413757,7.122716,6.1908774,5.983383,6.089017,6.221059,6.3153744,6.515323,6.398372,6.2097406,5.824933,5.4476705,5.6287565,5.8928404,6.1833324,6.360646,6.349328,6.149379,5.4891696,5.1345425,5.1760416,5.587258,6.2021956,6.089017,5.7909794,5.5570765,5.523123,5.7192993,5.353355,5.111907,5.0439997,4.991183,4.587512,3.9273026,3.2105038,2.5502944,2.0485353,1.7957695,1.5958204,1.4373702,1.3241913,1.2562841,1.20724,1.056335,0.935611,0.83752275,0.7696155,0.7582976,0.7469798,0.8563859,0.98465514,1.0601076,1.0374719,0.91297525,0.8337501,0.8563859,0.8601585,0.55080324,0.35462674,0.26031113,0.23390275,0.23013012,0.1659955,0.116951376,0.10186087,0.090543,0.08299775,0.07922512,0.08299775,0.06790725,0.06790725,0.08299775,0.090543,0.1056335,0.10186087,0.1056335,0.120724,0.10940613,0.1056335,0.14335975,0.14713238,0.120724,0.12826926,0.116951376,0.150905,0.15845025,0.13958712,0.1659955,0.14713238,0.1358145,0.120724,0.11317875,0.1358145,0.11317875,0.09808825,0.07922512,0.060362,0.06790725,0.07922512,0.10186087,0.1056335,0.090543,0.071679875,0.120724,0.08299775,0.056589376,0.08677038,0.16976812,0.23390275,0.29049212,0.28294688,0.24522063,0.29049212,0.362172,0.41876137,0.392353,0.33953625,0.45648763,0.52439487,0.7092535,0.73566186,0.5998474,0.5885295,0.6828451,0.84884065,1.1280149,1.4411428,1.5731846,1.2110126,1.1242423,1.1581959,1.2298758,1.3430545,0.9997456,1.0412445,1.0601076,0.8639311,0.49044126,0.56212115,0.76207024,1.0638802,1.2223305,0.784706,1.6222287,2.9803739,4.7836885,6.439871,6.8397694,6.881268,4.949684,2.9237845,1.8561316,1.9693103,2.987919,4.3913355,5.451443,5.87775,5.8098426,5.304311,9.265567,13.985121,16.146835,12.845788,16.35433,19.081938,17.1164,11.234878,6.888813,13.766309,12.687338,7.888559,3.4632697,3.3312278,9.861642,9.997457,7.8696957,6.0739264,5.6853456,3.3651814,3.4330888,4.1989317,4.6818275,4.6026025,2.9464202,3.0445085,2.3767538,0.86770374,0.8639311,0.72811663,0.73566186,0.6488915,0.5772116,0.935611,1.0827434,1.2600567,0.9922004,0.44894236,0.4678055,1.0223814,1.4034165,1.8599042,2.3390274,2.4974778,2.2560298,3.6783094,5.617439,6.9680386,6.670001,5.534441,6.5266414,6.9152217,6.0701537,5.485397,8.843033,8.805306,7.726336,7.3717093,8.918486,9.691874,9.5183325,9.771099,10.393582,9.910686,8.461998,8.975075,9.024119,8.409182,9.163706,9.420244,9.548513,10.284176,10.963248,9.525878,9.473062,9.280658,8.741172,7.9451485,7.284939,6.507778,6.802043,6.9491754,6.507778,5.8173876,5.3986263,5.3571277,5.824933,6.511551,6.700182,7.4169807,8.050782,9.22784,10.989656,12.811834,11.947904,11.510279,9.646602,6.255012,2.9728284,3.6594462,4.3686996,6.300284,7.7942433,4.353609,5.847569,5.4740787,5.8588867,7.9791017,11.1631975,6.8661776,4.5497856,3.7273536,4.1272516,5.674028,3.006782,2.5502944,2.6936543,2.686109,2.6483827,2.8521044,3.6292653,3.9122121,3.3576362,2.3880715,4.708236,4.08198,3.8178966,4.142342,2.1843498,3.3123648,2.8634224,3.3576362,6.3945994,12.642066,10.676529,10.650121,11.548005,13.162688,16.086473,17.89356,19.130981,19.198889,15.656394,4.2291126,6.5756855,10.197406,9.81637,5.5495315,2.8785129,8.284684,9.186342,7.805561,6.7756343,9.137298,5.96452,4.991183,6.7831798,9.186342,7.3415284,6.1720147,6.5568223,7.303802,7.4509344,6.2851934,6.507778,7.333983,9.35611,11.672502,11.883769,10.306811,9.688101,9.533423,9.937095,11.5857315,12.872196,13.27964,13.011784,12.294985,11.389555,9.748463,8.145098,7.960239,9.374973,11.370691,14.351066,18.919714,17.810562,12.151625,11.449917,13.905896,12.00072,10.872705,11.117926,8.812852,9.635284,9.748463,10.280403,11.223559,11.423509,7.7640624,6.9567204,7.9526935,8.669493,6.0022464,6.511551,4.8402777,4.255521,5.9682927,9.114662,8.967529,6.579458,5.2628117,6.0362,7.6131573,8.118689,8.216777,8.175279,7.7716074,6.307829,7.1076255,8.303548,9.639057,10.801025,11.423509,10.95193,11.329193,12.940104,15.396083,17.516298,20.915434,21.119154,19.236614,16.561823,14.603831,15.814844,15.384765,14.117163,12.759018,12.004493,8.314865,11.332966,12.774108,10.574668,8.89585,8.567632,8.118689,7.8923316,7.635793,6.530414,8.118689,9.386291,9.6201935,8.710991,7.141579,9.280658,9.593785,8.975075,8.688355,10.340765,10.287949,10.853842,11.249968,11.148107,10.691619,9.831461,11.046246,11.016065,9.484379,9.258021,8.477088,8.209232,8.741172,9.5183325,9.159933,8.846806,8.944894,8.5563135,7.7942433,7.7829256,7.4094353,6.5002327,7.4471617,9.386291,8.190369,7.515069,8.786444,11.208468,13.340002,13.0646,12.54775,13.023102,12.528888,11.415963,12.359119,11.740409,13.306048,15.109364,15.935568,15.339493,14.694374,14.494425,14.452927,14.068119,12.626976,11.7555,10.167224,8.45068,6.8435416,5.2062225,4.98741,5.100589,5.1081343,4.961002,4.9949555,5.1873593,5.311856,5.3458095,5.3458095,5.4363527,4.247976,3.9499383,4.3196554,4.82896,4.644101,3.983892,4.0178456,4.4139714,5.0175915,5.8513412,5.956975,6.5002327,7.7112455,9.352338,10.725573,11.3669195,11.604594,11.925267,12.377983,12.54775,13.109872,13.751218,14.452927,15.531898,17.644567,18.384,17.799244,17.855835,18.587723,18.104828,16.62973,16.324148,16.524097,17.014538,18.025602,18.218006,16.976812,15.99593,15.848798,16.007248,15.878979,15.196134,14.434063,14.222796,15.339493,15.83748,17.421982,19.002712,20.055275,20.594759,21.23988,20.492899,18.817854,17.350302,17.908651,17.765291,17.229578,17.399347,18.229324,18.557543,18.089737,18.33873,18.923487,19.304522,18.802763,17.45971,16.856089,16.765545,16.890041,16.874952,16.693865,16.603323,16.048746,14.977322,13.834216,13.079691,13.170234,13.317367,13.162688,12.740154,12.73261,12.974057,12.958967,12.830698,13.358865,14.667966,15.769572,16.746683,17.440845,17.429527,13.736128,14.2944765,14.875461,14.02662,12.140307,11.41219,10.8576145,10.642575,10.284176,9.963503,10.533169,11.363147,12.276122,12.642066,12.449662,12.31762,11.944131,12.261031,12.808062,13.12119,12.728837,13.041965,13.977575,14.705692,15.056546,15.524352,15.652621,15.501716,14.954685,14.362384,14.532151,13.860624,13.430545,13.336229,13.381501,13.057055,12.189351,11.355601,10.736891,10.167224,9.129752,9.005256,9.650374,10.125726,9.952185,9.103344,8.371455,7.699928,6.7077274,5.564622,4.991183,4.6818275,4.5007415,4.3347464,4.142342,3.953711,4.214022,4.2706113,4.266839,4.217795,4.0216184,4.025391,4.1083884,4.274384,4.534695,4.90064,4.8365054,4.772371,4.647874,4.4931965,4.4215164,4.447925,4.564876,4.5233774,4.3724723,4.4894238,4.5422406,4.5535583,4.617693,4.7572803,4.9044123,5.9192486,6.3116016,6.5568223,6.8246784,6.9869013,7.4773426,8.0206,8.439363,8.635539,8.560086,8.790216,8.748717,8.507269,7.9791017,6.937857,7.1679873,6.9567204,6.741681,6.8737226,7.624475,8.52236,9.382519,10.095545,10.555805,10.680302,11.114153,11.136789,11.065109,10.985884,10.7557535,10.79348,11.031156,11.3971,11.812089,12.181807,11.853588,11.363147,10.819888,10.657665,11.619685,12.174261,12.66093,12.932558,12.849561,12.291212,11.664956,11.034928,10.370946,9.563604,8.428044,8.062099,7.8017883,7.4169807,6.94163,6.6813188,6.5530496,6.5832305,6.8058157,7.066127,6.9982195,6.63982,6.48137,6.398372,6.3342376,6.2889657,6.2323766,6.6247296,7.020855,7.175533,7.0359454,6.356873,6.119198,6.3116016,6.851087,7.5905213,7.3188925,6.730363,6.2323766,5.983383,5.8664317,5.4891696,5.3344917,5.2967653,5.2288585,4.938366,4.4705606,3.7160356,2.8898308,2.1881225,1.7957695,1.5958204,1.4222796,1.2789198,1.1846043,1.177059,1.0601076,1.0789708,1.0223814,0.87902164,0.8186596,0.6752999,0.70170826,0.8639311,1.0601076,1.1091517,1.0714256,1.026154,1.0450171,1.0714256,0.90920264,0.6413463,0.43385187,0.34330887,0.33576363,0.2678564,0.19994913,0.15845025,0.12826926,0.1056335,0.09808825,0.120724,0.120724,0.124496624,0.12826926,0.10940613,0.10186087,0.08677038,0.090543,0.10940613,0.12826926,0.116951376,0.11317875,0.124496624,0.1358145,0.1358145,0.120724,0.13204187,0.14713238,0.16222288,0.1659955,0.14713238,0.12826926,0.11317875,0.10186087,0.09808825,0.08677038,0.090543,0.08677038,0.08299775,0.094315626,0.10186087,0.13204187,0.15467763,0.150905,0.124496624,0.11317875,0.1056335,0.10940613,0.150905,0.2565385,0.32821837,0.3169005,0.2565385,0.21881226,0.3055826,0.47535074,0.44894236,0.35085413,0.29049212,0.362172,0.55457586,0.83752275,0.84884065,0.5772116,0.35839936,0.30935526,0.3734899,0.43007925,0.6752999,1.6222287,0.98465514,1.1846043,1.2336484,0.9997456,1.1996948,0.7582976,0.6790725,0.7696155,0.7922512,0.4640329,0.5394854,0.59230214,0.65643674,0.73188925,0.784706,2.2673476,2.8256962,3.7801702,5.0666356,5.243949,4.7950063,3.3953626,2.5087957,2.3126192,1.6750455,2.1692593,3.7084904,5.2288585,5.855114,4.889322,6.3153744,13.671993,19.447882,21.130472,21.202152,21.017294,20.274086,20.02132,17.712475,7.201941,7.424526,6.549277,4.6931453,3.289729,5.070408,10.570895,9.869187,7.303802,5.1081343,3.4217708,3.3840446,4.293247,5.96452,7.5716586,7.624475,4.2819295,4.123479,3.3764994,1.5920477,1.6109109,1.2487389,1.3505998,1.1883769,0.90920264,1.5354583,1.4222796,1.2562841,0.94692886,0.67152727,0.87147635,1.8863125,1.8372684,1.5958204,1.6033657,1.8448136,2.4559789,4.447925,6.5756855,7.6848373,6.719045,6.2663302,7.020855,7.5792036,7.383027,6.7077274,8.858124,9.344792,8.786444,8.469543,10.325675,10.310584,10.186088,10.26154,10.427535,10.155907,7.91874,8.209232,8.318638,7.748972,8.201687,8.726082,8.820397,9.344792,9.955957,9.114662,9.288202,9.6201935,9.250477,8.254503,7.6697464,6.63982,6.1531515,6.1305156,5.9607477,4.4894238,4.3347464,4.315883,4.4894238,4.7950063,5.0553174,6.33801,7.462252,8.582722,9.963503,11.959221,12.208215,11.672502,9.039209,5.534441,4.9232755,5.613666,6.40969,6.2323766,5.243949,4.8440504,6.3719635,7.8244243,7.911195,6.6813188,5.534441,4.908185,6.360646,6.2399216,3.8971217,1.6863633,2.323937,3.31991,3.8669407,4.055572,4.90064,3.9650288,2.7200627,2.837014,3.4783602,1.2789198,3.3727267,2.6332922,2.9803739,4.3875628,2.886058,3.8858037,4.3083377,3.8141239,3.983892,8.314865,10.397354,7.1868505,3.7763977,2.9954643,5.3986263,7.8508325,9.578695,10.084227,9.103344,6.6134114,11.721546,14.25675,11.714001,5.983383,3.350091,12.645839,18.878216,17.47857,9.7220545,2.7389257,3.4557245,4.719554,5.692891,5.9720654,5.594803,6.722818,8.835487,9.635284,8.582722,6.862405,5.9909286,6.258785,8.439363,10.895341,9.559832,7.5037513,9.129752,10.20495,9.752235,10.016319,12.151625,12.359119,12.359119,12.332711,10.917976,8.99771,8.035691,8.499724,10.110635,11.834724,13.562587,16.908905,16.607096,12.487389,9.491924,12.268577,12.098808,11.996947,12.2270775,10.299266,7.745199,9.64283,10.253995,9.039209,10.646348,8.099826,7.032173,6.3116016,5.7570257,6.145606,9.786189,7.122716,4.195159,3.519859,4.1197066,9.454198,6.307829,4.183841,6.0550632,8.3525915,8.386545,8.194141,8.43559,8.707218,7.533932,6.7944975,6.881268,7.175533,7.9451485,10.374719,11.668729,13.317367,14.830189,16.192106,17.867151,20.387266,20.043957,18.617905,17.244669,16.418465,17.508753,16.161926,13.864397,11.102836,7.352846,3.7047176,8.884532,9.129752,3.350091,3.1199608,2.8634224,4.2328854,7.194396,9.857869,8.461998,5.172269,4.610148,5.617439,7.043491,7.756517,7.9451485,9.110889,9.7069645,9.378746,8.952439,10.435081,10.834979,10.77839,10.729345,10.982111,9.544742,10.506761,10.725573,9.812597,10.133271,7.9489207,7.8432875,8.605357,9.382519,9.688101,9.578695,9.22784,8.66572,8.107371,7.9451485,7.756517,6.5002327,6.990674,8.4544525,6.5266414,6.470052,9.906913,11.314102,10.510533,12.630749,11.446144,11.691365,10.838752,9.835234,13.109872,7.2887115,11.480098,15.222542,15.109364,14.811326,14.837734,14.215251,13.343775,12.321393,10.948157,9.793735,8.511042,7.2094865,5.956975,4.779916,4.6214657,4.696918,4.67051,4.436607,4.13857,4.776143,5.3684454,5.4250345,5.093044,5.149633,4.0517993,4.134797,4.346064,4.323428,4.3686996,3.7613072,3.6443558,3.9461658,4.7044635,6.0701537,6.33801,7.0548086,8.213005,9.439108,9.993684,10.250222,10.804798,11.544232,12.336484,13.008011,13.456953,14.086982,14.758509,15.603577,16.98813,18.674494,19.240387,19.17248,18.478317,16.690092,15.905387,16.290195,17.006994,17.810562,19.063074,19.104572,18.1086,17.501207,17.414436,16.667458,15.437581,15.184815,14.603831,13.645585,13.517315,14.950912,17.184307,19.289433,20.209951,18.742401,19.349794,18.278368,17.082445,16.678776,17.327667,17.37671,16.780636,16.856089,17.621931,17.795471,17.769064,18.104828,18.780127,19.398838,19.168707,17.184307,15.543215,15.184815,15.829934,15.984612,16.4826,16.260014,15.792209,15.086727,13.679539,12.928786,12.898605,12.974057,12.909923,12.853333,12.596795,12.781653,12.928786,12.81938,12.525115,12.894833,13.86817,15.116908,16.146835,16.309057,13.626721,14.320885,13.543724,12.242168,11.2801485,11.41219,11.7555,11.766817,11.170743,10.27663,10.008774,9.522105,9.922004,10.54826,11.133017,11.778135,12.15917,13.068373,13.920986,13.951167,12.193124,12.434572,12.936331,13.041965,12.740154,12.679792,12.253486,11.917723,11.7026825,11.796998,12.543978,12.261031,12.083718,12.106354,12.276122,12.37421,10.518079,10.008774,10.144588,10.167224,9.276885,8.99771,9.0807085,8.6732645,7.5905213,6.3342376,5.9418845,5.7909794,5.613666,5.3080835,4.927048,4.4630156,4.3309736,4.3309736,4.4441524,4.821415,5.2364035,5.304311,5.2062225,5.0854983,5.036454,5.1571784,5.3986263,5.594803,5.692891,5.7683434,5.6815734,5.6513925,5.572167,5.4476705,5.3873086,5.2137675,5.3382645,5.4891696,5.7079816,6.330465,6.013564,5.406172,4.8553686,4.561104,4.561104,5.292993,5.8437963,6.428553,7.145352,7.964011,8.514814,8.688355,8.790216,9.001483,9.352338,9.42779,9.473062,9.2844305,8.816625,8.194141,7.54525,7.356619,7.303802,7.3075747,7.5527954,8.273367,9.808825,11.234878,12.0724,12.268577,12.536433,12.759018,12.66093,12.223305,11.672502,11.661184,11.91395,12.189351,12.306303,12.147853,11.91395,12.23085,12.1101265,11.778135,12.694883,13.502225,14.143571,14.056801,13.343775,12.755245,12.449662,11.54046,10.540714,9.5032425,8.024373,7.756517,7.5716586,7.54525,7.6697464,7.828197,7.435844,6.907676,6.590776,6.5455046,6.5455046,6.6549106,7.039718,7.2660756,7.1302614,6.6662283,6.5228686,7.2094865,8.122461,8.661947,8.209232,7.2924843,7.322665,7.594294,7.624475,7.1264887,6.700182,6.4738245,6.1908774,5.8400235,5.6476197,5.7192993,5.802297,5.7079816,5.4250345,5.0968165,4.949684,4.447925,3.6594462,2.8445592,2.4408884,2.123988,1.7240896,1.3468271,1.0676528,0.94692886,0.83752275,0.83752275,0.8111144,0.7432071,0.73188925,0.55080324,0.5319401,0.76207024,1.1091517,1.2223305,1.3166461,1.3053282,1.4109617,1.5316857,1.2525115,0.8865669,0.6375736,0.49044126,0.42630664,0.42630664,0.32821837,0.29426476,0.24899325,0.1961765,0.24522063,0.3169005,0.29803738,0.26408374,0.23013012,0.18485862,0.1358145,0.11317875,0.1056335,0.1056335,0.090543,0.07922512,0.08677038,0.10940613,0.1358145,0.1358145,0.150905,0.150905,0.1659955,0.1659955,0.1056335,0.094315626,0.10186087,0.094315626,0.071679875,0.060362,0.060362,0.07922512,0.09808825,0.120724,0.1659955,0.15467763,0.14335975,0.13204187,0.1358145,0.19994913,0.1358145,0.20372175,0.28294688,0.3169005,0.3055826,0.3169005,0.32067314,0.31312788,0.3169005,0.36594462,0.58475685,0.47535074,0.32444575,0.26408374,0.29049212,0.422534,0.48666862,0.4678055,0.36971724,0.19994913,0.26031113,0.35839936,0.392353,0.48666862,0.97710985,1.20724,0.7432071,0.5998474,0.88279426,0.80734175,0.663982,0.73566186,0.8224323,0.7582976,0.42630664,0.6111652,0.6451189,0.60362,0.5885295,0.7469798,1.9579924,1.7354075,1.7014539,2.1051247,1.8636768,2.071171,2.3390274,2.384299,2.1013522,1.6033657,2.505023,3.8405323,4.5120597,4.376245,4.2404304,6.9755836,13.702174,18.780127,19.76101,17.380484,14.25675,12.083718,11.4838705,11.378237,8.971302,3.9310753,3.429316,4.146115,4.719554,5.7683434,8.4544525,8.786444,7.5527954,5.5080323,3.3727267,4.6554193,5.6061206,7.356619,9.307066,9.125979,4.878004,3.9989824,3.742444,3.31991,3.904667,2.7691069,2.5691576,1.9844007,1.0450171,1.1431054,1.1204696,0.6488915,0.3961256,0.5998474,1.0525624,1.6033657,1.6373192,1.6335466,1.7844516,2.0296721,2.5804756,4.666737,7.3453007,8.967529,7.17176,7.4018903,7.865923,8.047009,7.9300575,7.964011,10.272858,10.948157,10.582213,10.152134,11.031156,9.397609,10.076681,10.868933,10.816116,10.193633,8.288457,7.8395147,7.752744,7.6508837,7.858378,8.382772,8.367682,8.8618965,9.654147,9.261794,8.601585,9.235386,9.480607,8.963757,8.620448,6.9869013,5.945657,5.4740787,5.1232247,4.014073,3.8178966,4.032936,4.2404304,4.4101987,4.8968673,6.4738245,7.91874,8.914713,9.639057,10.789707,11.936585,10.216269,7.61693,6.009792,7.1566696,7.9262853,7.1000805,5.9984736,6.138061,9.261794,14.754736,11.276376,8.601585,8.412953,4.2894745,2.384299,6.221059,7.273621,3.9914372,1.7693611,2.3314822,2.5917933,2.8219235,3.9122121,7.352846,3.0709167,2.0636258,2.6785638,2.9992368,0.83752275,4.4177437,5.6287565,4.508287,2.1654868,0.8224323,5.621211,5.9682927,3.9612563,1.659955,1.0978339,1.9051756,1.5279131,1.1996948,1.9202662,4.4705606,8.047009,9.125979,8.009283,7.6131573,13.472044,17.391802,15.24895,11.5857315,8.722309,6.7454534,20.417446,32.89729,34.172436,22.77911,5.8136153,4.957229,6.2927384,5.5193505,3.410453,5.8136153,6.043745,7.624475,7.654656,6.047518,5.5080323,4.666737,5.8098426,7.032173,7.364164,6.790725,6.1305156,7.5301595,8.013056,7.5263867,8.941121,9.808825,9.639057,9.005256,8.986393,11.185833,8.926031,7.8017883,9.001483,11.725319,13.215506,12.479843,12.445889,13.079691,13.630494,12.604341,11.555551,10.038955,9.280658,9.639057,10.604849,7.9451485,9.110889,10.970794,11.427281,9.416472,9.035437,8.171506,7.0246277,5.9003854,5.2175403,6.085244,8.031919,8.201687,6.779407,6.9869013,3.2784111,2.2598023,1.9466745,1.9089483,3.2520027,1.358145,2.1579416,5.3080835,9.7069645,13.502225,5.6061206,4.044254,4.304565,4.708236,6.3945994,5.783434,7.643338,10.103089,11.631002,11.031156,10.435081,11.54046,14.177525,17.040947,17.701157,15.98084,14.441608,13.573905,11.84227,5.692891,4.459243,2.5502944,2.7200627,4.938366,6.379509,5.987156,7.1906233,8.646856,9.548513,9.597558,11.551778,11.993175,9.14107,5.243949,6.560595,7.7942433,7.835742,9.480607,11.348056,7.9036493,10.370946,11.434827,10.891568,9.884277,10.910432,9.971047,10.367173,10.18986,9.484379,10.253995,7.3000293,7.220804,8.360137,9.442881,9.552286,9.748463,9.4127,9.0957985,9.031664,9.156161,8.2507305,6.7341356,5.624984,4.779916,2.9011486,5.9494295,9.122208,10.823661,10.789707,10.054046,8.420499,12.525115,14.045483,13.257004,19.04421,8.726082,10.186088,13.634267,14.675511,14.298248,13.943622,12.728837,11.563096,10.510533,8.790216,8.031919,7.496206,6.828451,5.7909794,4.2404304,3.7537618,3.942393,4.4139714,4.7836885,4.7006907,5.0062733,5.191132,5.674028,6.066381,5.1873593,5.2137675,5.564622,5.342037,4.515832,3.9688015,3.3689542,3.2105038,3.3463185,3.7273536,4.4101987,4.9232755,5.873977,7.364164,8.967529,9.752235,10.299266,10.502988,10.770844,11.332966,12.238396,12.83447,13.837989,15.203679,16.682549,17.80679,19.002712,18.523588,17.554024,16.810818,16.55428,15.652621,15.297995,15.633758,16.546734,17.670975,18.670721,18.708447,18.43682,18.119919,17.670975,17.13149,16.795727,15.818617,14.381247,13.687083,15.00373,15.720529,16.244923,16.848543,17.655886,18.606586,17.542706,16.233604,15.679029,16.143063,16.58446,16.791954,17.003222,17.097536,16.648594,16.67123,16.724047,16.980585,17.301258,17.225805,15.897841,14.50197,14.539697,15.803526,16.388283,16.765545,16.74291,16.705183,16.437326,15.105591,13.849306,13.306048,13.087236,12.940104,12.755245,12.049765,12.257258,12.494934,12.366665,11.962994,11.668729,12.155397,13.091009,13.966258,14.0983,12.321393,14.226569,14.403882,13.973803,13.483362,12.913695,11.92904,11.570641,11.242422,10.7218,10.167224,10.020092,10.054046,10.182315,10.446399,10.985884,11.717773,12.419481,13.124963,13.336229,12.045992,12.162943,12.491161,12.479843,12.012038,11.434827,10.33322,10.465261,10.887795,11.216014,11.627231,11.563096,11.69891,11.778135,11.59705,11.031156,10.065364,9.646602,9.469289,9.178797,8.375228,7.0887623,6.48137,6.1041074,5.8136153,5.80607,5.7004366,5.9117036,6.149379,6.2625575,6.2361493,5.956975,5.6325293,5.349582,5.20245,5.2967653,5.4703064,5.59103,5.5004873,5.2854476,5.304311,5.492942,5.7381625,5.8173876,5.828706,6.19465,6.8699503,6.9567204,6.6020937,6.047518,5.6551647,5.3571277,5.270357,5.4288073,5.8136153,6.368191,6.4436436,6.7869525,7.201941,7.515069,7.564113,7.7225633,7.9791017,8.345046,8.748717,9.039209,9.374973,9.778644,10.231359,10.672756,11.027383,11.431054,11.449917,10.895341,9.895596,8.903395,7.914967,7.7037,7.865923,8.2507305,8.98262,10.287949,11.404645,12.106354,12.332711,12.193124,12.423254,12.536433,12.359119,11.981857,11.732863,11.838497,12.200669,12.543978,12.664702,12.427027,12.351574,12.781653,12.966512,12.958967,13.611631,14.290704,14.8339615,15.067864,14.822643,13.917213,13.132507,12.351574,11.7026825,11.065109,10.076681,9.623966,9.514561,9.49947,9.371201,8.975075,8.2507305,7.598067,7.1378064,6.952948,7.069899,7.250985,7.3868,7.707473,8.156415,8.412953,8.688355,9.201432,9.612649,9.695646,9.333474,9.167479,8.892077,8.707218,8.518587,7.9300575,7.84706,7.567886,7.1868505,6.820906,6.587003,6.5530496,6.356873,6.013564,5.5683947,5.1345425,5.0854983,4.708236,4.115934,3.4632697,2.9426475,2.516341,2.0900342,1.6373192,1.2261031,0.995973,0.8563859,0.8337501,0.84884065,0.8299775,0.7205714,0.6752999,0.7130261,0.84129536,1.0525624,1.3166461,1.4750963,1.5203679,1.5618668,1.5580941,1.3355093,1.1053791,0.9808825,0.8978847,0.8224323,0.7432071,0.6375736,0.5583485,0.45648763,0.392353,0.5357128,0.543258,0.38858038,0.271629,0.23767537,0.21881226,0.181086,0.17731337,0.181086,0.15845025,0.07922512,0.049044125,0.056589376,0.08677038,0.10940613,0.10186087,0.13204187,0.19240387,0.19240387,0.14713238,0.14335975,0.13958712,0.12826926,0.10186087,0.0754525,0.071679875,0.071679875,0.09808825,0.12826926,0.13958712,0.120724,0.14713238,0.12826926,0.1056335,0.10940613,0.150905,0.14713238,0.22258487,0.3169005,0.38480774,0.392353,0.46026024,0.4640329,0.45648763,0.44139713,0.35462674,0.42630664,0.41121614,0.3772625,0.34330887,0.29049212,0.3734899,0.41498876,0.44894236,0.44139713,0.30935526,0.20372175,0.32444575,0.4979865,0.66775465,0.9016574,0.80356914,0.56212115,0.48666862,0.6413463,0.88279426,0.66775465,0.694163,0.69793564,0.5998474,0.513077,0.5583485,0.68661773,0.7696155,0.88279426,1.2864652,1.3807807,2.0598533,2.1956677,1.7542707,1.8146327,1.5807298,1.5316857,2.033445,2.6219745,2.003264,3.1048703,3.9574835,4.315883,4.3875628,4.8402777,7.183078,9.903141,10.378491,9.012801,9.190115,6.221059,4.115934,3.1425967,3.4670424,5.1647234,2.848332,2.9011486,3.4217708,3.6330378,3.9122121,4.6252384,5.945657,6.4247804,5.704209,4.496969,6.247467,4.7648253,5.2250857,7.1340337,4.353609,2.2409391,1.7014539,1.7278622,1.901403,2.3805263,1.9579924,1.7882242,1.7995421,1.7731338,1.3656902,1.4071891,0.87147635,0.63002837,0.8299775,0.87147635,0.87147635,1.0072908,1.4071891,2.0900342,2.969056,3.4896781,6.0739264,9.22784,11.242422,10.197406,11.3971,11.41219,10.710483,10.601076,13.215506,13.841762,14.04171,12.970284,11.223559,10.823661,9.024119,9.348565,10.144588,10.325675,9.352338,8.880759,7.884786,7.326438,7.3000293,7.0284004,7.9715567,8.443134,8.756263,9.024119,9.152389,8.416726,9.25425,9.763554,9.491924,9.450426,8.458225,6.85486,5.613666,4.851596,3.8292143,4.093298,4.036709,3.9763467,4.2819295,5.3873086,6.620957,8.096053,9.171251,9.839006,10.763299,11.940358,9.937095,6.217286,3.2557755,4.5196047,7.6508837,8.692128,6.85486,4.353609,6.3945994,5.8136153,4.719554,4.2517486,4.779916,5.885295,3.006782,3.5274043,3.3538637,2.2673476,3.9310753,8.16396,9.020347,6.8737226,4.3875628,6.5002327,2.6936543,1.3468271,2.9200118,4.8968673,1.780679,2.505023,3.9159849,5.3684454,5.409944,1.7655885,3.731126,3.8178966,3.6971724,3.863168,3.6141748,2.848332,3.893349,4.6290107,4.055572,2.3088465,11.532914,11.559323,9.533423,8.937348,9.593785,13.551269,15.00373,13.053283,9.454198,8.646856,12.566614,24.556017,30.429993,23.95617,6.862405,10.646348,12.611885,10.914205,6.9567204,5.3986263,4.821415,5.462761,5.4476705,4.8968673,5.9117036,4.2404304,4.8100967,5.4967146,5.745708,6.5568223,5.0968165,5.8098426,6.752999,7.4509344,8.869441,10.242677,10.627484,10.084227,9.193887,9.035437,8.341274,8.054554,8.322411,9.688101,13.079691,14.260523,11.548005,10.401127,11.672502,11.615912,11.921495,11.68382,10.914205,10.137043,10.359629,8.850578,8.262049,8.13378,8.171506,8.254503,8.91094,7.707473,7.413208,9.265567,12.943876,6.5455046,7.805561,7.8508325,7.865923,19.108345,18.406637,9.050528,3.1576872,3.9197574,5.594803,2.8709676,4.745962,5.926794,5.511805,6.9869013,10.638803,8.024373,7.454707,10.159679,10.310584,12.445889,12.570387,11.69891,10.465261,9.114662,12.608112,16.561823,17.033401,15.441354,18.531134,16.690092,19.38752,16.795727,8.201687,1.9806281,5.7079816,5.9532022,6.519096,8.311093,9.333474,13.109872,7.5716586,5.6023483,8.601585,6.4738245,4.889322,4.7572803,7.020855,9.322156,6.013564,7.5188417,7.7602897,9.110889,10.974566,9.808825,9.431562,10.702937,11.072655,10.382264,10.861387,9.997457,10.26154,10.201178,9.740918,10.167224,7.0887623,7.0849895,8.375228,9.782416,10.770844,10.216269,9.148616,8.831716,9.393836,9.827688,8.122461,6.5945487,5.832478,5.824933,5.975838,7.277394,7.9828744,6.7341356,5.836251,11.2650585,8.650629,10.533169,11.200924,9.446653,8.582722,11.050018,9.846551,10.393582,12.985375,12.770335,12.81938,11.966766,10.831206,9.544742,7.7640624,7.564113,7.069899,6.273875,5.251494,4.1800685,3.682082,4.191386,4.745962,4.9723196,5.1043615,5.3571277,5.304311,5.4967146,5.726845,5.040227,5.0175915,4.7572803,4.689373,4.776143,4.52715,4.3422914,4.1008434,4.2064767,4.7120085,5.3382645,5.753253,6.6058664,7.4509344,8.182823,9.042982,9.57115,9.906913,10.378491,11.227332,12.626976,13.63804,14.388792,15.433809,16.65614,17.282394,17.67852,17.520071,16.780636,15.739391,14.943368,14.509516,14.894323,15.82239,16.976812,18.02183,18.38023,18.648085,18.557543,18.097282,17.497435,16.667458,16.31283,16.06761,15.573396,14.468017,13.864397,13.721037,14.358611,15.343266,15.494171,15.841252,15.848798,15.196134,14.437836,15.007503,16.052519,16.516552,16.486372,16.252468,16.331694,16.803272,16.863634,16.946632,16.976812,16.38451,15.629986,14.505743,14.071891,14.554788,15.324403,15.607349,15.388537,15.105591,14.618922,13.249459,12.404391,12.770335,13.20796,13.128735,12.47607,12.257258,12.483616,12.940104,13.340002,13.317367,13.181552,12.725064,12.487389,12.47607,12.170488,12.570387,13.264549,14.18507,14.445381,13.856852,12.913695,11.589504,10.906659,10.567122,10.374719,10.26154,10.378491,10.246449,10.253995,10.559577,11.072655,11.744182,12.053536,12.30253,12.393073,11.808316,11.891314,11.664956,11.351829,10.993429,10.419991,9.748463,9.97482,10.065364,9.831461,9.895596,10.499215,11.193378,11.332966,10.661438,9.303293,8.341274,7.7942433,7.564113,7.4169807,6.9869013,6.115425,5.485397,5.3080835,5.560849,5.9984736,6.017337,6.0512905,6.1229706,6.2323766,6.3229194,6.017337,5.753253,5.511805,5.3609,5.4363527,5.553304,5.4212623,5.089271,4.7308717,4.6554193,4.9459114,5.142088,5.3458095,5.6551647,6.1833324,6.571913,6.673774,6.507778,6.296511,6.462507,5.885295,5.66271,5.783434,6.2097406,6.900131,7.752744,8.367682,8.6732645,8.703445,8.616675,8.6732645,8.612903,8.59404,8.7600355,9.235386,10.269085,11.053791,11.495189,11.649866,11.710228,11.642321,11.223559,10.457717,9.537196,8.831716,8.571404,8.695901,8.98262,9.310839,9.65792,10.231359,11.091517,11.68382,11.959221,12.370438,12.728837,12.789199,12.491161,11.993175,11.676274,11.898859,11.91395,11.548005,11.019837,10.967021,11.231105,12.015811,12.759018,13.407909,14.434063,15.098045,15.230087,15.501716,15.875206,15.596032,14.898096,14.264296,13.690856,13.087236,12.264804,11.295239,10.838752,10.578441,10.246449,9.601331,8.809079,8.375228,8.103599,7.911195,7.816879,7.5792036,7.877241,8.514814,9.246704,9.767326,9.808825,10.186088,10.416218,10.461489,10.7557535,10.321902,9.789962,9.5032425,9.344792,8.718536,8.616675,8.409182,7.960239,7.3981175,7.1038527,6.9189944,6.6020937,6.247467,5.8588867,5.379763,4.8930945,4.6931453,4.459243,4.014073,3.2972744,2.837014,2.444661,2.0749438,1.7354075,1.4939595,1.4034165,1.237421,1.146878,1.1393328,1.056335,1.1846043,1.237421,1.3128735,1.4335974,1.5354583,1.720317,1.7240896,1.7165444,1.7278622,1.6524098,1.3619176,1.2147852,1.0902886,0.95447415,0.87902164,0.724344,0.6790725,0.58098423,0.4376245,0.42630664,0.38480774,0.33576363,0.331991,0.41498876,0.6149379,0.5394854,0.3734899,0.241448,0.18485862,0.120724,0.08677038,0.071679875,0.08299775,0.1056335,0.10186087,0.124496624,0.15845025,0.150905,0.116951376,0.14335975,0.120724,0.09808825,0.09808825,0.10940613,0.1056335,0.1056335,0.1358145,0.14713238,0.124496624,0.116951376,0.13958712,0.13204187,0.1358145,0.181086,0.27540162,0.2867195,0.35839936,0.43007925,0.47535074,0.5017591,0.58098423,0.59230214,0.543258,0.45648763,0.3772625,0.4074435,0.38103512,0.33576363,0.30181,0.30935526,0.331991,0.32821837,0.362172,0.40367088,0.3169005,0.22258487,0.44139713,0.60362,0.65643674,0.8563859,0.66775465,0.59607476,0.58098423,0.6488915,0.94692886,0.62625575,0.58475685,0.6111652,0.5998474,0.55080324,0.6073926,0.8111144,1.146878,1.4222796,1.3091009,1.0978339,3.2482302,3.8782585,2.6182017,2.6068838,2.4031622,1.8334957,1.8523588,2.372981,2.2899833,2.6446102,3.5575855,4.187614,4.429062,4.889322,6.696409,7.816879,7.0887623,4.9685473,3.561358,4.1272516,3.2557755,3.5462675,6.0550632,10.299266,8.933576,5.8513412,3.5538127,2.6936543,2.0862615,3.059599,4.274384,4.6290107,4.115934,3.8405323,4.9685473,3.1312788,3.5839937,5.553304,2.2258487,1.0827434,0.754525,0.8186596,1.0978339,1.6524098,1.3996439,1.5015048,1.7693611,1.9768555,1.8599042,1.5467763,1.2864652,1.2110126,1.1846043,0.7884786,0.995973,1.3091009,2.0673985,3.2369123,4.38379,4.6252384,7.032173,9.963503,12.012038,12.0082655,13.58145,13.951167,13.766309,14.034165,16.090246,16.380737,16.7995,15.339493,12.506252,11.302785,10.054046,9.58624,9.782416,9.876732,8.461998,9.159933,8.0206,7.326438,7.4584794,6.930312,7.533932,7.6584287,7.798016,8.14887,8.612903,7.745199,8.52236,9.129752,9.027891,8.918486,9.514561,8.114917,6.5266414,5.323174,3.8405323,4.164978,4.115934,3.92353,3.953711,4.7120085,5.764571,7.3151197,8.507269,9.024119,9.092027,11.016065,9.416472,5.624984,2.4182527,4.006528,6.851087,6.9454026,6.2361493,6.119198,7.432071,5.149633,4.606375,4.6252384,5.119452,7.118943,3.1161883,4.3083377,4.08198,1.7655885,2.6672459,9.5032425,9.25425,6.907676,6.221059,9.710737,4.772371,2.354118,3.2105038,4.9119577,1.8485862,2.4559789,2.584248,4.82896,7.492433,4.5799665,4.8402777,5.926794,5.5080323,3.863168,3.8669407,2.9992368,3.9989824,5.43258,5.8400235,3.7386713,6.7114997,8.586494,8.179051,6.8737226,8.631766,9.574923,10.672756,10.34831,9.167479,9.857869,10.310584,13.902123,15.267814,12.264804,5.96452,8.6732645,11.359374,13.079691,12.679792,8.809079,6.462507,5.3344917,4.949684,4.689373,3.8141239,5.492942,5.5382137,4.930821,4.4705606,4.7535076,4.82896,4.8440504,5.4288073,6.6850915,8.171506,8.36391,10.370946,11.4838705,10.672756,8.582722,7.7037,6.9491754,7.281166,9.031664,11.883769,13.324911,10.242677,9.7296,11.91395,9.967276,11.053791,12.73261,12.774108,11.219787,10.355856,10.378491,9.374973,8.688355,8.669493,8.68081,11.272603,9.258021,7.6282477,8.869441,12.943876,7.484888,9.631512,11.404645,11.204697,13.819125,17.274849,16.25624,12.185578,7.77538,7.0510364,4.2064767,5.3080835,6.537959,6.175787,4.568649,7.3113475,7.0812173,6.790725,7.062354,6.228604,8.695901,9.374973,9.759781,10.344538,10.612394,11.212241,13.12119,13.426772,12.438345,13.675766,13.815352,13.739901,10.231359,4.9044123,4.2027044,11.793225,10.4049,7.4999785,6.3945994,6.2625575,22.077402,12.068627,3.6066296,4.7648253,4.3083377,8.397863,5.873977,6.9491754,10.846297,5.828706,5.4174895,7.677292,9.0807085,9.280658,11.099063,9.95973,10.280403,10.710483,10.823661,11.114153,10.601076,10.567122,10.638803,10.570895,10.246449,7.3981175,6.9680386,7.907422,9.390063,10.812344,9.922004,9.152389,9.035437,9.333474,9.024119,7.5301595,7.5490227,6.983129,5.828706,6.156924,9.178797,6.673774,4.640329,6.1003346,11.099063,12.657157,10.982111,9.325929,8.280911,5.783434,9.446653,9.092027,9.507015,11.363147,11.227332,11.506506,11.212241,10.359629,9.163706,8.058327,7.7602897,7.0284004,6.0550632,5.070408,4.3385186,4.395108,4.696918,4.851596,4.9421387,5.515578,6.0362,5.8890676,5.775889,5.794752,5.455216,5.240176,4.817642,4.5460134,4.4894238,4.4215164,4.8063245,4.859141,4.8968673,5.0666356,5.3684454,6.175787,6.952948,7.4735703,7.7904706,8.20546,9.103344,10.159679,10.974566,11.548005,12.268577,13.189097,13.86817,14.577423,15.396083,16.218515,16.939087,17.222033,16.82968,15.841252,14.652876,14.456699,14.962231,15.811071,16.795727,17.829426,17.795471,18.048239,18.26705,18.350048,18.391546,16.950403,16.459963,16.520325,16.59955,16.03743,14.385019,13.819125,14.403882,15.39231,15.211224,15.00373,14.373701,13.50977,13.12119,14.422746,15.935568,15.99593,15.675257,15.562078,15.784663,15.99593,15.818617,16.222288,16.923996,16.395828,15.452672,14.203933,13.272095,13.053283,13.694629,14.743419,15.218769,15.049001,14.32843,13.343775,12.687338,13.204187,13.502225,13.106099,12.434572,12.510024,12.687338,13.12119,13.607859,13.592768,13.355092,13.230596,12.981603,12.623203,12.411936,12.83447,12.687338,13.275867,13.36641,12.668475,11.861133,10.782163,9.937095,9.507015,9.476834,9.616421,10.137043,10.325675,10.484125,10.7557535,11.102836,11.548005,11.578186,11.480098,11.423509,11.461235,11.336739,10.702937,10.133271,9.955957,10.246449,10.419991,10.487898,10.054046,9.333474,9.133525,10.050273,10.95193,10.993429,9.940866,8.152642,7.2887115,6.8397694,6.7152724,6.6586833,6.247467,5.745708,5.3609,5.402399,5.783434,6.013564,5.6363015,5.4740787,5.4174895,5.4288073,5.523123,5.3194013,5.194905,5.05909,4.908185,4.7874613,4.9534564,4.8553686,4.6931453,4.606375,4.6742826,4.8402777,4.889322,5.0175915,5.281675,5.583485,5.7909794,5.9682927,6.0701537,6.2021956,6.628502,6.375736,6.609639,7.0057645,7.454707,8.065872,8.718536,9.148616,9.348565,9.352338,9.246704,9.2995205,9.329701,9.208978,9.0543,9.25425,10.340765,11.114153,11.563096,11.668729,11.393328,11.102836,10.510533,9.8239155,9.21275,8.793989,9.208978,9.669238,9.884277,9.782416,9.507015,9.665465,10.27663,10.751981,11.046246,11.68382,12.049765,12.170488,11.951676,11.495189,11.121698,11.532914,11.348056,10.540714,9.703192,10.054046,10.7557535,11.649866,12.585477,13.532406,14.618922,14.626467,14.366156,14.735873,15.675257,16.18456,15.513034,14.841507,14.117163,13.336229,12.551523,11.551778,10.989656,10.695392,10.442626,9.910686,9.612649,9.525878,9.333474,8.956212,8.541223,8.160188,8.390318,9.125979,9.903141,9.899368,9.703192,10.250222,10.616167,10.801025,11.740409,10.872705,10.370946,10.106862,9.805053,9.024119,8.729855,8.548768,8.333729,8.080963,7.9225125,7.6697464,7.432071,7.039718,6.477597,5.881522,5.1571784,4.9459114,4.949684,4.749735,3.7952607,3.2972744,2.9086938,2.6219745,2.384299,2.1164427,2.2183034,2.033445,1.8976303,1.9202662,1.9768555,2.1013522,2.0108092,1.9353566,1.9391292,1.931584,2.0296721,2.0372176,2.0070364,1.9730829,1.9504471,1.5580941,1.4071891,1.2751472,1.0902886,0.9205205,0.7432071,0.7205714,0.6451189,0.482896,0.3734899,0.31312788,0.331991,0.47912338,0.70170826,0.8563859,0.65643674,0.4376245,0.27917424,0.19994913,0.1659955,0.12826926,0.10186087,0.090543,0.09808825,0.120724,0.1358145,0.13958712,0.12826926,0.120724,0.1358145,0.1056335,0.08299775,0.10186087,0.14335975,0.14713238,0.1659955,0.18863125,0.17731337,0.181086,0.32821837,0.2263575,0.18485862,0.2263575,0.33576363,0.4376245,0.42630664,0.47912338,0.5319401,0.59230214,0.76584285,0.754525,0.7696155,0.6413463,0.45648763,0.52062225,0.41498876,0.31312788,0.271629,0.29426476,0.331991,0.27540162,0.2565385,0.32067314,0.4074435,0.36594462,0.25276586,0.4376245,0.5357128,0.5055317,0.66775465,0.55457586,0.5885295,0.62248313,0.6752999,0.9507015,0.5885295,0.5357128,0.663982,0.9016574,1.2298758,0.95447415,0.98465514,1.2336484,1.3845534,0.87147635,1.1242423,3.006782,3.6443558,2.7125173,2.4220252,2.9539654,2.4786146,2.123988,2.2220762,2.323937,2.233394,3.429316,4.304565,4.715781,5.994701,6.700182,7.33021,7.466025,6.752999,4.8855495,3.9008942,3.097325,5.6400743,10.480352,12.344029,10.680302,6.571913,3.5802212,2.5691576,1.7240896,1.9466745,2.4597516,2.5314314,2.214531,2.354118,2.6672459,1.5165952,2.372981,4.1574326,1.2525115,0.6790725,0.43385187,0.422534,0.6488915,1.2223305,1.0940613,1.2600567,1.5505489,1.8372684,2.052308,1.7995421,1.7580433,1.6410918,1.358145,1.0186088,1.2449663,1.7429527,2.6483827,4.0216184,5.8437963,6.0512905,7.1906233,8.612903,10.306811,12.894833,14.1058445,14.4114275,14.762281,15.309312,15.414946,16.365646,17.471025,16.429781,13.577678,11.891314,11.18206,10.110635,9.756008,9.752235,8.29223,8.827943,7.835742,7.3453007,7.586749,7.001992,6.9152217,6.8246784,6.7454534,6.911449,7.7640624,7.2396674,7.586749,8.186596,8.544995,8.314865,9.842778,8.748717,7.2170315,6.017337,4.478106,4.5761943,4.6554193,4.4743333,4.217795,4.515832,5.2967653,7.0812173,8.6732645,9.310839,8.68081,10.729345,8.703445,4.938366,2.1579416,3.4745877,7.364164,5.4891696,4.644101,6.7379084,8.801534,6.617184,4.8327327,4.0216184,4.9232755,8.4544525,5.8437963,7.537705,7.594294,4.6931453,2.123988,7.360391,6.485142,4.6290107,4.738417,7.594294,4.104616,2.263575,2.3201644,2.9992368,1.5241405,2.546522,1.7580433,3.0407357,6.319147,7.564113,5.2137675,5.621211,5.036454,3.9273026,6.971811,4.7233267,3.731126,4.3800178,5.8664317,6.1908774,4.142342,6.356873,6.9265394,5.534441,7.4697976,7.020855,6.485142,6.0512905,6.319147,8.296002,8.458225,7.111398,5.3080835,4.104616,4.5724216,5.904158,7.360391,10.499215,13.468271,10.997202,7.6697464,5.43258,4.5007415,4.2517486,3.2331395,6.8397694,8.122461,6.9189944,4.610148,4.1612053,4.5460134,4.678055,5.0553174,5.945657,7.3717093,6.006019,8.126234,10.378491,10.510533,7.3679366,6.598321,5.7192993,6.6134114,8.809079,9.495697,9.601331,7.5301595,7.7414265,10.163452,10.216269,10.789707,10.906659,10.091772,8.7600355,8.22055,8.14887,7.2623034,7.5075235,8.816625,9.099571,11.223559,10.914205,9.408927,8.52236,10.627484,9.0543,9.7220545,12.562841,14.11339,7.515069,9.473062,12.736382,11.774363,7.164215,5.5797124,4.825187,9.073163,11.374464,10.253995,9.688101,11.940358,11.200924,7.6848373,4.123479,5.775889,5.330719,6.1116524,8.024373,10.555805,12.774108,9.307066,7.884786,7.997965,8.865668,9.446653,9.329701,7.5905213,4.7610526,2.8332415,5.247721,10.521852,13.547497,12.600568,9.107117,7.654656,18.157644,11.276376,6.1041074,7.798016,7.575431,8.548768,5.247721,5.089271,7.877241,5.798525,3.7801702,7.152897,8.729855,7.7942433,10.110635,9.933322,9.952185,10.238904,10.827434,11.725319,11.148107,10.86516,11.114153,11.423509,10.597303,8.284684,7.0963078,7.432071,8.816625,9.895596,9.435335,9.239159,9.024119,8.7600355,8.688355,7.828197,8.597813,7.786698,5.3873086,4.61392,7.9338303,5.1043615,4.647874,7.8621507,8.827943,13.490907,10.042727,7.484888,7.8395147,6.1606965,7.605612,8.190369,9.020347,9.861642,9.144843,9.933322,10.299266,9.884277,9.016574,8.741172,7.6622014,6.7756343,5.8211603,4.9157305,4.564876,4.8063245,4.8742313,4.8629136,4.98741,5.594803,6.1833324,6.307829,6.0776987,5.7306175,5.613666,5.2892203,4.9459114,4.7006907,4.61392,4.689373,5.240176,5.3910813,5.330719,5.3080835,5.6287565,6.375736,7.01331,7.3905725,7.5565677,7.748972,8.914713,10.246449,11.027383,11.216014,11.46878,11.996947,12.796744,13.626721,14.441608,15.388537,16.161926,16.403374,16.286423,15.773345,14.626467,14.562332,14.996184,15.7657995,16.897587,18.640541,18.048239,17.523844,17.346529,17.508753,17.72002,16.569368,16.218515,16.309057,16.452417,16.218515,14.78869,14.181297,14.219024,14.603831,14.909414,14.849052,13.932304,12.985375,12.792972,14.124708,15.467763,15.520579,15.214996,15.060319,15.124454,15.237633,15.015047,15.331948,15.946886,15.501716,14.592513,13.570132,12.653384,12.136535,12.408164,13.879487,14.667966,14.690601,14.120935,13.392818,12.770335,13.087236,13.234368,12.849561,12.310076,12.336484,12.562841,13.072145,13.660675,13.837989,13.547497,13.539951,13.272095,12.751472,12.559069,12.306303,12.510024,12.415709,11.898859,11.155652,10.714255,9.993684,9.190115,8.809079,8.858124,8.858124,9.654147,10.182315,10.359629,10.295494,10.284176,10.631257,10.661438,10.533169,10.502988,10.944386,10.47658,9.691874,8.99771,8.922258,10.095545,10.770844,10.653893,10.103089,9.529651,9.416472,10.03141,10.616167,10.49167,9.507015,8.013056,7.696155,7.537705,7.496206,7.326438,6.587003,5.9305663,5.6363015,5.643847,5.753253,5.6098933,4.636556,4.3800178,4.3347464,4.29702,4.357382,4.4630156,4.5196047,4.45547,4.2328854,3.8405323,3.99521,4.221567,4.5460134,4.9232755,5.2326307,5.149633,5.0439997,4.9421387,4.889322,4.9345937,5.3646727,5.6778007,5.915476,6.126743,6.3832817,6.8699503,7.828197,8.616675,9.0543,9.4127,9.239159,9.378746,9.714509,10.001229,9.876732,9.842778,10.099318,10.144588,9.835234,9.397609,9.861642,10.310584,10.808571,11.11038,10.661438,10.495442,10.121953,9.654147,9.175024,8.714764,9.469289,10.106862,10.178542,9.714509,9.21275,9.525878,9.857869,10.0276375,10.106862,10.438853,10.469034,10.687846,10.70671,10.465261,10.238904,10.710483,10.801025,10.340765,9.789962,10.227587,11.102836,11.7555,12.434572,13.189097,13.86817,13.162688,12.868423,13.377728,14.4152,15.0376835,14.324657,13.521088,12.619431,11.736636,11.106608,10.748209,10.533169,10.442626,10.374719,10.133271,10.442626,10.56335,10.340765,9.820143,9.246704,9.133525,9.114662,9.631512,10.159679,9.246704,9.216523,10.121953,10.61994,10.744436,11.883769,11.18206,10.921749,10.544487,9.857869,9.027891,8.60913,8.458225,8.612903,8.944894,9.148616,8.959985,8.956212,8.526133,7.647111,6.8850408,6.2135134,5.8702044,5.915476,5.8626595,4.6856003,3.9989824,3.5123138,3.1840954,2.9426475,2.6974268,3.0256453,3.0445085,2.987919,3.0369632,3.2972744,3.2935016,2.9766011,2.6483827,2.4672968,2.4522061,2.3880715,2.4182527,2.3767538,2.2409391,2.11267,1.720317,1.6033657,1.5015048,1.2902378,0.9922004,0.8262049,0.7582976,0.6790725,0.5696664,0.4979865,0.43007925,0.40367088,0.5885295,0.8526133,0.7432071,0.47535074,0.4074435,0.35839936,0.27540162,0.21881226,0.21881226,0.23013012,0.21503963,0.181086,0.17354076,0.181086,0.15845025,0.14335975,0.14713238,0.13204187,0.13204187,0.12826926,0.1358145,0.16222288,0.19994913,0.24899325,0.2565385,0.26031113,0.362172,0.7432071,0.543258,0.41121614,0.46026024,0.6187105,0.63002837,0.58098423,0.6790725,0.7696155,0.8903395,1.2525115,1.0223814,0.9808825,0.80356914,0.55457586,0.69039035,0.4074435,0.271629,0.27540162,0.34330887,0.331991,0.23390275,0.241448,0.32821837,0.43385187,0.46026024,0.3055826,0.35085413,0.39989826,0.4074435,0.4640329,0.41876137,0.4678055,0.5093044,0.5885295,0.8903395,0.5772116,0.5998474,0.8337501,1.327964,2.2975287,1.5882751,1.2751472,1.1317875,0.95447415,0.5772116,1.4939595,1.5618668,1.6146835,1.7089992,1.1506506,2.5238862,2.8634224,2.6710186,2.354118,2.233394,2.282438,3.7386713,4.708236,5.4212623,8.216777,7.6622014,7.3717093,8.122461,9.250477,8.643084,3.199186,2.3126192,6.1795597,10.695392,7.4584794,5.5985756,3.7990334,2.8219235,2.595566,2.2258487,0.8639311,0.66020936,0.80734175,0.90920264,0.98842776,0.9280658,0.6488915,1.5958204,2.7804246,0.784706,0.73566186,0.4376245,0.3055826,0.49044126,0.87147635,0.91674787,0.965792,1.2336484,1.629774,1.7580433,2.0372176,2.1353056,1.8636768,1.448688,1.50905,1.4675511,2.0145817,2.795515,4.08198,6.749226,7.122716,6.862405,6.5568223,7.677292,12.611885,12.887287,12.879742,13.347548,13.702174,11.996947,13.487134,15.531898,15.762027,13.973803,12.113899,11.887542,10.393582,9.631512,9.688101,8.726082,8.07719,7.303802,7.062354,7.201941,6.7756343,6.2135134,6.1720147,5.8928404,5.643847,6.7039547,7.020855,6.907676,7.4207535,8.348819,8.209232,9.665465,8.733627,7.5226145,6.7114997,5.564622,5.5193505,5.643847,5.50426,5.2364035,5.5306683,5.926794,7.84706,9.88805,10.9594755,10.26154,11.766817,8.805306,4.851596,2.3767538,2.8332415,8.246958,5.311856,3.1765501,5.1571784,8.741172,6.6624556,3.2444575,1.6863633,3.6028569,9.001483,10.570895,10.050273,9.997457,9.476834,4.0480266,4.561104,3.6066296,2.071171,1.0412445,1.8334957,1.1732863,1.327964,1.388326,1.2223305,1.4901869,2.7087448,1.8523588,1.961765,4.738417,10.555805,4.4630156,2.7011995,2.7841973,4.6856003,10.842525,7.032173,3.8669407,3.1954134,5.1269975,8.024373,6.1305156,6.4511886,6.330465,5.323174,5.194905,5.715527,4.4441524,3.187868,3.308592,5.723072,5.50426,5.0553174,4.8742313,4.9157305,4.564876,5.6891184,4.561104,5.50426,8.703445,10.231359,7.9753294,5.9720654,4.991183,5.032682,5.3194013,8.318638,10.687846,9.186342,5.138315,4.447925,3.9989824,5.028909,5.50426,5.3194013,6.296511,4.3007927,5.13077,7.1679873,8.216777,5.511805,5.666483,5.2854476,6.326692,8.20546,7.805561,5.9305663,6.187105,6.356873,6.7831798,10.374719,10.080454,7.5301595,5.1798143,4.255521,4.7346444,4.168751,3.7235808,5.0062733,7.635793,9.250477,8.903395,11.2801485,11.646093,9.559832,8.858124,11.276376,8.582722,9.95973,13.664448,7.01331,4.044254,3.029418,3.3048196,3.983892,3.9688015,5.87775,12.943876,15.562078,13.570132,16.237377,19.851553,17.342756,10.212496,4.112161,8.835487,5.9305663,5.8928404,7.405663,9.593785,12.015811,7.2887115,4.8666863,4.3611546,5.330719,7.284939,5.0741806,4.538468,3.3576362,2.1390784,4.4139714,4.678055,13.045737,16.754227,13.555041,11.725319,5.089271,5.4174895,9.533423,13.257004,11.393328,3.338773,2.7841973,5.643847,7.7904706,5.032682,3.7273536,6.651138,8.269594,7.533932,7.8923316,8.892077,9.616421,10.061591,10.661438,12.30253,11.431054,11.121698,11.52537,11.966766,10.917976,9.216523,7.383027,7.0963078,8.179051,8.582722,9.031664,9.186342,8.586494,7.9300575,9.065618,8.495952,8.443134,7.281166,4.9949555,3.1954134,4.8365054,3.742444,5.0515447,7.9300575,5.5683947,9.899368,7.960239,6.688864,7.6320205,6.952948,7.383027,7.654656,8.416726,8.986393,7.3717093,8.333729,9.156161,9.190115,8.778898,9.25425,7.394345,6.379509,5.523123,4.798779,4.8629136,4.8138695,4.7535076,4.8855495,5.2062225,5.4740787,5.904158,6.2851934,6.043745,5.379763,5.27413,5.1647234,5.040227,5.062863,5.240176,5.4212623,5.6363015,5.617439,5.50426,5.5570765,6.168242,6.5266414,6.934085,7.1076255,7.118943,7.394345,8.620448,9.7069645,10.18986,10.216269,10.536942,10.702937,11.619685,12.73261,13.747445,14.6302395,14.973549,14.800008,14.739646,14.758509,14.173752,14.2944765,14.766054,15.667711,17.267305,20.013775,18.995167,17.452164,16.41092,16.075155,15.833707,15.418718,15.32063,15.350811,15.328176,15.101818,14.6151495,14.147344,13.426772,12.96274,14.037937,14.57365,14.226569,13.604086,13.29473,13.849306,14.592513,15.131999,15.17727,14.826416,14.562332,14.886778,14.871688,14.709465,14.422746,13.8719425,13.226823,12.823153,12.404391,12.0233555,12.064855,13.268322,13.920986,14.1058445,13.79649,12.875969,12.181807,12.438345,12.898605,13.087236,12.792972,12.400619,12.58925,13.117417,13.698401,14.045483,13.8870325,13.505998,13.045737,12.630749,12.355347,10.940613,11.514051,12.691111,12.687338,11.506506,10.970794,10.140816,9.567377,9.567377,9.933322,9.933322,10.103089,9.771099,9.118435,8.405409,7.964011,8.6732645,9.005256,9.190115,9.480607,10.163452,9.590013,8.548768,7.8395147,7.677292,7.6923823,7.7376537,7.7225633,7.8961043,8.367682,9.125979,9.125979,9.107117,9.076936,9.001483,8.820397,9.186342,9.031664,8.797762,8.503497,7.7225633,6.8925858,6.096562,5.43258,5.0477724,5.1571784,4.436607,3.9008942,3.6066296,3.5274043,3.5387223,3.9688015,4.3309736,4.353609,4.1083884,3.9989824,3.85185,4.134797,4.4177437,4.5120597,4.485651,4.4630156,4.4743333,4.515832,4.738417,5.4476705,5.983383,6.3116016,6.511551,6.7756343,7.3868,7.8621507,8.646856,9.205205,9.473062,9.88805,10.340765,10.56335,10.653893,10.514306,9.842778,9.65792,9.25425,9.288202,9.665465,9.567377,10.227587,10.740664,11.012292,11.000975,10.695392,10.121953,9.952185,9.42779,8.458225,7.6282477,8.959985,9.65792,9.876732,9.922004,10.238904,10.140816,10.216269,10.182315,10.084227,10.314357,9.544742,9.710737,9.80128,9.616421,9.752235,9.676784,10.56335,11.223559,11.106608,10.299266,10.435081,10.759526,11.200924,11.68382,12.147853,12.585477,12.943876,13.264549,13.302276,12.498707,12.264804,11.593277,10.868933,10.374719,10.299266,10.812344,11.151879,11.09529,10.740664,10.499215,10.352083,10.223814,10.303039,10.442626,10.163452,10.272858,10.54826,10.770844,10.589758,9.491924,10.223814,11.185833,11.16697,10.518079,11.140562,11.823407,11.646093,10.740664,9.699419,9.552286,9.367428,9.525878,9.597558,9.661693,10.284176,10.26154,10.510533,10.344538,9.64283,8.850578,7.9828744,7.7376537,7.7640624,7.492433,6.149379,4.927048,4.2102494,3.6141748,3.150142,3.2331395,3.5651307,3.9499383,4.032936,3.9688015,4.4101987,4.4818783,4.1272516,3.6066296,3.1463692,2.916239,2.8030603,2.6672459,2.5880208,2.4899325,2.1353056,1.9881734,1.8259505,1.629774,1.418507,1.237421,1.0902886,0.8865669,0.73566186,0.65643674,0.59607476,0.5093044,0.3961256,0.3734899,0.41498876,0.36594462,0.4376245,0.59607476,0.62625575,0.5017591,0.36594462,0.513077,0.66775465,0.694163,0.55080324,0.32067314,0.26031113,0.18863125,0.14713238,0.13204187,0.1056335,0.20372175,0.24899325,0.21503963,0.17354076,0.26031113,0.30935526,0.3470815,0.43385187,0.66020936,1.1581959,1.2826926,1.0450171,0.9922004,1.1317875,0.9620194,0.91297525,1.2562841,1.5430037,1.690136,1.9844007,1.3845534,1.1544232,1.0450171,0.8978847,0.6413463,0.4074435,0.46026024,0.44894236,0.30935526,0.26031113,0.26031113,0.29426476,0.29049212,0.29049212,0.47157812,0.47157812,0.49044126,0.5772116,0.6828451,0.67152727,0.40367088,0.33576363,0.29803738,0.35462674,0.7922512,0.5998474,0.7884786,1.0072908,1.3958713,2.5804756,2.3088465,1.8863125,1.5015048,1.3468271,1.6033657,2.2258487,1.6675003,1.1431054,0.9318384,0.38103512,1.2864652,2.5616124,2.8445592,2.2447119,2.3805263,2.5276587,3.9914372,5.304311,6.688864,10.069136,9.314611,5.938112,3.712263,3.1237335,1.4034165,1.3807807,4.67051,5.7381625,3.2369123,0.0,0.21881226,0.7130261,0.9016574,0.784706,0.9318384,0.7582976,0.5357128,0.4376245,0.52439487,0.73188925,1.1091517,1.1695137,1.3392819,1.5052774,0.9922004,1.3807807,0.8941121,0.5998474,0.724344,0.62625575,0.62625575,0.845068,1.3468271,1.7316349,1.1581959,1.7316349,2.2258487,2.2673476,1.9730829,1.9391292,2.1202152,2.3390274,2.7879698,3.893349,6.349328,6.4926877,7.043491,7.5075235,8.228095,10.374719,9.608876,10.578441,11.283921,10.676529,8.650629,8.639311,11.68382,13.6682205,13.200415,11.627231,12.445889,10.076681,8.563859,8.846806,8.7751255,7.5792036,6.7944975,6.2436943,5.8966126,5.8588867,5.7872066,5.3458095,5.0553174,5.13077,5.5080323,6.7039547,6.8397694,7.2283497,8.073418,8.4544525,9.733373,9.031664,8.114917,7.4697976,6.2851934,6.8359966,6.6624556,6.387054,6.541732,7.567886,7.7037,8.990166,10.834979,12.347801,12.359119,13.936077,11.69891,7.6848373,4.2404304,4.044254,5.764571,4.7836885,3.5575855,3.9688015,7.322665,4.357382,1.6373192,1.7957695,4.508287,6.485142,12.917468,6.560595,5.353355,10.759526,7.7829256,5.7683434,3.2218218,1.6109109,2.0296721,5.20245,2.1503963,2.8709676,3.9461658,3.783943,2.625747,4.515832,3.5877664,5.3759904,10.555805,14.939595,5.560849,3.4557245,4.115934,5.13077,6.1795597,5.583485,4.06689,4.5422406,7.001992,8.514814,6.696409,5.855114,4.52715,2.9464202,3.0822346,3.742444,4.327201,5.247721,6.519096,7.752744,3.6254926,3.289729,6.006019,9.156161,8.239413,7.84706,6.0211096,4.2328854,4.2517486,8.13378,9.74469,9.21275,9.876732,11.117926,8.345046,11.631002,9.337247,5.6023483,2.9200118,2.1503963,3.4330888,5.292993,5.492942,4.221567,4.074435,3.6707642,4.61392,5.492942,5.7570257,5.7079816,6.620957,6.228604,5.692891,6.549277,10.710483,8.073418,12.762791,12.755245,6.700182,3.9084394,4.9685473,7.5301595,7.4584794,4.8063245,3.8292143,6.820906,7.5490227,7.145352,7.284939,10.178542,9.469289,9.484379,10.393582,10.846297,7.964011,14.007756,11.042474,7.213259,6.670001,9.552286,9.465516,7.375482,6.790725,8.3525915,9.842778,10.197406,5.4703064,5.093044,9.1825695,8.560086,5.3382645,9.4013815,9.152389,3.8292143,3.5236318,6.881268,6.907676,5.9984736,5.142088,3.92353,2.897376,5.4401255,5.111907,2.2069857,3.7688525,2.7313805,1.7127718,1.1091517,2.2560298,7.432071,12.0082655,6.5530496,2.8558772,4.0103,4.425289,5.0968165,4.3385186,3.3161373,2.4710693,1.5430037,2.2975287,8.409182,20.862616,27.283625,1.9693103,5.20245,7.515069,8.793989,9.016574,8.209232,7.9300575,9.288202,10.555805,11.227332,12.0082655,11.653639,11.695138,12.064855,12.102581,10.529396,9.099571,7.405663,6.7114997,7.152897,7.752744,8.68081,8.718536,7.9941926,7.4207535,8.710991,7.1264887,5.4665337,4.847823,5.040227,4.4403796,6.198423,3.6254926,2.3616633,3.6368105,4.274384,6.349328,9.0543,9.895596,8.601585,7.111398,8.820397,8.284684,8.620448,9.691874,8.118689,7.250985,7.786698,8.107371,8.156415,9.416472,8.156415,6.571913,5.4363527,5.081726,5.3873086,5.300538,4.949684,5.010046,5.5004873,5.7683434,6.255012,5.9117036,5.379763,4.991183,4.7610526,5.492942,5.704209,5.666483,5.617439,5.753253,5.4967146,5.485397,5.481624,5.5193505,5.934339,6.802043,6.8925858,6.462507,5.9796104,6.089017,7.432071,8.635539,9.344792,9.58624,9.782416,10.061591,10.710483,11.197151,11.649866,12.849561,13.249459,13.113645,12.777881,12.600568,12.955194,13.539951,14.290704,15.339493,16.950403,19.500698,19.24416,17.980331,16.920223,16.429781,16.052519,14.709465,14.264296,14.332202,14.637785,15.015047,14.747191,14.222796,13.426772,12.830698,13.36641,13.792717,13.800262,13.532406,13.249459,13.336229,13.920986,14.637785,15.064092,14.988639,14.403882,14.649103,14.792462,14.7170105,14.335975,13.5663595,12.50248,12.411936,12.381755,12.321393,12.970284,13.702174,14.920732,15.30554,14.426518,12.740154,11.910177,12.830698,14.252977,15.32063,15.562078,14.524607,14.064346,13.856852,13.630494,13.151371,13.287186,12.974057,12.996693,13.419228,13.5663595,9.220296,9.989911,10.93684,11.864905,12.525115,12.642066,12.51757,11.370691,10.733118,11.031156,11.604594,11.872451,11.193378,10.3634,9.81637,9.601331,9.556059,9.371201,8.990166,8.461998,7.964011,7.61693,7.326438,7.1604424,7.149124,7.3000293,7.5829763,7.748972,7.91874,8.035691,7.9036493,7.6886096,7.756517,8.013056,8.2507305,8.137552,8.503497,8.567632,8.314865,7.7942433,7.111398,6.25124,5.7494807,5.485397,5.3458095,5.2288585,4.3649273,4.3913355,4.636556,4.7610526,4.772371,4.817642,4.889322,4.7874613,4.496969,4.191386,4.085753,4.2781568,4.429062,4.357382,4.0216184,3.7348988,3.731126,3.8858037,4.217795,4.8968673,5.7570257,6.2436943,6.4210076,6.5040054,6.858632,7.6584287,8.284684,8.763808,9.031664,8.948667,9.25425,9.782416,10.253995,10.627484,11.087745,10.250222,9.58624,9.522105,9.910686,10.069136,9.710737,9.35611,9.276885,9.393836,9.25425,9.0543,8.661947,8.326183,8.194141,8.311093,9.303293,9.556059,9.552286,9.431562,9.016574,9.25425,9.397609,9.461743,9.574923,9.97482,9.623966,9.578695,9.635284,9.669238,9.616421,9.650374,10.186088,10.789707,11.080199,10.714255,10.691619,11.1782875,11.691365,12.027128,12.257258,12.449662,12.411936,12.012038,11.521597,11.604594,11.978085,11.59705,11.249968,11.223559,11.32542,11.114153,10.774617,10.650121,10.899114,11.476325,11.710228,11.59705,11.415963,11.438599,11.921495,12.54775,12.709973,12.725064,12.619431,12.113899,11.725319,11.593277,11.442371,11.32542,11.615912,11.548005,11.355601,10.699164,9.937095,10.163452,10.106862,9.81637,9.514561,9.276885,9.039209,9.533423,10.321902,10.714255,10.54826,10.20495,10.314357,10.212496,10.076681,9.74469,8.710991,7.3151197,6.0286546,5.089271,4.557331,4.3083377,4.5309224,4.82896,5.05909,5.1760416,5.2628117,4.938366,4.4931965,4.032936,3.663219,3.4896781,3.6896272,3.6443558,3.4783602,3.2331395,2.8822856,2.4031622,2.1051247,1.8900851,1.7429527,1.7240896,1.5769572,1.4637785,1.3355093,1.177059,1.0110635,0.8563859,0.69793564,0.633801,0.7432071,1.086516,1.2751472,1.3241913,1.2638294,1.1317875,0.9393836,0.88279426,0.83752275,0.875249,0.9393836,0.8941121,0.49044126,0.33576363,0.30181,0.3055826,0.29049212,0.32067314,0.33576363,0.38480774,0.47535074,0.5885295,0.724344,0.69039035,0.80734175,1.1280149,1.4524606,1.5354583,1.3204187,1.3204187,1.4864142,1.2185578,1.3920987,1.7278622,2.0258996,2.2409391,2.4823873,2.1013522,1.7844516,1.4449154,1.1091517,0.9205205,0.69793564,0.6526641,0.633801,0.5470306,0.331991,0.2263575,0.26408374,0.331991,0.39989826,0.5357128,0.513077,0.5281675,0.6149379,0.66020936,0.40367088,0.30181,0.39989826,0.4979865,0.5470306,0.633801,0.7432071,0.8601585,1.3619176,2.233394,3.0671442,2.3692086,1.4713237,0.8903395,0.80734175,1.0525624,1.871222,1.20724,0.58098423,0.52062225,0.5772116,1.0902886,2.4899325,3.3312278,3.308592,3.2482302,3.3727267,4.063117,5.0025005,5.994701,6.983129,6.217286,4.3611546,2.7691069,2.1051247,2.354118,1.2751472,3.5689032,3.5462675,1.5128226,3.7952607,2.1805773,1.5769572,1.1280149,0.63002837,0.55080324,0.6149379,0.573439,0.5281675,0.55080324,0.66020936,0.9318384,1.5920477,1.8334957,1.5731846,1.4298248,1.1657411,0.69793564,0.44139713,0.4074435,0.22258487,0.211267,0.49044126,0.83752275,1.0789708,1.0638802,0.94315624,1.0487897,1.358145,1.8070874,2.2786655,2.5993385,2.625747,2.4559789,3.1727777,6.8359966,7.937603,8.873214,8.963757,8.473316,8.616675,5.300538,6.2399216,7.0585814,6.530414,6.6134114,6.8058157,8.854351,10.989656,11.838497,10.419991,11.283921,9.691874,8.477088,8.303548,7.6622014,6.379509,5.726845,5.251494,5.0138187,5.6023483,5.9192486,5.3458095,5.0515447,5.119452,4.5309224,5.885295,6.058836,6.2814207,6.8661776,7.194396,8.114917,7.798016,7.624475,7.6207023,6.458734,6.5002327,6.9680386,7.24344,7.3981175,8.179051,8.224322,8.488406,8.986393,10.038955,12.249713,13.9888935,13.381501,9.7069645,4.5233774,1.6524098,3.6858547,4.2781568,3.4255435,2.8332415,5.8966126,3.0860074,1.6146835,1.6373192,3.108643,5.7909794,6.0701537,5.3684454,7.3981175,10.808571,9.186342,6.1078796,3.4783602,1.871222,2.867195,9.046755,4.881777,2.7540162,4.606375,7.8998766,5.6287565,4.346064,5.772116,7.2396674,7.7037,7.748972,8.959985,6.688864,4.851596,4.406426,3.3350005,5.2175403,5.304311,4.538468,4.0706625,5.2779026,5.523123,6.6624556,7.356619,7.8923316,10.186088,10.680302,5.8928404,4.0706625,7.364164,11.84227,8.612903,8.130007,10.7218,13.336229,9.510788,6.8435416,6.3719635,6.2097406,6.1003346,7.413208,8.83926,8.084735,7.2094865,7.413208,9.065618,14.283158,10.525623,5.4740787,2.9803739,3.0897799,2.7502437,5.3194013,6.217286,4.7044635,3.8556228,3.8707132,5.511805,6.722818,7.039718,7.586749,8.09228,7.001992,5.6363015,5.3986263,7.7829256,6.971811,9.420244,10.499215,8.22055,3.2482302,4.8553686,7.4094353,6.911449,3.5651307,1.7655885,4.6327834,9.216523,10.038955,7.7150183,8.967529,10.974566,10.257768,9.982366,10.272858,8.171506,10.514306,11.778135,10.001229,6.760544,7.1604424,7.043491,7.7150183,8.013056,8.371455,10.819888,8.458225,4.8742313,10.748209,19.18757,5.753253,6.043745,8.812852,10.061591,7.99042,2.9992368,5.7419353,7.9338303,10.461489,11.461235,6.3153744,5.80607,4.6290107,3.6783094,2.9539654,1.5467763,1.3694628,1.2449663,2.3314822,4.5724216,6.7114997,8.243186,8.858124,8.337502,6.79827,4.6931453,5.560849,7.0284004,7.043491,5.3571277,3.531177,1.9730829,4.9723196,11.664956,14.950912,1.5279131,5.010046,7.0057645,7.443389,6.983129,7.0246277,8.76758,9.654147,10.416218,11.16697,11.423509,11.498961,11.476325,11.581959,11.370691,9.748463,8.963757,7.598067,6.809588,6.8963585,7.2887115,7.911195,7.6282477,7.1076255,6.8359966,7.115171,6.25124,4.821415,3.651901,4.1272516,8.175279,9.778644,6.0286546,3.1199608,4.6856003,11.8045435,7.541477,5.764571,7.6320205,10.393582,7.3792543,11.099063,9.786189,8.688355,8.952439,7.643338,6.7944975,7.2170315,7.699928,7.8961043,8.303548,7.575431,6.507778,5.6363015,5.2967653,5.6287565,5.20245,5.485397,5.726845,5.572167,5.05909,6.006019,5.8136153,5.560849,5.5193505,5.138315,5.4703064,6.1305156,6.4210076,6.273875,6.25124,6.300284,6.2135134,5.934339,5.6589375,5.836251,6.3719635,6.670001,6.620957,6.466279,6.820906,7.960239,8.59404,8.850578,8.967529,9.280658,9.250477,9.525878,10.231359,11.046246,11.189606,10.955703,10.921749,11.02361,11.306557,11.955449,12.521342,13.264549,14.219024,15.611122,17.889788,19.127209,18.26705,16.882498,15.746937,14.830189,13.732355,13.283413,13.27964,13.50977,13.721037,12.913695,12.649611,12.864652,13.087236,12.464753,13.2607765,13.4644985,13.124963,12.713746,13.091009,13.920986,14.2077055,13.981348,13.313594,12.31762,12.385528,12.73261,12.947649,12.955194,13.015556,12.713746,12.762791,12.917468,13.196642,13.8719425,14.694374,15.052773,14.720782,13.721037,12.351574,12.019584,13.011784,14.373701,15.098045,14.109617,12.898605,13.192869,13.407909,13.113645,13.019329,12.830698,12.970284,13.268322,13.456953,13.174006,9.895596,10.751981,11.076427,11.710228,12.653384,13.053283,13.241914,12.359119,11.861133,12.128989,12.479843,12.0724,11.02361,10.186088,9.9257765,10.11818,10.114408,10.182315,10.159679,9.861642,9.0807085,9.303293,9.310839,9.488152,9.880505,10.231359,10.499215,10.0465,9.2844305,8.5563135,8.156415,8.20546,8.5563135,8.990166,9.2844305,9.239159,9.333474,9.009028,8.601585,8.216777,7.752744,6.9680386,6.304056,5.832478,5.4250345,4.727099,4.504514,4.7535076,5.0553174,5.160951,4.991183,4.7874613,4.678055,4.4101987,3.9499383,3.5085413,3.4481792,3.731126,3.8254418,3.6028569,3.31991,3.3463185,3.4972234,3.821669,4.353609,5.089271,5.8626595,6.4511886,6.749226,6.851087,7.0774446,7.435844,7.7376537,8.031919,8.201687,7.9715567,8.152642,8.880759,9.439108,9.756008,10.382264,9.623966,9.073163,8.926031,9.016574,8.820397,8.488406,8.114917,7.967784,7.9828744,7.7602897,8.156415,8.318638,8.469543,8.797762,9.435335,10.140816,10.140816,9.899368,9.552286,8.933576,9.220296,9.386291,9.461743,9.612649,10.11818,10.325675,10.419991,10.442626,10.352083,10.020092,10.970794,11.378237,11.627231,11.8045435,11.714001,11.00852,11.219787,11.548005,11.732863,12.027128,11.921495,12.068627,11.812089,11.348056,11.740409,11.680047,11.442371,11.219787,11.200924,11.581959,11.615912,11.7026825,11.823407,12.128989,12.909923,13.268322,13.106099,12.970284,13.166461,13.743673,14.498198,15.098045,15.490398,15.418718,14.43029,12.849561,11.936585,11.378237,11.080199,11.155652,10.974566,11.1631975,10.963248,10.469034,10.627484,10.593531,10.287949,10.125726,10.069136,9.578695,9.680555,10.125726,10.559577,10.846297,11.038701,11.691365,11.529142,11.1782875,10.827434,10.231359,8.548768,7.3453007,6.33801,5.572167,5.409944,5.553304,5.7004366,5.723072,5.59103,5.349582,5.0854983,4.889322,4.5120597,4.032936,3.8971217,3.9725742,4.032936,3.8895764,3.5802212,3.3425457,3.0369632,2.8407867,2.7087448,2.6144292,2.5427492,2.3503454,2.1768045,2.082489,2.0258996,1.8825399,1.4939595,1.177059,1.0450171,1.1695137,1.5958204,1.7995421,1.9957186,2.0145817,1.8259505,1.569412,1.4373702,1.2298758,1.1732863,1.2449663,1.1581959,0.845068,0.59607476,0.513077,0.5772116,0.6375736,0.663982,0.8111144,0.98465514,1.1355602,1.2562841,1.5845025,1.3807807,1.4222796,1.7882242,1.8561316,1.9579924,2.0070364,2.0258996,1.9730829,1.7316349,1.690136,2.0862615,2.6521554,3.0633714,2.9652832,2.5276587,2.173032,1.750498,1.3053282,1.0827434,0.87147635,0.7507524,0.63002837,0.48666862,0.3772625,0.271629,0.34330887,0.452715,0.5772116,0.77716076,0.6073926,0.4678055,0.422534,0.46026024,0.5017591,0.513077,0.6451189,0.77338815,0.8903395,1.0789708,1.2185578,1.2336484,1.8485862,3.0105548,3.8556228,2.6785638,1.5128226,0.88279426,0.79602385,0.7696155,1.116697,0.8941121,0.7205714,0.8224323,1.0299267,1.5543215,3.1840954,3.99521,3.6971724,3.6028569,3.731126,5.081726,5.938112,5.975838,6.255012,4.323428,2.546522,1.5241405,1.4562333,2.1277604,4.90064,5.221313,3.2935016,1.4939595,4.3875628,2.5917933,1.9278114,1.3128735,0.55457586,0.33953625,0.4678055,0.55080324,0.5885295,0.6111652,0.66020936,0.66020936,1.1431054,1.6109109,1.720317,1.2864652,0.8337501,0.543258,0.4074435,0.331991,0.1056335,0.06790725,0.27540162,0.52439487,0.73188925,0.91674787,0.72811663,0.784706,0.84884065,1.0035182,1.6524098,2.2673476,2.3578906,2.2069857,3.0105548,6.8774953,8.68081,9.408927,9.22784,8.820397,9.405154,6.330465,5.8173876,6.1418333,6.319147,6.1418333,6.1003346,6.851087,8.299775,9.601331,9.1825695,9.167479,8.394091,7.805561,7.413208,6.2851934,5.6778007,5.451443,4.8855495,4.327201,5.1835866,5.8400235,5.4250345,5.2364035,5.2967653,4.3800178,5.142088,5.1571784,5.3986263,5.885295,5.692891,6.7567716,6.7114997,6.8397694,7.250985,6.911449,6.4738245,7.141579,7.643338,7.8319697,8.695901,8.854351,8.544995,8.469543,9.144843,10.914205,12.034674,13.249459,10.367173,4.29702,1.0336993,2.2748928,3.3651814,3.8141239,3.8707132,4.5422406,2.6710186,2.757789,2.5767028,1.9957186,2.9803739,3.8103511,9.612649,12.321393,9.948412,6.571913,5.1534057,5.270357,3.9310753,2.897376,8.68081,5.0213637,3.2784111,5.4288073,8.36391,3.8782585,2.4484336,3.500996,4.5799665,4.5196047,3.4594972,4.8666863,5.142088,4.587512,3.531177,2.3126192,6.2814207,7.91874,5.824933,2.8596497,6.145606,5.3571277,4.715781,4.459243,5.5683947,9.782416,12.351574,9.699419,7.2698483,6.971811,7.2057137,6.802043,7.624475,9.1976595,9.978593,7.3377557,6.7152724,8.299775,9.25425,8.733627,7.8810134,7.828197,7.232122,6.221059,6.1041074,9.382519,17.942604,16.837225,10.401127,3.802806,3.0709167,4.7346444,7.586749,9.205205,8.360137,4.991183,4.7950063,5.9720654,7.364164,8.122461,7.7187905,7.4999785,6.270103,5.934339,6.688864,7.0510364,6.900131,7.17176,6.8246784,5.281675,2.4220252,3.3123648,5.3156285,6.6058664,5.7192993,1.5354583,3.1312788,6.9982195,9.367428,8.892077,6.6360474,11.012292,10.853842,10.446399,10.93684,10.367173,9.001483,9.329701,9.420244,8.76758,8.29223,7.1302614,7.6584287,7.835742,7.6923823,9.359882,7.2887115,4.217795,10.155907,20.258997,14.818871,11.861133,9.95973,9.039209,8.428044,6.8699503,7.032173,6.436098,7.145352,8.099826,5.1269975,4.4101987,3.4972234,2.8747404,2.4710693,1.6788181,1.5467763,1.961765,4.606375,7.635793,5.6891184,6.0626082,7.3868,7.277394,5.9532022,6.2436943,6.515323,6.888813,7.111398,6.3945994,3.4066803,2.8445592,5.3458095,7.575431,7.194396,2.837014,3.0030096,3.7537618,4.3309736,4.561104,4.851596,6.858632,8.8769865,10.250222,10.917976,11.423509,11.050018,10.8576145,10.831206,10.502988,8.956212,8.801534,7.6810646,7.009537,7.1302614,7.3188925,7.567886,6.907676,6.4549613,6.4247804,6.126743,5.670255,4.859141,4.093298,5.062863,10.7218,11.102836,8.307321,6.205968,6.096562,6.6850915,4.346064,7.643338,12.015811,14.377474,13.12119,12.0082655,8.763808,7.183078,7.665974,7.220804,6.488915,6.749226,7.1868505,7.4999785,7.914967,7.069899,6.730363,6.247467,5.6363015,5.583485,5.089271,5.7607985,6.439871,6.428553,5.4778514,5.764571,5.6400743,5.553304,5.696664,5.994701,5.8588867,6.319147,6.760544,7.001992,7.284939,6.960493,6.620957,6.25124,6.0776987,6.5643673,6.7454534,6.832224,6.9189944,7.020855,7.032173,7.443389,7.91874,8.303548,8.737399,9.65792,9.533423,9.220296,9.224068,9.514561,9.510788,9.725827,9.967276,10.076681,10.144588,10.47658,11.102836,11.7555,12.698656,14.268067,16.874952,18.79899,17.452164,15.652621,14.622695,14.015302,13.283413,12.815607,12.626976,12.54775,12.196897,12.261031,12.1101265,12.272349,12.593022,12.2270775,12.377983,12.377983,12.030901,11.593277,11.759273,12.585477,12.996693,12.925014,12.381755,11.476325,11.77059,12.200669,12.543978,12.838243,13.355092,13.185325,13.35132,13.539951,13.713491,14.124708,14.977322,15.064092,14.351066,13.223051,12.498707,12.781653,13.8870325,14.807553,14.7736,13.245687,11.759273,12.272349,12.808062,12.770335,12.940104,12.992921,13.275867,13.456953,13.385274,13.113645,9.793735,10.076681,10.310584,10.917976,11.857361,12.626976,13.011784,12.898605,13.158916,13.830443,14.079436,12.54775,11.18206,10.423763,10.31813,10.484125,10.86516,11.442371,11.747954,11.642321,11.310329,11.996947,12.045992,12.012038,12.091263,12.136535,11.955449,11.32542,10.559577,9.940866,9.714509,9.97482,10.11818,10.197406,10.250222,10.299266,10.269085,9.582467,9.009028,8.763808,8.499724,7.5263867,6.7680893,6.047518,5.27413,4.432834,4.466788,4.708236,4.919503,4.919503,4.587512,4.266839,4.0593443,3.682082,3.2482302,3.289729,3.218049,3.3689542,3.4745877,3.4142256,3.2218218,3.338773,3.610402,4.036709,4.5724216,5.1571784,5.907931,6.462507,6.7379084,6.8133607,6.911449,6.9944468,7.220804,7.4207535,7.466025,7.273621,7.4282985,8.141325,8.684583,8.98262,9.612649,9.092027,8.620448,8.329956,8.197914,8.050782,7.6395655,7.4094353,7.3188925,7.333983,7.424526,8.050782,8.322411,8.695901,9.258021,9.748463,10.061591,9.978593,9.812597,9.556059,8.907167,9.288202,9.680555,10.008774,10.265312,10.487898,11.480098,11.544232,11.45369,11.461235,11.310329,12.0233555,12.102581,12.076173,12.189351,12.400619,11.853588,11.8045435,11.872451,11.959221,12.245941,12.0082655,11.940358,11.706455,11.32542,11.148107,10.61994,10.759526,11.087745,11.544232,12.528888,13.313594,13.924759,14.094527,13.996439,14.226569,14.641558,14.811326,14.973549,15.188588,15.365902,15.83748,16.395828,16.546734,16.044973,14.898096,13.460726,12.381755,11.359374,10.559577,10.601076,10.56335,10.944386,11.117926,11.057564,11.348056,11.1782875,10.985884,11.314102,11.812089,11.249968,10.676529,10.502988,10.604849,10.891568,11.32542,12.14408,11.778135,11.261286,10.982111,10.665211,9.390063,8.477088,7.61693,6.79827,6.3455553,6.25124,6.258785,6.0739264,5.6551647,5.2326307,5.191132,5.2288585,4.957229,4.447925,4.2328854,4.3121104,4.398881,4.2706113,3.9273026,3.591539,3.4972234,3.4029078,3.3123648,3.240685,3.218049,3.0520537,2.8332415,2.7502437,2.7653341,2.625747,2.142851,1.7957695,1.750498,1.9994912,2.354118,2.4899325,2.8143783,2.9313297,2.7389257,2.4408884,2.2598023,2.0447628,1.9693103,1.9957186,1.8599042,1.6675003,1.3694628,1.2411937,1.3317367,1.4675511,1.6184561,1.9278114,2.233394,2.463524,2.625747,2.9124665,2.757789,2.71629,2.7879698,2.4371157,2.6031113,2.7200627,2.7200627,2.595566,2.4333432,2.04099,2.354118,2.9954643,3.5085413,3.350091,3.059599,2.6634734,2.1654868,1.6825907,1.4260522,1.0940613,0.9695646,0.814887,0.60362,0.52439487,0.46026024,0.5281675,0.5998474,0.66020936,0.77716076,0.48666862,0.5017591,0.44139713,0.32444575,0.56589377,0.56589377,0.79602385,1.1355602,1.4449154,1.5618668,1.4826416,1.7052265,2.463524,3.451952,3.8141239,2.7313805,1.5769572,0.9242931,0.8299775,0.84884065,1.0299267,1.2185578,1.5505489,1.9164935,1.961765,2.5201135,4.0404816,4.8063245,4.429062,3.8443048,4.847823,6.5568223,6.9491754,5.994701,5.670255,3.3651814,1.539231,1.0902886,1.8297231,2.4974778,6.258785,6.2889657,4.0706625,2.0258996,3.5236318,2.1164427,2.071171,1.6448646,0.66020936,0.47912338,0.633801,0.7809334,0.7997965,0.724344,0.7130261,0.513077,0.59230214,1.1695137,1.7580433,1.1808317,0.6187105,0.44894236,0.41876137,0.33953625,0.08677038,0.05281675,0.16976812,0.4074435,0.62248313,0.5696664,0.58098423,0.7696155,0.7092535,0.58475685,1.20724,2.1315331,2.3880715,2.203213,2.4408884,4.610148,7.383027,7.707473,7.069899,7.115171,9.691874,7.914967,7.0887623,6.549277,6.1229706,6.1041074,6.2663302,5.9682927,6.4549613,7.6018395,7.8998766,7.6093845,7.1679873,6.5530496,5.7381625,4.7120085,4.82896,4.878004,4.4215164,3.7688525,3.9725742,4.776143,4.7836885,4.6554193,4.534695,4.063117,4.2027044,4.2328854,4.5912848,5.0553174,4.715781,5.6476197,5.8098426,6.2021956,6.9755836,7.435844,6.647365,7.111398,7.564113,7.8923316,9.129752,10.499215,9.250477,8.262049,8.571404,9.367428,10.808571,12.619431,10.435081,4.825187,1.2789198,2.173032,2.6106565,3.0369632,3.8782585,5.5306683,3.640583,3.1425967,3.4934506,3.4594972,1.1280149,2.5012503,8.582722,10.170997,6.273875,4.093298,3.4255435,5.798525,5.50426,3.7613072,8.707218,4.821415,3.3651814,4.768598,6.511551,3.138824,1.7731338,2.5012503,3.1425967,3.2255943,3.9989824,3.4029078,4.8855495,5.0025005,3.7575345,4.5950575,6.058836,7.5112963,5.7872066,3.6594462,9.861642,9.016574,5.4703064,2.6031113,2.4220252,5.5797124,15.056546,17.014538,14.354838,9.405154,3.8971217,8.424272,10.008774,9.325929,7.360391,5.413717,7.326438,10.427535,13.189097,14.071891,11.532914,8.952439,7.8734684,6.862405,6.085244,7.3151197,14.019074,18.89708,14.7736,4.961002,3.240685,5.062863,8.703445,11.329193,10.782163,5.5759397,4.7912335,5.243949,6.300284,7.039718,6.221059,6.3455553,5.1458607,6.096562,8.91094,9.525878,7.9489207,5.9305663,4.2102494,2.9841464,1.9164935,2.3616633,4.5761943,7.175533,7.9036493,3.6330378,3.8065786,5.1571784,7.9413757,10.197406,7.756517,11.446144,11.2650585,10.699164,10.906659,10.7218,9.631512,8.744945,8.646856,9.046755,8.797762,7.533932,9.152389,9.473062,8.273367,9.291975,10.106862,7.5490227,8.480861,12.857106,13.777626,10.125726,7.745199,6.8397694,7.0472636,7.4509344,7.7942433,7.2623034,7.043491,7.01331,5.7419353,4.6290107,3.9348478,3.7198083,3.519859,2.3616633,3.218049,4.0480266,6.2097406,8.246958,5.8966126,6.3908267,6.228604,5.594803,5.5797124,8.152642,8.424272,7.2057137,6.2323766,5.4665337,3.0897799,3.5877664,4.983638,4.606375,2.8106055,2.9615107,6.398372,9.989911,8.122461,3.4557245,6.9227667,6.0512905,8.001738,9.756008,10.3634,10.933067,10.79348,10.631257,10.56335,10.325675,9.261794,9.039209,8.114917,7.466025,7.405663,7.575431,7.6282477,6.6813188,6.1644692,6.2889657,6.0362,5.541986,4.9723196,4.6554193,5.832478,10.691619,9.593785,8.816625,9.382519,9.442881,4.315883,2.8785129,10.461489,17.120173,17.923742,12.928786,13.389046,8.341274,5.73439,6.952948,6.85486,6.3153744,6.458734,6.741681,6.964266,7.281166,6.5040054,6.72659,6.647365,5.9984736,5.5457587,5.6853456,6.1003346,6.5530496,6.6662283,5.9418845,5.281675,5.43258,5.692891,5.9418845,6.647365,6.255012,6.4021444,6.7341356,7.1302614,7.6923823,7.3113475,6.862405,6.48137,6.368191,6.7831798,6.779407,6.8359966,7.0585814,7.3000293,7.1604424,7.533932,7.8734684,8.307321,8.929804,9.786189,9.778644,9.26934,8.805306,8.605357,8.563859,8.75249,8.922258,9.009028,9.114662,9.507015,10.186088,10.695392,11.4838705,12.928786,15.335721,17.63325,16.652367,15.184815,14.392565,13.807808,13.038192,12.434572,12.174261,12.121444,11.830952,12.287439,12.053536,11.947904,12.174261,12.321393,12.0233555,11.6008215,11.189606,10.929295,10.989656,11.593277,12.1101265,12.166716,11.649866,10.70671,11.031156,11.529142,12.019584,12.498707,13.128735,13.124963,13.498452,13.81158,13.981348,14.260523,14.735873,14.7736,14.18507,13.445636,13.6833105,14.128481,14.849052,15.105591,14.434063,12.645839,11.25374,11.646093,12.106354,12.185578,12.691111,13.041965,13.415455,13.547497,13.381501,13.0646,8.484633,8.050782,8.616675,9.64283,10.782163,11.898859,12.453435,12.966512,13.93985,15.173498,15.762027,13.675766,12.245941,11.551778,11.348056,11.0613365,11.744182,12.313848,12.362892,12.068627,12.200669,12.894833,12.943876,12.562841,12.049765,11.793225,11.25374,11.02361,11.174516,11.487643,11.457462,11.506506,11.012292,10.480352,10.220041,10.352083,10.472807,9.978593,9.439108,9.125979,8.990166,7.6508837,7.001992,6.258785,5.281675,4.587512,4.2592936,4.3347464,4.436607,4.3196554,3.8707132,3.5651307,3.308592,2.9652832,2.8143783,3.5462675,3.5575855,3.451952,3.5349495,3.7198083,3.5538127,3.591539,3.9725742,4.3724723,4.6931453,5.0553174,5.7796617,6.168242,6.326692,6.375736,6.4210076,6.56814,6.900131,7.0774446,7.0472636,7.0585814,7.281166,7.7376537,8.137552,8.473316,9.046755,8.654402,8.186596,7.8319697,7.77538,8.167733,7.54525,7.333983,7.2924843,7.435844,8.031919,8.52236,8.52236,8.778898,9.21275,8.952439,8.82417,8.914713,9.163706,9.25425,8.590267,9.016574,9.759781,10.495442,10.917976,10.748209,12.291212,12.3289385,12.242168,12.551523,12.921241,12.445889,12.106354,12.019584,12.196897,12.559069,12.728837,12.611885,12.453435,12.396846,12.47607,12.310076,11.766817,11.378237,11.083972,10.235131,9.748463,10.393582,11.589504,12.985375,14.449154,15.648849,16.146835,15.961976,15.39231,15.015047,15.558306,16.131744,16.467508,16.493916,16.343012,16.24115,16.101564,15.4074,14.339747,13.773854,13.396591,12.54775,11.400873,10.412445,10.329447,10.38981,10.736891,11.155652,11.581959,12.128989,11.966766,11.887542,12.468526,13.257004,12.751472,11.978085,11.476325,11.1782875,11.117926,11.415963,12.098808,11.657412,11.16697,11.00852,10.861387,10.442626,9.680555,8.922258,8.194141,7.224577,6.628502,6.458734,6.1795597,5.674028,5.2552667,5.4174895,5.5268955,5.3684454,4.9760923,4.640329,4.8553686,4.878004,4.719554,4.38379,3.8480775,3.7613072,3.6481283,3.5538127,3.519859,3.5764484,3.4783602,3.31991,3.2670932,3.2859564,3.127506,2.806833,2.6144292,2.757789,3.150142,3.4029078,3.4557245,3.7009451,3.8065786,3.6707642,3.429316,3.2633207,3.1840954,3.1727777,3.1765501,3.1048703,2.987919,2.7426984,2.6936543,2.886058,3.0709167,3.3689542,3.7650797,4.164978,4.4743333,4.606375,4.6818275,4.817642,4.7044635,4.217795,3.3764994,3.5123138,3.3764994,3.2369123,3.1840954,3.138824,2.5087957,2.6521554,3.1312788,3.572676,3.6481283,3.712263,3.2633207,2.7011995,2.2296214,1.8674494,1.3958713,1.3166461,1.1883769,0.91297525,0.72811663,0.7205714,0.7922512,0.80734175,0.754525,0.7432071,0.27917424,0.573439,0.63002837,0.35085413,0.51684964,0.513077,0.8526133,1.4562333,1.991946,1.8599042,1.7240896,2.2371666,3.0520537,3.6292653,3.229367,2.6332922,1.6750455,1.0299267,0.98842776,1.4600059,2.1390784,2.463524,2.9501927,3.4444065,3.127506,3.942393,5.0062733,5.764571,5.73439,4.5120597,6.9227667,7.492433,6.7379084,5.4250345,4.5724216,2.8143783,1.5203679,1.5354583,2.5804756,3.2557755,4.115934,6.0248823,5.160951,2.3013012,2.806833,1.720317,2.535204,2.2711203,0.77716076,0.7469798,1.1053791,1.3392819,1.2902378,1.0148361,0.77716076,0.5017591,0.31312788,0.814887,1.6373192,1.4109617,0.6187105,0.4376245,0.43385187,0.35462674,0.14335975,0.14335975,0.2263575,0.4678055,0.6488915,0.271629,0.38103512,0.6375736,0.7167987,0.7582976,1.3505998,2.4786146,2.916239,2.4710693,1.5958204,1.4034165,4.6214657,4.7874613,3.9084394,4.3347464,8.737399,8.409182,8.213005,6.911449,5.2062225,5.764571,6.436098,5.80607,5.564622,6.1116524,6.5756855,6.700182,6.175787,5.1458607,4.0782075,3.7386713,3.7952607,3.7688525,3.6292653,3.2746384,2.5238862,3.1350515,3.6028569,3.5877664,3.270866,3.308592,3.3236825,3.663219,4.1272516,4.4705606,4.3875628,4.821415,5.172269,5.855114,6.828451,7.5716586,6.820906,7.0359454,7.360391,7.779153,9.129752,12.15917,10.56335,8.612903,8.073418,8.209232,10.567122,11.955449,10.306811,5.994701,1.8448136,3.0445085,2.5427492,1.7354075,2.41448,6.8058157,4.779916,2.4559789,3.350091,5.4250345,1.0789708,1.1129243,2.6672459,2.897376,2.0447628,3.4557245,2.5578396,4.508287,5.0666356,4.821415,9.193887,5.0477724,3.1350515,3.1312788,4.0404816,4.1536603,2.4484336,3.731126,4.6026025,4.847823,7.435844,7.1038527,7.9828744,7.598067,6.673774,9.103344,4.768598,5.462761,5.594803,5.7872066,12.902377,14.351066,9.435335,4.183841,1.7844516,2.565385,16.448645,21.036158,18.912169,12.804289,5.5985756,13.936077,15.1395445,12.355347,8.299775,5.2665844,8.654402,12.570387,16.90136,19.90437,18.18028,12.344029,9.948412,8.646856,6.9869013,4.4139714,4.772371,13.59654,13.985121,5.3759904,3.5349495,3.3538637,7.84706,11.212241,10.480352,5.523123,3.874486,3.7198083,4.183841,4.52715,4.142342,5.511805,4.4177437,5.904158,10.174769,12.619431,8.937348,5.43258,3.6556737,3.3953626,2.6597006,3.180323,5.794752,8.122461,8.60913,6.5455046,6.620957,5.855114,7.914967,11.664956,11.174516,12.004493,11.378237,10.842525,10.487898,8.937348,10.744436,10.4049,9.156161,8.118689,8.288457,7.8696957,10.921749,11.7894535,9.955957,10.035183,13.287186,11.747954,7.5490227,3.4179983,2.6710186,2.6031113,3.9688015,5.5457587,6.168242,4.7346444,6.9189944,9.208978,10.110635,9.310839,7.677292,6.458734,5.270357,5.240176,5.534441,3.3915899,5.4288073,6.6058664,6.937857,6.8058157,6.9454026,7.9941926,6.85486,6.0512905,6.7379084,8.695901,9.861642,8.280911,5.9230213,4.187614,3.893349,4.0970707,3.3878171,2.203213,1.358145,2.071171,11.374464,19.195116,14.70192,4.0103,10.163452,7.073672,7.232122,8.397863,9.352338,9.922004,10.725573,10.77839,10.759526,10.782163,10.397354,9.597558,8.899622,8.20546,7.7037,7.8810134,8.0206,6.9755836,6.356873,6.5002327,6.4738245,5.7192993,5.0968165,4.7120085,5.511805,9.265567,7.254758,8.492179,10.650121,11.185833,7.333983,3.8480775,10.33322,17.84829,19.123436,8.52236,15.641303,9.276885,5.1269975,6.9567204,6.5832305,6.273875,6.360646,6.4474163,6.3644185,6.187105,5.855114,6.3417826,6.628502,6.319147,5.643847,6.571913,6.466279,6.247467,6.1795597,5.885295,4.8629136,5.3458095,5.975838,6.3644185,7.073672,6.6360474,6.519096,6.6020937,6.8661776,7.3792543,7.4697976,7.092535,6.692637,6.48137,6.4436436,6.360646,6.673774,7.0774446,7.3679366,7.443389,8.273367,8.420499,8.699674,9.22784,9.416472,9.540969,9.352338,9.020347,8.646856,8.235641,7.858378,7.7187905,7.854605,8.265821,8.937348,9.540969,10.038955,10.695392,11.717773,13.238141,15.611122,16.063837,15.814844,15.290449,14.143571,12.989148,12.257258,12.027128,12.162943,12.298758,12.385528,12.193124,11.993175,11.996947,12.344029,12.185578,11.536687,10.944386,10.672756,10.695392,11.129244,11.457462,11.302785,10.627484,9.725827,10.103089,10.7557535,11.374464,11.830952,12.166716,12.47607,13.019329,13.528633,13.902123,14.2077055,14.068119,13.992666,13.902123,14.132254,15.403628,15.524352,15.482853,15.143317,14.226569,12.298758,11.332966,11.442371,11.570641,11.619685,12.46098,12.781653,13.094781,13.328684,13.340002,12.909923,8.299775,8.582722,8.726082,9.49947,10.774617,11.521597,12.095036,12.174261,12.619431,13.626721,14.724555,14.347293,13.445636,12.664702,12.162943,11.61214,12.08749,11.099063,10.140816,9.661693,9.065618,9.016574,9.295748,9.608876,10.050273,11.125471,11.551778,11.329193,11.419736,11.774363,11.321648,10.49167,9.782416,9.34102,9.205205,9.276885,9.691874,10.382264,10.33322,9.673011,9.673011,8.296002,7.7112455,7.1679873,6.247467,4.8666863,4.304565,4.112161,4.006528,3.7348988,3.0520537,2.8936033,2.6144292,2.5427492,2.727608,2.9615107,3.4972234,3.6141748,3.4594972,3.2255943,3.127506,3.8480775,4.5233774,4.8138695,4.9232755,5.5683947,5.617439,5.8211603,6.1418333,6.507778,6.8359966,6.8359966,6.8925858,6.8661776,6.900131,7.4018903,7.7301087,7.7376537,7.6282477,7.4999785,7.3377557,6.9869013,6.760544,6.802043,7.1566696,7.7678347,7.865923,7.696155,7.586749,7.677292,7.9338303,8.52236,9.205205,9.42779,8.914713,7.707473,7.364164,8.065872,8.809079,8.98262,8.345046,8.273367,9.107117,9.880505,10.246449,10.469034,11.348056,12.196897,12.717519,12.970284,13.396591,13.128735,12.943876,12.864652,12.826925,12.679792,12.166716,12.076173,11.778135,11.242422,11.046246,10.997202,11.042474,11.144334,11.310329,11.566868,11.725319,12.404391,13.917213,15.731846,16.463736,16.501461,15.777118,14.928277,14.5132885,15.015047,15.8676605,15.826162,15.528125,15.475307,16.03743,15.328176,14.558559,13.65313,12.932558,13.091009,12.468526,11.506506,11.136789,11.159425,10.269085,10.121953,10.725573,11.495189,12.042219,12.178034,12.83447,12.872196,12.513797,12.102581,12.113899,12.543978,12.50248,12.245941,12.015811,12.038446,12.370438,12.479843,12.37421,12.264804,12.559069,12.178034,11.140562,10.001229,9.0807085,8.469543,7.1000805,6.477597,6.1229706,5.80607,5.523123,5.7909794,5.915476,5.828706,5.583485,5.3269467,5.2288585,5.149633,4.9949555,4.749735,4.4705606,4.191386,3.9084394,3.8971217,4.0178456,3.7235808,3.5764484,3.5953116,3.7047176,3.7990334,3.7386713,3.7386713,3.8103511,3.9461658,4.134797,4.3800178,4.4403796,4.3007927,4.146115,4.0782075,4.0895257,4.1762958,4.2328854,4.2328854,4.2291126,4.3649273,4.5120597,4.4818783,4.82896,5.4740787,5.7079816,5.938112,6.2436943,6.620957,6.888813,6.6662283,6.8133607,7.1981683,7.0170827,6.1078796,4.9760923,4.7308717,4.183841,3.651901,3.380272,3.5387223,2.9916916,3.2105038,3.6330378,3.9159849,3.953711,4.134797,3.6481283,3.1539145,2.746471,1.9542197,1.6486372,1.5807298,1.3619176,0.9695646,0.76207024,0.8865669,1.0902886,1.1883769,1.2298758,1.50905,0.52062225,0.3772625,0.44139713,0.4678055,0.56589377,0.94315624,1.0827434,1.4675511,2.022127,2.1051247,2.886058,2.9539654,3.31991,3.9612563,3.8141239,3.0822346,2.2598023,1.7655885,1.8976303,2.837014,4.436607,4.727099,4.715781,4.606375,3.7990334,5.873977,6.5568223,6.907676,7.062354,6.255012,9.088254,6.3719635,3.893349,3.6556737,3.874486,1.8863125,1.7919968,1.9089483,1.780679,2.1805773,1.9881734,6.2663302,6.058836,1.8787673,3.7235808,2.686109,4.093298,3.2972744,0.45648763,0.5017591,1.5543215,2.071171,2.1277604,1.7165444,0.77716076,0.47157812,0.3055826,0.6790725,1.4449154,1.9240388,0.7997965,0.5281675,0.47912338,0.39989826,0.41121614,0.46026024,0.5998474,0.6752999,0.663982,0.68661773,0.4074435,0.30935526,0.44139713,0.8865669,1.7391801,2.886058,3.4859054,2.8936033,1.720317,1.8297231,2.8822856,3.610402,3.8367596,4.587512,8.103599,9.2995205,7.748972,6.4474163,6.0324273,4.776143,5.1043615,5.270357,4.9534564,4.561104,5.2326307,5.1232247,4.768598,4.4630156,4.447925,4.8968673,3.138824,2.7389257,2.7917426,2.7804246,2.546522,2.4861598,3.0407357,3.5387223,3.4896781,2.565385,3.270866,4.1083884,4.504514,4.3875628,4.1800685,4.353609,4.9345937,5.6476197,6.2663302,6.6058664,6.7152724,7.33021,7.752744,7.835742,7.9791017,10.921749,12.351574,11.053791,8.246958,7.598067,9.076936,10.884023,10.008774,6.326692,2.5804756,3.5802212,3.682082,2.8596497,1.8146327,1.9844007,3.1425967,1.9957186,1.2147852,1.4713237,1.4335974,1.2034674,3.361409,4.353609,3.6858547,3.904667,5.2854476,3.1048703,1.8599042,3.1539145,5.692891,4.983638,3.8895764,3.2029586,2.9954643,2.6408374,1.7844516,3.3651814,6.5530496,9.231613,8.009283,10.891568,12.491161,13.728582,14.203933,12.193124,5.5495315,8.944894,10.231359,7.5792036,9.461743,14.25675,12.178034,7.2170315,3.8480775,7.032173,5.534441,6.9152217,8.575176,9.371201,9.627739,14.011529,14.475562,12.875969,10.137043,6.255012,10.797253,15.731846,18.350048,19.87796,25.480309,16.022339,12.091263,10.638803,9.175024,5.7683434,3.3123648,4.112161,4.429062,3.3274553,2.655928,3.169005,6.7643166,9.231613,8.880759,6.560595,3.742444,2.9615107,3.4029078,3.99521,3.4330888,5.251494,4.5799665,5.406172,8.235641,10.11818,7.432071,5.221313,4.696918,5.564622,6.043745,6.092789,6.828451,7.816879,8.20546,6.730363,9.989911,9.156161,10.804798,13.932304,9.978593,10.272858,11.012292,12.166716,12.234623,8.254503,8.83926,10.012547,10.751981,10.691619,10.133271,9.544742,8.484633,9.288202,10.450171,6.590776,6.1531515,6.4738245,5.873977,4.353609,3.5839937,5.4891696,7.33021,8.544995,8.484633,6.40969,5.1647234,5.0439997,5.251494,5.2137675,4.5761943,3.9914372,4.3121104,4.4630156,4.610148,6.149379,6.330465,7.6584287,8.103599,7.3000293,6.530414,7.484888,8.141325,8.2507305,7.466025,5.342037,7.488661,7.432071,6.515323,5.8966126,6.530414,5.492942,4.115934,3.2557755,3.1576872,3.4632697,3.0369632,6.0626082,7.17176,5.2062225,3.2067313,7.537705,5.9192486,5.3910813,7.7112455,9.382519,10.325675,10.438853,10.616167,10.948157,10.725573,9.895596,9.590013,9.110889,8.431817,8.16396,8.616675,7.7225633,7.1340337,7.0963078,6.4247804,5.775889,5.6778007,4.5497856,4.274384,10.193633,8.692128,10.816116,8.2507305,2.6483827,5.5985756,2.535204,3.7462165,9.963503,16.7995,14.784918,17.70493,9.937095,5.3344917,6.8397694,6.485142,6.349328,6.417235,6.307829,5.8702044,5.172269,5.221313,5.772116,6.379509,6.5568223,5.8136153,6.205968,6.4474163,6.4738245,6.1418333,5.2628117,5.3759904,5.6400743,6.092789,6.8058157,7.9036493,7.3792543,6.8359966,6.8435416,7.2698483,7.2924843,7.8432875,7.484888,6.971811,6.7152724,6.7756343,6.40969,6.8397694,7.364164,7.6886096,7.91874,8.114917,8.265821,8.567632,8.975075,9.171251,9.073163,9.333474,9.318384,8.726082,7.5527954,7.515069,7.54525,7.6282477,7.6886096,7.567886,7.8131065,8.7600355,9.880505,10.8576145,11.627231,13.336229,14.962231,16.22606,16.475054,14.694374,13.460726,12.943876,12.600568,12.151625,11.566868,11.857361,12.498707,12.3289385,11.574413,11.857361,11.989402,11.940358,11.057564,9.65792,9.046755,9.842778,9.748463,9.273112,8.907167,9.14107,10.627484,11.59705,12.083718,12.095036,11.581959,11.898859,12.2270775,12.694883,13.185325,13.306048,13.000465,12.521342,12.864652,14.252977,16.158154,15.988385,15.580941,15.131999,14.362384,12.479843,11.747954,11.61214,11.714001,12.034674,12.864652,12.570387,12.223305,12.385528,12.872196,12.725064,7.9338303,8.058327,8.311093,9.359882,10.899114,11.653639,12.249713,12.721292,13.113645,13.192869,12.464753,11.465008,10.985884,10.861387,10.95193,11.125471,11.02361,10.336992,9.688101,9.303293,9.027891,9.152389,9.81637,10.49167,11.125471,12.098808,13.192869,12.423254,10.9594755,9.714509,9.367428,9.224068,9.378746,9.759781,10.435081,11.634775,11.785681,11.449917,10.555805,9.552286,9.405154,8.201687,7.515069,7.250985,6.9755836,5.9305663,5.455216,4.6742826,3.8480775,3.2067313,2.9539654,3.0897799,2.927557,2.7238352,2.6710186,2.9124665,3.2444575,3.4783602,3.5500402,3.5538127,3.7386713,4.164978,4.8629136,5.2854476,5.5457587,6.387054,6.964266,6.779407,6.3832817,6.145606,6.2625575,6.2927384,6.2889657,6.360646,6.6322746,7.24344,7.092535,6.651138,6.2021956,6.006019,6.326692,6.6360474,7.141579,7.352846,7.2924843,7.4735703,7.2962565,7.356619,7.8206515,8.382772,8.239413,8.98262,9.450426,9.276885,8.590267,8.047009,8.016829,8.571404,8.993938,9.159933,9.529651,9.963503,10.970794,11.691365,11.947904,12.238396,12.706201,13.65313,14.547242,14.943368,14.483108,14.6151495,14.667966,14.339747,13.63804,12.875969,12.381755,11.996947,11.472552,10.872705,10.559577,11.046246,11.415963,11.812089,12.185578,12.287439,12.427027,12.370438,12.83447,13.50977,13.072145,14.083209,14.988639,15.24895,15.120681,15.660167,15.55076,14.992412,14.947141,15.494171,15.841252,15.339493,14.93205,14.237886,13.313594,12.653384,12.664702,12.264804,12.234623,12.845788,13.86817,12.785426,12.864652,13.204187,13.2607765,12.849561,12.600568,12.751472,12.623203,12.287439,12.593022,12.853333,13.04951,13.200415,13.268322,13.174006,13.249459,13.158916,13.272095,13.8719425,15.120681,15.173498,14.286931,13.011784,11.555551,9.763554,7.9941926,6.952948,6.221059,5.643847,5.353355,5.1534057,5.1798143,5.142088,4.98741,4.8855495,4.7572803,4.708236,4.5497856,4.2592936,3.9574835,3.874486,3.874486,3.9650288,4.0291634,3.832987,4.036709,4.327201,4.4139714,4.2404304,3.99521,3.9273026,4.0706625,4.3083377,4.644101,5.2099953,5.20245,5.3156285,5.2250857,5.05909,5.3948536,5.2967653,5.0213637,4.8327327,4.745962,4.561104,5.194905,5.8513412,6.485142,6.9793563,7.17176,7.375482,7.9941926,8.582722,8.831716,8.582722,7.8810134,7.7678347,7.647111,7.062354,5.6815734,5.409944,4.8629136,4.4139714,4.1989317,4.112161,4.568649,4.3686996,4.164978,4.1536603,4.074435,4.38379,3.9801195,3.451952,2.9501927,2.1956677,1.6486372,1.5845025,1.7316349,1.8599042,1.7995421,1.4147344,1.0601076,1.0827434,1.3732355,1.3392819,0.6526641,0.5017591,0.5885295,0.80356914,1.2223305,1.3770081,1.086516,1.2525115,1.9164935,2.2748928,2.8030603,3.1652324,3.6141748,4.172523,4.6214657,3.5575855,3.3651814,3.7499893,4.4215164,5.1081343,6.598321,5.9192486,5.300538,5.2779026,4.678055,5.3382645,7.066127,8.307321,8.60913,8.624221,10.627484,9.152389,7.1906233,5.59103,3.0445085,1.3996439,1.3091009,2.6219745,5.534441,10.604849,5.4891696,5.515578,4.745962,2.5993385,3.8443048,3.802806,2.7879698,1.6184561,0.8978847,1.0148361,2.0560806,2.4408884,2.354118,1.871222,0.9507015,0.7507524,0.55080324,0.7809334,1.3392819,1.5807298,1.2110126,0.84884065,0.52062225,0.331991,0.47157812,0.8941121,1.0827434,0.90543,0.58098423,0.663982,0.34330887,0.23390275,0.39989826,1.1016065,2.8143783,3.4444065,3.8254418,3.0520537,1.7127718,1.8938577,2.2484846,3.0445085,3.6028569,4.1197066,5.66271,6.40969,6.511551,6.1833324,5.353355,3.6669915,4.1612053,4.7610526,4.7006907,4.1197066,4.085753,3.6934,3.4330888,3.2218218,3.2557755,4.032936,3.7273536,3.7273536,3.6254926,3.4029078,3.4142256,3.2670932,3.591539,3.863168,3.9273026,4.0178456,4.6931453,5.2892203,5.6476197,5.775889,5.8513412,5.5080323,6.039973,6.511551,6.670001,6.971811,7.1906233,7.567886,8.216777,8.846806,8.748717,10.978339,12.921241,12.468526,10.140816,9.076936,8.669493,10.295494,10.269085,7.564113,3.8367596,3.5877664,5.2250857,6.115425,5.4476705,4.2404304,4.9232755,2.9539654,1.1996948,0.7696155,1.0072908,5.070408,8.296002,7.3151197,3.6934,3.942393,4.617693,4.6629643,4.557331,4.323428,3.531177,4.561104,7.858378,8.235641,5.775889,5.802297,5.6891184,6.643593,7.6395655,8.929804,12.015811,16.720274,15.856343,15.399856,16.388283,14.901869,14.128481,12.883514,9.64283,6.0362,6.8133607,6.4549613,4.7572803,3.3689542,3.1652324,4.2517486,6.5002327,4.9949555,4.044254,4.6214657,4.3800178,5.1081343,5.994701,6.7039547,6.7152724,5.304311,9.522105,12.178034,16.565596,21.711456,22.394302,15.82239,11.61214,10.487898,10.906659,9.061845,5.7306175,6.6813188,6.330465,3.772625,2.7879698,5.353355,7.3981175,8.5563135,8.409182,6.5002327,4.304565,2.6219745,2.837014,4.0103,2.8822856,5.670255,4.183841,3.3840446,4.8855495,6.9793563,6.7454534,6.0776987,5.3571277,5.089271,5.8966126,8.4544525,8.043237,7.8998766,8.744945,8.790216,9.510788,10.095545,10.193633,10.220041,11.321648,11.144334,11.208468,11.604594,11.717773,10.220041,10.065364,10.714255,10.763299,10.18986,10.352083,10.850069,10.080454,10.9594755,13.302276,13.819125,11.336739,8.986393,7.2170315,6.187105,5.772116,6.934085,6.1795597,6.149379,7.5527954,9.178797,9.21275,8.805306,8.8618965,8.933576,7.213259,6.4926877,7.2170315,7.360391,6.9152217,7.907422,7.6810646,8.254503,7.8923316,6.692637,6.56814,6.5530496,6.5455046,7.3717093,8.461998,7.8319697,8.367682,7.3717093,6.221059,5.617439,5.5797124,5.938112,4.821415,3.399135,2.7011995,3.610402,7.303802,5.828706,6.7379084,9.963503,7.7942433,4.1197066,2.1579416,3.169005,6.462507,9.397609,9.371201,9.87296,10.827434,11.46878,10.359629,10.095545,9.548513,9.307066,9.239159,8.480861,8.228095,7.907422,7.6584287,7.3415284,6.5341864,5.485397,5.010046,3.9989824,2.9086938,3.7613072,9.797507,9.95973,8.375228,7.0887623,6.089017,3.8065786,4.0782075,5.983383,8.582722,10.902886,11.566868,6.8246784,5.1081343,7.333983,6.900131,6.043745,6.1342883,6.360646,6.168242,5.247721,5.138315,5.3458095,5.5268955,5.775889,6.5945487,6.349328,6.5228686,6.3644185,5.8098426,5.4967146,5.5382137,5.4401255,6.1041074,7.4735703,8.552541,8.552541,8.186596,7.7150183,7.33021,7.1604424,7.3868,7.3377557,6.952948,6.5643673,6.907676,7.01331,7.2358947,7.273621,7.1981683,7.466025,7.605612,7.7829256,8.2507305,8.952439,9.537196,9.261794,8.446907,7.9300575,7.756517,7.164215,7.164215,7.3868,7.073672,6.3153744,6.006019,7.039718,7.5565677,8.084735,8.850578,9.797507,10.917976,11.944131,13.309821,14.649103,14.781145,14.93205,14.622695,13.826671,12.759018,11.857361,11.419736,10.816116,10.616167,11.159425,12.551523,11.876224,11.808316,11.529142,10.589758,8.914713,9.239159,9.042982,8.83926,8.91094,9.2995205,9.820143,10.819888,11.589504,11.774363,11.348056,11.529142,11.133017,11.204697,11.857361,12.279895,13.060828,13.445636,13.645585,14.109617,15.535669,15.599804,14.735873,14.25675,14.079436,12.736382,11.574413,10.9594755,10.657665,10.808571,11.910177,12.057309,11.283921,11.2801485,12.30253,13.189097,9.125979,8.967529,8.91094,9.616421,10.850069,11.461235,12.298758,13.600313,13.81158,12.593022,10.819888,10.246449,9.87296,9.789962,9.967276,10.269085,9.880505,9.933322,9.805053,9.371201,9.046755,9.522105,10.54826,11.136789,11.068882,10.906659,11.16697,10.269085,9.276885,8.756263,8.7600355,9.393836,10.061591,10.744436,11.415963,12.030901,11.208468,10.174769,9.220296,8.695901,9.016574,8.458225,7.8696957,7.752744,7.828197,7.0548086,6.0701537,5.0175915,4.112161,3.482133,3.2029586,3.1048703,2.9501927,2.837014,2.8219235,2.9351022,3.2444575,3.519859,3.8292143,4.1498876,4.38379,4.689373,5.119452,5.5985756,6.198423,7.141579,7.2698483,6.971811,6.579458,6.277648,6.0814714,6.009792,6.0512905,6.1003346,6.330465,7.183078,7.4735703,7.194396,6.700182,6.307829,6.330465,6.696409,7.152897,7.3151197,7.111398,6.7680893,6.8171334,7.3151197,8.00551,8.669493,9.148616,9.476834,9.81637,10.001229,9.986138,9.835234,9.929549,10.159679,10.518079,11.042474,11.812089,12.872196,13.79649,14.535924,14.977322,14.924504,15.384765,15.701665,16.026112,16.173243,15.652621,15.679029,15.603577,15.369675,14.867915,13.920986,12.90615,12.0233555,11.197151,10.578441,10.529396,11.099063,11.661184,12.193124,12.468526,12.045992,11.917723,11.729091,12.064855,12.657157,12.415709,13.943622,15.475307,16.075155,15.882751,16.116653,15.799753,15.690348,16.03743,16.678776,17.037174,16.42601,16.033657,15.324403,14.611377,15.041456,14.320885,14.249205,14.505743,14.611377,13.936077,13.79649,13.422999,13.234368,13.219278,12.932558,13.336229,13.392818,13.36641,13.324911,13.132507,13.249459,13.445636,13.679539,13.875714,13.951167,13.905896,13.79649,14.139798,14.924504,15.607349,15.697892,15.049001,13.898351,12.396846,10.589758,9.133525,7.9262853,6.9567204,6.255012,5.904158,5.4250345,5.119452,4.8553686,4.6516466,4.6931453,4.610148,4.496969,4.3196554,4.063117,3.731126,3.6783094,3.6594462,3.802806,4.0291634,4.063117,3.8292143,3.9612563,4.183841,4.217795,3.7462165,4.014073,3.8971217,3.8707132,4.2517486,5.168496,5.643847,6.115425,6.119198,5.824933,6.043745,5.8966126,5.704209,5.73439,5.915476,5.8513412,6.477597,7.152897,7.7187905,8.126234,8.461998,8.722309,9.514561,10.280403,10.585986,10.11818,9.35611,8.6732645,8.424272,8.194141,6.7831798,6.0626082,5.4476705,4.961002,4.640329,4.5309224,4.696918,4.7421894,4.776143,4.7912335,4.67051,4.9345937,4.436607,3.7914882,3.2255943,2.6068838,2.003264,1.6071383,1.7089992,2.071171,1.9504471,1.7316349,1.7467253,1.9278114,2.033445,1.6825907,1.0186088,0.8337501,0.7884786,0.84129536,1.2223305,1.7957695,1.6335466,1.7995421,2.3692086,2.4371157,2.5804756,3.0897799,3.5424948,3.85185,4.2819295,4.1612053,4.104616,4.3913355,4.9987283,5.621211,6.25124,4.881777,3.942393,4.346064,5.5004873,6.1795597,7.394345,8.903395,10.321902,11.121698,11.019837,8.650629,5.783434,3.5160866,2.2786655,2.5389767,1.9089483,2.2258487,4.919503,10.989656,7.726336,7.1340337,5.4665337,2.7917426,2.9954643,3.4670424,1.9089483,0.9280658,1.1053791,0.9997456,2.3428001,2.9313297,2.7841973,2.1843498,1.6788181,1.3543724,0.9205205,0.72811663,0.8299775,0.9808825,1.1204696,0.8903395,0.5583485,0.32067314,0.2867195,0.6526641,0.87902164,0.7696155,0.49044126,0.56589377,0.271629,0.47912338,1.0223814,1.6825907,2.1654868,1.9730829,2.1466236,1.8976303,1.297783,1.2940104,1.5505489,1.841041,3.1840954,5.0477724,5.342037,5.624984,5.8966126,5.2175403,3.62172,2.0975795,3.4632697,4.2819295,4.115934,3.4670424,3.7801702,3.0105548,2.9049213,2.8143783,2.8219235,3.7499893,3.5349495,3.99521,4.1083884,3.7914882,3.92353,4.2819295,4.1008434,4.146115,4.561104,4.8742313,5.492942,5.9607477,6.2814207,6.651138,7.435844,7.1264887,7.333983,7.9300575,8.469543,8.190369,8.141325,8.254503,8.529905,9.280658,11.129244,11.736636,11.321648,10.95193,11.299012,12.630749,9.439108,11.004747,12.185578,10.412445,5.6778007,4.3121104,4.22534,5.2628117,6.296511,5.247721,5.983383,5.8400235,4.508287,2.595566,1.6033657,4.395108,5.9192486,5.172269,3.7348988,5.764571,6.4474163,6.85486,6.2436943,4.719554,3.229367,5.7419353,8.36391,7.7338815,4.9119577,5.402399,6.3908267,8.190369,8.843033,8.175279,7.798016,10.367173,10.246449,10.220041,10.250222,7.5037513,8.397863,8.473316,9.125979,10.533169,11.631002,8.627994,6.270103,5.0251365,4.357382,2.7238352,5.0439997,5.13077,5.2099953,6.25124,7.964011,8.880759,9.242931,8.465771,6.9189944,5.926794,9.024119,10.567122,12.838243,15.660167,16.38451,11.891314,10.140816,10.382264,11.631002,12.653384,9.473062,9.865415,8.235641,4.1989317,2.5578396,4.3649273,6.33801,7.6207023,8.073418,8.288457,6.617184,3.8782585,3.772625,5.221313,2.4069347,5.692891,4.266839,3.138824,4.5120597,7.786698,7.654656,7.405663,7.8432875,8.035691,5.311856,8.348819,9.186342,9.57115,10.042727,9.948412,10.699164,11.193378,10.533169,9.661693,11.363147,11.306557,11.480098,11.099063,10.310584,10.197406,10.310584,10.570895,10.70671,10.582213,10.178542,9.839006,9.424017,9.635284,10.714255,12.419481,10.808571,9.559832,8.390318,7.1906233,6.043745,7.062354,7.0812173,7.020855,7.33021,7.967784,8.050782,8.175279,8.495952,8.66572,7.816879,8.439363,9.103344,9.159933,8.688355,8.511042,8.8618965,8.329956,7.3113475,6.790725,8.3525915,9.597558,9.261794,8.827943,8.710991,8.231868,7.3415284,6.4436436,6.221059,6.4474163,5.9984736,6.1305156,5.9909286,4.938366,3.308592,2.4031622,5.6778007,5.070408,5.1081343,7.8244243,12.766563,3.591539,1.1581959,2.7087448,6.009792,9.390063,8.888305,9.567377,10.691619,11.257513,9.993684,9.725827,9.510788,9.540969,9.5183325,8.669493,8.190369,8.239413,8.114917,7.6282477,7.092535,5.745708,4.7874613,3.9348478,3.2746384,3.240685,7.1264887,9.186342,10.838752,11.321648,7.673519,4.2027044,4.353609,5.6891184,6.8171334,7.3981175,6.907676,5.100589,5.4891696,7.647111,7.1868505,5.9796104,5.5985756,5.8400235,6.0701537,5.2099953,5.040227,5.040227,5.138315,5.5268955,6.670001,6.3342376,6.270103,5.7683434,5.1081343,5.5457587,5.6853456,6.0248823,6.7077274,7.6886096,8.710991,9.103344,8.971302,8.488406,7.84706,7.24344,7.2660756,7.443389,7.4282985,7.220804,7.1793056,7.284939,7.2962565,7.17176,6.964266,6.8435416,7.2057137,7.6282477,8.058327,8.529905,9.171251,9.118435,8.103599,7.2170315,6.851087,6.7077274,6.4926877,6.7831798,6.63982,6.066381,5.9909286,6.4549613,6.851087,7.213259,7.7640624,8.937348,9.737145,10.235131,11.019837,12.076173,12.770335,14.426518,14.852824,14.124708,12.838243,12.08749,11.427281,10.401127,9.910686,10.529396,12.487389,11.544232,11.1631975,11.140562,11.027383,10.133271,9.903141,9.774872,9.812597,9.929549,9.895596,9.937095,10.533169,11.200924,11.5857315,11.4838705,11.491416,11.053791,11.053791,11.54046,11.747954,12.1252165,12.683565,12.600568,12.411936,14.02662,14.837734,13.928532,13.124963,12.860879,12.189351,11.717773,11.072655,10.401127,10.125726,10.978339,11.7894535,11.6008215,11.400873,11.608367,12.049765,10.642575,9.778644,9.752235,10.216269,10.770844,10.948157,11.502733,12.623203,12.577931,11.11038,9.454198,9.6051035,9.408927,9.231613,9.261794,9.537196,9.450426,9.8239155,9.95973,9.676784,9.314611,9.567377,10.008774,10.227587,10.050273,9.559832,9.224068,8.529905,8.27714,8.646856,9.190115,10.0276375,10.355856,10.465261,10.555805,10.748209,9.7220545,8.782671,8.390318,8.488406,8.52236,8.446907,8.254503,8.213005,8.175279,7.564113,6.2097406,5.292993,4.515832,3.832987,3.4179983,3.150142,3.1237335,3.1425967,3.1727777,3.3463185,3.5802212,3.8065786,4.093298,4.4101987,4.5988297,4.8968673,5.1269975,5.5004873,6.0362,6.5568223,6.730363,6.587003,6.300284,6.013564,5.836251,6.0286546,6.119198,6.138061,6.3116016,7.0812173,7.5829763,7.454707,7.069899,6.7152724,6.587003,6.673774,6.903904,7.0548086,6.9793563,6.587003,6.888813,7.4773426,8.084735,8.771353,9.940866,9.703192,9.865415,10.295494,10.718028,10.710483,11.065109,11.476325,12.00072,12.623203,13.230596,14.196388,14.84528,15.596032,16.35433,16.509007,17.078674,16.950403,16.70141,16.542961,16.35433,16.335466,16.029884,15.792209,15.543215,14.796235,13.290957,12.15917,11.246195,10.657665,10.759526,11.193378,11.627231,12.091263,12.419481,12.234623,11.895086,11.830952,12.272349,12.90615,12.883514,13.788944,15.264041,15.988385,15.984612,16.622187,16.018566,16.097792,16.724047,17.463482,17.57666,16.791954,16.580687,16.278877,16.158154,17.429527,15.890297,15.645076,15.860115,15.369675,12.672247,13.45318,13.404137,13.181552,13.185325,13.585222,14.48688,14.43029,14.50197,14.815099,14.509516,14.234114,14.068119,14.147344,14.403882,14.569878,14.2944765,14.385019,14.807553,15.30554,15.39231,15.411173,14.984866,14.120935,12.928786,11.634775,10.257768,8.941121,7.854605,7.1302614,6.851087,6.3832817,5.885295,5.342037,4.8666863,4.7006907,4.606375,4.504514,4.3724723,4.187614,3.9197574,3.8707132,3.7499893,3.783943,3.9914372,4.1536603,3.6594462,3.5651307,3.904667,4.376245,4.357382,4.432834,4.2064767,4.1197066,4.5460134,5.7796617,7.141579,7.5037513,7.326438,7.115171,7.4094353,7.111398,6.72659,6.598321,6.688864,6.598321,7.3188925,7.888559,8.333729,8.722309,9.159933,9.876732,10.827434,11.548005,11.800771,11.532914,10.774617,10.152134,10.152134,10.076681,8.035691,7.0057645,6.039973,5.3194013,4.919503,4.817642,4.798779,5.010046,5.251494,5.379763,5.311856,5.353355,4.534695,3.7235808,3.270866,3.0105548,2.5314314,1.9693103,1.841041,1.9957186,1.6071383,1.8561316,2.2371666,2.4559789,2.3692086,1.9994912,1.4901869,1.2826926,1.20724,1.1846043,1.2411937,1.9730829,2.1277604,2.3616633,2.6823363,2.463524,2.4220252,3.0369632,3.4896781,3.610402,3.8858037,4.647874,4.8629136,4.927048,5.0213637,5.149633,4.5233774,3.289729,3.0935526,4.357382,6.2889657,7.0510364,8.0206,9.488152,11.125471,11.970539,9.152389,6.300284,3.904667,2.3692086,1.9881734,5.3571277,5.1835866,3.5689032,3.5160866,8.922258,9.820143,9.024119,6.511551,3.6254926,3.0407357,2.6898816,1.4335974,0.69039035,0.724344,0.62625575,1.991946,2.565385,2.3993895,1.8448136,1.539231,1.1996948,0.814887,0.49044126,0.35839936,0.55457586,1.0035182,0.9280658,0.6488915,0.3734899,0.18863125,0.3470815,0.4979865,0.49044126,0.392353,0.49044126,0.52062225,1.2713746,1.7882242,1.6825907,1.1544232,0.724344,0.7507524,0.79602385,0.70170826,0.6149379,1.0487897,1.0978339,2.625747,4.817642,4.1612053,4.6856003,4.7308717,3.9499383,2.7200627,2.1466236,3.289729,3.610402,3.3236825,3.029418,3.7009451,2.9841464,2.9954643,3.0746894,3.127506,3.640583,3.270866,3.942393,4.45547,4.406426,4.1800685,4.8025517,4.3800178,4.093298,4.466788,5.406172,5.907931,6.5002327,6.8435416,7.1566696,8.179051,8.197914,8.069645,8.431817,9.242931,9.767326,10.054046,10.167224,9.846551,10.001229,12.672247,12.347801,10.465261,9.914458,11.54046,14.132254,10.982111,12.664702,13.721037,11.736636,7.3377557,4.8327327,3.4934506,3.9763467,5.587258,6.25124,6.858632,7.273621,6.1908774,4.376245,4.6516466,5.6363015,5.451443,4.991183,5.342037,7.7716074,8.314865,8.43559,7.3717093,5.383536,3.7537618,5.2665844,5.692891,4.666737,3.4481792,4.938366,6.696409,8.345046,8.684583,7.5075235,5.6061206,4.9949555,7.092535,8.311093,6.934085,3.1539145,4.425289,5.59103,9.333474,14.535924,16.24115,12.404391,9.820143,7.4169807,5.0213637,3.3878171,4.2630663,4.6818275,5.783434,7.6093845,9.088254,9.8239155,9.948412,8.8618965,7.152897,6.571913,7.575431,9.258021,10.137043,10.401127,11.921495,11.174516,10.419991,10.616167,11.827179,13.20796,12.4307995,11.174516,8.103599,4.187614,2.674791,3.0860074,4.919503,8.224322,11.234878,10.370946,6.771862,4.587512,4.538468,5.142088,2.704972,4.715781,4.293247,4.0706625,5.5759397,9.258021,7.907422,7.748972,8.258276,8.412953,6.677546,9.601331,10.985884,11.136789,10.680302,10.570895,11.314102,11.732863,11.227332,10.295494,10.529396,10.661438,11.076427,10.438853,9.276885,9.97482,9.57115,9.552286,10.03141,10.695392,10.804798,9.424017,9.035437,9.261794,9.876732,10.789707,9.899368,9.371201,9.020347,8.480861,7.194396,7.360391,8.284684,8.548768,8.09228,8.20546,8.126234,8.167733,8.322411,8.567632,8.873214,10.8576145,11.393328,11.004747,10.0465,8.729855,9.291975,8.050782,6.964266,7.1000805,8.616675,10.280403,10.438853,9.435335,7.997965,7.2623034,6.0739264,5.9117036,6.3153744,6.719045,6.428553,6.2889657,5.9117036,5.300538,4.38379,3.0105548,4.112161,4.214022,3.5236318,4.06689,9.691874,2.8181508,1.3091009,2.9539654,6.0248823,9.25425,9.005256,9.64283,10.453944,10.695392,9.608876,8.918486,9.027891,9.484379,9.752235,9.201432,8.699674,8.975075,8.782671,7.9225125,7.24344,6.039973,5.032682,4.172523,3.5651307,3.4481792,4.8063245,8.254503,11.234878,11.574413,7.4811153,4.61392,4.4101987,5.670255,6.930312,6.458734,5.089271,4.821415,6.1644692,7.9451485,7.2962565,6.1041074,5.621211,5.8966126,6.2851934,5.455216,4.7836885,4.8365054,5.100589,5.4891696,6.349328,6.3417826,6.1720147,5.6061206,5.0968165,5.764571,5.753253,6.436098,7.3415284,8.213005,9.005256,9.34102,9.175024,8.786444,8.29223,7.6282477,7.6207023,7.798016,7.8621507,7.745199,7.6131573,7.665974,7.492433,7.2396674,6.9755836,6.677546,6.7567716,7.224577,7.8017883,8.341274,8.816625,8.812852,7.6886096,6.541732,5.9909286,6.156924,5.956975,6.3908267,6.7152724,6.719045,6.700182,6.1041074,6.33801,6.72659,7.122716,7.9225125,9.0807085,9.548513,9.929549,10.469034,11.053791,13.287186,14.279386,14.068119,13.174006,12.570387,11.974312,10.955703,10.178542,10.31813,12.061082,11.608367,11.189606,11.151879,11.404645,11.404645,10.714255,10.585986,10.7218,10.816116,10.567122,10.725573,11.268831,11.819634,12.079946,11.84227,11.517824,11.129244,11.080199,11.321648,11.359374,11.431054,11.823407,11.615912,11.208468,12.321393,13.513543,13.370183,12.73261,12.136535,11.796998,11.966766,11.442371,10.533169,9.793735,10.038955,10.9594755,11.423509,11.4838705,11.2650585,10.978339,11.283921,9.718282,9.993684,10.484125,10.518079,10.355856,10.174769,10.174769,9.9257765,9.291975,8.43559,8.89585,9.009028,8.892077,8.843033,9.333474,9.725827,9.789962,9.850324,9.918231,9.7069645,9.22784,8.405409,8.084735,8.345046,8.537451,8.412953,8.09228,8.322411,9.122208,9.797507,10.253995,9.752235,9.020347,8.597813,8.869441,8.529905,8.280911,8.552541,8.967529,8.348819,8.341274,8.431817,8.390318,8.09228,7.5112963,6.1833324,5.5457587,4.8930945,4.0970707,3.6028569,3.3576362,3.4557245,3.5123138,3.531177,3.904667,4.044254,4.1498876,4.195159,4.247976,4.4818783,4.7044635,4.8327327,4.979865,5.1232247,5.1232247,5.915476,6.1342883,5.975838,5.73439,5.7909794,6.300284,6.3455553,6.3116016,6.432326,6.749226,6.9265394,6.79827,6.643593,6.6058664,6.700182,6.6020937,6.8397694,7.0812173,7.164215,7.0887623,7.488661,7.7904706,8.084735,8.6732645,10.061591,9.718282,9.759781,10.125726,10.585986,10.736891,11.332966,12.189351,12.940104,13.381501,13.494679,13.758763,14.173752,14.898096,15.7657995,16.31283,16.976812,17.010767,16.644821,16.248695,16.343012,16.644821,16.222288,15.841252,15.671484,15.271586,13.558814,12.513797,11.796998,11.374464,11.536687,11.740409,11.766817,11.962994,12.396846,12.838243,12.54775,12.721292,13.053283,13.257004,13.068373,13.283413,14.57365,15.237633,15.335721,16.675003,15.924251,15.777118,16.4411,17.30503,16.954176,16.260014,16.388283,16.724047,17.225805,18.395319,16.961721,16.275105,16.086473,15.339493,12.174261,13.13628,13.736128,13.822898,13.834216,14.777372,15.486626,15.396083,15.554533,16.105335,16.29774,15.456445,14.750964,14.577423,14.84528,14.977322,14.664193,14.999957,15.343266,15.437581,15.418718,15.279131,15.049001,14.581196,13.879487,13.079691,11.359374,9.835234,8.6732645,7.9526935,7.696155,7.424526,6.964266,6.2663302,5.4778514,4.9421387,4.67051,4.5837393,4.485651,4.327201,4.191386,4.172523,4.055572,3.983892,4.0216184,4.1612053,3.85185,3.7273536,4.085753,4.8629136,5.624984,5.383536,5.172269,5.2062225,5.753253,7.145352,8.959985,8.790216,8.341274,8.469543,9.186342,8.83926,8.016829,7.273621,6.828451,6.5455046,7.4169807,8.062099,8.529905,8.903395,9.314611,10.574668,11.6875925,12.313848,12.468526,12.555296,11.7894535,11.736636,12.151625,11.936585,9.125979,8.080963,6.907676,6.270103,6.1342883,5.723072,5.723072,5.745708,5.8098426,5.828706,5.624984,5.4401255,4.236658,3.2972744,3.1124156,3.3915899,3.078462,2.6182017,2.3201644,2.0749438,1.3770081,1.8938577,2.2409391,2.3692086,2.3013012,2.1277604,1.9089483,1.7919968,1.8599042,1.9579924,1.6939086,2.1390784,2.5314314,2.7426984,2.6898816,2.354118,2.3880715,3.0520537,3.4972234,3.572676,3.8178966,4.647874,5.3646727,5.5570765,5.1647234,4.4931965,2.938875,2.6823363,3.85185,5.802297,7.092535,8.20546,9.295748,9.839006,9.910686,10.201178,6.304056,4.0216184,3.2746384,3.1539145,1.9240388,7.356619,8.477088,5.9230213,3.1765501,6.530414,10.544487,9.767326,7.118943,4.7610526,4.0970707,2.0485353,1.1129243,0.5055317,0.049044125,0.19240387,1.0827434,1.3732355,1.2525115,0.90920264,0.5583485,0.38858038,0.3055826,0.1961765,0.1358145,0.41876137,0.9997456,0.98465514,0.7394345,0.48666862,0.29426476,0.30935526,0.35462674,0.5696664,0.8526133,0.8526133,1.4826416,2.2899833,2.11267,1.0714256,0.58098423,0.5093044,0.44139713,0.3470815,0.24899325,0.21503963,0.7130261,0.9205205,1.9429018,3.2255943,2.535204,3.4670424,3.4330888,3.3123648,3.4481792,3.6594462,3.5085413,3.1350515,3.0181,3.2821836,3.7047176,3.308592,3.4859054,3.7952607,3.9688015,3.9159849,3.561358,4.036709,4.8553686,5.3194013,4.504514,4.938366,4.6026025,3.9273026,3.8669407,5.885295,6.3832817,7.1604424,7.484888,7.496206,8.201687,8.526133,8.14887,7.8923316,8.484633,10.533169,11.883769,12.540206,12.117672,11.415963,12.404391,12.668475,11.68382,11.012292,11.559323,13.5663595,12.472299,13.573905,13.340002,10.948157,8.280911,5.0741806,3.942393,3.6783094,4.195159,6.5002327,7.183078,6.7680893,5.7419353,5.6853456,9.258021,9.382519,8.692128,7.997965,8.016829,9.371201,9.171251,8.741172,7.7037,6.0739264,4.2894745,3.2670932,2.2409391,2.022127,2.916239,4.6931453,6.6586833,6.8737226,6.8850408,7.2698483,7.635793,4.9459114,8.035691,9.710737,7.6207023,4.2706113,5.455216,5.5683947,8.224322,12.777881,14.32843,11.785681,9.937095,6.960493,4.08198,5.5683947,4.919503,3.519859,4.1083884,6.013564,5.1345425,6.356873,6.828451,6.7756343,6.5002327,6.3945994,5.674028,7.805561,8.903395,8.529905,9.688101,12.513797,10.650121,9.80128,10.997202,10.601076,13.3626375,11.223559,7.8206515,5.100589,3.2821836,3.1652324,4.5988297,9.80128,15.199906,11.419736,5.2364035,5.13077,5.27413,4.0404816,4.0480266,3.8895764,4.3875628,4.9987283,6.168242,9.34102,8.348819,8.13378,6.809588,5.9418845,10.514306,12.08749,12.162943,11.664956,11.208468,11.121698,11.204697,11.472552,11.249968,10.525623,9.944639,9.842778,9.989911,9.439108,8.714764,9.80128,8.258276,8.031919,8.718536,9.906913,11.208468,9.8239155,9.171251,9.922004,11.299012,11.068882,10.095545,9.201432,9.035437,9.359882,9.039209,8.016829,8.650629,8.99771,8.918486,10.087999,10.035183,9.514561,9.224068,9.612649,10.887795,13.155144,13.389046,12.415709,10.850069,9.110889,8.820397,7.303802,6.8774953,7.7716074,8.16396,8.601585,9.307066,8.846806,7.33021,6.428553,5.772116,6.1078796,6.3116016,6.1833324,6.4474163,6.5530496,4.8666863,4.266839,5.119452,5.300538,4.5724216,3.6556737,2.7087448,1.9051756,1.4373702,1.7882242,1.961765,3.5538127,6.530414,9.224068,9.548513,9.895596,10.201178,10.182315,9.325929,8.171506,8.235641,9.065618,9.97482,10.072908,9.590013,9.839006,9.450426,8.239413,7.2283497,6.3945994,5.643847,4.6931453,3.6481283,2.9615107,4.1989317,7.6848373,9.673011,8.7600355,5.8890676,5.3948536,4.6290107,4.9987283,6.349328,6.983129,5.643847,5.617439,6.8850408,8.243186,7.2962565,6.436098,6.2436943,6.5040054,6.6813188,5.9192486,4.4931965,4.727099,5.191132,5.4476705,6.0626082,6.3719635,6.187105,5.8173876,5.6287565,6.0324273,5.975838,6.647365,7.8017883,8.971302,9.480607,9.510788,9.190115,8.748717,8.329956,7.99042,8.141325,8.20546,8.152642,8.058327,8.103599,8.062099,7.7678347,7.4018903,7.1378064,7.118943,6.6322746,6.8359966,7.492433,8.228095,8.526133,8.337502,7.1378064,5.987156,5.455216,5.624984,5.666483,6.258785,6.952948,7.383027,7.2585306,6.3153744,6.3417826,6.6624556,6.851087,6.72659,8.371455,9.216523,9.695646,10.061591,10.374719,12.0082655,13.023102,13.460726,13.422999,13.094781,12.694883,11.849815,10.95193,10.585986,11.555551,11.996947,12.012038,11.932813,11.951676,12.106354,11.099063,10.8576145,10.978339,11.125471,11.016065,11.438599,12.200669,12.736382,12.728837,12.083718,11.570641,11.197151,11.057564,11.091517,11.091517,11.246195,11.332966,11.159425,10.823661,10.714255,11.627231,12.570387,12.672247,12.030901,11.732863,12.079946,11.589504,10.650121,9.752235,9.473062,10.057818,10.838752,11.476325,11.563096,10.627484,9.842778,8.76758,8.737399,9.144843,9.646602,10.148361,9.695646,9.216523,9.016574,8.91094,8.239413,7.960239,8.209232,8.379,8.646856,9.978593,9.895596,9.480607,9.4127,9.718282,9.782416,8.937348,7.647111,6.63982,6.330465,6.8058157,7.111398,7.0585814,8.224322,9.918231,9.186342,9.318384,8.703445,8.446907,8.624221,8.269594,8.280911,8.458225,8.616675,8.812852,9.337247,9.107117,8.43559,8.228095,8.36391,7.707473,6.5455046,5.753253,5.172269,4.6742826,4.1498876,3.772625,3.5123138,3.4255435,3.5387223,3.8292143,4.146115,4.134797,4.036709,4.1272516,4.715781,4.447925,4.315883,4.2592936,4.4177437,5.111907,5.794752,6.4436436,6.900131,7.069899,6.911449,6.692637,6.5002327,6.273875,6.0550632,5.983383,5.7872066,5.873977,6.119198,6.40969,6.651138,7.043491,7.745199,8.043237,7.84706,7.673519,8.103599,8.273367,8.122461,8.084735,9.110889,9.940866,10.257768,10.740664,11.566868,12.419481,12.566614,12.996693,13.717264,14.324657,14.007756,14.007756,14.656648,15.339493,15.565851,14.969776,15.75071,16.505234,16.45619,15.792209,15.671484,16.697638,16.429781,16.16947,16.222288,15.931795,14.2077055,13.29473,12.894833,12.955194,13.626721,13.502225,13.13628,12.932558,12.864652,12.434572,12.543978,13.151371,12.925014,11.955449,11.747954,14.045483,15.826162,15.758255,14.562332,15.015047,15.55076,15.686575,16.124199,16.67123,16.218515,16.28265,16.361876,16.55428,17.01831,17.942604,18.248188,17.591751,16.840998,16.0412,14.418973,15.324403,15.256495,15.1395445,15.264041,15.290449,15.7657995,15.70921,15.814844,16.28265,16.84477,15.724301,14.800008,14.441608,14.611377,14.894323,15.577168,15.83748,16.060064,16.275105,16.188334,15.580941,15.580941,15.648849,15.399856,14.618922,12.653384,10.733118,9.4013815,8.624221,7.7829256,7.586749,7.1981683,6.571913,5.881522,5.5382137,4.8327327,4.4818783,4.1612053,3.8367596,3.7386713,3.7499893,3.9273026,4.146115,4.3309736,4.4403796,4.3196554,4.52715,4.878004,5.292993,5.783434,6.820906,6.228604,5.9796104,6.752999,7.9489207,8.231868,7.786698,7.647111,8.231868,9.367428,9.733373,8.967529,7.7942433,6.888813,6.851087,7.194396,8.186596,8.888305,9.118435,9.461743,10.38981,11.619685,12.58925,12.909923,12.359119,12.140307,12.23085,12.261031,11.664956,9.673011,8.661947,8.443134,9.348565,10.27663,8.726082,7.7376537,7.435844,7.0887623,6.356873,5.292993,5.2099953,3.9801195,3.059599,3.0860074,3.8895764,3.500996,3.1463692,2.9615107,2.7691069,2.0598533,2.0108092,2.0900342,2.3163917,2.505023,2.2748928,2.1164427,2.305074,2.595566,2.7917426,2.7313805,2.9992368,3.3878171,3.3123648,2.7540162,2.2447119,2.3654358,2.8898308,3.2444575,3.3764994,3.7688525,3.6707642,4.6629643,5.4438977,5.372218,4.45547,3.4179983,4.447925,5.938112,7.1038527,7.9941926,11.510279,11.476325,8.710991,5.515578,5.66271,6.149379,4.2291126,3.0746894,2.9501927,1.20724,3.5123138,4.8666863,5.0025005,4.0404816,2.5012503,6.3116016,8.654402,7.4697976,4.353609,4.561104,1.6825907,0.49421388,0.116951376,0.033953626,0.1056335,0.21503963,0.39989826,0.44139713,0.32821837,0.23013012,0.20372175,0.150905,0.10940613,0.150905,0.38103512,0.95447415,0.84129536,0.663982,0.62625575,0.5017591,0.62625575,0.784706,1.7844516,3.0030096,2.3805263,3.6141748,2.6295197,1.3543724,0.72811663,0.70170826,0.69039035,0.5017591,0.38103512,0.35085413,0.23013012,0.21503963,0.41498876,1.116697,2.4371157,4.3196554,3.9989824,4.014073,4.768598,5.5004873,4.255521,3.561358,3.8254418,4.45547,4.7912335,4.1197066,3.4594972,4.1272516,4.745962,4.9534564,5.4174895,4.9157305,4.82896,5.485397,6.2361493,5.43258,5.6400743,5.270357,4.398881,4.1272516,6.590776,7.5792036,8.073418,8.062099,7.9300575,8.469543,8.737399,8.107371,7.515069,7.594294,8.66572,11.072655,13.083464,14.079436,13.490907,10.819888,13.2607765,14.7321005,14.132254,12.909923,15.045229,12.642066,10.638803,10.008774,10.012547,8.194141,5.7872066,4.5912848,3.5236318,2.655928,3.2029586,5.696664,6.749226,7.118943,8.246958,12.238396,10.321902,9.997457,9.574923,9.224068,10.970794,9.382519,7.677292,6.3116016,5.300538,4.22534,3.2746384,2.505023,2.7917426,3.350091,1.7391801,3.5462675,2.9539654,4.357382,7.6093845,8.024373,5.7570257,4.9232755,4.353609,3.5236318,2.546522,1.8787673,1.1959221,1.0487897,1.267602,0.9620194,3.1840954,2.584248,1.2864652,1.7844516,6.971811,5.4363527,4.0178456,3.1614597,2.7653341,2.1654868,10.819888,11.631002,9.261794,6.700182,5.2326307,6.039973,6.9454026,7.062354,6.541732,6.5756855,6.6247296,4.485651,4.859141,7.635793,7.9036493,11.895086,13.717264,13.196642,10.069136,3.9688015,5.040227,6.937857,9.393836,11.223559,10.344538,6.8171334,8.424272,7.907422,4.9647746,6.270103,6.1116524,5.311856,4.1612053,3.99521,7.2170315,12.90615,12.064855,7.8244243,6.0739264,15.471535,11.747954,9.42779,10.9594755,14.151116,12.162943,12.332711,10.661438,9.137298,9.14107,11.457462,10.212496,8.967529,7.9262853,7.5188417,8.424272,7.1906233,6.779407,7.3000293,8.171506,8.13378,8.571404,7.8131065,7.835742,8.82417,9.14107,9.016574,9.454198,8.6732645,7.3075747,8.394091,7.914967,7.6697464,7.515069,7.643338,8.560086,8.499724,8.646856,8.809079,9.582467,12.3893,13.13628,12.276122,11.306557,10.710483,9.978593,7.7338815,5.715527,6.477597,9.639057,11.887542,10.899114,10.155907,9.559832,8.929804,8.024373,7.194396,6.4474163,5.9984736,6.009792,6.6058664,6.9869013,5.111907,3.9574835,4.5196047,5.8136153,5.0062733,3.772625,2.867195,2.474842,2.1805773,3.5839937,3.4594972,4.859141,7.914967,9.857869,10.016319,9.782416,9.895596,10.155907,9.397609,8.360137,7.854605,8.428044,9.793735,10.819888,10.355856,10.038955,9.42779,8.643084,8.360137,7.3717093,6.3832817,5.6513925,5.062863,4.134797,3.9159849,8.76758,10.79348,8.4544525,6.560595,6.3908267,5.9532022,5.2288585,4.5422406,4.5761943,6.2851934,6.7039547,7.4811153,8.394091,7.3717093,7.0774446,6.7114997,6.4474163,6.300284,6.1041074,4.5761943,4.7006907,5.040227,5.3156285,6.379509,6.221059,5.7494807,5.3759904,5.349582,5.753253,6.888813,7.5565677,8.265821,9.0807085,9.627739,9.774872,9.812597,9.016574,7.7829256,7.598067,8.062099,8.269594,8.616675,8.922258,8.424272,7.8244243,7.5188417,7.3113475,7.2924843,7.828197,7.7301087,7.586749,7.356619,7.232122,7.6584287,7.488661,6.9227667,6.326692,5.832478,5.3571277,5.3684454,5.828706,6.25124,6.488915,6.7454534,7.696155,7.8244243,7.647111,7.273621,6.40969,7.164215,8.160188,9.050528,9.627739,9.812597,10.216269,10.691619,11.336739,12.128989,12.925014,12.777881,12.098808,11.314102,10.850069,11.155652,11.936585,12.679792,12.947649,12.706201,12.313848,11.042474,10.691619,10.853842,11.114153,11.016065,10.819888,11.129244,11.623458,11.940358,11.657412,11.815862,11.812089,11.717773,11.555551,11.261286,10.868933,10.570895,10.284176,9.861642,9.0807085,9.348565,10.310584,11.106608,11.389555,11.351829,11.778135,11.080199,10.367173,10.095545,10.069136,10.899114,11.747954,12.543978,12.604341,10.650121,10.7218,8.552541,8.058327,8.175279,8.337502,8.473316,7.9451485,7.7338815,7.9413757,8.367682,8.507269,8.412953,8.5563135,8.620448,8.654402,9.076936,9.359882,9.34102,8.91094,8.156415,7.3415284,7.484888,7.326438,7.0359454,6.8058157,6.8435416,6.990674,7.2962565,8.518587,9.876732,9.027891,7.726336,7.77538,8.231868,8.654402,9.099571,8.820397,8.865668,8.8618965,9.024119,10.144588,9.971047,9.431562,9.397609,9.65792,8.888305,6.722818,6.228604,6.0550632,5.50426,4.52715,4.745962,4.776143,4.561104,4.1989317,3.9159849,3.9008942,3.9876647,4.08198,4.123479,4.104616,4.1083884,4.063117,3.9612563,3.8820312,3.953711,4.98741,5.613666,5.726845,5.6023483,5.8626595,5.643847,5.5759397,5.560849,5.613666,5.885295,6.2663302,6.387054,6.6850915,7.1378064,7.273621,7.911195,8.7600355,9.344792,9.333474,8.578949,8.273367,8.416726,8.620448,8.869441,9.510788,10.7218,11.216014,11.351829,11.532914,12.2119875,13.140053,14.351066,15.113135,15.011275,13.970031,13.717264,13.834216,14.068119,14.245432,14.260523,15.041456,15.245177,14.762281,14.068119,14.230342,14.796235,14.34352,14.086982,14.464244,15.150862,14.385019,13.905896,13.905896,14.403882,15.260268,15.169725,14.683057,14.139798,13.539951,12.543978,12.019584,12.223305,12.238396,11.823407,11.431054,12.51757,13.943622,14.7736,14.962231,15.354584,15.347038,16.275105,17.384256,18.052011,17.795471,18.040693,18.240643,18.659403,19.251705,19.640285,18.919714,17.282394,16.878725,17.538933,16.761772,17.022083,17.022083,16.927769,16.712729,16.131744,15.973294,15.384765,15.211224,15.543215,15.735619,14.837734,14.535924,14.50197,14.539697,14.57365,14.720782,15.082954,15.513034,15.878979,16.056292,15.845025,16.063837,16.407146,16.38451,15.339493,13.732355,11.766817,10.103089,9.0543,8.563859,7.7225633,7.01331,6.537959,6.224831,5.8437963,5.5570765,5.3986263,5.1873593,4.938366,4.8629136,4.715781,4.666737,4.6554193,4.7233267,4.991183,4.908185,4.817642,4.979865,5.3646727,5.6363015,6.138061,6.039973,5.9607477,6.387054,7.6810646,7.152897,6.960493,7.1076255,7.564113,8.269594,8.578949,8.284684,7.7678347,7.2094865,6.5945487,6.6322746,7.424526,8.333729,8.914713,8.922258,9.948412,10.593531,11.532914,12.438345,12.004493,11.491416,11.306557,11.057564,10.465261,9.344792,8.175279,8.028146,8.07719,7.964011,7.8017883,7.7112455,7.997965,7.6018395,6.387054,5.149633,4.67051,4.29702,3.7009451,3.1840954,3.6594462,3.4745877,3.229367,2.916239,2.686109,2.867195,2.3767538,2.033445,2.3390274,3.0218725,3.006782,2.5729303,2.8634224,3.0520537,2.916239,2.8181508,3.2029586,3.429316,3.218049,2.4710693,1.267602,1.4864142,2.474842,3.1954134,3.2821836,3.0369632,3.4859054,4.1008434,4.3347464,4.0404816,3.4670424,3.904667,5.1571784,7.0774446,9.21275,10.816116,11.1782875,8.416726,5.198677,3.440634,4.3309736,3.108643,5.7004366,7.0887623,6.326692,6.515323,4.3007927,3.572676,3.3840446,3.1237335,2.5012503,8.224322,6.6813188,3.9801195,2.886058,2.8294687,1.0714256,0.32444575,0.08299775,0.03772625,0.071679875,0.090543,0.17354076,0.21503963,0.18863125,0.120724,0.211267,0.13204187,0.09808825,0.17354076,0.26031113,0.5583485,0.8186596,0.77716076,0.51684964,0.45648763,1.7882242,2.7389257,3.1350515,2.938875,2.2598023,3.1576872,3.127506,2.6408374,1.8938577,0.7884786,0.8337501,0.7922512,0.62248313,0.38858038,0.27917424,0.62625575,0.5583485,0.8526133,1.8146327,3.2557755,3.2821836,3.7877154,4.214022,4.2027044,3.610402,3.0407357,3.3953626,3.6594462,3.640583,3.983892,4.115934,4.1272516,4.5120597,5.1081343,5.062863,5.956975,5.6476197,5.4665337,5.873977,6.4436436,6.40969,6.175787,5.372218,4.825187,6.579458,7.7942433,8.477088,9.039209,9.740918,10.676529,11.004747,10.069136,8.858124,8.028146,7.911195,9.865415,10.484125,11.155652,12.140307,12.562841,11.197151,11.9064045,11.529142,10.789707,14.313339,13.898351,10.653893,8.873214,9.310839,9.1825695,7.2170315,5.6400743,3.7047176,2.3880715,4.398881,6.881268,9.344792,11.129244,11.989402,12.102581,9.933322,9.955957,9.8239155,9.246704,9.993684,9.714509,9.246704,8.009283,6.405917,5.802297,4.749735,3.078462,3.8480775,6.115425,4.9119577,6.017337,3.9612563,4.534695,7.2887115,5.534441,4.406426,3.4217708,2.5314314,2.1277604,3.0369632,2.6182017,1.8259505,3.187868,5.8136153,5.379763,4.6931453,3.4481792,3.1312788,3.9273026,4.689373,2.7426984,5.7683434,9.533423,10.265312,4.6554193,9.552286,12.46098,13.641812,13.008011,10.1294985,9.469289,9.64283,10.623712,11.8045435,11.996947,8.801534,8.043237,6.696409,4.6214657,4.5460134,5.481624,7.6622014,7.91874,5.515578,2.1353056,4.881777,9.224068,11.465008,10.359629,7.149124,8.054554,9.876732,9.148616,6.40969,6.221059,5.8588867,6.0626082,6.2851934,6.1229706,5.311856,6.217286,7.828197,7.164215,5.772116,9.7220545,10.110635,9.276885,8.959985,9.65792,10.646348,11.442371,10.970794,9.771099,8.677037,8.797762,8.36391,8.375228,7.8395147,6.9567204,7.115171,6.900131,6.9869013,7.3453007,7.809334,8.096053,9.540969,9.397609,8.831716,8.311093,7.6131573,8.07719,9.684328,9.563604,7.8998766,7.9413757,8.488406,8.661947,8.933576,9.250477,9.024119,8.631766,9.201432,9.767326,10.518079,12.815607,13.7851715,13.000465,11.823407,10.729345,9.295748,8.035691,7.2698483,7.33021,8.273367,9.884277,9.8239155,8.990166,8.2507305,7.8923316,7.624475,7.009537,6.145606,5.938112,6.4964604,7.145352,6.477597,6.4738245,6.126743,5.292993,4.7044635,5.2137675,3.9122121,2.7087448,2.6823363,4.0970707,4.6818275,5.062863,6.519096,8.790216,10.076681,10.080454,10.186088,10.242677,10.042727,9.325929,8.865668,9.235386,10.03141,10.910432,11.563096,11.204697,10.291721,9.261794,8.458225,8.130007,7.5716586,6.368191,5.27413,4.4743333,3.5839937,3.240685,5.481624,7.122716,7.0849895,6.4021444,4.67051,6.6247296,10.834979,13.011784,6.006019,7.303802,7.907422,8.028146,7.756517,7.0510364,7.2660756,6.990674,6.6850915,6.5756855,6.651138,5.4401255,5.3986263,5.5457587,5.696664,6.477597,6.277648,5.994701,5.9305663,6.1531515,6.4964604,6.9982195,7.360391,7.8998766,8.60913,9.175024,9.009028,9.246704,9.1825695,8.669493,8.122461,8.586494,8.597813,8.548768,8.544995,8.386545,7.6886096,7.322665,7.2094865,7.326438,7.707473,8.047009,8.167733,7.997965,7.7301087,7.805561,7.1566696,6.85486,6.722818,6.5530496,6.089017,5.564622,5.6325293,6.1229706,6.7454534,7.1000805,7.9715567,8.009283,7.7640624,7.5716586,7.54525,7.383027,7.7904706,8.371455,9.001483,9.797507,9.948412,10.148361,10.657665,11.41219,12.019584,12.313848,11.9064045,11.589504,11.619685,11.740409,12.1101265,12.585477,13.083464,13.245687,12.434572,11.099063,10.397354,10.223814,10.487898,11.102836,11.8045435,12.242168,12.54775,12.593022,12.00072,11.570641,11.359374,11.502733,11.691365,11.1631975,10.401127,10.016319,9.612649,9.0957985,8.677037,9.042982,9.337247,9.763554,10.367173,11.02361,11.646093,11.495189,11.1782875,11.0613365,11.242422,11.476325,12.155397,12.54775,12.298758,11.419736,9.58624,8.243186,7.5075235,7.232122,7.2094865,7.1793056,7.54525,7.61693,7.635793,7.6923823,7.696155,7.624475,7.696155,7.779153,7.9489207,8.503497,8.793989,8.590267,8.114917,7.4697976,6.6360474,6.858632,7.0849895,7.2170315,7.2396674,7.2283497,6.971811,7.3981175,8.412953,9.201432,8.228095,7.5565677,7.7187905,8.016829,8.054554,7.7338815,8.303548,8.43559,8.382772,8.560086,9.567377,9.914458,9.963503,10.042727,9.929549,8.820397,7.858378,7.3981175,7.175533,6.862405,6.0324273,5.8928404,5.515578,4.957229,4.3913355,4.1008434,4.1197066,4.104616,4.036709,3.9348478,3.85185,3.92353,3.7537618,3.5877664,3.482133,3.2972744,3.9876647,4.5422406,4.8742313,5.081726,5.462761,5.7570257,5.8136153,5.80607,5.881522,6.1720147,6.1833324,6.3116016,6.6662283,7.1264887,7.3377557,8.175279,8.571404,8.650629,8.66572,8.967529,8.831716,8.959985,9.163706,9.465516,10.125726,10.767072,11.427281,11.921495,12.30253,12.849561,13.86817,14.64533,14.992412,14.667966,13.36641,13.0646,13.174006,13.419228,13.570132,13.434318,13.328684,13.223051,13.185325,13.147598,12.909923,12.921241,12.823153,12.864652,13.2607765,14.166207,14.313339,14.18507,14.037937,14.162435,14.883006,15.222542,15.316857,14.988639,14.136025,12.736382,11.446144,11.057564,10.948157,10.891568,11.0613365,11.827179,12.657157,13.502225,14.264296,14.818871,15.471535,16.724047,18.002966,18.693357,18.135008,17.38803,17.180534,17.520071,18.270823,19.149845,18.391546,17.667202,18.244415,19.417702,18.51227,18.097282,17.731337,17.263533,16.648594,15.939341,15.792209,15.150862,15.011275,15.494171,15.841252,15.290449,14.762281,14.543469,14.600059,14.569878,14.558559,14.728328,15.041456,15.4074,15.663939,16.105335,16.429781,16.848543,17.04472,16.16947,14.901869,13.226823,11.45369,9.940866,9.061845,8.213005,7.54525,7.213259,7.141579,7.001992,6.7680893,6.511551,6.2436943,5.983383,5.7570257,5.5495315,5.4174895,5.3458095,5.3269467,5.383536,5.4212623,5.3609,5.342037,5.379763,5.342037,5.4174895,5.617439,5.783434,6.0211096,6.7077274,6.730363,6.7454534,7.0284004,7.5905213,8.197914,8.416726,8.382772,7.997965,7.3075747,6.5228686,6.3455553,7.17176,8.29223,8.993938,8.567632,9.06939,10.03141,11.09529,11.834724,11.77059,10.95193,10.680302,10.431308,9.854096,8.7751255,8.258276,8.130007,7.8696957,7.4169807,7.175533,6.9265394,7.333983,7.322665,6.462507,4.9760923,4.2706113,4.0895257,3.9273026,3.712263,3.8405323,3.5085413,3.2557755,3.059599,3.048281,3.5160866,3.0143273,2.4371157,2.4182527,2.8332415,2.795515,2.7502437,3.0181,3.078462,2.9501927,3.187868,3.5047686,3.7877154,3.1916409,1.8900851,1.0676528,1.2751472,2.11267,2.5012503,2.444661,3.0369632,3.9876647,4.8100967,5.1156793,5.0175915,5.1232247,6.828451,7.798016,8.850578,9.952185,10.201178,8.544995,5.9607477,4.587512,4.2027044,2.2296214,1.5656394,3.9122121,5.885295,5.9909286,4.6214657,4.353609,3.3236825,3.4557245,4.776143,5.43258,6.541732,4.123479,2.04099,1.6184561,1.6373192,0.5319401,0.150905,0.056589376,0.030181,0.060362,0.060362,0.08299775,0.1056335,0.10186087,0.056589376,0.13204187,0.18863125,0.271629,0.32444575,0.18485862,0.43007925,0.965792,1.3430545,1.4901869,1.6976813,2.7011995,3.5349495,3.0746894,1.9504471,2.565385,3.3840446,3.1161883,2.6898816,2.3390274,1.6033657,1.5845025,1.2751472,0.97333723,0.7809334,0.63002837,0.6451189,0.6752999,0.7432071,1.1657411,2.5691576,3.3915899,4.0895257,3.99521,3.240685,2.7615614,2.6634734,2.8219235,3.078462,3.500996,4.398881,4.878004,4.6856003,4.957229,5.6325293,5.4703064,6.2323766,5.881522,5.59103,5.994701,7.164215,7.073672,6.6549106,5.7192993,5.119452,6.730363,7.77538,8.5563135,9.246704,10.005001,10.982111,11.77059,11.6875925,10.7218,9.310839,8.3525915,8.703445,8.899622,9.2995205,10.291721,12.276122,10.450171,10.227587,10.095545,10.174769,12.234623,14.50197,11.457462,8.635539,8.243186,9.137298,8.337502,7.020855,5.300538,4.1008434,5.149633,6.983129,9.088254,10.978339,12.336484,13.023102,11.46878,10.589758,9.752235,9.031664,9.201432,9.110889,8.733627,7.786698,6.692637,6.571913,5.907931,3.85185,3.9763467,5.458988,3.108643,4.3724723,3.4330888,4.67051,6.937857,3.5575855,6.722818,5.247721,3.3764994,3.4972234,6.1418333,6.719045,6.519096,7.816879,10.11818,10.182315,8.175279,6.115425,5.413717,5.7004366,4.825187,3.3010468,7.9225125,13.7700815,15.067864,5.2062225,6.6058664,7.4282985,7.6622014,7.118943,5.4212623,6.519096,7.2396674,10.110635,14.622695,17.206944,14.279386,15.350811,14.369928,9.9257765,5.2628117,5.726845,5.4363527,5.040227,4.5196047,3.2067313,7.696155,11.400873,12.306303,10.050273,5.9192486,6.379509,8.028146,7.7716074,6.0814714,6.971811,6.862405,5.8890676,6.187105,7.594294,7.665974,5.462761,5.613666,5.2854476,4.459243,5.934339,8.507269,9.273112,9.175024,9.337247,11.083972,11.295239,10.646348,9.857869,9.092027,7.9300575,7.7376537,7.699928,7.213259,6.5341864,6.771862,6.5002327,6.8661776,7.6131573,8.27714,8.152642,8.345046,8.443134,8.394091,8.273367,8.296002,8.239413,9.578695,10.11818,9.344792,8.424272,7.997965,8.175279,8.60913,9.156161,9.846551,10.057818,10.269085,10.642575,11.472552,13.200415,13.513543,12.543978,11.514051,10.650121,9.208978,7.99042,7.6093845,7.7829256,8.213005,8.597813,8.937348,8.416726,7.726336,7.356619,7.567886,7.5263867,6.7643166,6.2927384,6.4247804,6.7756343,5.4438977,5.6476197,5.904158,5.7192993,5.5797124,5.292993,4.29702,3.4783602,3.5877664,5.2288585,5.87775,6.2097406,7.2094865,8.741172,9.563604,9.906913,10.035183,9.967276,9.756008,9.5183325,9.6051035,10.34831,11.027383,11.438599,11.9064045,11.61214,11.087745,9.906913,8.473316,8.009283,7.6584287,6.85486,5.881522,5.010046,4.5120597,4.06689,3.9688015,5.081726,6.771862,6.911449,4.063117,6.7114997,12.181807,15.403628,8.918486,8.590267,8.235641,7.8734684,7.4773426,6.964266,7.2472124,6.9944468,6.6850915,6.5530496,6.587003,6.119198,6.485142,6.5568223,6.270103,6.620957,6.477597,6.1833324,5.9494295,6.009792,6.609639,6.862405,6.9189944,7.2962565,8.096053,9.001483,8.756263,8.944894,9.058073,8.831716,8.228095,8.341274,8.416726,8.488406,8.480861,8.194141,7.6131573,7.073672,6.8963585,7.152897,7.647111,7.7338815,7.9526935,7.960239,7.7602897,7.7414265,7.654656,7.4169807,6.990674,6.4738245,6.1078796,5.7683434,5.783434,6.3342376,7.1076255,7.2887115,7.7678347,8.065872,8.360137,8.465771,7.828197,7.1000805,7.3075747,7.707473,8.024373,8.45068,8.786444,9.125979,9.540969,10.035183,10.559577,10.872705,11.140562,11.302785,11.438599,11.729091,12.196897,12.917468,13.558814,13.664448,12.630749,11.642321,10.774617,10.155907,9.97482,10.484125,11.189606,11.649866,11.7894535,11.514051,10.702937,10.559577,10.544487,10.914205,11.472552,11.559323,10.589758,10.242677,9.884277,9.1976595,8.171506,8.511042,8.446907,8.888305,9.789962,10.170997,10.740664,10.891568,11.02361,11.283921,11.581959,11.668729,12.306303,12.740154,12.743927,12.638294,8.578949,8.235641,7.647111,7.1340337,6.771862,6.4021444,7.0472636,7.24344,7.0585814,6.6813188,6.428553,6.375736,6.4511886,6.63982,6.990674,7.654656,7.91874,7.7338815,7.4999785,7.326438,7.0472636,7.122716,7.250985,7.413208,7.4773426,7.2283497,7.164215,7.6093845,8.394091,8.820397,7.6584287,7.375482,7.3075747,7.364164,7.2698483,6.56814,7.1566696,7.5226145,7.745199,8.058327,8.827943,9.469289,9.906913,9.876732,9.239159,7.9941926,8.080963,7.7678347,7.541477,7.33021,6.5266414,6.0626082,5.6400743,5.2326307,4.851596,4.534695,4.5988297,4.4818783,4.217795,3.9310753,3.8556228,3.99521,3.7914882,3.6594462,3.6934,3.682082,3.942393,4.2064767,4.5007415,4.821415,5.1345425,5.621211,5.6476197,5.666483,5.873977,6.19465,5.753253,6.0248823,6.4436436,6.79827,7.2358947,7.6697464,7.914967,8.265821,8.918486,9.982366,9.865415,9.665465,9.529651,9.593785,9.97482,10.49167,11.25374,12.019584,12.630749,13.000465,13.641812,14.219024,14.392565,13.936077,12.736382,12.279895,12.513797,12.947649,13.215506,13.091009,12.415709,12.170488,12.31762,12.506252,12.0724,12.178034,12.427027,12.755245,13.226823,14.037937,14.558559,14.524607,14.203933,14.003984,14.479335,14.720782,14.962231,14.656648,13.626721,12.049765,10.729345,10.144588,9.948412,10.065364,10.710483,11.653639,12.279895,13.068373,14.083209,14.984866,16.044973,16.67123,17.342756,17.80679,17.048492,16.373192,16.158154,16.478827,17.338985,18.666948,18.327412,18.451908,19.625195,20.88148,19.700647,18.810308,18.025602,17.252214,16.4826,15.833707,15.720529,15.422491,15.565851,16.116653,16.38451,15.814844,15.060319,14.592513,14.524607,14.592513,14.554788,14.596286,14.811326,15.120681,15.279131,15.984612,16.38451,16.822134,17.191853,16.939087,15.705438,14.234114,12.3893,10.495442,9.318384,8.624221,8.14887,7.9413757,7.9489207,8.013056,7.9262853,7.564113,7.1264887,6.670001,6.1078796,5.9796104,5.8437963,5.670255,5.4778514,5.323174,5.3571277,5.3759904,5.2967653,5.1232247,4.9421387,4.908185,5.160951,5.4438977,5.643847,5.80607,6.0512905,6.149379,6.620957,7.484888,8.2507305,8.492179,8.431817,7.964011,7.2170315,6.541732,6.466279,7.213259,8.190369,8.7751255,8.299775,8.216777,9.510788,10.56335,10.7557535,10.457717,10.186088,10.076681,10.020092,9.673011,8.439363,7.9715567,8.126234,8.039464,7.5112963,7.009537,6.470052,7.0170827,7.4094353,7.020855,5.8400235,4.617693,4.236658,4.1612053,4.0970707,4.0103,3.4859054,3.0709167,3.0143273,3.3161373,3.7160356,3.3274553,2.969056,2.776652,2.7540162,2.776652,3.308592,3.2633207,3.0935526,3.0860074,3.3463185,3.863168,4.123479,3.440634,2.173032,1.7278622,1.6524098,2.1956677,2.354118,2.2069857,2.9200118,4.044254,5.247721,5.945657,6.3719635,7.594294,9.684328,9.854096,9.061845,8.235641,8.265821,6.3945994,4.5460134,4.0895257,4.3649273,2.6634734,3.8480775,3.2821836,3.591539,4.266839,1.659955,3.0030096,2.957738,3.5877664,4.9987283,5.311856,3.7009451,2.0975795,1.1129243,0.8224323,0.7394345,0.20749438,0.06790725,0.0452715,0.02263575,0.049044125,0.05281675,0.049044125,0.0452715,0.0452715,0.041498873,0.20749438,0.3169005,0.43007925,0.48666862,0.3169005,1.7354075,2.4182527,2.6144292,2.7125173,3.2482302,3.572676,3.5236318,2.9351022,2.5880208,4.195159,4.402653,3.0671442,2.3277097,2.4899325,2.033445,2.1541688,1.6071383,1.2185578,1.1846043,1.0789708,0.6488915,0.6149379,0.5583485,0.76207024,2.203213,3.451952,4.1989317,3.8895764,2.8558772,2.305074,2.425798,2.3956168,2.9086938,3.8707132,4.395108,5.534441,5.594803,5.4438977,5.515578,5.7872066,6.273875,6.3832817,6.5455046,6.934085,7.466025,7.432071,7.0963078,6.590776,6.488915,7.7829256,8.541223,8.869441,9.061845,9.374973,10.038955,10.751981,10.906659,10.265312,9.291975,9.171251,8.76758,8.601585,8.386545,8.627994,10.631257,10.891568,10.948157,11.004747,11.189606,11.52537,14.120935,12.377983,9.491924,7.7602897,8.567632,9.578695,8.465771,6.9491754,6.0512905,6.089017,7.24344,8.473316,9.578695,10.748209,12.562841,11.830952,10.310584,9.076936,8.5563135,8.537451,8.00551,7.443389,6.8058157,6.3342376,6.5455046,6.40969,4.689373,4.7421894,5.624984,2.082489,3.4368613,3.6745367,4.346064,4.825187,2.3088465,6.7114997,6.5455046,4.7610526,3.832987,5.7419353,6.609639,7.1038527,8.122461,9.8239155,11.631002,9.993684,7.5112963,5.904158,5.323174,4.349837,4.402653,9.718282,14.0907545,13.309821,5.1760416,6.4247804,6.085244,5.032682,3.8707132,2.9426475,5.270357,5.907931,8.235641,12.619431,16.395828,16.056292,19.36111,20.036411,17.01831,14.449154,14.603831,8.552541,4.8553686,5.8437963,7.594294,9.231613,10.472807,10.159679,8.443134,6.7944975,4.7572803,6.4021444,6.790725,5.4891696,6.598321,7.443389,5.8966126,5.3382645,6.670001,8.337502,6.7567716,5.100589,4.6931453,5.221313,4.7120085,7.1378064,9.099571,9.820143,9.80128,10.816116,10.891568,9.7220545,8.835487,8.488406,7.6923823,8.069645,7.9753294,7.4396167,6.8246784,6.8435416,6.8133607,7.0812173,7.779153,8.461998,8.114917,7.424526,7.699928,7.7904706,7.605612,8.111144,8.186596,9.042982,9.740918,9.812597,9.265567,7.877241,7.956466,8.484633,9.107117,10.106862,10.597303,10.661438,10.982111,11.774363,12.7477,12.604341,11.631002,10.895341,10.453944,9.34102,7.9715567,7.6093845,7.9451485,8.43559,8.311093,8.371455,7.865923,7.3151197,7.115171,7.515069,7.6508837,7.092535,6.617184,6.488915,6.462507,5.221313,5.1647234,5.3080835,5.3759904,5.798525,5.1571784,4.9345937,4.727099,4.772371,5.9720654,6.700182,6.9265394,7.466025,8.458225,9.367428,9.699419,9.748463,9.665465,9.601331,9.74469,10.438853,11.234878,11.721546,11.921495,12.291212,11.619685,11.619685,10.627484,8.801534,8.137552,7.5188417,7.3679366,6.63982,5.3910813,4.8138695,5.342037,4.8440504,4.889322,5.617439,5.753253,3.6179473,5.138315,11.144334,16.471281,9.97482,10.012547,8.650629,7.635793,7.3905725,6.9869013,7.3113475,7.201941,6.8699503,6.5266414,6.356873,6.3229194,6.8435416,6.9793563,6.7341356,7.066127,7.2396674,6.888813,6.2399216,5.798525,6.3342376,6.7152724,6.72659,6.990674,7.699928,8.627994,8.43559,8.533678,8.544995,8.318638,7.9338303,8.058327,8.269594,8.488406,8.533678,8.152642,7.4471617,6.8246784,6.6322746,6.888813,7.2585306,7.2660756,7.5490227,7.828197,7.9300575,7.809334,7.8696957,7.696155,7.17176,6.511551,6.258785,6.356873,6.2663302,6.63982,7.424526,7.865923,8.231868,8.511042,8.918486,9.201432,8.620448,7.635793,7.3981175,7.360391,7.2924843,7.277394,7.809334,8.182823,8.582722,9.031664,9.431562,9.582467,9.97482,10.552032,11.133017,11.378237,11.7894535,12.966512,13.728582,13.494679,12.30253,11.6875925,10.861387,10.18986,9.891823,10.042727,10.47658,11.0613365,11.212241,10.789707,10.11818,10.11818,10.035183,10.306811,10.982111,11.747954,10.816116,10.502988,10.170997,9.431562,8.137552,8.088508,8.107371,8.597813,9.344792,9.5183325,9.986138,10.223814,10.480352,10.816116,11.125471,11.472552,12.128989,12.593022,12.845788,13.358865,8.379,8.375228,8.062099,7.5075235,6.809588,6.0701537,6.2625575,6.4474163,6.349328,6.0286546,5.885295,5.7796617,5.704209,5.836251,6.19465,6.651138,6.9189944,6.9869013,7.0057645,7.111398,7.424526,7.564113,7.5603404,7.4999785,7.2924843,6.6586833,7.3000293,7.8696957,8.5563135,8.850578,7.54525,6.802043,6.3644185,6.3229194,6.458734,6.217286,6.1342883,6.722818,7.4207535,8.058327,8.865668,9.337247,9.5032425,9.076936,8.156415,7.220804,7.496206,7.54525,7.413208,6.930312,5.745708,5.251494,5.2250857,5.402399,5.5193505,5.292993,5.20245,5.040227,4.7308717,4.4101987,4.429062,4.647874,4.5422406,4.5120597,4.6856003,4.9421387,4.8063245,4.5422406,4.346064,4.3347464,4.5535583,4.817642,4.7912335,4.9949555,5.5306683,6.0814714,5.485397,5.692891,6.0550632,6.40969,7.0812173,7.0812173,7.7187905,8.952439,10.374719,11.208468,10.653893,10.065364,9.684328,9.556059,9.540969,10.657665,11.423509,11.996947,12.434572,12.679792,12.796744,13.588995,13.894578,13.340002,12.37421,11.589504,11.785681,12.340257,12.811834,12.955194,12.336484,11.996947,11.883769,11.868678,11.781908,12.528888,12.864652,13.230596,13.788944,14.418973,14.901869,15.026365,15.0905,15.222542,15.373446,14.909414,14.437836,13.751218,12.743927,11.415963,10.570895,10.084227,9.831461,9.88805,10.540714,11.793225,12.664702,13.505998,14.396337,15.147089,15.98084,15.890297,15.90916,16.127972,15.686575,16.305285,16.652367,16.863634,17.274849,18.43682,18.500954,18.297232,19.127209,20.432537,19.779873,19.255478,18.365139,17.372938,16.520325,16.0412,16.01102,16.21097,16.580687,16.878725,16.675003,15.788436,15.188588,14.70192,14.377474,14.5132885,14.407655,14.441608,14.649103,14.886778,14.830189,15.4074,15.863888,16.324148,16.840998,17.37671,16.203424,14.652876,12.668475,10.638803,9.390063,8.786444,8.529905,8.416726,8.371455,8.4544525,8.544995,8.152642,7.5603404,6.8661776,5.975838,5.9192486,5.8702044,5.6325293,5.2779026,5.1081343,5.0854983,5.13077,5.081726,4.949684,4.8930945,4.938366,5.093044,5.406172,5.80607,6.085244,5.885295,5.8173876,6.379509,7.5188417,8.624221,8.952439,8.741172,8.179051,7.4018903,6.511551,6.749226,7.213259,7.726336,8.043237,7.835742,7.8432875,9.06939,9.767326,9.4013815,8.6581745,9.435335,9.435335,9.454198,9.435335,8.477088,7.281166,7.8017883,8.209232,7.8734684,7.3490734,6.6850915,7.5075235,8.2507305,8.126234,7.149124,5.2779026,4.696918,4.485651,4.255521,4.142342,3.5349495,2.9652832,2.9351022,3.3538637,3.5462675,3.127506,3.229367,3.1199608,2.8332415,3.1539145,3.9763467,3.5424948,3.240685,3.4368613,3.4859054,4.3875628,4.719554,4.285702,3.4557245,3.1350515,2.3428001,2.674791,2.9954643,2.8558772,2.5087957,3.4368613,5.0062733,6.217286,7.2472124,9.424017,11.41219,10.306811,7.492433,5.138315,6.2097406,5.1571784,3.8480775,3.3878171,3.983892,4.9421387,6.8737226,4.3347464,2.7011995,2.7728794,0.77338815,1.237421,3.0030096,4.1272516,3.8593953,2.6634734,1.5731846,1.086516,0.80734175,0.5093044,0.12826926,0.120724,0.08677038,0.06790725,0.06790725,0.06413463,0.05281675,0.05281675,0.05281675,0.07922512,0.15845025,0.42630664,0.5281675,0.58475685,0.8111144,1.5241405,4.5460134,4.708236,4.1197066,4.014073,4.708236,4.8025517,4.715781,4.67051,5.1835866,7.0963078,5.5457587,3.2859564,2.4861598,2.8785129,1.7693611,2.2786655,1.7052265,1.3091009,1.3656902,1.1657411,0.6451189,0.392353,0.32821837,0.7205714,2.2069857,3.150142,3.9763467,3.9310753,3.1237335,2.5540671,2.5012503,2.4559789,3.1916409,4.327201,4.3121104,6.0512905,6.375736,5.7004366,5.0439997,6.0248823,6.379509,7.33021,8.22055,8.511042,7.786698,7.8131065,7.937603,8.412953,9.190115,9.910686,10.510533,10.016319,9.205205,8.677037,8.854351,9.088254,8.714764,8.190369,8.216777,9.733373,9.552286,8.854351,7.986647,7.6697464,9.005256,11.589504,12.917468,13.238141,12.898605,12.362892,12.830698,12.940104,11.272603,8.620448,7.99042,10.159679,9.367428,8.043237,7.33021,7.066127,7.726336,8.22055,8.36391,8.710991,10.593531,10.510533,9.21275,8.322411,8.182823,7.8621507,6.673774,6.0550632,5.6853456,5.5457587,5.9305663,6.1644692,5.353355,5.617439,6.1795597,3.3651814,4.3686996,4.5724216,3.6443558,2.2673476,2.1541688,3.6707642,5.7306175,5.6400743,3.7084904,3.2331395,3.380272,4.006528,4.9647746,6.4247804,8.888305,8.420499,6.8435416,4.9949555,3.5802212,3.218049,5.5797124,9.74469,10.27663,7.1566696,5.80607,11.189606,11.936585,9.854096,7.118943,6.2399216,8.737399,8.707218,8.284684,9.058073,12.061082,13.743673,18.059555,20.700394,23.118647,32.531345,30.260225,15.79598,6.432326,7.2057137,10.906659,7.3981175,6.7567716,6.1908774,5.847569,8.83926,4.927048,5.855114,6.700182,5.9607477,5.59103,7.0548086,6.228604,4.991183,4.689373,6.145606,7.250985,5.726845,6.0512905,7.865923,5.975838,6.530414,8.952439,10.133271,9.514561,9.103344,9.676784,8.756263,7.6207023,7.009537,7.1264887,8.209232,8.793989,8.578949,7.7716074,7.0812173,7.4999785,7.3868,7.533932,7.914967,7.7112455,7.492433,7.937603,7.696155,6.828451,6.809588,7.805561,8.661947,9.088254,9.193887,9.491924,7.914967,7.9300575,8.669493,9.522105,10.133271,10.27663,10.601076,11.0613365,11.480098,11.555551,11.589504,10.963248,10.382264,9.971047,9.258021,8.254503,7.8923316,7.956466,8.182823,8.262049,7.809334,7.175533,7.224577,7.8998766,8.239413,7.4697976,6.8397694,6.6586833,6.760544,6.488915,5.670255,5.5495315,5.2590394,4.8365054,5.221313,5.194905,5.6853456,5.8966126,5.9305663,6.79827,7.1793056,7.3151197,7.6923823,8.484633,9.578695,9.49947,9.608876,9.650374,9.669238,10.03141,11.212241,11.868678,12.117672,12.204442,12.483616,11.446144,11.619685,10.993429,9.4013815,8.514814,7.4018903,7.6622014,7.069899,5.3571277,4.195159,5.9117036,6.56814,5.9117036,4.52715,3.8707132,3.6330378,3.4142256,8.971302,16.177015,11.027383,10.8576145,8.990166,7.6810646,7.454707,7.1038527,7.5301595,7.541477,7.2094865,6.688864,6.187105,6.145606,6.48137,6.79827,7.0774446,7.6584287,8.16396,7.7301087,6.79827,5.9682927,5.9984736,6.549277,6.8850408,7.2283497,7.6697464,8.137552,7.997965,8.058327,7.9941926,7.748972,7.533932,7.9753294,8.2507305,8.446907,8.507269,8.201687,7.2887115,6.8359966,6.7680893,6.862405,6.7643166,6.9152217,7.213259,7.7112455,8.156415,7.986647,7.598067,7.4697976,7.1981683,6.7680893,6.5266414,6.952948,6.7869525,6.9189944,7.586749,8.401636,9.1825695,9.273112,9.454198,9.967276,10.499215,9.0957985,7.9941926,7.3000293,6.94163,6.6662283,7.0284004,7.303802,7.8432875,8.537451,8.801534,8.820397,8.865668,9.623966,10.740664,10.823661,11.189606,12.54775,13.283413,12.83447,11.668729,11.212241,10.612394,10.186088,9.982366,9.778644,10.091772,10.819888,11.065109,10.687846,10.336992,10.174769,9.899368,9.993684,10.601076,11.52537,10.895341,10.627484,10.280403,9.616421,8.575176,7.748972,7.967784,8.469543,8.91094,9.35611,9.846551,9.940866,9.891823,9.87296,9.986138,10.834979,11.54046,11.91395,12.23085,13.219278,8.209232,7.9413757,7.333983,6.7944975,6.398372,5.873977,6.25124,6.5228686,6.858632,7.3113475,7.8131065,7.2887115,6.405917,5.8626595,5.904158,6.3342376,6.405917,6.25124,6.0286546,5.9230213,6.119198,6.7152724,7.141579,7.020855,6.428553,5.8890676,6.696409,7.8206515,8.620448,8.60913,7.462252,6.5228686,5.7570257,5.4401255,5.4967146,5.5080323,6.3153744,6.900131,7.7716074,9.024119,10.329447,10.38981,9.337247,8.280911,7.7338815,7.598067,8.197914,8.620448,8.333729,7.164215,5.292993,4.636556,4.534695,4.8629136,5.511805,6.379509,5.8890676,5.613666,5.4703064,5.587258,6.270103,6.4436436,6.349328,6.304056,6.349328,6.224831,5.3344917,4.4441524,3.7047176,3.3463185,3.663219,3.904667,4.2404304,4.847823,5.726845,6.730363,6.1908774,5.2779026,5.2062225,6.043745,6.7152724,7.9451485,9.0957985,9.963503,10.47658,10.695392,9.669238,9.488152,9.774872,10.26154,10.789707,12.351574,13.023102,12.992921,12.777881,13.230596,13.132507,13.445636,13.615403,13.290957,12.313848,11.216014,11.004747,11.427281,11.966766,11.857361,11.344283,10.785934,10.718028,11.197151,11.793225,12.785426,12.985375,13.008011,13.185325,13.5663595,14.358611,15.497944,17.172989,18.632996,18.218006,17.206944,15.47908,14.313339,13.966258,13.687083,12.491161,11.5857315,10.899114,10.529396,10.770844,12.151625,13.211733,13.754991,13.547497,12.313848,12.974057,14.317112,15.369675,15.916705,16.539188,17.73511,18.629223,17.96524,16.444872,16.739138,16.810818,14.826416,14.27184,15.875206,17.610613,19.379974,19.025349,17.497435,15.98084,15.8676605,16.648594,17.112627,17.127718,16.735365,16.11288,15.245177,15.120681,14.969776,14.588741,14.34352,14.064346,13.909668,14.019074,14.1926155,13.902123,14.596286,15.007503,15.482853,16.192106,17.120173,16.961721,15.109364,12.90615,11.000975,9.352338,8.778898,8.729855,8.692128,8.526133,8.4544525,8.186596,7.7150183,7.194396,6.609639,5.7683434,5.485397,5.7079816,5.783434,5.6098933,5.643847,5.8173876,5.934339,5.8702044,5.7872066,6.1041074,5.934339,6.0550632,6.6020937,7.6093845,9.001483,8.684583,8.039464,8.073418,9.076936,10.589758,10.8576145,10.785934,10.163452,8.744945,6.255012,6.560595,6.719045,6.8737226,6.9567204,6.7152724,8.397863,9.205205,9.076936,8.548768,8.744945,9.49947,8.91094,8.345046,8.356364,8.695901,7.062354,7.3377557,8.311093,8.888305,8.118689,7.1906233,8.175279,9.461743,9.469289,6.6360474,4.745962,4.5120597,4.6327834,4.5799665,4.5912848,4.006528,3.7047176,3.519859,3.410453,3.4481792,2.6295197,2.746471,2.6182017,2.323937,3.2029586,3.5462675,3.2557755,3.3764994,4.0480266,4.485651,5.342037,6.477597,6.1720147,4.82896,4.991183,2.8898308,3.078462,3.7198083,3.6330378,2.2899833,2.8747404,4.798779,6.56814,7.8621507,9.522105,12.427027,9.654147,5.907931,3.8895764,4.3196554,2.916239,2.7841973,4.6327834,6.6247296,4.3800178,2.1202152,3.6971724,4.0782075,2.4220252,2.1051247,1.6788181,5.692891,7.352846,5.485397,4.5309224,1.4675511,0.9507015,0.875249,0.422534,0.030181,0.18863125,0.10186087,0.124496624,0.271629,0.19994913,0.10186087,0.150905,0.23390275,0.34330887,0.55080324,0.52439487,0.83752275,0.94315624,1.6939086,5.3571277,7.8319697,5.7607985,4.689373,5.8702044,6.270103,6.990674,10.797253,10.819888,7.8395147,10.269085,5.349582,3.9197574,4.2102494,4.1498876,1.3430545,2.2220762,1.7655885,1.3732355,1.2034674,0.150905,0.23767537,0.1961765,0.32821837,1.0223814,2.7313805,2.7087448,3.874486,4.4215164,3.9688015,3.5538127,3.2482302,3.410453,3.821669,4.5196047,5.8136153,6.5455046,6.300284,5.80607,5.80607,7.0510364,6.571913,8.213005,9.733373,10.035183,9.156161,9.0957985,9.665465,10.899114,12.276122,12.740154,13.498452,12.672247,10.767072,8.903395,8.820397,9.344792,9.144843,8.756263,8.718536,9.597558,8.854351,7.9262853,7.3868,7.7602897,9.507015,10.801025,12.608112,13.5663595,13.290957,12.37421,11.091517,12.868423,13.472044,11.408418,7.9036493,8.062099,8.778898,8.756263,7.8621507,7.141579,7.3000293,7.284939,7.303802,7.7602897,9.261794,9.578695,9.073163,8.83926,8.654402,6.9567204,5.2137675,4.640329,4.4931965,4.5497856,5.111907,5.3080835,5.511805,3.9499383,2.0108092,4.255521,4.636556,3.6141748,3.169005,3.6179473,3.6330378,2.1805773,3.5085413,6.0739264,8.088508,7.5527954,6.7831798,6.2814207,6.8850408,7.2887115,4.044254,3.640583,5.5985756,5.666483,3.8405323,4.3800178,8.601585,5.934339,3.6556737,4.817642,8.224322,20.836208,22.413166,16.59955,9.684328,10.574668,14.86037,15.580941,14.136025,12.853333,15.015047,13.562587,14.479335,18.21046,29.211435,55.966892,47.00691,23.254461,7.605612,5.304311,3.9386206,2.263575,3.8707132,4.4931965,4.727099,10.023865,7.4018903,4.564876,5.50426,8.643084,6.8359966,6.300284,6.0626082,6.168242,6.0739264,4.67051,5.119452,6.700182,8.167733,8.918486,8.941121,7.5263867,9.533423,10.352083,8.797762,7.1264887,7.5527954,8.82417,8.639311,6.858632,5.4778514,6.1116524,8.27714,9.352338,8.669493,7.5226145,7.0585814,6.63982,6.609639,6.809588,6.5756855,7.5301595,7.967784,8.201687,8.065872,6.94163,8.175279,9.673011,10.069136,9.125979,7.7225633,6.2436943,6.187105,7.435844,9.495697,11.476325,11.314102,11.744182,11.872451,11.3971,10.604849,11.2650585,11.25374,10.27663,8.880759,8.4544525,8.990166,8.831716,8.009283,6.9793563,6.6360474,6.477597,6.587003,8.533678,11.378237,11.657412,8.2507305,6.6322746,6.368191,6.6850915,6.439871,5.1835866,5.3156285,5.572167,5.6476197,6.2097406,6.270103,6.25124,6.349328,6.8737226,8.239413,7.835742,7.5527954,8.137552,9.224068,9.322156,9.21275,9.771099,9.948412,9.835234,10.665211,11.729091,12.15917,11.925267,11.446144,11.581959,11.472552,11.32542,10.884023,10.076681,9.001483,7.9300575,7.7150183,7.062354,5.6476197,4.134797,4.5007415,5.455216,6.673774,7.213259,5.492942,5.6778007,5.6287565,6.2851934,9.710737,19.134754,9.820143,7.9791017,8.122461,7.7640624,7.3868,7.7640624,7.4094353,7.220804,7.1302614,6.1041074,6.092789,6.5266414,7.0963078,7.575431,7.8432875,8.013056,7.352846,6.7944975,6.5341864,5.9984736,6.1305156,7.1000805,7.9941926,8.360137,8.16396,7.8961043,7.9753294,8.235641,8.303548,7.5829763,7.8395147,7.986647,8.122461,8.179051,7.9338303,7.4697976,7.5829763,7.748972,7.61693,7.020855,6.7643166,6.862405,7.2283497,7.6697464,7.888559,7.5603404,7.201941,6.8850408,6.5530496,6.0286546,6.4436436,6.7643166,7.175533,7.54525,7.462252,9.122208,9.703192,10.514306,11.9064045,13.2607765,10.378491,8.284684,7.1679873,6.6662283,5.8588867,5.383536,5.885295,6.858632,7.77538,8.118689,8.216777,8.552541,8.990166,9.495697,10.11818,11.41219,11.981857,12.276122,12.3289385,11.778135,11.155652,10.917976,10.352083,9.424017,8.790216,9.374973,9.88805,9.978593,9.639057,9.201432,9.273112,9.574923,10.242677,11.000975,11.185833,11.050018,10.978339,10.748209,10.137043,8.941121,7.111398,6.8737226,7.5263867,8.537451,9.552286,10.344538,10.005001,9.363655,8.82417,8.360137,9.631512,10.469034,10.853842,11.219787,12.449662,7.4509344,7.183078,6.7379084,6.319147,6.0512905,5.983383,6.2851934,6.7680893,7.4509344,8.175279,8.616675,8.152642,7.8923316,7.6584287,7.3981175,7.1981683,7.3000293,6.858632,6.387054,6.1342883,6.092789,6.2625575,6.651138,6.7944975,6.696409,6.8435416,6.7379084,7.2924843,7.5188417,7.01331,5.9720654,6.058836,6.273875,6.439871,6.5002327,6.5228686,6.9567204,6.651138,6.820906,7.567886,7.888559,8.194141,8.013056,7.673519,7.3868,7.232122,7.8395147,7.8923316,7.4396167,6.609639,5.5985756,5.458988,5.3910813,5.8136153,6.72659,7.707473,7.9338303,8.126234,8.409182,8.412953,7.2585306,6.9152217,6.470052,6.187105,6.013564,5.5797124,5.7607985,5.372218,4.9723196,4.776143,4.6742826,4.938366,5.5797124,6.1795597,6.5228686,6.5945487,6.741681,7.1566696,7.443389,7.5037513,7.5301595,7.9753294,9.21275,10.223814,10.521852,10.133271,9.763554,9.627739,9.918231,10.555805,11.1782875,12.261031,12.823153,13.0646,13.275867,13.864397,13.58145,13.52486,13.264549,12.706201,12.128989,11.589504,11.781908,11.996947,11.944131,11.747954,10.687846,10.212496,10.284176,10.774617,11.442371,12.204442,12.47607,12.611885,13.019329,14.139798,14.920732,15.935568,17.139036,18.135008,18.168962,16.882498,15.871433,15.0376835,14.649103,15.335721,14.286931,12.679792,11.18206,10.378491,10.759526,11.231105,11.725319,11.883769,11.6875925,11.472552,12.061082,13.185325,14.1926155,15.052773,16.36942,17.23335,17.716248,17.222033,16.222288,16.252468,17.086218,17.142809,17.312576,18.085964,19.538425,20.839981,20.175999,17.976559,15.618668,15.441354,16.55428,17.142809,17.1164,16.625957,16.052519,16.271332,16.539188,16.331694,15.716756,15.343266,14.524607,14.056801,13.736128,13.547497,13.656902,14.117163,14.852824,15.279131,15.55076,16.546734,16.33924,15.207452,13.604086,11.872451,10.231359,9.258021,9.031664,8.7751255,8.322411,8.122461,8.273367,8.152642,7.8432875,7.375482,6.7077274,6.330465,6.1229706,5.8211603,5.4778514,5.4740787,5.5004873,5.7381625,6.19465,6.741681,7.115171,7.5112963,7.5565677,7.6622014,8.231868,9.673011,8.827943,8.284684,9.084481,10.744436,11.272603,11.434827,11.461235,11.151879,10.186088,8.137552,8.058327,8.190369,7.91874,7.2698483,6.8963585,8.024373,8.661947,8.710991,8.348819,8.047009,9.125979,8.9788475,8.684583,8.76758,9.186342,9.442881,8.914713,9.390063,10.487898,9.631512,8.45068,8.07719,8.050782,7.6395655,5.832478,4.2819295,3.8669407,4.063117,4.432834,4.640329,4.142342,3.8707132,3.742444,3.7348988,3.9008942,3.4745877,3.8405323,4.183841,4.3385186,4.779916,4.436607,4.5196047,3.92353,3.8065786,7.586749,6.907676,5.66271,4.5196047,3.8669407,3.8292143,4.3385186,5.0025005,5.05909,4.5535583,4.349837,5.0553174,6.530414,7.7376537,8.514814,9.559832,10.167224,6.1078796,3.2029586,2.8558772,2.022127,2.463524,3.138824,2.886058,1.7919968,1.20724,2.082489,2.3692086,1.9391292,2.1390784,5.8173876,6.8133607,7.5301595,6.119198,3.0746894,1.2223305,1.3807807,1.0336993,0.5357128,0.1659955,0.116951376,0.20749438,0.1358145,0.35085413,0.66775465,0.271629,0.30935526,0.51684964,0.58475685,0.49044126,0.513077,0.935611,1.1355602,2.1692593,4.45547,7.786698,8.7600355,6.8661776,6.1531515,7.5188417,8.710991,9.314611,11.332966,11.3820095,9.884277,11.076427,6.8661776,5.3571277,5.172269,4.6554193,1.8674494,2.795515,1.5958204,0.663982,0.58475685,0.13958712,0.362172,0.633801,1.2147852,2.0560806,2.7804246,3.8480775,5.0779533,5.13077,4.2328854,4.142342,4.217795,4.255521,4.610148,5.3571277,6.2889657,6.7077274,6.590776,6.470052,6.779407,7.816879,7.537705,8.3525915,9.061845,9.590013,10.985884,11.608367,10.63503,10.170997,10.789707,11.544232,13.875714,12.860879,10.989656,9.756008,9.661693,12.336484,12.989148,11.815862,10.148361,10.438853,9.842778,9.171251,8.854351,9.171251,10.26154,10.453944,11.332966,12.113899,12.566614,13.008011,12.479843,13.249459,14.822643,15.441354,12.113899,9.314611,8.126234,7.654656,7.5226145,7.884786,7.594294,7.533932,7.673519,8.043237,8.710991,8.816625,8.605357,8.790216,9.167479,8.643084,6.428553,4.7836885,3.904667,3.9122121,4.8440504,5.27413,5.221313,5.73439,6.3455553,5.0854983,7.194396,6.3342376,4.2706113,3.2255943,5.8664317,2.8030603,1.9994912,2.1088974,2.6483827,4.025391,6.643593,6.5341864,6.1041074,5.379763,2.0183544,2.191895,5.9796104,6.6322746,4.745962,8.262049,8.627994,8.009283,7.5792036,7.5792036,7.333983,14.943368,13.441863,8.986393,6.9755836,12.027128,11.057564,15.82239,20.311813,21.869907,21.179516,17.255987,16.135517,16.165699,20.677757,38.00165,29.479292,14.053028,4.9760923,4.3724723,3.240685,4.4403796,5.6551647,4.8063245,3.108643,5.1043615,4.8063245,4.6742826,5.281675,6.7077274,8.533678,7.752744,6.4436436,7.9791017,11.393328,11.393328,6.9454026,8.22055,8.948667,7.854605,8.646856,7.5075235,8.197914,8.805306,8.575176,7.907422,8.179051,7.696155,6.990674,6.571913,6.930312,8.27714,9.001483,8.375228,7.213259,7.8508325,7.066127,6.56814,6.330465,6.4021444,6.8925858,6.9755836,6.6662283,6.5945487,6.628502,5.855114,6.1795597,8.111144,9.21275,8.782671,7.865923,5.9909286,5.553304,6.2663302,7.828197,9.910686,10.174769,10.054046,9.608876,8.990166,8.420499,9.322156,9.850324,9.469289,8.488406,8.050782,8.567632,8.809079,8.529905,7.9036493,7.492433,6.934085,6.7039547,7.3151197,8.707218,10.27663,8.258276,6.9567204,6.587003,6.8246784,6.8058157,6.2814207,5.485397,5.0515447,5.2326307,5.8928404,6.4436436,6.741681,7.4396167,8.473316,9.06939,8.130007,7.9451485,8.843033,10.084227,9.861642,9.439108,9.522105,9.891823,10.536942,11.680047,11.872451,11.793225,11.578186,11.351829,11.204697,10.359629,9.556059,9.495697,9.7069645,8.526133,7.4811153,6.888813,6.247467,5.66271,5.8211603,5.3269467,5.251494,5.828706,6.187105,4.357382,5.723072,5.5985756,5.8136153,7.854605,12.883514,7.84706,7.937603,8.835487,8.707218,8.190369,7.4169807,6.8397694,7.0359454,7.4471617,6.3832817,6.2436943,6.48137,7.0284004,7.6320205,7.8432875,7.5829763,7.4735703,7.2170315,6.779407,6.398372,6.7077274,7.4207535,8.22055,8.907167,9.382519,8.8618965,8.590267,8.326183,7.964011,7.54525,8.341274,8.956212,8.873214,8.145098,7.4207535,7.33021,7.145352,7.0812173,7.069899,6.7756343,6.6549106,6.8699503,6.8058157,6.643593,7.352846,7.303802,7.069899,6.741681,6.349328,5.8437963,5.4891696,5.6325293,6.0814714,6.579458,6.828451,8.07719,9.439108,10.687846,11.7555,12.759018,10.114408,8.503497,7.756517,7.2585306,5.945657,4.991183,5.1043615,5.5306683,6.096562,7.1906233,7.5527954,7.9225125,8.288457,8.797762,9.763554,11.465008,12.0082655,12.128989,12.049765,11.461235,11.065109,11.189606,10.774617,9.876732,9.691874,9.329701,9.26934,9.258021,9.246704,9.382519,9.631512,9.627739,9.756008,10.035183,10.110635,10.570895,10.650121,10.325675,9.680555,8.903395,6.760544,6.4738245,7.1906233,8.307321,9.465516,10.231359,9.846551,9.446653,9.393836,9.239159,9.835234,10.33322,10.502988,10.33322,10.023865,6.779407,6.4210076,6.33801,6.198423,5.9494295,5.836251,5.824933,6.3116016,7.213259,8.209232,8.744945,8.186596,7.9036493,7.7716074,7.7376537,7.835742,7.7640624,7.432071,6.907676,6.398372,6.2436943,6.149379,6.5832305,6.9227667,6.9755836,6.971811,6.3342376,6.3455553,6.5530496,6.488915,5.6815734,6.009792,6.719045,7.1793056,7.0887623,6.4926877,6.217286,6.1418333,6.4436436,6.8435416,6.571913,6.692637,6.730363,6.72659,6.790725,7.122716,7.5490227,7.5037513,7.4018903,7.466025,7.7376537,7.5188417,7.2887115,7.462252,8.175279,9.276885,10.001229,10.34831,10.518079,10.133271,8.265821,7.914967,7.5527954,7.0057645,6.4210076,6.270103,6.4134626,6.398372,6.145606,5.783434,5.643847,5.873977,6.1041074,6.439871,6.858632,7.2094865,8.394091,9.310839,9.661693,9.525878,9.382519,9.495697,9.865415,10.03141,9.820143,9.371201,9.529651,9.673011,9.884277,10.269085,10.93684,11.676274,12.359119,12.970284,13.536179,14.151116,13.9888935,13.86817,13.58145,13.113645,12.653384,12.351574,12.291212,12.128989,11.796998,11.491416,11.042474,11.200924,12.012038,13.204187,14.2077055,14.962231,15.562078,15.69412,15.633758,16.260014,17.882242,18.395319,18.523588,18.376457,17.463482,17.557796,16.675003,15.890297,15.660167,15.818617,14.894323,13.347548,11.763044,10.601076,10.216269,10.38981,10.751981,11.050018,11.283921,11.710228,12.494934,13.494679,14.400109,15.207452,16.244923,17.063583,17.769064,17.908651,17.72002,18.12369,18.746174,18.97253,18.708447,18.399092,19.040438,20.258997,19.757236,18.572634,17.274849,15.958203,16.516552,17.214487,17.425755,17.08999,16.705183,16.569368,16.15438,15.546988,14.84528,14.120935,13.272095,12.932558,12.770335,12.657157,12.691111,12.909923,13.445636,14.0983,14.830189,15.799753,15.520579,14.735873,13.396591,11.751727,10.340765,9.597558,9.484379,9.276885,8.846806,8.646856,8.858124,8.333729,7.8395147,7.624475,7.4169807,7.213259,6.983129,6.6134114,6.1531515,5.836251,5.926794,6.149379,6.387054,6.5228686,6.4738245,6.937857,7.1793056,7.149124,7.1679873,7.911195,7.5565677,7.8395147,9.020347,10.7557535,12.113899,12.702429,12.1252165,11.1631975,10.26154,9.529651,9.273112,9.024119,8.684583,8.197914,7.5829763,8.103599,8.548768,8.816625,8.827943,8.52236,9.14107,9.159933,8.918486,8.865668,9.556059,10.646348,9.771099,9.680555,10.797253,11.234878,10.9594755,10.152134,9.363655,8.597813,7.3075747,5.2779026,4.006528,4.055572,4.9044123,4.957229,4.7346444,4.4403796,4.1612053,4.074435,4.4630156,5.0175915,5.5268955,5.692891,5.5382137,5.383536,5.1798143,5.775889,6.221059,6.432326,7.17176,5.824933,4.2706113,3.6292653,3.9273026,4.0970707,5.6098933,6.25124,6.0248823,5.492942,5.783434,6.1720147,7.6207023,9.159933,9.771099,8.379,6.8473144,3.6179473,2.1881225,2.637065,1.6146835,2.5616124,3.5085413,2.5540671,0.3772625,0.21881226,0.9205205,1.2562841,1.1242423,2.0787163,7.3377557,9.258021,6.719045,3.5764484,1.6184561,0.55080324,1.780679,1.1883769,0.39989826,0.13958712,0.21881226,0.14713238,0.35462674,0.7092535,0.8941121,0.38103512,0.36594462,0.5055317,0.58098423,0.62625575,0.9242931,1.7995421,2.3277097,3.9763467,6.5945487,8.420499,8.080963,7.854605,8.096053,8.718536,9.224068,10.446399,11.027383,10.502988,9.574923,10.133271,8.2507305,6.903904,6.56814,6.156924,3.0520537,4.3121104,2.595566,1.086516,0.76207024,0.41121614,0.97710985,1.780679,2.1994405,2.3654358,3.150142,3.8178966,4.429062,4.432834,4.0178456,4.112161,4.6818275,4.6214657,4.8138695,5.624984,6.8850408,6.971811,7.0359454,6.964266,7.164215,8.578949,9.084481,8.865668,8.397863,8.5563135,10.601076,11.52537,10.729345,9.737145,9.669238,11.25374,14.117163,13.739901,12.064855,10.672756,10.789707,13.5663595,14.479335,13.174006,11.042474,11.227332,10.657665,10.374719,10.367173,10.676529,11.385782,11.080199,11.125471,11.449917,12.128989,13.377728,13.958713,14.313339,14.78869,15.546988,16.55428,13.981348,11.057564,9.159933,8.4544525,7.888559,7.748972,7.911195,8.031919,8.118689,8.537451,8.639311,8.303548,8.099826,8.243186,8.597813,6.8661776,5.281675,4.398881,4.304565,4.610148,5.311856,5.2779026,5.726845,6.6360474,6.730363,7.220804,5.240176,4.002755,4.466788,5.3269467,4.266839,5.070408,4.214022,1.9202662,2.1353056,3.663219,3.8065786,3.8405323,4.0404816,3.7084904,2.8747404,3.6594462,3.731126,3.380272,5.4778514,6.7114997,7.6923823,9.027891,10.208723,9.590013,10.650121,8.137552,5.696664,5.3684454,7.594294,8.130007,11.174516,17.610613,23.058285,17.904879,13.845533,16.810818,15.705438,12.132762,20.353312,17.28994,8.956212,4.5196047,4.979865,3.1576872,4.9421387,5.775889,5.0062733,3.561358,3.9499383,4.221567,7.009537,8.13378,7.066127,6.907676,7.6018395,7.33021,10.56335,15.513034,14.147344,8.194141,7.6584287,7.5226145,6.6020937,7.567886,8.13378,7.8810134,7.8131065,8.299775,9.073163,8.975075,8.586494,7.8508325,7.281166,7.9791017,9.065618,9.337247,7.914967,5.873977,6.25124,5.6476197,5.772116,5.8702044,5.855114,6.304056,7.01331,7.213259,6.7944975,6.1305156,6.0701537,6.511551,7.598067,8.280911,8.243186,7.9036493,6.089017,5.0968165,5.311856,6.752999,9.099571,9.525878,8.816625,8.001738,7.6622014,7.9451485,7.7829256,8.054554,8.228095,8.152642,8.043237,8.473316,8.412953,8.431817,8.4544525,7.779153,7.4584794,7.4169807,7.3981175,7.5829763,8.586494,7.997965,7.3981175,6.903904,6.590776,6.4926877,5.7419353,5.3759904,5.458988,5.975838,6.828451,7.8961043,8.043237,8.356364,9.024119,9.333474,8.492179,8.575176,9.688101,11.050018,10.963248,10.499215,10.227587,10.386037,10.944386,11.631002,11.502733,11.189606,10.95193,10.714255,10.0465,8.941121,8.239413,8.382772,8.748717,7.6584287,6.903904,6.5568223,6.0362,5.4703064,5.692891,6.2361493,6.8925858,7.33021,7.1378064,5.8211603,5.975838,5.59103,5.062863,5.142088,6.9189944,6.907676,8.035691,9.009028,9.186342,8.582722,7.443389,7.0057645,7.2962565,7.6395655,6.6360474,6.349328,6.519096,6.809588,6.9944468,6.964266,6.692637,7.039718,7.3000293,7.2623034,7.2057137,7.537705,7.6848373,8.00551,8.514814,8.884532,8.567632,8.612903,8.624221,8.386545,7.877241,8.424272,8.790216,8.718536,8.201687,7.4773426,7.3377557,7.122716,6.8359966,6.48137,6.0739264,5.9418845,6.5228686,6.79827,6.670001,6.952948,6.7341356,6.6662283,6.549277,6.33801,6.145606,5.904158,5.80607,5.938112,6.149379,6.0550632,6.587003,7.3868,8.714764,10.174769,10.740664,8.8769865,7.605612,7.17176,7.1000805,6.187105,5.2892203,5.028909,5.1458607,5.5797124,6.48137,6.9227667,7.3188925,7.7678347,8.446907,9.639057,11.276376,11.812089,12.0082655,12.091263,11.759273,11.344283,10.804798,10.167224,9.661693,9.725827,9.231613,9.231613,9.4013815,9.420244,8.990166,9.291975,9.57115,10.023865,10.416218,10.099318,10.144588,10.137043,10.080454,9.933322,9.582467,7.3075747,6.530414,6.6850915,7.3717093,8.356364,9.099571,9.548513,9.673011,9.593785,9.578695,9.971047,9.929549,10.005001,10.170997,9.827688,6.1795597,5.9607477,6.19465,6.2323766,5.945657,5.7419353,5.3194013,5.73439,6.651138,7.6810646,8.394091,7.888559,7.4282985,7.2358947,7.3679366,7.696155,7.6923823,7.360391,6.7152724,6.0626082,5.987156,6.138061,6.6813188,7.0548086,7.0585814,6.8435416,6.379509,6.187105,6.379509,6.617184,6.1041074,6.2927384,6.964266,7.3792543,7.1566696,6.2851934,5.975838,6.1342883,6.3531003,6.326692,5.8588867,6.145606,6.405917,6.7379084,7.220804,7.911195,7.809334,7.624475,7.9300575,8.797762,9.793735,9.952185,9.805053,9.627739,9.869187,11.144334,11.578186,11.706455,11.517824,10.831206,9.288202,9.016574,8.575176,8.088508,7.7150183,7.635793,7.643338,7.4773426,6.8774953,6.047518,5.643847,5.9418845,6.255012,6.7869525,7.5301595,8.280911,9.631512,10.725573,11.223559,11.223559,11.287694,10.759526,10.257768,9.759781,9.329701,9.103344,9.288202,9.416472,9.6201935,9.971047,10.472807,11.3669195,12.102581,12.872196,13.622949,14.053028,13.815352,13.739901,13.713491,13.585222,13.185325,12.838243,12.698656,12.615658,12.581704,12.717519,13.13628,13.890805,15.256495,16.98813,18.323639,19.040438,19.553514,19.70442,19.572378,19.462973,20.06282,19.994913,19.798737,19.447882,18.342503,19.108345,18.874443,18.259504,17.50498,16.486372,15.905387,14.826416,13.449409,12.106354,11.234878,10.974566,11.11038,11.442371,11.91395,12.619431,13.215506,14.053028,15.022593,16.146835,17.580433,18.402864,18.500954,18.49718,18.700903,19.093256,18.946123,18.829172,18.350048,17.746428,17.897333,18.666948,18.704676,18.685812,18.376457,16.622187,16.62973,17.048492,17.255987,17.05981,16.716501,16.22606,15.358356,14.535924,13.890805,13.253232,12.468526,12.151625,12.132762,12.200669,12.083718,12.140307,12.408164,13.155144,14.219024,15.01882,14.837734,14.335975,13.20796,11.608367,10.170997,9.646602,9.273112,8.926031,8.654402,8.6581745,8.620448,7.9338303,7.4094353,7.352846,7.5527954,7.5905213,7.3905725,7.1000805,6.779407,6.4210076,6.477597,6.560595,6.4134626,6.0248823,5.6287565,5.9682927,6.349328,6.530414,6.6020937,6.9869013,7.2170315,8.16396,9.665465,11.593277,13.894578,14.9358225,14.283158,12.864652,11.604594,11.434827,11.348056,10.597303,9.842778,9.235386,8.443134,8.616675,8.993938,9.397609,9.6201935,9.416472,8.854351,8.809079,8.831716,9.039209,10.11818,11.363147,10.593531,10.170997,10.744436,11.249968,12.185578,11.902632,11.227332,10.484125,9.476834,7.1906233,4.8553686,4.22534,5.062863,5.119452,5.036454,4.9119577,4.5950575,4.3121104,4.6742826,5.696664,6.017337,6.066381,5.9682927,5.560849,5.59103,6.4021444,7.3151197,7.394345,5.462761,4.036709,3.0633714,3.2105038,4.236658,4.9760923,6.2399216,6.4436436,6.4247804,6.4511886,6.228604,6.458734,8.83926,10.751981,10.212496,5.873977,3.9386206,2.173032,2.003264,2.9766011,2.7540162,2.6785638,3.1048703,2.1466236,0.23013012,0.10940613,0.8978847,1.1242423,1.4449154,2.9124665,6.960493,8.016829,5.7192993,3.1425967,1.6976813,1.0940613,1.4901869,1.0186088,0.482896,0.25276586,0.27917424,0.3055826,0.6828451,0.935611,0.8337501,0.392353,0.36971724,0.52062225,0.80356914,1.2449663,1.961765,3.3878171,3.863168,4.9987283,6.9454026,8.401636,7.383027,8.756263,10.397354,11.057564,10.355856,9.948412,10.450171,10.072908,8.986393,9.307066,9.042982,7.3717093,6.643593,6.319147,3.0105548,3.904667,3.3764994,2.2748928,1.327964,1.1129243,1.6486372,2.3805263,2.637065,2.5729303,3.1539145,2.727608,2.7615614,3.2029586,3.8178966,4.22534,5.4703064,5.7570257,5.945657,6.571913,7.8621507,7.9753294,8.526133,8.443134,8.039464,8.986393,9.740918,8.948667,7.907422,7.805561,9.748463,10.144588,10.33322,9.952185,9.771099,11.676274,13.170234,13.434318,12.664702,11.608367,11.551778,12.898605,13.324911,12.706201,11.800771,12.245941,11.781908,11.506506,11.34051,11.336739,11.7026825,11.314102,10.997202,10.970794,11.389555,12.321393,13.758763,14.7170105,14.588741,14.509516,17.380484,17.28994,14.50197,11.747954,9.963503,8.303548,7.956466,8.09228,7.9262853,7.598067,8.186596,9.118435,8.98262,8.299775,7.7037,7.9300575,7.0548086,5.907931,5.2590394,5.1647234,4.9534564,5.594803,5.583485,5.6363015,6.2814207,7.865923,6.9755836,4.708236,4.587512,6.168242,5.0439997,5.583485,6.6134114,5.9003854,3.7990334,3.218049,3.1840954,3.8707132,4.859141,6.0626082,7.7225633,4.821415,2.6521554,2.1956677,3.199186,4.172523,7.0510364,8.258276,9.031664,9.918231,10.789707,10.49167,8.179051,6.56814,6.643593,7.6697464,9.367428,9.352338,14.0907545,20.443855,15.690348,13.577678,19.074392,16.81459,7.575431,8.262049,8.941121,5.6551647,4.1762958,5.194905,4.285702,5.0515447,5.413717,5.27413,4.8440504,4.6554193,3.832987,6.888813,8.529905,7.3113475,5.6551647,6.9793563,7.194396,10.340765,14.992412,14.234114,10.1294985,7.8206515,6.4474163,5.8664317,6.6586833,7.6508837,7.575431,7.2924843,7.5490227,8.967529,8.552541,8.91094,8.843033,8.477088,9.273112,9.156161,8.959985,7.6282477,5.704209,5.3344917,4.779916,5.2137675,5.583485,5.6551647,5.994701,6.4511886,7.303802,7.224577,6.40969,6.587003,7.020855,7.484888,7.6848373,7.6093845,7.54525,6.0776987,4.979865,4.949684,6.228604,8.567632,8.937348,8.13378,7.2924843,7.0963078,7.7829256,7.115171,7.164215,7.575431,7.9338303,7.752744,8.001738,7.9338303,8.099826,8.303548,7.6093845,7.7942433,8.156415,8.612903,8.850578,8.318638,8.552541,8.424272,7.699928,6.7077274,6.360646,5.587258,5.7381625,6.2663302,6.8774953,7.5490227,9.031664,9.220296,9.076936,9.005256,8.869441,8.52236,8.744945,9.35611,10.193633,11.091517,11.283921,11.046246,11.012292,11.2650585,11.348056,11.00852,10.54826,10.114408,9.650374,8.873214,7.7150183,7.2962565,7.4396167,7.6697464,7.2283497,6.458734,6.25124,5.975838,5.5004873,5.191132,5.7570257,6.470052,6.8473144,6.7869525,6.598321,5.96452,5.6363015,4.881777,4.08198,4.727099,7.1264887,8.118689,8.899622,9.556059,9.065618,7.9791017,7.4094353,7.4811153,7.7225633,7.0812173,7.039718,7.356619,7.4999785,7.2698483,6.79827,6.63982,6.911449,7.3490734,7.8319697,8.375228,8.284684,8.14887,8.114917,8.171506,8.137552,8.22055,8.314865,8.329956,8.201687,7.8961043,8.27714,8.439363,8.631766,8.714764,8.152642,7.564113,7.213259,6.752999,6.224831,6.043745,5.904158,6.2021956,6.515323,6.670001,6.749226,6.4738245,6.466279,6.3417826,6.1342883,6.300284,6.5832305,6.4436436,6.598321,6.930312,6.4926877,5.975838,5.7683434,6.832224,8.714764,9.537196,8.333729,7.284939,6.7756343,6.6247296,6.0512905,5.5985756,5.2175403,5.142088,5.3873086,5.7570257,6.047518,6.428553,7.1000805,8.099826,9.333474,10.725573,11.45369,11.808316,11.944131,11.887542,11.574413,10.61994,9.80128,9.450426,9.42779,8.944894,8.858124,8.869441,8.756263,8.360137,8.763808,9.623966,10.687846,11.449917,11.148107,10.378491,9.993684,9.876732,9.81637,9.522105,7.6622014,6.673774,6.439871,6.779407,7.4282985,8.013056,8.918486,9.442881,9.522105,9.703192,9.9257765,9.548513,9.537196,9.906913,9.7296,5.8098426,6.0211096,6.3719635,6.40969,6.1078796,5.881522,5.281675,5.643847,6.360646,7.0963078,7.8017883,7.5527954,7.092535,6.8850408,7.020855,7.201941,7.4773426,7.0812173,6.2927384,5.624984,5.855114,6.4964604,7.0812173,7.3113475,7.2057137,7.141579,7.0510364,6.8435416,6.7756343,6.8058157,6.6058664,6.7114997,7.0510364,7.254758,7.17176,6.8661776,7.2094865,7.1264887,6.7077274,6.126743,5.643847,6.2663302,7.020855,7.8508325,8.597813,8.98262,8.567632,8.367682,8.914713,10.103089,11.204697,11.846043,11.838497,11.41219,11.268831,12.581704,12.253486,11.996947,11.532914,10.827434,10.099318,9.767326,9.242931,9.137298,9.337247,8.986393,8.8769865,8.239413,7.1868505,6.0739264,5.5193505,6.115425,6.85486,7.748972,8.66572,9.322156,10.012547,11.087745,11.725319,11.830952,12.049765,10.940613,10.231359,9.756008,9.457971,9.378746,9.352338,9.49947,9.869187,10.367173,10.7557535,11.649866,12.083718,12.664702,13.385274,13.630494,13.158916,13.109872,13.475817,13.879487,13.607859,13.472044,13.845533,14.385019,14.999957,15.826162,16.592005,17.391802,18.48209,19.866644,21.311558,21.300241,21.292696,21.696367,22.209444,21.82841,20.462717,20.285404,20.549488,20.730574,20.519308,20.85507,21.394556,21.09652,19.764782,18.078419,17.784155,17.157898,16.052519,14.78869,14.147344,13.313594,12.800517,12.702429,13.0646,13.917213,14.0907545,14.8339615,15.965749,17.467255,19.493153,20.187317,19.4592,18.904623,18.923487,18.731083,17.595524,17.23335,17.033401,16.848543,16.991903,17.05981,17.584206,18.033148,17.938831,16.893814,16.77309,16.58446,16.407146,16.25624,16.075155,15.784663,15.207452,14.581196,14.064346,13.721037,12.713746,12.083718,11.955449,12.162943,12.245941,12.223305,12.385528,13.060828,14.086982,14.815099,14.796235,14.5132885,13.494679,11.819634,10.106862,9.390063,8.409182,7.756517,7.6622014,8.016829,7.699928,7.194396,6.8737226,6.9265394,7.360391,7.635793,7.4094353,7.1566696,7.020855,6.8397694,6.858632,6.809588,6.4738245,5.915476,5.4703064,5.692891,6.1229706,6.72659,7.432071,8.13378,8.737399,9.87296,11.461235,13.502225,16.071383,17.105082,16.878725,15.569623,13.985121,13.5663595,13.675766,12.543978,11.136789,9.978593,9.175024,9.152389,9.442881,9.782416,9.948412,9.759781,8.175279,8.001738,8.529905,9.495697,11.083972,11.883769,11.548005,11.185833,10.948157,10.020092,11.868678,12.487389,12.528888,12.249713,11.498961,9.012801,5.855114,4.323428,4.67051,5.1081343,4.8553686,4.847823,4.7120085,4.4931965,4.659192,5.27413,5.2665844,5.6589375,6.356873,6.1644692,5.828706,6.2399216,6.398372,5.6287565,3.5500402,2.727608,2.8294687,3.7763977,5.1269975,6.1116524,6.304056,5.9192486,6.3153744,7.0170827,5.73439,6.907676,10.676529,12.034674,9.137298,3.2972744,2.4522061,1.8523588,2.1768045,3.2746384,4.1536603,2.5804756,2.2560298,1.4826416,0.23390275,0.15845025,2.7426984,2.3805263,2.7841973,4.8855495,6.8171334,5.6853456,6.017337,5.040227,2.7691069,1.9730829,0.7696155,0.7809334,0.7582976,0.392353,0.3169005,0.6413463,0.9997456,0.98842776,0.6451189,0.4376245,0.55457586,0.9695646,1.6109109,2.3767538,3.1237335,5.270357,5.281675,5.3269467,6.4247804,8.446907,7.5037513,9.650374,12.00072,12.925014,12.057309,9.348565,10.201178,10.386037,9.178797,9.352338,9.442881,6.809588,5.281675,4.930821,2.0862615,1.8033148,3.1614597,3.1916409,1.8448136,2.0108092,2.0673985,2.2371666,2.6144292,2.987919,2.837014,1.5354583,1.3392819,2.354118,3.9499383,4.7836885,6.7454534,7.624475,7.858378,7.9791017,8.616675,9.06939,10.227587,10.544487,9.763554,8.880759,9.027891,8.016829,7.2170315,7.5603404,9.559832,9.084481,10.34831,11.544232,12.344029,13.898351,12.370438,12.223305,12.540206,12.777881,12.770335,11.491416,11.087745,11.551778,12.46098,12.970284,12.468526,11.91395,11.355601,10.970794,11.072655,10.93684,10.668983,10.453944,10.378491,10.38981,12.091263,13.898351,14.320885,13.849306,14.954685,17.25976,16.32792,14.003984,11.570641,9.733373,8.865668,8.699674,8.024373,7.149124,7.8810134,9.6201935,10.001229,9.265567,8.054554,7.4018903,7.118943,6.4210076,6.039973,6.039973,5.836251,5.9607477,5.983383,6.085244,6.571913,7.8810134,7.360391,6.168242,6.360646,7.352846,5.9230213,5.9230213,4.991183,4.727099,5.3382645,5.6476197,5.670255,6.9491754,8.258276,9.367428,11.012292,7.0284004,3.9989824,3.4972234,5.081726,6.330465,9.556059,10.238904,8.854351,7.3188925,8.993938,11.502733,10.042727,8.639311,9.25425,11.785681,13.332457,12.019584,12.872196,15.977067,16.490145,16.407146,21.424738,18.915941,8.816625,3.6179473,4.8930945,4.315883,3.8707132,4.5837393,6.519096,5.3458095,5.081726,5.221313,5.342037,5.111907,3.410453,4.357382,5.764571,6.5530496,6.771862,8.394091,7.6093845,8.130007,10.597303,12.581704,11.657412,8.635539,6.3455553,5.881522,6.6247296,6.515323,7.224577,7.2283497,6.7869525,7.91874,7.3377557,8.114917,8.8618965,9.359882,10.56335,9.193887,8.284684,7.405663,6.5040054,5.934339,4.889322,4.9987283,5.3194013,5.560849,6.0776987,5.564622,6.4964604,7.2057137,7.213259,7.2283497,7.3905725,7.6584287,7.5263867,7.020855,6.677546,6.009792,5.3344917,5.3759904,6.417235,8.314865,8.431817,7.8206515,7.175533,6.903904,7.164215,6.983129,7.1566696,7.492433,7.677292,7.277394,7.2962565,7.643338,7.9715567,8.00551,7.5301595,7.9300575,8.329956,9.695646,11.034928,9.416472,9.461743,9.291975,8.465771,7.303802,6.903904,6.4134626,6.6360474,7.1302614,7.54525,7.6320205,9.159933,9.7296,9.544742,8.944894,8.394091,8.465771,8.548768,8.333729,8.461998,10.518079,11.59705,11.61214,11.419736,11.336739,11.155652,10.499215,9.940866,9.2995205,8.605357,8.099826,6.9869013,6.6813188,6.6549106,6.7680893,7.24344,6.296511,5.8588867,5.80607,5.753253,5.0553174,4.4177437,4.1762958,4.38379,4.991183,5.836251,5.7381625,5.772116,5.3571277,4.9534564,6.058836,7.6584287,7.986647,8.6732645,9.714509,9.473062,8.741172,7.809334,7.4094353,7.54525,7.454707,8.035691,8.60913,8.865668,8.616675,7.816879,7.5792036,7.326438,7.4471617,8.145098,9.405154,8.884532,8.741172,8.586494,8.265821,7.8621507,8.114917,7.8432875,7.4811153,7.3415284,7.598067,8.088508,8.2507305,8.7600355,9.408927,9.092027,7.9715567,7.2962565,6.719045,6.3229194,6.6360474,6.56814,6.096562,6.0512905,6.515323,6.8133607,6.4964604,6.4134626,6.175787,5.934339,6.387054,7.1604424,7.3792543,7.9753294,8.846806,8.884532,8.371455,7.0057645,6.6247296,7.726336,9.461743,8.809079,8.084735,7.352846,6.628502,5.8400235,5.764571,5.4250345,5.1873593,5.168496,5.2099953,5.43258,5.6098933,6.3342376,7.5829763,8.737399,9.759781,10.834979,11.446144,11.544232,11.570641,11.566868,10.804798,9.929549,9.2844305,8.941121,8.643084,8.235641,7.77538,7.5037513,7.835742,8.405409,9.740918,11.219787,12.287439,12.434572,11.216014,10.325675,9.665465,9.144843,8.677037,7.7112455,6.9793563,6.677546,6.7869525,7.069899,7.4999785,8.152642,8.82417,9.382519,9.797507,10.005001,9.631512,9.42779,9.5032425,9.329701,5.9796104,6.7379084,6.9567204,6.9189944,6.7341356,6.3342376,6.319147,6.6850915,7.032173,7.2057137,7.277394,7.24344,7.1868505,7.383027,7.726336,7.752744,7.9941926,8.058327,7.4697976,6.771862,7.492433,8.00551,8.288457,8.2507305,8.167733,8.66572,7.77538,7.141579,6.628502,6.300284,6.4247804,6.9491754,7.1793056,7.515069,8.197914,9.307066,9.989911,9.318384,8.137552,7.009537,6.2399216,6.1908774,7.624475,9.046755,9.480607,8.469543,9.224068,9.789962,10.423763,11.348056,12.740154,12.253486,11.619685,11.216014,11.314102,12.068627,11.751727,11.415963,11.0613365,10.684074,10.269085,9.695646,10.008774,10.242677,10.023865,9.597558,8.597813,7.9791017,7.4509344,7.194396,7.888559,9.0957985,9.0957985,9.231613,9.725827,9.688101,10.152134,10.801025,11.00852,10.684074,10.269085,10.133271,10.291721,10.336992,10.084227,9.597558,10.061591,11.423509,12.166716,12.294985,13.321139,12.355347,11.895086,11.970539,12.445889,13.030646,12.774108,12.664702,13.355092,14.426518,14.388792,15.769572,17.267305,18.531134,19.413929,19.987368,19.915688,19.787418,19.225298,18.795218,20.006231,17.452164,17.135263,18.297232,19.764782,19.972277,20.277859,21.24365,21.4436,20.922977,21.179516,21.534143,21.088974,20.930523,21.130472,20.75321,19.87419,19.232841,18.365139,17.493662,17.516298,16.712729,14.999957,13.913441,14.124708,15.441354,15.916705,16.98813,18.006739,18.629223,18.79899,19.078165,20.028866,20.504217,20.160908,19.440336,17.37671,16.724047,16.45619,16.21097,16.29774,16.429781,16.603323,16.625957,16.516552,16.478827,16.603323,15.954432,15.294222,15.211224,16.11288,16.271332,16.422237,16.346785,15.882751,14.894323,13.038192,11.887542,11.4838705,11.830952,12.894833,12.81938,13.057055,13.79649,14.973549,16.28265,16.086473,15.633758,14.252977,12.15917,10.438853,8.948667,7.7225633,7.0887623,7.149124,7.798016,7.673519,6.903904,6.617184,7.0812173,7.6886096,8.239413,8.073418,7.605612,7.0849895,6.6058664,7.0963078,7.1981683,6.990674,6.620957,6.300284,6.5228686,7.17176,8.118689,9.25425,10.514306,11.634775,12.740154,13.528633,14.460471,16.754227,16.840998,16.28265,15.260268,14.313339,14.373701,13.8870325,12.774108,11.389555,10.140816,9.507015,8.89585,8.650629,8.616675,8.601585,8.394091,7.598067,7.5188417,8.4544525,10.303039,12.574159,12.083718,12.310076,12.385528,11.7026825,9.933322,12.0082655,12.721292,13.219278,13.671993,13.245687,9.265567,5.9909286,4.2328854,4.1574326,5.2779026,4.5460134,3.8782585,4.025391,4.8063245,5.111907,4.8666863,4.991183,6.2851934,8.103599,8.360137,6.3945994,5.583485,4.847823,3.5236318,1.388326,2.3163917,4.3800178,6.6322746,8.065872,7.6131573,6.417235,5.715527,5.983383,6.379509,4.745962,9.250477,13.313594,12.117672,6.5568223,3.2331395,2.9313297,2.8445592,2.637065,2.5804756,3.5538127,2.323937,2.4069347,1.7165444,0.27917424,0.24522063,5.6513925,5.062863,5.0854983,7.8319697,10.895341,8.465771,8.13378,6.2851934,3.1539145,2.837014,1.3128735,1.3619176,1.146878,0.40367088,0.42630664,0.7809334,1.116697,1.0676528,0.77716076,0.9016574,1.3015556,2.2258487,3.138824,3.5877664,3.2331395,6.300284,6.2323766,6.5228686,8.009283,8.850578,8.533678,10.695392,10.899114,9.495697,11.642321,12.155397,10.929295,10.121953,10.197406,9.903141,10.291721,6.5002327,4.002755,3.893349,2.867195,1.3430545,1.8221779,2.1164427,1.8523588,2.4861598,2.0372176,2.2258487,2.969056,3.6179473,2.9615107,2.0560806,1.8674494,2.8332415,4.52715,5.6778007,8.009283,8.892077,8.771353,8.167733,7.6923823,8.288457,9.590013,11.385782,11.993175,8.269594,7.488661,5.6815734,5.413717,7.4094353,10.559577,10.291721,12.181807,15.599804,19.074392,20.29295,15.448899,12.543978,12.513797,14.675511,16.739138,11.808316,11.1782875,12.106354,12.725064,12.053536,10.759526,10.310584,10.182315,10.167224,10.374719,10.876478,10.552032,10.0276375,9.718282,9.842778,11.174516,12.0724,12.981603,13.792717,13.856852,14.698147,15.301767,14.622695,13.019329,12.238396,11.6008215,11.32542,10.133271,8.503497,8.650629,8.797762,9.265567,9.224068,8.465771,7.4169807,6.779407,6.5568223,6.5455046,6.6058664,6.6662283,5.9230213,6.2323766,6.590776,6.6850915,6.8661776,7.9300575,8.09228,7.7640624,7.24344,6.730363,4.6290107,3.0331905,2.2899833,2.7691069,4.8666863,6.6850915,7.7187905,7.462252,6.971811,8.865668,8.36391,5.775889,5.3571277,7.3075747,7.7829256,9.846551,11.404645,10.023865,6.4436436,4.561104,5.1835866,4.983638,6.149379,8.318638,8.575176,13.8719425,14.784918,12.113899,9.556059,13.717264,11.996947,18.248188,20.873934,15.494171,4.957229,7.533932,7.575431,5.492942,4.187614,9.031664,5.7117543,4.6252384,3.904667,3.059599,2.9766011,4.3422914,4.1800685,3.953711,5.406172,10.544487,15.731846,13.238141,9.125979,7.3453007,9.752235,9.322156,7.175533,5.8928404,6.3945994,7.91874,7.4169807,7.7150183,7.673519,7.394345,8.224322,7.564113,7.6848373,8.073418,8.843033,10.710483,9.808825,8.484633,7.3490734,6.8133607,7.0812173,4.8327327,4.38379,4.398881,4.5761943,5.613666,6.0776987,6.2135134,6.971811,8.194141,8.620448,9.133525,8.529905,7.6093845,6.63982,5.372218,6.432326,6.277648,6.5756855,7.7187905,8.805306,8.499724,7.3981175,6.7454534,6.6247296,5.96452,6.247467,6.673774,6.907676,7.009537,7.462252,7.364164,7.786698,8.503497,9.009028,8.544995,8.09228,7.33021,8.288457,10.306811,10.023865,8.744945,8.039464,7.7829256,7.8810134,8.269594,7.3792543,7.4207535,7.884786,8.194141,7.707473,8.511042,9.416472,9.691874,9.416472,9.491924,9.224068,8.8618965,8.91094,9.684328,11.321648,12.189351,12.038446,11.314102,10.642575,10.850069,9.8239155,9.310839,8.884532,8.356364,7.7829256,6.8661776,6.40969,6.1342883,6.1342883,6.8661776,6.462507,5.621211,5.4401255,5.7909794,5.3269467,4.7648253,4.285702,4.2781568,4.715781,5.142088,5.8626595,6.043745,5.8211603,5.7796617,6.9265394,6.670001,7.375482,8.390318,9.107117,8.971302,9.031664,8.179051,7.24344,6.771862,7.001992,8.137552,8.790216,9.35611,9.74469,9.352338,8.511042,7.914967,7.4811153,7.635793,9.307066,9.540969,9.058073,8.714764,8.59404,7.9941926,7.654656,7.201941,6.937857,7.062354,7.6584287,8.062099,7.9526935,8.428044,9.382519,9.507015,8.394091,7.4207535,6.7567716,6.488915,6.620957,6.730363,6.2097406,6.300284,7.032173,7.201941,6.115425,5.926794,6.126743,6.5228686,7.2170315,7.997965,9.144843,10.061591,11.057564,13.36641,16.712729,13.736128,9.020347,6.3644185,8.805306,9.291975,9.424017,9.125979,8.269594,6.6850915,6.156924,5.587258,5.168496,5.0741806,5.4778514,6.3945994,5.8890676,5.8890676,6.907676,8.043237,8.371455,9.699419,10.86516,11.299012,11.031156,11.363147,10.868933,9.774872,8.575176,8.024373,8.782671,8.469543,7.8810134,7.5527954,7.7376537,8.394091,9.612649,10.914205,11.9064045,12.298758,11.932813,10.77839,9.5032425,8.601585,8.409182,8.322411,7.960239,7.383027,6.851087,6.851087,7.5226145,7.8734684,8.563859,9.514561,9.918231,10.917976,10.785934,10.182315,9.718282,9.963503,6.1644692,6.930312,7.333983,7.4396167,7.3981175,7.454707,7.696155,7.5527954,7.5037513,7.533932,7.118943,7.533932,7.8961043,7.9753294,7.9225125,8.288457,8.601585,8.548768,7.960239,7.2887115,7.5792036,7.496206,7.6810646,7.6848373,7.466025,7.4094353,7.5226145,7.6886096,7.6886096,7.6508837,8.047009,9.020347,9.797507,10.461489,11.072655,11.676274,10.933067,9.4013815,8.035691,7.3113475,7.2170315,7.352846,8.635539,9.97482,10.797253,11.042474,10.989656,11.016065,11.355601,12.189351,13.619176,13.63804,13.189097,13.04951,13.196642,12.789199,12.140307,11.317875,10.819888,10.782163,11.000975,11.246195,10.676529,9.756008,9.016574,9.046755,9.035437,8.75249,8.714764,9.129752,9.914458,10.499215,9.910686,9.454198,9.465516,9.322156,10.148361,10.601076,10.650121,10.378491,9.963503,10.306811,10.827434,10.910432,10.7218,11.208468,11.291467,11.883769,12.5326605,12.777881,12.162943,12.064855,12.370438,12.366665,12.253486,13.140053,13.5663595,15.143317,16.539188,17.108854,16.91645,18.863125,19.270569,19.08571,18.787672,18.414183,17.180534,17.346529,17.071129,16.380737,17.16167,16.493916,17.040947,17.95015,18.881989,20.04773,21.719002,22.439573,22.266033,21.375692,20.081682,21.900087,21.251196,20.764528,21.417192,22.53389,22.115128,22.548979,21.28515,18.881989,18.995167,18.18028,16.81459,15.841252,15.731846,16.505234,17.780382,18.670721,19.025349,19.029121,19.18757,18.953669,20.315586,21.541689,21.70391,20.673985,19.281887,18.463226,18.101055,18.033148,18.040693,17.199398,16.708956,16.607096,16.478827,15.452672,15.01882,14.6151495,14.151116,13.970031,14.84528,15.452672,16.109108,16.429781,16.24115,15.562078,14.803781,13.7700815,12.73261,12.049765,12.174261,12.147853,12.581704,13.43809,14.68683,16.305285,16.550507,16.324148,15.456445,14.003984,12.242168,10.3634,8.756263,7.828197,7.537705,7.394345,7.2623034,6.620957,6.387054,6.85486,7.677292,8.695901,8.809079,8.345046,7.707473,7.3868,7.4773426,7.4811153,7.413208,7.284939,7.0812173,7.009537,7.383027,8.043237,8.812852,9.461743,9.442881,10.642575,12.359119,14.215251,16.16947,16.36942,16.678776,16.143063,14.875461,14.056801,13.215506,11.6875925,9.955957,8.646856,8.529905,8.729855,8.865668,8.8769865,8.533678,7.4282985,8.156415,7.960239,8.635539,10.514306,12.464753,13.147598,13.181552,12.215759,10.763299,10.212496,11.566868,11.834724,12.623203,13.615403,12.574159,9.767326,7.699928,6.330465,5.73439,6.085244,5.1269975,4.0593443,4.2781568,5.6098933,6.296511,5.3080835,5.383536,6.458734,7.7150183,7.5792036,6.2889657,4.538468,3.482133,3.1161883,2.2673476,3.0407357,5.6778007,8.458225,9.7296,7.9300575,5.515578,5.613666,5.783434,5.764571,7.4811153,13.788944,11.461235,7.0849895,3.99521,2.2447119,1.7731338,1.8976303,3.097325,4.315883,2.957738,2.757789,2.033445,1.0827434,0.36594462,0.52439487,4.7421894,6.820906,7.254758,6.0626082,2.7917426,4.678055,5.168496,4.8063245,4.214022,4.0706625,3.180323,1.901403,0.9205205,0.573439,0.84129536,0.9016574,1.2261031,1.4147344,1.4260522,1.5467763,2.5767028,3.1010978,3.338773,3.8971217,5.7607985,5.983383,5.3156285,6.277648,8.401636,8.239413,8.99771,12.140307,12.864652,10.31813,7.6018395,10.47658,8.605357,8.126234,9.171251,5.8626595,7.484888,5.975838,4.055572,2.9803739,2.5502944,2.003264,1.7655885,1.4147344,1.2185578,2.1466236,2.6597006,2.6068838,2.9124665,3.5764484,3.6669915,3.7801702,3.5462675,3.9688015,5.172269,6.40969,7.7150183,8.0206,8.228095,8.601585,8.790216,7.405663,7.654656,8.941121,10.235131,10.065364,10.367173,9.110889,7.3377557,7.2283497,12.083718,13.985121,13.370183,14.132254,17.731337,23.19787,17.991648,13.611631,12.381755,13.736128,14.237886,11.393328,11.125471,12.15917,12.694883,10.431308,9.80128,9.839006,10.069136,10.250222,10.352083,10.167224,9.763554,9.582467,9.891823,10.7557535,11.627231,11.732863,11.7894535,12.385528,13.9888935,14.226569,14.079436,13.928532,14.539697,17.05981,18.289686,17.312576,14.354838,11.34051,11.887542,11.555551,10.114408,9.118435,8.729855,7.7225633,6.9869013,6.530414,6.530414,6.771862,6.620957,6.205968,7.073672,7.5301595,7.277394,7.3905725,8.91094,9.544742,9.808825,9.846551,9.4013815,7.496206,7.122716,6.8435416,6.326692,6.356873,5.8890676,5.492942,5.20245,4.938366,4.496969,7.01331,8.00551,7.232122,5.6061206,5.1835866,8.692128,9.740918,11.197151,11.672502,5.515578,5.0741806,5.160951,8.069645,11.091517,6.511551,12.015811,13.558814,13.970031,14.750964,16.060064,11.751727,13.445636,16.52787,15.792209,5.4703064,6.8774953,5.772116,4.7120085,4.779916,5.6023483,6.1795597,5.2250857,3.9763467,3.3953626,4.1612053,4.9119577,8.197914,8.431817,7.7187905,15.863888,18.757492,11.144334,6.013564,7.009537,8.420499,7.8961043,6.930312,6.2851934,6.2851934,6.8435416,7.4773426,7.462252,7.533932,8.035691,8.933576,7.77538,8.114917,8.465771,8.2507305,7.7942433,8.160188,8.567632,8.103599,7.164215,7.4207535,4.979865,4.244203,4.255521,4.4441524,4.6629643,5.6551647,6.6322746,7.3151197,7.7037,8.073418,8.458225,8.544995,8.190369,7.1868505,5.2628117,6.432326,6.360646,6.507778,7.183078,7.54525,7.7187905,7.4396167,6.7831798,6.2399216,6.722818,7.032173,6.851087,6.56814,6.620957,7.5112963,7.352846,8.175279,10.069136,11.551778,9.533423,8.477088,8.16396,8.89585,10.31813,11.404645,11.11038,9.880505,8.741172,8.096053,7.7338815,6.881268,6.802043,7.2396674,8.047009,9.171251,9.359882,9.703192,9.97482,10.005001,9.688101,8.744945,8.480861,9.0957985,10.393582,11.785681,12.506252,11.996947,11.133017,10.412445,9.944639,9.291975,8.914713,8.627994,8.20546,7.3679366,6.7454534,6.168242,5.8588867,5.8664317,6.0739264,6.3719635,6.270103,6.126743,5.9305663,5.300538,4.45547,3.7009451,4.006528,5.081726,5.3759904,6.387054,7.454707,7.624475,7.2094865,7.7678347,6.6549106,7.0548086,8.009283,8.726082,8.582722,8.699674,8.563859,7.914967,7.0812173,6.990674,7.9526935,8.650629,9.337247,9.80128,9.4013815,8.7751255,8.299775,7.752744,7.564113,8.809079,8.480861,8.096053,7.9338303,7.8206515,7.115171,6.560595,6.911449,7.5226145,7.8734684,7.575431,8.379,8.586494,8.620448,8.650629,8.627994,8.152642,7.7037,7.3075747,6.900131,6.3417826,6.0512905,6.628502,6.9454026,6.6813188,6.3342376,6.56814,7.220804,7.183078,6.700182,7.375482,8.273367,9.310839,10.589758,12.608112,16.271332,18.150099,13.705947,8.560086,6.1833324,7.8998766,8.692128,8.993938,8.620448,7.937603,7.8432875,6.730363,6.485142,6.096562,5.3156285,4.636556,5.511805,5.775889,5.873977,6.145606,6.820906,7.111398,8.013056,9.231613,10.442626,11.287694,11.1782875,10.880251,9.906913,8.586494,8.073418,8.382772,7.605612,7.1000805,7.281166,7.6018395,7.4396167,8.307321,9.6201935,10.910432,11.796998,12.340257,12.264804,10.884023,8.793989,7.84706,8.103599,8.209232,8.0206,7.61693,7.303802,7.6622014,7.9489207,8.669493,9.556059,9.590013,9.740918,10.140816,10.585986,10.95193,11.197151,6.1833324,6.651138,6.809588,7.069899,7.541477,8.058327,8.2507305,8.084735,7.786698,7.462252,7.0812173,7.745199,8.186596,8.360137,8.428044,8.7600355,9.148616,9.137298,9.016574,8.880759,8.624221,8.465771,8.443134,8.560086,8.688355,8.560086,8.699674,8.873214,8.975075,9.0543,9.314611,10.472807,11.574413,12.306303,12.47607,12.019584,10.86516,9.491924,8.409182,7.9715567,8.367682,9.231613,10.38981,11.589504,12.600568,13.200415,12.721292,12.178034,11.891314,12.140307,13.162688,13.36641,13.241914,12.97783,12.619431,12.064855,11.676274,11.283921,11.276376,11.563096,11.59705,11.11038,10.087999,9.084481,8.677037,9.469289,10.287949,10.272858,10.148361,10.321902,10.906659,10.668983,10.336992,10.076681,10.020092,10.265312,10.808571,11.121698,11.446144,11.763044,11.800771,11.92904,11.623458,11.136789,10.79348,10.989656,11.102836,11.223559,11.634775,12.106354,11.917723,12.325166,12.766563,12.974057,13.158916,14.019074,14.030393,15.339493,16.94286,17.659658,16.146835,17.18808,17.282394,17.595524,18.30855,18.606586,16.735365,17.244669,17.580433,17.338985,18.251959,18.561316,18.976303,19.636513,20.345766,20.568352,21.21347,21.503962,21.617142,21.651094,21.598278,23.41291,22.77911,22.03213,22.367893,23.850534,24.005213,23.775084,22.303759,20.179771,19.436563,18.663176,17.603067,16.38451,15.588487,16.229834,18.319866,19.534653,20.081682,20.23636,20.330677,20.602304,21.639776,22.375439,22.416937,22.024584,21.439827,20.632486,20.16468,20.100546,20.017548,18.342503,17.37671,17.274849,17.437073,16.497688,15.505488,14.943368,14.418973,13.958713,13.966258,14.5132885,15.471535,16.180788,16.260014,15.641303,15.01882,13.902123,12.596795,11.566868,11.434827,11.446144,11.7026825,12.404391,13.592768,15.158407,15.543215,15.629986,15.301767,14.5132885,13.264549,11.506506,10.001229,8.748717,7.798016,7.220804,7.1378064,6.5832305,6.4134626,6.8774953,7.6395655,8.465771,8.571404,8.130007,7.435844,6.907676,6.8359966,6.9152217,6.8774953,6.617184,6.198423,6.1606965,6.5530496,7.1566696,7.77538,8.201687,8.307321,8.914713,10.110635,11.774363,13.577678,14.864142,15.70921,16.403374,16.908905,16.859861,15.999702,14.241659,11.778135,9.408927,8.552541,8.756263,9.084481,9.258021,9.152389,8.778898,9.450426,9.171251,9.537196,11.00852,12.913695,13.505998,12.883514,11.548005,10.329447,10.386037,10.831206,10.921749,11.442371,12.113899,11.6008215,10.272858,9.34102,8.337502,7.0963078,5.783434,5.1873593,4.06689,4.187614,5.670255,6.9869013,5.828706,5.956975,6.651138,7.3113475,7.466025,6.6360474,4.666737,3.2633207,3.006782,3.338773,3.8820312,5.194905,7.164215,8.507269,6.7756343,4.7912335,5.111907,5.191132,5.873977,11.378237,11.657412,7.0246277,3.5953116,2.7426984,1.1016065,1.2110126,4.063117,6.1833324,5.6400743,2.022127,2.9086938,2.1881225,1.3015556,1.2525115,2.6182017,5.8400235,7.986647,7.643338,5.251494,3.078462,3.9876647,4.217795,4.538468,5.111907,5.4967146,3.2029586,1.5316857,0.95824677,1.3392819,1.9164935,1.7882242,2.123988,2.0749438,1.7052265,2.003264,2.7540162,3.7462165,4.2781568,4.5988297,5.9192486,5.560849,5.4967146,8.028146,12.019584,12.902377,11.415963,13.536179,14.475562,12.00072,6.436098,9.559832,8.118689,7.322665,7.575431,4.485651,5.9532022,5.5457587,4.293247,3.0746894,2.5729303,1.9164935,1.901403,2.3126192,2.8634224,3.2029586,2.9426475,2.8407867,3.338773,4.304565,5.0175915,4.357382,3.6934,3.7084904,4.557331,5.8966126,6.960493,6.802043,6.6662283,7.141579,8.14887,6.971811,7.4169807,8.544995,9.442881,9.205205,10.789707,9.884277,8.103599,7.54525,10.774617,13.630494,13.072145,12.249713,13.747445,19.595015,16.429781,12.736382,11.208468,11.898859,12.2270775,10.978339,10.838752,10.921749,10.536942,9.175024,9.756008,9.97482,9.95973,9.74469,9.246704,8.8618965,8.801534,9.110889,9.861642,11.170743,12.4307995,12.777881,12.687338,12.883514,14.324657,14.490653,14.468017,14.4114275,14.777372,16.305285,17.20317,17.1164,15.445127,13.0646,12.321393,11.083972,9.092027,8.416726,8.899622,8.16396,7.333983,6.7756343,6.6662283,6.934085,7.2472124,6.9755836,7.4509344,7.4396167,6.9265394,7.0849895,9.099571,10.608622,11.189606,11.057564,11.042474,10.080454,9.122208,8.846806,9.231613,9.556059,9.310839,7.665974,6.4964604,6.085244,5.1345425,6.25124,7.254758,8.386545,8.514814,5.1345425,6.560595,8.499724,11.657412,14.320885,12.381755,11.853588,10.257768,11.3820095,12.491161,4.293247,7.960239,10.570895,12.740154,14.551015,15.565851,10.993429,10.484125,10.808571,9.563604,5.1798143,5.0968165,4.172523,3.5839937,3.6330378,3.7575345,6.1720147,5.80607,5.5268955,5.8928404,5.1798143,4.496969,7.352846,8.333729,7.865923,12.2270775,11.819634,8.526133,7.1378064,8.2507305,8.262049,7.33021,7.0170827,7.250985,7.5301595,6.934085,7.4396167,7.009537,7.5188417,9.0807085,10.035183,8.933576,8.439363,8.27714,8.13378,7.6584287,7.748972,8.084735,7.8206515,7.0585814,6.828451,4.983638,4.346064,4.459243,4.8440504,5.0025005,5.624984,6.2927384,6.7341356,7.0284004,7.586749,7.6320205,8.122461,8.36391,8.028146,7.1302614,7.496206,7.3113475,7.322665,7.424526,6.6549106,6.85486,7.201941,6.8359966,6.0626082,6.3531003,7.4018903,7.254758,6.590776,6.168242,6.828451,6.9265394,8.001738,10.11818,11.721546,9.623966,8.59404,8.631766,8.654402,8.8618965,10.740664,10.589758,9.8239155,8.846806,8.099826,8.047009,7.496206,7.141579,7.3113475,8.099826,9.352338,9.529651,9.529651,9.590013,9.552286,8.865668,8.45068,8.903395,9.869187,11.148107,12.698656,12.853333,11.895086,10.989656,10.408672,9.510788,9.540969,9.480607,9.1825695,8.503497,7.3075747,6.560595,6.0776987,5.7683434,5.613666,5.674028,6.149379,6.2851934,6.0701537,5.6778007,5.458988,4.5950575,3.9801195,3.8103511,4.036709,4.3875628,5.7306175,6.9227667,7.2396674,6.8850408,6.990674,6.270103,7.0774446,8.314865,9.107117,8.812852,8.786444,8.695901,8.45068,8.171506,8.197914,8.586494,9.14107,9.593785,9.782416,9.635284,9.076936,8.835487,8.529905,8.341274,9.031664,8.748717,8.431817,8.239413,8.099826,7.7112455,7.2698483,7.2887115,7.6923823,8.16396,8.130007,8.899622,8.816625,8.646856,8.59404,8.307321,7.907422,7.6093845,7.3905725,7.1038527,6.4738245,6.462507,6.9454026,7.149124,6.9152217,6.6850915,7.073672,7.8131065,8.122461,7.91874,7.828197,8.431817,8.537451,8.782671,9.6051035,11.257513,12.253486,9.748463,7.3679366,6.590776,6.760544,7.786698,8.952439,9.265567,8.639311,7.8961043,7.250985,6.722818,6.4134626,6.1041074,5.247721,5.1345425,5.372218,5.7004366,5.8966126,5.7570257,6.3644185,7.322665,8.160188,8.9788475,10.438853,10.34831,10.265312,9.891823,9.26934,8.790216,8.643084,8.337502,8.035691,7.8621507,7.907422,7.7301087,8.303548,9.14107,9.971047,10.7557535,11.657412,12.400619,11.763044,9.789962,7.798016,8.050782,8.944894,9.64283,9.646602,8.790216,8.103599,8.035691,8.797762,10.155907,11.419736,10.612394,9.982366,10.144588,10.974566,11.604594,5.987156,6.2889657,6.326692,6.7454534,7.6508837,8.601585,8.75249,8.714764,8.394091,7.964011,7.9036493,8.616675,8.929804,9.156161,9.4127,9.6051035,10.012547,10.287949,10.702937,10.974566,10.291721,10.359629,10.56335,10.940613,11.291467,11.170743,10.970794,10.506761,10.174769,10.133271,10.303039,11.09529,12.196897,12.966512,13.008011,12.166716,11.404645,10.484125,9.752235,9.601331,10.435081,11.589504,12.344029,13.057055,13.788944,14.27184,13.577678,12.925014,12.457208,12.264804,12.381755,12.057309,11.695138,11.566868,11.574413,11.257513,11.159425,11.174516,11.359374,11.498961,11.076427,10.050273,9.450426,9.442881,10.137043,11.581959,12.1252165,12.2270775,11.981857,11.642321,11.608367,11.102836,11.027383,11.034928,11.053791,11.314102,11.570641,11.936585,12.347801,12.672247,12.740154,12.58925,11.846043,11.117926,10.691619,10.536942,10.838752,11.000975,11.2650585,11.676274,12.057309,12.740154,13.321139,13.626721,13.792717,14.283158,14.407655,14.84528,16.075155,17.150352,15.701665,16.36942,16.874952,18.029375,19.38752,19.240387,18.248188,19.010258,19.281887,18.976303,20.130728,19.798737,19.960958,20.700394,21.31533,20.30804,20.017548,20.296722,20.934296,21.805773,22.877197,24.054256,23.55627,22.586706,22.232079,23.4695,23.997667,23.45441,22.17549,20.673985,19.625195,18.599041,17.738882,16.761772,16.056292,16.724047,19.323385,20.711712,21.436056,21.888771,22.277351,22.035902,22.005722,21.918951,21.67373,21.322876,20.934296,20.304268,19.923233,19.896824,19.923233,18.331184,17.516298,17.60684,18.03692,17.512526,16.195879,15.686575,15.645076,15.603577,14.969776,14.852824,15.546988,15.954432,15.671484,14.999957,13.860624,12.917468,11.996947,11.204697,10.891568,11.00852,11.336739,12.091263,13.223051,14.43029,14.743419,14.679284,14.354838,13.807808,12.989148,11.664956,10.56335,9.359882,8.145098,7.4584794,7.2698483,6.7454534,6.5756855,6.9491754,7.5603404,8.258276,8.265821,7.8621507,7.3151197,6.858632,6.8246784,6.9189944,6.888813,6.617184,6.089017,6.006019,6.296511,6.7680893,7.284939,7.756517,8.258276,8.394091,8.782671,9.703192,11.106608,13.075918,14.407655,15.433809,16.199652,16.459963,16.754227,16.373192,14.468017,11.5857315,9.639057,9.152389,9.280658,9.737145,10.269085,10.63503,11.185833,10.782163,10.808571,11.581959,12.340257,13.038192,12.325166,11.378237,10.812344,10.672756,9.989911,9.725827,9.948412,10.419991,10.56335,10.450171,9.944639,9.201432,8.028146,5.8928404,5.564622,4.606375,4.606375,5.8211603,7.164215,6.375736,6.5266414,6.7643166,6.94163,7.6131573,6.8133607,5.304311,4.063117,3.8405323,5.1647234,5.4174895,5.6891184,6.4738245,7.2283497,6.3531003,5.4665337,5.1873593,5.7117543,7.835742,12.951422,8.062099,4.164978,2.505023,2.3465726,0.9620194,1.9579924,6.94163,8.986393,6.930312,5.353355,4.825187,2.9539654,3.289729,5.7079816,6.3832817,7.175533,7.2358947,6.092789,4.504514,4.447925,4.402653,3.8820312,4.032936,4.6290107,4.074435,2.0900342,1.177059,1.4637785,2.546522,3.4896781,3.289729,2.886058,2.3201644,1.961765,2.5012503,3.127506,4.3422914,5.13077,5.0968165,4.478106,5.349582,5.6287565,9.442881,15.452672,16.874952,12.774108,12.253486,12.574159,11.3820095,6.6813188,8.213005,7.7225633,6.9793563,6.187105,4.002755,5.3382645,5.383536,4.6818275,3.7499893,3.0860074,2.033445,2.4069347,3.2029586,3.7801702,3.8707132,2.9011486,2.7389257,3.4029078,4.557331,5.5306683,4.4894238,3.7650797,3.3764994,3.5236318,4.5761943,5.50426,5.726845,5.670255,5.9003854,7.122716,6.620957,7.2924843,8.013056,8.080963,7.201941,9.680555,9.318384,8.307321,8.175279,9.820143,12.611885,12.015811,10.499215,11.038701,17.093763,16.573141,13.091009,11.140562,11.5857315,11.661184,11.076427,10.544487,9.654147,8.820397,9.26934,10.518079,10.616167,10.238904,9.680555,8.850578,8.480861,8.59404,9.159933,10.072908,11.121698,12.31762,12.781653,12.755245,12.725064,13.385274,14.358611,15.022593,14.803781,13.856852,13.053283,13.773854,14.905642,14.664193,13.075918,11.955449,10.306811,8.892077,8.699674,9.288202,8.786444,7.8696957,7.462252,7.273621,7.2924843,7.809334,7.586749,7.5829763,7.224577,6.7341356,7.115171,8.8618965,10.887795,11.868678,11.706455,11.548005,11.566868,10.18986,9.7220545,10.616167,11.476325,11.642321,10.612394,9.363655,8.167733,6.590776,6.8058157,7.0887623,9.397609,11.951676,9.220296,6.937857,8.16396,10.691619,13.087236,14.713238,15.863888,16.622187,16.422237,13.381501,4.285702,7.220804,9.507015,11.068882,11.898859,12.038446,8.348819,7.956466,7.1868505,5.4703064,5.3609,4.142342,3.2331395,3.7537618,5.2137675,5.5193505,6.771862,6.4738245,6.3908267,7.073672,7.828197,5.160951,5.9192486,6.990674,7.3113475,7.8810134,6.760544,7.0548086,7.624475,7.9715567,8.231868,7.326438,8.597813,9.971047,10.016319,7.99042,7.798016,6.7643166,7.5301595,9.891823,10.77839,10.495442,9.242931,8.224322,7.8998766,7.9791017,7.61693,7.364164,7.1679873,6.8699503,6.2135134,5.0251365,4.466788,4.5120597,4.961002,5.4401255,5.8890676,6.25124,6.3908267,6.439871,6.7643166,6.8925858,7.6131573,8.080963,8.122461,8.231868,8.137552,7.7301087,7.492433,7.352846,6.6850915,6.4738245,6.85486,6.9454026,6.6624556,6.72659,7.6622014,7.541477,6.760544,6.0248823,6.319147,7.001992,8.3525915,10.201178,11.25374,9.110889,8.4544525,8.82417,8.469543,7.911195,9.9257765,10.091772,9.7069645,8.944894,8.209232,8.152642,7.7301087,7.4396167,7.598067,8.243186,9.114662,9.540969,9.424017,9.103344,8.646856,7.865923,8.356364,9.186342,10.314357,11.781908,13.698401,13.694629,12.00072,10.702937,10.246449,9.454198,9.805053,9.778644,9.431562,8.737399,7.5603404,6.541732,5.9909286,5.7079816,5.5683947,5.5193505,5.8890676,6.228604,6.0739264,5.523123,5.251494,4.745962,4.1800685,3.4896781,2.969056,3.2670932,4.7535076,5.9909286,6.330465,5.915476,5.66271,5.8626595,6.8473144,8.0206,8.888305,9.06939,9.159933,8.8769865,8.699674,8.786444,8.9788475,9.107117,9.537196,9.737145,9.714509,9.993684,9.767326,9.4127,9.224068,9.273112,9.420244,9.167479,8.888305,8.575176,8.258276,8.016829,8.167733,8.028146,7.9338303,8.039464,8.329956,8.967529,8.228095,7.654656,7.677292,7.647111,7.699928,7.699928,7.54525,7.284939,7.118943,7.152897,7.1906233,7.2057137,7.1868505,7.1302614,7.5112963,7.9715567,8.45068,8.643084,7.986647,8.088508,7.6093845,7.183078,7.1264887,7.424526,8.737399,8.692128,8.405409,8.062099,6.930312,8.8769865,10.069136,10.065364,9.118435,8.156415,7.484888,6.749226,6.387054,6.2889657,5.8173876,5.2175403,5.149633,5.379763,5.455216,4.7233267,5.3684454,6.5756855,7.454707,7.967784,8.952439,9.691874,9.835234,9.759781,9.597558,9.261794,8.7751255,9.012801,9.016574,8.639311,8.552541,8.179051,8.296002,8.688355,9.231613,9.884277,10.816116,11.970539,12.2270775,11.027383,8.390318,8.360137,9.352338,10.329447,10.665211,10.11818,9.016574,8.677037,9.231613,10.638803,12.694883,12.083718,10.499215,9.861642,10.574668,11.54046,5.7570257,6.145606,6.3455553,6.8661776,7.8508325,9.06939,9.454198,9.548513,9.390063,9.242931,9.601331,10.291721,10.450171,10.627484,10.921749,10.955703,11.283921,11.910177,12.596795,12.894833,12.147853,12.464753,13.238141,13.853079,14.019074,13.751218,12.992921,11.876224,11.076427,10.86516,11.106608,11.461235,12.385528,13.155144,13.340002,12.800517,12.67602,12.185578,11.6875925,11.680047,12.800517,13.585222,13.641812,13.705947,13.9888935,14.177525,13.189097,12.762791,12.555296,12.291212,11.732863,10.759526,9.993684,10.186088,10.974566,10.861387,10.725573,10.763299,10.804798,10.653893,10.084227,9.314611,9.695646,10.963248,12.66093,14.136025,13.977575,14.147344,13.951167,13.27964,12.630749,12.415709,12.102581,11.947904,11.966766,11.932813,12.095036,12.649611,12.883514,12.596795,12.113899,11.7894535,11.336739,10.925522,10.646348,10.514306,10.895341,11.400873,11.7026825,11.921495,12.642066,13.4644985,14.279386,14.535924,14.27184,14.1058445,14.826416,14.769827,15.573396,17.014538,16.999449,17.886015,19.017803,20.413673,21.05502,18.863125,19.553514,20.602304,20.304268,19.217752,20.160908,18.908396,18.946123,19.794964,20.421219,19.21398,18.923487,19.413929,20.455173,21.760502,22.982832,23.511,23.43932,22.673477,21.941587,22.813063,23.103556,22.93756,22.100037,20.828663,19.810055,18.685812,17.969013,17.655886,17.738882,18.172735,20.564579,21.737865,22.258488,22.696112,23.620405,22.013268,20.689075,20.213724,20.232588,19.455427,18.678267,18.070873,17.957695,18.221779,18.312323,17.28994,16.920223,17.1164,17.538933,17.587978,16.320375,16.063837,16.837225,17.844517,17.486116,16.716501,16.52787,16.056292,15.169725,14.452927,12.940104,12.287439,11.951676,11.574413,10.982111,11.291467,11.932813,12.853333,13.837989,14.50197,14.520834,14.064346,13.479589,12.887287,12.170488,11.261286,10.552032,9.646602,8.605357,7.9526935,7.594294,7.115171,6.8774953,7.0170827,7.435844,8.209232,8.228095,7.9753294,7.699928,7.4471617,7.492433,7.4509344,7.4169807,7.33021,6.9793563,6.6586833,6.688864,6.964266,7.424526,8.058327,8.722309,8.89585,8.91094,9.152389,10.065364,12.2270775,13.992666,14.400109,13.800262,13.853079,15.531898,16.74291,16.033657,13.50977,10.853842,9.703192,9.178797,9.857869,11.234878,11.721546,12.513797,12.00072,11.717773,11.815862,11.076427,12.2119875,12.106354,11.834724,11.676274,11.136789,9.393836,8.367682,8.341274,9.016574,9.525878,10.197406,9.669238,9.14107,8.605357,6.8397694,6.609639,5.9003854,5.832478,6.537959,7.17176,6.8925858,6.8850408,6.587003,6.4134626,7.752744,7.443389,6.4738245,5.6325293,5.692891,7.4282985,7.997965,7.6018395,7.073672,6.79827,6.7114997,7.232122,6.4134626,8.09228,11.465008,11.091517,5.458988,3.5877664,2.886058,2.516341,3.3915899,5.5004873,9.7296,10.065364,7.635793,10.733118,7.2396674,3.5651307,4.9949555,9.631512,8.390318,6.63982,5.2892203,4.2706113,3.802806,4.38379,4.5233774,3.5274043,3.0030096,2.8030603,1.0223814,1.0751982,1.4826416,2.704972,4.376245,5.311856,5.0968165,3.5274043,2.5804756,2.8445592,3.5160866,4.142342,5.3646727,6.039973,5.3382645,2.7238352,5.451443,5.534441,9.718282,17.074902,18.99894,12.536433,9.1976595,9.246704,10.487898,8.27714,6.9793563,7.360391,7.0585814,5.455216,3.651901,5.6098933,6.017337,5.7004366,5.100589,4.2592936,2.8030603,3.2859564,3.6028569,3.2859564,3.4745877,2.4823873,2.1541688,2.686109,3.7914882,4.715781,4.4743333,3.9763467,3.1614597,2.5616124,3.2821836,3.8971217,4.9345937,5.4778514,5.6023483,6.368191,6.217286,6.6850915,6.7341356,6.1833324,5.7117543,8.624221,9.065618,8.850578,9.076936,10.11818,11.729091,10.687846,9.314611,10.431308,17.384256,19.047983,15.192361,12.672247,13.019329,12.453435,11.808316,10.767072,9.495697,8.858124,10.419991,11.359374,11.216014,10.718028,10.201178,9.6051035,9.314611,9.314611,9.793735,10.480352,10.631257,11.068882,11.302785,11.408418,11.415963,11.317875,13.211733,14.656648,14.335975,12.336484,10.148361,11.800771,13.664448,13.687083,12.215759,11.970539,11.336739,10.823661,10.461489,10.178542,9.782416,8.590267,8.201687,7.8206515,7.3717093,7.4811153,7.496206,7.443389,7.1793056,7.009537,7.6886096,8.624221,10.442626,11.830952,12.166716,11.506506,12.0233555,10.967021,10.272858,10.593531,11.310329,11.348056,12.162943,11.736636,9.81637,7.8998766,8.416726,8.360137,9.914458,12.679792,13.690856,9.548513,8.948667,9.288202,9.691874,11.027383,13.230596,18.365139,18.817854,13.189097,6.2625575,9.933322,10.967021,10.3634,9.190115,8.586494,5.583485,7.3377557,8.786444,8.567632,9.042982,5.907931,3.440634,5.1760416,9.314611,8.695901,7.118943,6.888813,6.270103,6.0512905,9.522105,6.398372,5.624984,6.1116524,6.741681,6.356873,6.749226,6.692637,6.6134114,7.0812173,8.82417,9.167479,15.475307,18.38023,15.067864,9.2844305,8.152642,6.8737226,7.6093845,9.906913,10.70671,11.419736,10.38981,8.926031,7.9338303,7.907422,7.4094353,6.749226,6.598321,6.7379084,6.0550632,5.2099953,4.6252384,4.38379,4.5988297,5.4212623,6.1003346,6.4021444,6.326692,6.009792,5.7381625,6.066381,6.9793563,7.537705,7.6320205,7.9791017,8.114917,7.5716586,7.0774446,6.9491754,7.111398,6.511551,6.4926877,6.85486,7.3453007,7.6584287,7.6923823,7.4207535,6.8473144,6.2889657,6.3945994,7.4396167,8.899622,10.223814,10.502988,8.465771,8.280911,8.8618965,8.661947,8.145098,9.759781,10.374719,10.084227,9.322156,8.431817,7.654656,7.1340337,7.1981683,7.643338,8.235641,8.741172,9.242931,9.216523,8.6581745,7.828197,7.2283497,8.303548,8.99771,10.18986,12.038446,13.9888935,13.600313,11.548005,10.155907,9.903141,9.431562,9.74469,9.446653,9.06939,8.707218,8.031919,6.851087,6.0286546,5.692891,5.674028,5.4891696,5.73439,6.1833324,6.221059,5.692891,4.9119577,4.8629136,4.2027044,3.2972744,2.6295197,2.7804246,4.0895257,5.27413,5.4891696,4.859141,4.429062,5.5457587,6.3342376,7.1076255,8.031919,9.125979,9.405154,9.009028,8.646856,8.639311,8.914713,9.2844305,9.597558,9.767326,9.963503,10.597303,10.676529,9.948412,9.608876,9.827688,9.737145,9.280658,8.937348,8.518587,8.016829,7.6093845,8.337502,8.488406,8.107371,7.6282477,7.8621507,8.360137,7.122716,6.156924,6.255012,6.990674,7.647111,7.9715567,7.77538,7.435844,7.8734684,7.677292,7.4773426,7.322665,7.254758,7.273621,7.9941926,8.179051,8.397863,8.563859,7.914967,7.6810646,7.2962565,7.0963078,7.322665,8.141325,10.321902,12.483616,13.008011,11.604594,9.2844305,12.283667,12.106354,10.408672,8.7751255,8.748717,7.5905213,6.851087,6.224831,5.7494807,5.8098426,5.6098933,5.3269467,5.160951,4.961002,4.22534,4.353609,5.59103,6.9265394,7.7112455,7.677292,9.344792,9.782416,9.714509,9.537196,9.310839,8.684583,9.148616,9.5032425,9.390063,9.25425,8.394091,8.031919,8.254503,8.854351,9.337247,10.080454,11.32542,12.336484,12.136535,9.510788,8.993938,9.205205,9.710737,10.238904,10.691619,10.103089,9.74469,9.952185,10.868933,12.438345,13.053283,11.532914,10.246449,10.212496,11.140562,5.904158,6.428553,6.85486,7.2887115,7.911195,8.971302,10.11818,10.352083,10.4049,10.725573,11.442371,12.310076,12.528888,12.691111,12.883514,12.664702,12.785426,13.347548,13.781399,13.856852,13.687083,13.894578,14.852824,15.297995,14.898096,14.252977,12.419481,11.714001,11.544232,11.59705,11.84227,12.913695,13.898351,14.381247,14.2077055,13.472044,13.27964,13.328684,12.96274,12.543978,13.472044,13.766309,13.117417,13.030646,13.58145,13.396591,11.676274,11.072655,10.7557535,10.585986,11.125471,10.940613,11.09529,11.02361,10.665211,10.484125,9.861642,9.767326,10.148361,10.691619,10.86516,10.642575,11.506506,12.713746,13.671993,13.917213,14.939595,15.433809,15.271586,14.7170105,14.449154,14.351066,13.147598,12.128989,11.872451,12.238396,12.272349,12.90615,13.166461,12.672247,11.61214,10.929295,10.61994,10.608622,10.710483,10.63503,10.684074,11.246195,11.7026825,12.336484,14.313339,15.214996,15.871433,16.275105,16.203424,15.226315,15.313085,15.728074,17.18808,19.040438,19.270569,19.063074,20.074137,20.862616,19.960958,15.882751,16.652367,18.41041,18.361366,16.618414,16.203424,17.180534,16.822134,16.874952,17.738882,18.433046,18.248188,18.157644,19.24416,21.322876,22.933788,23.190327,24.242887,24.895552,25.0955,25.92548,24.899324,24.393793,23.726038,22.311304,19.700647,19.893051,19.364883,19.232841,19.455427,18.844261,19.821371,20.560806,20.628714,20.485353,21.4851,20.043957,18.21046,18.429274,20.258997,20.372175,19.417702,18.070873,18.13878,19.191343,18.568861,17.01831,16.28265,15.852571,15.841252,17.014538,16.195879,15.754482,16.490145,18.135008,19.31584,19.183798,17.769064,16.72782,16.392056,15.746937,15.309312,14.347293,13.570132,13.083464,12.37421,12.887287,13.4644985,14.019074,14.43029,14.524607,13.93985,13.830443,13.837989,13.611631,12.815607,11.827179,11.042474,10.084227,8.990166,8.209232,8.024373,7.7602897,7.432071,7.1793056,7.277394,7.865923,8.2507305,8.439363,8.265821,7.3868,7.273621,7.020855,6.8737226,6.881268,6.881268,6.296511,6.270103,6.620957,7.213259,7.9338303,8.52236,9.190115,9.559832,9.869187,10.955703,14.007756,15.833707,16.21097,16.048746,17.380484,17.916197,16.74291,14.849052,12.706201,10.253995,9.789962,8.265821,8.729855,10.929295,11.306557,12.049765,11.604594,11.11038,11.076427,11.3820095,12.113899,12.528888,12.166716,11.45369,11.672502,9.548513,7.360391,6.7379084,7.647111,8.394091,9.639057,9.80128,9.631512,9.205205,7.9489207,8.167733,7.7225633,7.624475,7.9300575,7.7225633,7.2924843,6.7756343,5.772116,5.300538,7.7678347,10.4049,8.873214,7.598067,8.088508,8.941121,11.736636,9.046755,6.6058664,6.2097406,5.723072,8.284684,8.98262,12.344029,15.275358,7.0510364,3.5462675,2.5502944,2.003264,3.1124156,10.374719,14.075664,13.230596,9.461743,6.277648,9.110889,5.5570765,2.425798,1.3958713,2.0560806,1.9089483,1.81086,4.908185,5.670255,3.9914372,5.1873593,3.5538127,3.289729,2.3088465,0.91297525,1.8146327,1.9240388,2.8407867,5.0251365,7.3377557,7.0359454,6.741681,5.0213637,4.432834,5.3080835,5.7381625,5.406172,7.567886,8.099826,5.8136153,2.4559789,5.726845,5.9796104,9.593785,17.048492,22.918697,12.67602,8.854351,11.827179,16.550507,12.574159,8.141325,8.646856,8.216777,5.5080323,3.6783094,7.069899,8.311093,8.367682,7.7037,6.2851934,4.1762958,4.3611546,4.1536603,2.9954643,2.4710693,1.569412,0.9393836,1.177059,2.1654868,3.0671442,4.214022,3.31991,2.11267,1.8297231,3.218049,3.4745877,4.217795,5.0062733,5.5759397,5.8437963,5.8702044,5.983383,5.666483,5.372218,6.530414,9.850324,11.083972,10.967021,10.359629,10.238904,9.21275,9.359882,8.98262,9.65792,16.252468,19.289433,16.90136,14.649103,14.237886,13.502225,12.917468,12.321393,11.480098,10.736891,11.016065,10.944386,10.77839,10.627484,10.559577,10.61994,10.435081,10.419991,10.56335,10.54826,9.703192,9.495697,9.884277,10.386037,10.536942,9.903141,10.967021,12.657157,12.736382,11.189606,10.223814,13.445636,15.203679,14.622695,12.789199,12.740154,15.475307,14.822643,13.117417,11.819634,11.491416,9.450426,8.035691,6.937857,6.0286546,5.3571277,6.270103,6.7643166,7.001992,7.2887115,8.058327,8.8618965,9.778644,11.11038,12.351574,12.193124,12.37421,11.5857315,10.702937,10.26154,10.469034,10.650121,11.619685,11.476325,10.525623,11.306557,9.842778,9.239159,8.646856,8.296002,9.491924,10.370946,10.819888,10.140816,8.8769865,8.805306,5.9117036,7.33021,9.461743,9.88805,7.3868,10.838752,12.479843,10.785934,8.296002,11.627231,7.598067,12.96274,18.387774,20.319359,20.979568,12.253486,5.300538,6.1003346,11.027383,6.851087,4.398881,6.273875,6.7077274,4.5535583,3.2972744,5.1156793,5.6325293,5.80607,6.089017,6.4549613,6.270103,5.704209,7.254758,10.499215,12.083718,15.746937,34.093212,39.19003,25.431265,9.552286,7.220804,7.224577,7.9451485,8.68081,9.64283,10.182315,11.046246,10.914205,9.6051035,8.103599,7.3717093,6.6020937,6.3644185,6.5568223,6.40969,5.553304,5.0477724,4.4931965,4.1612053,5.0062733,5.66271,5.5193505,5.4740787,5.613666,5.1873593,4.5912848,5.7683434,7.164215,7.9300575,7.9036493,8.439363,8.152642,7.726336,7.2698483,6.3153744,6.2436943,6.115425,6.006019,6.1418333,6.911449,6.937857,6.651138,6.5832305,6.809588,6.94163,7.039718,7.8998766,8.465771,8.4544525,8.329956,8.488406,8.903395,8.967529,8.941121,9.978593,10.076681,10.182315,9.695646,8.473316,6.8359966,6.3342376,6.458734,7.0359454,7.7150183,7.9338303,7.8131065,8.039464,7.99042,7.567886,7.201941,7.9451485,8.646856,9.940866,11.559323,12.3289385,9.25425,8.714764,9.2995205,9.725827,8.835487,9.469289,8.99771,8.567632,8.567632,8.605357,7.5792036,6.590776,5.926794,5.624984,5.4778514,5.8702044,5.7381625,5.87775,6.145606,5.462761,5.3156285,4.8138695,3.9348478,3.1463692,3.4029078,4.146115,4.4630156,4.236658,3.7198083,3.5236318,5.2099953,6.043745,6.779407,7.805561,9.125979,8.820397,8.567632,8.397863,8.412953,8.805306,9.58624,9.559832,10.072908,11.197151,11.732863,11.099063,10.382264,9.808825,9.616421,10.054046,9.322156,8.699674,8.29223,7.9753294,7.4018903,7.5716586,7.6886096,7.4735703,7.0812173,7.0812173,7.322665,6.507778,6.0550632,6.587003,7.91874,7.9791017,7.877241,7.5603404,7.322665,7.8131065,7.960239,7.9941926,7.6282477,7.149124,7.432071,8.846806,9.137298,8.918486,8.586494,8.314865,8.473316,8.386545,8.601585,9.446653,11.046246,12.721292,18.184053,20.911661,18.772581,14.022847,16.35433,13.822898,10.038955,7.699928,8.590267,8.114917,7.145352,6.089017,5.4212623,5.6778007,6.043745,5.8513412,5.5570765,5.3948536,5.372218,4.5535583,5.070408,6.4134626,7.726336,7.8131065,8.763808,9.661693,10.137043,10.054046,9.507015,8.967529,9.431562,10.095545,10.303039,9.522105,8.692128,8.337502,8.59404,9.046755,8.729855,9.06939,10.382264,12.113899,12.955194,10.819888,9.695646,8.884532,8.963757,9.789962,10.499215,10.582213,10.419991,10.653893,11.231105,11.41219,12.770335,12.559069,11.283921,10.005001,10.344538,6.1116524,6.8737226,7.3113475,7.84706,8.835487,10.570895,11.378237,11.434827,11.646093,12.185578,12.494934,12.940104,12.438345,11.736636,11.299012,11.272603,12.08749,12.759018,13.347548,13.815352,14.015302,13.9888935,13.9888935,14.000212,13.698401,12.457208,13.185325,12.996693,12.6345215,12.438345,12.3289385,12.377983,12.408164,12.721292,13.298503,13.815352,14.743419,14.811326,14.332202,13.747445,13.619176,13.913441,13.649357,13.751218,14.022847,13.177779,11.389555,10.465261,10.250222,10.502988,10.902886,10.8576145,11.317875,11.77059,11.902632,11.593277,10.9594755,10.646348,10.812344,11.404645,12.181807,13.837989,14.060574,13.788944,13.604086,13.732355,14.992412,14.66042,14.188843,14.2944765,14.973549,13.694629,12.868423,12.415709,12.419481,13.128735,12.570387,12.174261,11.631002,10.93684,10.38981,9.982366,10.291721,10.472807,10.4049,10.672756,10.906659,11.646093,12.279895,12.649611,13.057055,13.792717,14.735873,15.188588,14.849052,13.81158,14.569878,15.16218,15.958203,16.882498,17.41821,18.28214,19.334703,19.481836,18.68204,17.935059,16.965494,17.206944,17.670975,18.229324,19.610106,20.255224,21.160654,20.243906,18.233097,18.678267,18.85558,19.074392,19.164934,19.391293,20.455173,21.085201,21.349285,21.877453,22.862108,24.091984,22.413166,22.01704,21.288923,19.817598,18.406637,18.316093,18.025602,18.0671,18.199142,17.40312,15.882751,16.044973,16.94286,18.278368,20.4099,19.349794,18.293459,18.757492,20.30804,20.564579,19.146072,18.357594,18.617905,19.334703,18.900852,18.53868,17.25976,16.724047,17.546478,19.296976,17.659658,16.21097,15.150862,14.826416,15.777118,16.84477,17.384256,16.91645,15.875206,15.599804,16.029884,15.848798,15.471535,14.943368,13.962485,14.211478,14.539697,15.414946,16.618414,17.225805,15.818617,14.769827,14.464244,14.84528,15.430037,14.928277,13.091009,11.038701,9.424017,8.428044,7.854605,7.405663,6.952948,6.5945487,6.643593,7.4735703,8.028146,8.341274,8.390318,8.118689,8.299775,7.6923823,7.0472636,6.9265394,7.699928,7.2396674,7.250985,7.3000293,7.2396674,7.2283497,7.432071,7.911195,8.492179,9.2844305,10.661438,12.47607,14.305794,15.524352,15.961976,15.916705,15.347038,16.659912,16.708956,14.667966,12.00072,9.144843,8.050782,8.6581745,9.891823,9.695646,8.058327,7.4999785,7.9262853,9.06939,10.469034,10.352083,11.091517,11.091517,10.295494,10.182315,7.326438,5.7683434,5.8211603,6.94163,7.745199,9.167479,9.469289,9.133525,8.4544525,7.5603404,7.6810646,7.4999785,8.013056,8.7600355,7.8319697,7.8319697,7.707473,6.6813188,6.0324273,9.073163,10.106862,9.103344,8.646856,9.193887,9.050528,8.59404,7.4735703,6.9944468,7.4018903,7.8696957,12.525115,17.372938,20.613623,17.980331,2.7389257,2.3428001,1.8146327,4.236658,7.624475,4.957229,15.626213,9.87296,9.899368,15.460217,3.8593953,2.6031113,1.9881734,1.3958713,1.5845025,4.678055,4.2781568,3.2331395,2.4786146,2.5276587,3.4896781,1.2110126,1.8334957,2.8521044,3.350091,3.9876647,4.4705606,6.0324273,8.903395,11.574413,10.819888,9.129752,6.7454534,6.375736,7.3981175,5.8211603,7.2623034,9.027891,7.858378,4.4403796,3.3953626,9.793735,12.113899,13.924759,16.52787,18.964987,17.557796,16.81459,15.467763,13.664448,12.97783,7.0887623,6.7756343,7.6697464,7.164215,4.398881,7.1378064,8.397863,9.333474,9.940866,9.0807085,5.564622,6.9944468,6.0550632,2.1051247,1.1921495,1.750498,1.3958713,1.0450171,1.2751472,2.2862108,3.3463185,2.8030603,2.0108092,1.9844007,3.4142256,3.7688525,3.6254926,4.349837,6.013564,7.394345,7.537705,6.971811,6.7379084,7.3151197,8.643084,9.922004,9.839006,9.899368,10.680302,11.838497,12.423254,12.253486,10.974566,9.993684,12.50248,13.521088,13.936077,13.93985,13.460726,12.174261,13.011784,13.381501,13.204187,12.396846,10.868933,10.544487,10.514306,10.604849,10.823661,11.351829,10.906659,10.061591,10.005001,10.638803,10.559577,10.33322,10.744436,10.789707,10.438853,10.63503,10.446399,11.710228,12.713746,12.943876,13.102326,14.539697,14.649103,14.279386,14.200161,15.098045,18.58395,16.908905,14.083209,12.570387,13.29473,10.661438,8.8618965,7.6131573,6.700182,5.9909286,6.749226,7.073672,6.881268,6.590776,7.115171,8.224322,8.360137,9.061845,10.593531,11.959221,12.31762,11.751727,10.435081,9.2844305,9.940866,9.989911,9.820143,9.869187,10.382264,11.427281,10.412445,9.005256,8.314865,8.477088,8.650629,7.624475,7.9828744,8.333729,8.850578,11.306557,14.830189,12.777881,11.476325,12.540206,12.879742,14.290704,16.060064,15.758255,14.354838,16.192106,7.7414265,9.993684,18.221779,23.835445,14.388792,9.224068,4.115934,5.855114,11.378237,7.7904706,3.4330888,3.4142256,4.266839,3.9688015,1.9278114,1.961765,2.4559789,3.127506,4.168751,6.2851934,7.2057137,9.22784,12.796744,17.886015,23.98635,39.970963,68.084564,67.424355,35.790894,9.688101,7.1000805,6.4549613,7.4094353,8.782671,8.544995,9.208978,11.140562,11.385782,9.756008,8.82417,7.9941926,7.3377557,6.79827,6.4021444,6.273875,4.9232755,4.304565,3.9461658,3.8820312,4.6742826,5.5683947,5.4212623,5.3571277,5.6853456,5.934339,5.5495315,6.1795597,7.1378064,7.854605,7.8810134,7.6923823,7.835742,8.197914,8.107371,6.3153744,5.832478,6.326692,6.7341356,6.903904,7.594294,7.0548086,6.5002327,6.477597,6.881268,6.9680386,6.8397694,6.8435416,6.828451,6.858632,7.194396,8.360137,8.631766,8.371455,8.14887,8.7600355,8.661947,9.318384,9.242931,8.126234,6.858632,6.6813188,6.7454534,6.903904,7.0887623,7.3000293,7.118943,6.964266,7.1264887,7.5075235,7.6282477,8.130007,8.480861,9.125979,9.5032425,8.058327,9.220296,8.778898,8.941121,9.793735,9.322156,9.665465,8.956212,8.062099,7.696155,8.446907,7.8017883,7.1378064,6.617184,6.224831,5.745708,6.3229194,5.8136153,5.142088,4.9345937,5.511805,5.160951,4.5988297,3.7877154,3.1727777,3.682082,3.4330888,3.2784111,3.3538637,3.5387223,3.451952,4.666737,5.8098426,6.6549106,7.424526,8.771353,8.620448,8.646856,8.646856,8.646856,8.903395,9.869187,9.993684,10.1294985,10.748209,11.940358,11.434827,10.834979,9.842778,8.944894,9.431562,9.835234,9.216523,8.20546,7.3377557,7.0472636,6.8058157,6.4549613,6.628502,7.17176,7.141579,6.9454026,6.349328,6.1606965,6.72659,7.91874,8.575176,8.00551,7.3377557,7.1604424,7.5301595,7.6018395,8.167733,8.103599,7.5565677,7.9451485,8.82417,9.899368,9.963503,8.907167,7.7301087,10.242677,10.963248,12.223305,14.4152,15.954432,20.723028,35.36836,40.740578,31.018522,13.679539,9.371201,8.382772,8.186596,7.828197,7.907422,7.5301595,7.250985,6.6586833,5.794752,5.1647234,5.8928404,6.149379,6.009792,5.6061206,5.1043615,4.52715,5.1760416,6.149379,6.900131,7.201941,7.9791017,8.661947,9.446653,9.88805,8.918486,7.9828744,9.009028,10.329447,10.684074,9.22784,8.778898,8.13378,7.9941926,8.265821,8.043237,7.9451485,9.118435,11.027383,12.619431,12.321393,10.336992,9.06939,8.899622,9.616421,10.412445,10.265312,10.20495,10.227587,10.359629,10.668983,11.868678,13.015556,12.81938,11.570641,11.151879,6.8774953,7.284939,8.284684,9.567377,10.884023,12.034674,12.079946,11.310329,11.434827,12.510024,12.958967,12.785426,12.012038,11.151879,10.699164,11.125471,12.3289385,12.845788,13.158916,13.415455,13.430545,13.7851715,13.27964,13.060828,13.170234,12.540206,13.475817,13.309821,13.283413,13.570132,13.29473,12.498707,12.73261,13.63804,14.566105,14.558559,14.618922,14.618922,14.0907545,13.166461,12.577931,12.992921,13.053283,13.057055,13.177779,13.45318,11.917723,11.1631975,11.125471,11.419736,11.363147,11.408418,11.653639,11.947904,12.106354,11.879996,12.064855,11.891314,11.84227,12.004493,12.053536,12.721292,13.4644985,14.0983,14.418973,14.219024,13.977575,13.226823,12.849561,13.060828,13.411682,13.008011,12.875969,13.124963,13.5663595,13.736128,12.411936,11.517824,11.004747,10.770844,10.661438,10.695392,11.355601,11.446144,10.944386,11.019837,10.884023,11.072655,11.083972,10.895341,10.974566,11.348056,12.200669,12.894833,13.234368,13.468271,14.196388,14.667966,14.992412,15.365902,16.063837,16.380737,17.723793,18.304777,18.221779,19.462973,18.61036,18.874443,19.579924,20.258997,20.655123,20.323132,20.474035,19.753464,18.319866,17.84829,17.384256,17.599297,17.546478,16.969267,16.286423,16.45619,16.765545,17.429527,18.376457,19.270569,18.934805,18.62545,18.063328,17.252214,16.471281,16.546734,16.24115,15.920478,15.667711,15.294222,13.966258,14.230342,15.154634,16.18456,17.165443,17.659658,18.414183,18.99894,19.225298,19.123436,18.168962,17.961468,18.406637,18.878216,18.221779,17.897333,16.920223,16.429781,16.999449,18.659403,17.629477,16.592005,15.331948,14.094527,13.5663595,14.169979,14.728328,14.890551,14.611377,14.128481,14.758509,14.818871,14.815099,14.739646,14.083209,14.479335,14.841507,15.890297,17.395575,18.16519,16.927769,16.044973,15.826162,16.086473,16.15438,15.052773,12.860879,10.804798,9.439108,8.631766,7.8131065,7.488661,7.273621,7.0510364,6.971811,7.877241,8.0206,7.699928,7.3679366,7.643338,8.088508,7.7037,7.2887115,7.3075747,7.865923,7.624475,7.8319697,8.047009,8.035691,7.7829256,7.605612,7.9941926,8.692128,9.616421,10.819888,12.083718,13.35132,14.181297,14.6151495,15.181043,14.1926155,14.66042,14.939595,14.366156,13.27964,10.27663,8.926031,8.884532,9.235386,8.469543,6.6662283,6.8850408,7.7376537,8.831716,10.797253,10.725573,11.287694,10.872705,9.616421,9.390063,7.039718,5.7607985,5.8400235,6.8058157,7.4169807,8.684583,8.854351,8.575176,8.243186,7.9941926,8.235641,8.36391,8.590267,8.718536,8.141325,8.171506,8.744945,8.560086,8.356364,10.917976,10.227587,9.159933,8.345046,8.080963,8.329956,6.9265394,6.6058664,7.284939,8.518587,9.469289,13.604086,17.508753,18.772581,14.535924,1.50905,1.388326,1.4713237,4.1612053,7.7942433,6.6020937,9.665465,5.138315,7.6207023,14.320885,5.0666356,2.1994405,2.8181508,2.5125682,1.1921495,3.0935526,2.3503454,1.4147344,0.90920264,1.0110635,1.4449154,1.9730829,3.229367,4.889322,6.3229194,6.609639,8.582722,9.710737,11.25374,12.479843,10.646348,9.940866,8.035691,7.4811153,7.9941926,6.477597,8.75249,9.21275,7.624475,6.149379,9.314611,12.951422,12.928786,12.925014,14.581196,17.516298,32.297443,34.530838,26.87618,15.328176,9.231613,11.925267,9.978593,8.575176,8.552541,6.398372,8.031919,7.594294,6.6813188,6.519096,7.960239,5.149633,6.258785,5.010046,1.2789198,1.0789708,2.323937,1.9466745,1.3015556,1.237421,2.0900342,2.7313805,2.2786655,1.871222,2.1843498,3.4179983,3.99521,4.5309224,5.5382137,7.069899,8.744945,9.4127,9.280658,8.66572,8.235641,8.986393,9.333474,10.080454,10.95193,11.725319,12.272349,12.925014,12.37421,11.506506,11.140562,12.015811,12.057309,13.20796,14.7321005,15.324403,13.075918,12.830698,13.117417,13.057055,12.185578,10.457717,10.536942,10.578441,10.729345,11.140562,11.993175,11.510279,8.816625,8.314865,10.321902,11.083972,11.593277,11.61214,11.068882,10.325675,10.186088,10.469034,11.61214,13.053283,14.2944765,14.93205,15.414946,15.380992,15.773345,16.920223,18.568861,21.175745,18.632996,14.800008,12.276122,12.400619,10.016319,8.499724,7.3717093,6.5568223,6.379509,6.8699503,7.232122,7.4282985,7.3792543,6.964266,7.254758,7.0246277,7.8319697,9.680555,11.031156,10.725573,10.638803,9.922004,9.016574,9.639057,9.416472,9.386291,9.876732,11.00852,12.706201,11.536687,10.084227,9.0807085,8.60913,8.088508,8.778898,8.231868,7.6923823,7.9451485,9.314611,12.083718,11.966766,11.529142,11.876224,12.668475,13.72481,14.426518,14.3095665,15.618668,23.292187,12.37421,8.99771,11.197151,13.675766,7.805561,5.1081343,4.4630156,7.405663,10.770844,6.688864,4.0517993,4.3724723,6.013564,6.6813188,3.399135,1.5279131,1.5203679,2.474842,4.06689,6.598321,8.944894,12.061082,15.999702,21.68505,30.92798,46.05998,71.10266,67.405495,34.244118,8.812852,7.605612,6.6662283,6.7944975,7.7037,7.9941926,8.948667,10.891568,10.978339,9.420244,9.469289,8.827943,7.8810134,7.0284004,6.511551,6.4436436,5.2062225,4.353609,3.6783094,3.380272,4.0895257,5.2250857,5.6778007,5.8626595,5.975838,6.009792,5.692891,6.3417826,7.4094353,8.356364,8.643084,8.069645,7.9036493,7.7904706,7.352846,6.217286,5.5193505,6.330465,6.960493,7.092535,7.756517,7.0510364,6.2889657,6.0022464,6.168242,6.205968,6.730363,6.809588,6.4964604,6.247467,6.911449,7.7942433,8.130007,8.039464,7.865923,8.197914,7.624475,8.778898,9.424017,8.733627,7.2698483,7.1038527,6.8246784,6.6247296,6.6322746,6.9227667,6.6247296,6.571913,6.8963585,7.4169807,7.6622014,8.182823,8.341274,8.099826,8.103599,9.688101,8.386545,8.107371,8.899622,9.9257765,9.461743,9.329701,8.52236,7.6622014,7.3151197,7.986647,7.745199,7.2396674,6.911449,6.7680893,6.3908267,6.5530496,6.1078796,5.413717,4.9345937,5.240176,5.070408,4.436607,3.7084904,3.2482302,3.440634,3.270866,3.180323,3.259548,3.4330888,3.451952,4.2706113,5.3382645,5.987156,6.470052,7.9489207,8.2507305,8.582722,8.518587,8.231868,8.488406,9.639057,10.103089,10.227587,10.416218,11.133017,10.438853,10.216269,9.699419,9.001483,9.110889,9.314611,9.06939,8.60913,7.960239,6.9491754,6.9793563,6.2625575,6.0776987,6.530414,6.560595,6.696409,6.673774,6.8397694,7.2057137,7.435844,8.084735,8.001738,7.6886096,7.5603404,7.937603,8.167733,8.480861,8.82417,9.175024,9.510788,9.552286,11.649866,12.577931,11.400873,9.469289,11.566868,13.517315,16.535416,20.115637,22.050993,38.922173,63.82904,62.493534,36.258698,22.035902,17.399347,11.321648,7.8206515,7.488661,7.5075235,7.2057137,7.115171,6.7454534,5.907931,4.7233267,5.160951,5.836251,5.956975,5.5306683,5.3458095,4.8930945,5.2590394,5.907931,6.417235,6.507778,7.066127,7.5490227,8.367682,9.178797,8.91094,8.495952,9.148616,9.929549,10.170997,9.476834,8.843033,8.16396,8.088508,8.379,7.8923316,7.4207535,7.9489207,9.439108,11.065109,11.23865,9.789962,8.729855,8.446907,9.107117,10.665211,11.000975,10.442626,9.854096,9.733373,10.246449,11.593277,13.0646,13.664448,13.147598,12.038446,7.250985,7.5301595,8.990166,10.963248,12.789199,13.788944,12.593022,11.714001,11.876224,12.755245,12.992921,12.279895,11.400873,10.725573,10.608622,11.408418,12.468526,13.211733,13.754991,14.053028,13.924759,14.019074,13.196642,12.672247,12.770335,12.936331,13.72481,13.830443,14.166207,14.781145,14.867915,14.260523,14.48688,15.033911,15.23386,14.249205,13.936077,13.830443,13.419228,12.766563,12.513797,12.830698,12.759018,12.543978,12.479843,12.932558,11.887542,11.6875925,11.823407,11.876224,11.521597,11.570641,11.672502,11.8045435,11.864905,11.68382,11.808316,11.61214,11.766817,12.257258,12.377983,12.038446,12.434572,13.189097,13.79649,13.626721,12.510024,12.102581,12.015811,12.042219,12.155397,12.630749,12.645839,12.777881,13.091009,13.113645,11.857361,10.748209,10.231359,10.314357,10.521852,10.642575,11.299012,11.529142,11.219787,11.125471,10.804798,10.480352,10.012547,9.525878,9.405154,9.857869,10.861387,12.034674,13.132507,14.045483,14.449154,14.554788,14.649103,14.777372,14.750964,14.354838,15.365902,16.335466,16.98813,18.206688,18.316093,19.074392,19.794964,19.998686,19.398838,18.938578,18.51227,18.052011,17.36162,16.097792,15.282904,15.358356,15.328176,14.735873,13.671993,13.634267,14.177525,15.271586,16.4411,16.791954,17.14658,17.010767,16.407146,15.543215,14.803781,15.030138,14.694374,14.162435,13.736128,13.634267,12.966512,13.200415,13.754991,14.166207,14.109617,15.131999,16.580687,17.452164,17.591751,17.663431,17.20317,17.327667,18.025602,18.859352,18.934805,18.074646,17.229578,16.478827,16.078928,16.475054,16.399601,16.637276,15.973294,14.279386,12.5326605,12.249713,12.045992,12.438345,13.113645,12.913695,13.094781,13.045737,13.091009,13.223051,13.12119,13.875714,14.766054,16.22606,17.727566,17.742655,17.086218,16.244923,16.033657,16.31283,15.973294,13.970031,11.815862,10.325675,9.57115,8.873214,7.937603,7.6697464,7.5490227,7.424526,7.4999785,7.7376537,7.413208,6.8774953,6.5643673,7.001992,7.4584794,7.17176,7.0774446,7.4018903,7.635793,7.6207023,7.8244243,8.171506,8.461998,8.405409,8.254503,8.733627,9.480607,10.231359,10.831206,11.634775,12.449662,12.96274,13.385274,14.43029,13.404137,12.725064,12.90615,13.588995,13.536179,10.891568,9.574923,8.952439,8.511042,7.8696957,6.952948,7.726336,8.790216,9.906913,12.015811,12.2270775,11.974312,10.834979,9.397609,9.261794,7.360391,6.2851934,6.304056,7.069899,7.6093845,8.854351,8.918486,8.899622,9.035437,8.710991,9.06939,9.042982,8.8618965,8.733627,8.83926,8.710991,9.1976595,9.461743,10.001229,12.645839,11.125471,9.22784,7.4396167,6.8473144,9.133525,7.673519,7.567886,7.7716074,8.069645,9.046755,11.966766,12.4307995,11.691365,9.024119,1.7165444,1.2713746,1.8070874,5.2062225,9.016574,6.4210076,4.6290107,3.9574835,7.3113475,11.140562,5.4401255,4.006528,3.9612563,2.8106055,1.0299267,2.0296721,0.8601585,0.814887,1.0940613,1.6071383,3.0030096,5.0553174,6.8133607,8.495952,9.740918,9.593785,11.431054,11.627231,12.061082,12.551523,10.861387,10.672756,9.510788,9.005256,9.046755,7.7829256,9.793735,7.964011,7.24344,9.359882,12.800517,12.279895,11.827179,12.483616,15.271586,21.221016,46.79564,57.177906,44.20762,19.1008,12.442118,20.77962,15.679029,9.684328,7.7225633,7.1000805,6.9454026,5.6853456,4.244203,3.832987,5.956975,3.7462165,4.825187,4.1197066,1.388326,1.2336484,3.218049,2.6483827,1.7580433,1.5845025,1.9806281,2.5993385,2.5427492,2.4333432,2.686109,3.5274043,4.534695,5.674028,6.488915,7.141579,8.401636,9.650374,10.042727,9.457971,8.612903,9.012801,9.2844305,10.612394,12.061082,12.943876,12.811834,13.087236,11.766817,11.068882,11.717773,12.943876,13.109872,14.381247,16.135517,16.746683,13.585222,12.581704,12.604341,12.419481,11.536687,10.231359,10.785934,10.740664,10.785934,11.072655,11.212241,9.87296,7.914967,8.028146,10.0465,10.955703,11.548005,11.8045435,11.672502,11.23865,10.729345,11.329193,12.393073,13.879487,15.448899,16.45619,16.350557,16.071383,16.418465,17.384256,18.168962,19.595015,17.618158,14.188843,11.317875,11.09529,9.318384,8.088508,7.17176,6.647365,6.903904,7.2698483,7.4396167,7.816879,8.07719,7.1906233,6.85486,6.620957,7.2698483,8.575176,9.310839,8.548768,8.707218,8.707218,8.52236,9.175024,8.959985,9.242931,10.035183,11.317875,13.008011,11.827179,10.676529,9.740918,9.031664,8.375228,9.884277,9.175024,8.465771,8.130007,6.6586833,8.235641,10.182315,11.45369,11.91395,12.336484,13.551269,14.056801,13.381501,13.766309,20.183544,13.219278,9.922004,10.310584,11.502733,7.7338815,3.4481792,4.617693,7.7602897,9.012801,4.1272516,3.3953626,5.100589,7.6697464,8.850578,5.7117543,3.0822346,2.5578396,3.3651814,4.9723196,7.0849895,10.744436,15.071637,18.5085,22.07363,29.32084,38.34496,49.88542,45.365814,25.001186,7.816879,7.4811153,6.85486,6.643593,7.066127,7.8734684,8.639311,10.186088,10.555805,9.869187,10.291721,9.416472,8.262049,7.352846,6.888813,6.7643166,5.9192486,4.749735,3.821669,3.5387223,4.112161,5.1798143,6.1116524,6.6624556,6.7567716,6.4738245,6.085244,6.466279,7.303802,8.09228,8.141325,7.8206515,7.745199,7.3377557,6.609639,6.1606965,6.0550632,6.832224,7.326438,7.435844,8.137552,7.4094353,6.590776,6.089017,5.9607477,5.9003854,6.722818,6.9227667,6.4738245,6.058836,7.0585814,7.364164,7.533932,7.413208,7.1604424,7.2698483,6.8699503,7.91874,9.005256,9.156161,7.8508325,7.537705,7.1868505,6.8661776,6.6247296,6.462507,6.138061,6.300284,6.7039547,7.141579,7.4811153,7.964011,8.073418,7.4471617,7.0849895,9.329701,7.4282985,7.7414265,8.831716,9.635284,9.480607,8.967529,8.114917,7.4811153,7.326438,7.6584287,7.6093845,7.1981683,7.092535,7.2924843,7.1302614,6.488915,6.1305156,5.624984,5.1043615,5.2326307,5.292993,4.6554193,3.9386206,3.4481792,3.1727777,3.2670932,3.2029586,3.187868,3.3123648,3.5538127,3.7650797,4.538468,5.2062225,5.8173876,7.1566696,7.5301595,8.024373,8.07719,7.809334,8.024373,8.812852,9.424017,9.767326,9.95973,10.325675,9.831461,9.582467,9.480607,9.371201,9.031664,8.578949,8.397863,8.371455,8.126234,7.039718,7.443389,6.7152724,6.228604,6.296511,6.156924,6.356873,6.9680386,7.5112963,7.6697464,7.3000293,7.6395655,8.001738,8.265821,8.446907,8.695901,9.073163,9.050528,9.325929,9.967276,10.393582,10.446399,12.728837,14.241659,13.985121,12.989148,14.124708,16.086473,19.644058,23.895807,26.265015,45.580856,69.49175,65.48522,42.51371,50.968163,53.59391,29.558517,10.691619,7.1076255,7.2396674,6.930312,6.960493,6.7039547,5.938112,4.8402777,4.6554193,5.342037,5.7607985,5.666483,5.6815734,5.4967146,5.6400743,5.8966126,6.0362,5.80607,6.349328,6.8058157,7.3490734,8.07719,9.046755,9.246704,9.420244,9.476834,9.416472,9.348565,8.733627,8.2507305,8.480861,8.967529,8.216777,7.5037513,7.5527954,8.597813,10.023865,10.355856,9.782416,8.7751255,8.209232,8.582722,10.020092,11.25374,10.974566,9.846551,8.914713,9.6051035,11.427281,12.755245,13.822898,14.339747,13.45318,6.930312,7.598067,9.363655,11.876224,14.403882,15.811071,13.234368,12.623203,12.67602,12.672247,12.487389,11.993175,11.23865,10.725573,10.827434,11.819634,12.585477,13.743673,14.803781,15.422491,15.396083,14.754736,13.758763,12.898605,12.600568,13.215506,14.151116,14.84528,15.335721,15.712983,16.105335,16.452417,16.109108,15.441354,14.551015,13.302276,13.619176,13.411682,13.181552,13.230596,13.6682205,13.72481,13.321139,12.762791,12.189351,11.578186,11.00852,11.370691,11.536687,11.204697,10.880251,10.880251,11.057564,11.193378,11.189606,11.080199,10.627484,10.521852,11.23865,12.581704,13.694629,12.985375,12.0724,11.646093,11.766817,11.864905,11.136789,11.46878,11.732863,11.631002,11.729091,12.106354,11.763044,11.291467,11.091517,11.378237,11.080199,10.20495,9.593785,9.559832,9.880505,9.665465,10.0465,10.589758,10.989656,11.042474,10.967021,10.54826,10.144588,9.846551,9.457971,10.197406,11.491416,13.091009,14.524607,15.082954,14.93205,14.807553,15.045229,15.165953,13.902123,13.158916,13.302276,14.128481,15.045229,15.101818,15.920478,16.999449,17.67852,17.655886,16.984358,17.301258,17.040947,16.467508,15.588487,14.169979,13.7700815,13.815352,13.728582,13.494679,13.622949,13.634267,14.347293,15.848798,17.342756,17.150352,16.822134,16.731592,16.022339,14.784918,14.04171,14.252977,13.736128,13.091009,12.664702,12.536433,12.0233555,11.978085,12.185578,12.359119,12.140307,12.510024,13.43809,14.634012,15.826162,16.77309,16.65614,16.803272,17.674747,19.15739,20.575897,19.229069,18.157644,16.920223,15.516807,14.388792,14.652876,15.811071,15.7657995,14.102073,12.08749,11.295239,10.495442,10.661438,11.642321,12.178034,11.785681,11.6008215,11.517824,11.544232,11.815862,12.728837,14.169979,16.029884,17.4333,16.77309,16.82968,16.022339,15.79598,16.135517,15.569623,12.974057,11.012292,10.091772,9.846551,9.125979,8.171506,7.7301087,7.4282985,7.273621,7.6584287,6.964266,6.4436436,6.2625575,6.417235,6.7152724,6.9227667,6.515323,6.56814,7.1302614,7.213259,7.405663,7.4169807,7.6584287,8.137552,8.469543,8.83926,9.57115,10.321902,10.748209,10.502988,10.876478,11.578186,12.287439,12.909923,13.600313,12.691111,11.785681,12.00072,12.97783,12.894833,10.559577,9.846551,9.073163,8.013056,7.914967,8.035691,8.929804,10.087999,11.378237,13.011784,13.102326,11.936585,10.529396,9.601331,9.593785,7.84706,6.8171334,6.8171334,7.5301595,8.043237,9.480607,9.718282,10.008774,10.340765,9.461743,9.673011,9.133525,8.816625,9.122208,9.861642,9.35611,8.858124,8.933576,10.114408,12.917468,11.657412,8.771353,6.270103,6.228604,10.797253,9.771099,9.676784,8.443134,6.6586833,7.5565677,9.759781,7.254758,5.523123,5.2137675,2.1466236,1.5241405,2.0108092,5.9418845,9.525878,2.8294687,3.8405323,5.994701,8.296002,8.526133,3.2331395,5.8966126,4.255521,1.8900851,1.0638802,2.6898816,1.3317367,1.9768555,3.2935016,5.0439997,8.084735,9.42779,11.106608,12.468526,13.068373,12.687338,13.060828,12.370438,12.37421,13.000465,12.359119,11.710228,11.046246,10.861387,10.736891,9.318384,9.763554,5.9192486,6.598321,11.529142,11.3669195,8.695901,10.227587,13.12119,17.316349,25.555761,49.115807,66.91882,53.020473,20.145817,19.666695,28.256962,19.1008,8.82417,4.8629136,5.455216,4.1536603,3.5236318,3.3350005,3.5538127,4.327201,2.4823873,3.9348478,4.085753,2.142851,1.1280149,3.9310753,3.4066803,2.41448,2.123988,2.003264,2.7728794,3.2935016,3.4557245,3.4783602,3.8895764,5.243949,6.349328,6.549277,6.224831,6.7869525,8.14887,8.737399,8.820397,8.797762,9.201432,9.774872,10.612394,11.962994,13.347548,13.577678,13.996439,11.944131,10.914205,12.083718,14.302021,14.800008,15.807299,16.490145,15.920478,13.057055,12.543978,12.332711,11.962994,11.272603,10.397354,11.034928,10.861387,10.834979,10.665211,8.809079,6.7944975,7.707473,8.790216,9.265567,10.33322,10.287949,11.314102,12.272349,12.58925,12.279895,12.796744,13.951167,15.414946,16.90136,18.199142,17.263533,16.056292,15.482853,15.30554,14.124708,15.079182,14.9358225,12.936331,10.352083,10.49167,9.318384,8.224322,7.4584794,7.1793056,7.435844,7.884786,7.7942433,8.145098,8.805306,8.548768,8.088508,7.7376537,7.533932,7.4999785,7.635793,7.1340337,7.2660756,7.594294,8.028146,8.850578,8.646856,8.843033,9.590013,10.789707,12.140307,11.302785,10.597303,10.076681,9.684328,9.246704,9.80128,9.35611,9.559832,9.612649,6.2814207,7.6810646,9.601331,11.6875925,13.332457,13.645585,14.283158,15.23386,13.962485,11.117926,10.525623,9.442881,11.09529,15.743164,19.289433,13.275867,5.8098426,4.402653,5.7419353,6.300284,2.354118,1.81086,4.063117,7.069899,8.820397,7.3188925,4.881777,4.112161,4.6214657,5.881522,7.2283497,11.449917,17.493662,20.368402,19.859098,20.519308,23.1941,20.432537,17.052265,13.804035,7.3679366,6.828451,6.63982,6.6624556,6.9454026,7.7640624,8.194141,9.371201,10.412445,10.891568,10.868933,9.390063,8.3525915,7.6622014,7.2358947,6.9982195,6.587003,5.138315,4.187614,4.2706113,4.908185,5.560849,6.3945994,7.1302614,7.5075235,7.273621,6.8661776,6.820906,7.118943,7.3415284,6.670001,6.771862,7.1981683,7.1378064,6.530414,6.0512905,6.7944975,7.432071,7.7150183,7.8810134,8.654402,7.9941926,7.2170315,6.6813188,6.477597,6.4021444,6.8171334,6.8850408,6.4549613,6.1229706,7.254758,7.1264887,7.0170827,6.647365,6.1795597,6.228604,6.507778,6.8473144,7.8206515,8.835487,8.111144,7.6508837,7.5188417,7.3415284,6.8925858,6.0814714,5.726845,6.0022464,6.4021444,6.7643166,7.2698483,7.5716586,7.567886,7.0849895,6.3417826,5.9494295,6.9755836,7.9489207,8.627994,9.050528,9.552286,8.873214,7.9828744,7.54525,7.6395655,7.756517,7.756517,7.4169807,7.4018903,7.7225633,7.7150183,6.3455553,5.881522,5.481624,5.13077,5.6513925,5.726845,5.1647234,4.466788,3.8443048,3.2029586,3.2935016,3.048281,2.9237845,3.127506,3.6292653,3.270866,3.6669915,4.5120597,5.5382137,6.519096,6.688864,7.118943,7.4018903,7.484888,7.647111,7.7829256,8.243186,8.763808,9.26934,9.869187,10.012547,9.590013,9.58624,9.854096,9.099571,8.231868,7.677292,7.413208,7.3453007,7.3000293,7.745199,7.273621,6.8699503,6.7680893,6.4474163,6.273875,7.201941,7.8961043,7.956466,7.8961043,8.054554,8.326183,8.820397,9.276885,9.06939,9.484379,9.5032425,9.522105,9.80128,10.47658,11.227332,12.875969,14.400109,15.456445,16.376965,16.905132,18.025602,21.209698,25.751938,28.811537,38.348732,49.9156,49.677925,48.840405,83.63532,94.20622,50.15705,14.120935,6.832224,7.1906233,6.790725,6.964266,6.7039547,5.9003854,5.3458095,4.5799665,4.8553686,5.4438977,5.824933,5.6778007,5.9003854,6.0701537,6.115425,5.975838,5.5985756,6.145606,6.6058664,6.7077274,6.983129,8.75249,9.439108,9.563604,9.34102,8.986393,8.692128,8.533678,8.390318,8.865668,9.5032425,8.76758,8.114917,8.024373,8.703445,9.812597,10.469034,10.495442,9.242931,8.246958,8.099826,8.465771,10.525623,11.608367,10.536942,8.461998,8.858124,10.850069,11.830952,13.162688,14.781145,15.169725,6.270103,7.6018395,10.069136,13.487134,16.70141,17.591751,14.286931,12.268577,11.125471,10.695392,11.046246,12.623203,12.657157,11.91395,11.442371,12.58925,13.88326,14.600059,15.116908,15.531898,15.641303,15.373446,14.524607,13.690856,13.385274,14.068119,14.750964,15.754482,16.214743,15.848798,14.969776,15.675257,14.894323,14.037937,13.777626,14.022847,14.475562,14.230342,13.932304,13.936077,14.32843,14.460471,14.385019,13.200415,11.348056,10.589758,10.076681,10.352083,10.193633,9.525878,9.416472,9.416472,9.57115,9.563604,9.495697,9.87296,10.789707,11.921495,13.034419,14.075664,15.196134,13.20796,11.849815,11.080199,10.729345,10.499215,10.314357,10.725573,11.332966,11.581959,10.789707,10.18986,9.940866,9.944639,9.986138,9.703192,10.374719,10.782163,10.70671,10.382264,10.469034,9.880505,9.955957,10.3634,10.899114,11.457462,11.763044,11.695138,11.763044,12.0082655,12.0082655,12.14408,13.026875,14.396337,15.629986,15.777118,14.581196,15.067864,16.052519,16.35433,14.815099,13.694629,13.521088,13.7851715,14.11339,14.298248,14.369928,15.396083,16.263786,16.376965,15.656394,16.252468,15.845025,15.00373,14.120935,13.411682,13.864397,14.252977,14.245432,14.147344,14.894323,14.173752,15.128226,16.35433,16.84477,15.992157,14.830189,14.102073,13.95494,14.249205,14.543469,14.724555,13.377728,11.921495,11.121698,11.11038,10.533169,10.529396,10.834979,11.065109,10.710483,11.091517,12.264804,13.290957,14.196388,15.992157,16.637276,16.682549,17.225805,18.485863,19.806282,18.68204,17.659658,16.31283,14.890551,14.32843,13.449409,13.275867,13.196642,12.66093,11.185833,10.63503,10.167224,9.989911,10.197406,10.774617,10.725573,10.831206,11.038701,11.242422,11.291467,11.498961,12.393073,13.72481,15.196134,16.478827,17.40689,18.104828,18.41041,17.7917,15.350811,12.860879,11.065109,10.133271,9.771099,9.246704,8.345046,7.5792036,7.0359454,6.8171334,7.0510364,6.696409,6.405917,6.296511,6.4247804,6.790725,6.7039547,6.462507,6.579458,6.934085,6.7756343,7.152897,7.164215,7.194396,7.443389,7.91874,9.092027,10.080454,10.831206,11.016065,10.038955,10.529396,11.246195,12.196897,13.087236,13.306048,12.525115,11.725319,11.59705,12.038446,12.162943,10.744436,10.740664,10.1294985,8.771353,8.394091,9.088254,10.352083,11.393328,11.876224,11.902632,10.827434,9.899368,9.748463,10.144588,10.008774,8.937348,7.356619,7.0774446,7.9715567,7.9941926,9.510788,10.382264,10.7557535,10.70671,10.253995,9.80128,9.110889,8.922258,9.559832,10.925522,9.510788,8.001738,8.001738,9.26934,9.718282,9.1825695,6.511551,4.7421894,5.621211,9.612649,10.148361,10.431308,8.98262,7.0057645,8.360137,10.827434,9.175024,7.696155,6.6020937,1.9994912,0.6073926,0.16976812,0.10186087,0.38858038,1.5731846,5.5004873,5.6325293,4.5233774,3.4142256,2.2447119,3.953711,2.3465726,0.88279426,1.0902886,2.5804756,2.003264,4.617693,7.9262853,10.623712,12.58925,13.7851715,13.807808,14.290704,15.324403,15.471535,16.41092,15.354584,14.317112,13.762536,12.604341,12.336484,11.812089,11.627231,11.480098,10.163452,7.4999785,4.52715,5.621211,9.144843,7.462252,6.937857,7.564113,9.989911,14.056801,18.829172,25.446356,32.89729,26.280106,11.231105,13.917213,25.427492,13.245687,2.8747404,2.293756,1.9542197,3.0030096,3.0256453,2.776652,2.6182017,2.5314314,2.837014,3.399135,3.218049,2.093807,0.6413463,3.5236318,3.9763467,3.4557245,2.9086938,2.7615614,2.7011995,3.1048703,3.7047176,4.2404304,4.485651,5.462761,6.4210076,6.462507,5.8966126,6.224831,6.541732,7.2094865,8.160188,9.016574,9.0807085,9.6051035,9.661693,10.182315,11.54046,13.5663595,15.467763,13.875714,13.075918,14.351066,15.961976,15.181043,14.490653,13.373956,12.325166,12.864652,13.083464,12.204442,11.672502,11.631002,10.910432,10.921749,10.906659,11.193378,10.453944,5.7079816,6.2323766,7.6622014,7.3453007,6.428553,9.857869,9.7220545,10.823661,11.747954,12.132762,12.694883,14.0983,16.078928,17.96524,19.417702,20.432537,17.72002,15.350811,14.196388,13.70972,11.902632,13.743673,15.082954,13.502225,10.310584,10.529396,9.699419,8.959985,8.186596,7.5075235,7.322665,7.960239,8.29223,9.42779,11.355601,12.955194,12.174261,10.714255,9.110889,7.9300575,7.7829256,8.209232,8.473316,8.635539,8.91094,9.64283,8.473316,8.186596,8.461998,9.454198,11.812089,11.3820095,11.249968,10.819888,10.087999,9.612649,10.186088,8.2507305,8.533678,10.868933,10.223814,8.635539,9.303293,11.272603,13.43809,14.509516,12.5326605,12.030901,11.09529,10.646348,14.418973,7.643338,9.22784,14.867915,19.270569,16.143063,11.774363,5.1873593,1.9844007,3.1954134,5.292993,2.8785129,2.2296214,4.1612053,7.111398,7.111398,4.1574326,3.5387223,4.349837,5.613666,6.2851934,9.484379,16.950403,19.994913,16.478827,10.804798,9.035437,7.997965,7.752744,7.964011,7.9036493,7.111398,6.25124,5.7419353,5.8966126,6.9567204,8.179051,9.261794,10.257768,10.797253,10.103089,8.4544525,7.865923,7.4471617,6.9491754,6.790725,6.741681,5.2628117,4.255521,4.5535583,5.9192486,6.0550632,6.043745,6.3342376,6.907676,7.2623034,7.2623034,7.6923823,8.114917,8.024373,6.8661776,6.3531003,6.571913,6.934085,6.809588,5.5382137,5.6853456,6.590776,7.250985,7.5792036,8.424272,8.043237,7.1981683,6.730363,6.85486,7.17176,7.001992,6.9680386,6.802043,6.6662283,7.1566696,6.6058664,6.790725,6.6020937,6.119198,6.6058664,6.888813,6.3908267,6.7680893,7.7829256,7.2924843,6.85486,6.72659,6.7944975,6.8133607,6.4247804,5.715527,5.9418845,6.307829,6.609639,7.232122,7.33021,6.7680893,6.2625575,5.9494295,5.3873086,7.643338,8.246958,8.43559,8.903395,9.797507,9.137298,8.186596,7.8319697,8.160188,8.4544525,8.695901,8.401636,8.039464,7.8734684,7.9338303,6.6020937,5.8513412,5.4288073,5.4212623,6.224831,5.9192486,5.458988,5.0062733,4.508287,3.6783094,3.4934506,3.108643,2.8294687,2.8709676,3.3727267,3.2859564,3.3312278,3.8895764,4.8968673,5.798525,6.349328,6.5228686,6.6058664,6.7944975,7.17176,7.4018903,7.6282477,7.865923,8.329956,9.431562,10.038955,10.47658,10.70671,10.453944,9.186342,8.661947,7.7150183,6.7077274,6.360646,7.752744,7.643338,7.2585306,7.164215,7.435844,7.643338,7.364164,7.816879,8.024373,8.07719,9.14107,9.835234,9.495697,9.208978,9.020347,7.9338303,8.337502,8.967529,9.703192,10.465261,11.246195,11.917723,13.211733,14.48688,15.486626,16.343012,16.18456,18.029375,22.413166,28.321096,33.217964,34.315796,34.327114,35.71167,45.32809,74.4188,78.54605,40.310497,10.989656,6.541732,7.6886096,7.164215,7.2623034,6.7379084,5.66271,5.43258,4.52715,4.3309736,4.6856003,5.13077,4.8968673,5.3609,5.7607985,6.360646,6.94163,6.820906,6.771862,6.7944975,6.6247296,6.530414,7.322665,8.75249,9.495697,9.714509,9.352338,8.118689,8.5563135,8.7600355,9.061845,9.367428,9.110889,9.073163,8.880759,8.880759,9.333474,10.4049,10.540714,9.303293,8.073418,7.4509344,7.232122,9.367428,12.136535,12.276122,9.95973,8.7751255,9.359882,9.74469,11.3820095,14.132254,16.28265,7.5301595,9.258021,12.396846,15.30554,16.271332,13.479589,11.559323,10.589758,10.642575,11.314102,11.766817,12.219532,12.049765,11.84227,12.068627,13.087236,14.196388,14.905642,15.0905,15.045229,15.456445,15.267814,14.988639,14.800008,14.667966,14.373701,14.694374,15.00373,14.886778,14.48688,14.456699,15.154634,14.754736,14.456699,14.558559,14.460471,14.279386,13.951167,13.841762,14.003984,14.181297,14.366156,13.736128,12.67602,11.695138,11.457462,10.834979,10.016319,9.333474,9.156161,9.865415,10.208723,10.295494,10.336992,10.359629,10.201178,11.216014,11.710228,12.543978,13.592768,13.70972,12.67602,12.332711,11.91395,11.046246,9.7296,9.34102,9.835234,10.789707,11.5857315,11.385782,11.16697,10.770844,10.540714,10.582213,10.77839,11.227332,11.751727,12.279895,12.479843,11.785681,11.649866,11.593277,11.876224,12.393073,12.679792,13.230596,12.955194,12.883514,13.177779,13.166461,12.883514,13.060828,13.287186,13.645585,14.739646,14.196388,14.709465,15.682802,16.392056,15.988385,14.739646,13.788944,13.445636,13.36641,12.562841,12.423254,13.158916,13.773854,14.045483,14.558559,14.920732,14.803781,14.381247,13.81158,13.230596,13.826671,13.140053,12.540206,12.6345215,13.234368,12.766563,13.58145,13.909668,13.381501,13.026875,13.389046,13.407909,13.253232,13.011784,12.66093,12.826925,11.781908,10.386037,9.435335,9.654147,9.22784,9.163706,9.333474,9.525878,9.454198,9.688101,10.808571,12.034674,12.96274,13.573905,15.599804,17.267305,17.923742,17.723793,17.644567,16.59955,16.109108,15.316857,14.1926155,13.521088,13.4644985,13.106099,12.777881,12.204442,10.502988,9.386291,9.273112,9.654147,10.269085,11.125471,11.615912,11.891314,12.193124,12.396846,12.034674,11.940358,12.540206,13.460726,14.547242,15.8676605,16.746683,18.795218,19.372429,17.554024,14.166207,12.0082655,11.197151,10.914205,10.612394,10.0276375,8.880759,8.088508,7.5037513,7.1604424,7.2924843,7.0170827,6.33801,5.9720654,6.058836,6.1418333,6.488915,6.405917,6.541732,6.903904,6.8737226,7.1038527,7.33021,7.699928,8.288457,9.065618,10.325675,11.2650585,11.932813,12.004493,10.770844,10.050273,10.201178,11.012292,12.140307,13.109872,12.875969,11.736636,10.714255,10.125726,9.574923,8.099826,7.7640624,8.13378,8.718536,8.952439,11.034928,11.883769,11.680047,10.989656,10.77839,10.506761,10.137043,10.993429,12.506252,12.208215,11.317875,8.967529,7.7150183,8.031919,8.299775,9.129752,9.812597,10.340765,10.589758,10.314357,10.167224,9.374973,9.0807085,9.578695,10.340765,7.7338815,7.333983,8.737399,10.77839,11.502733,7.9262853,6.5266414,7.001992,8.311093,8.661947,9.793735,10.106862,9.156161,8.107371,9.718282,6.741681,5.240176,4.5950575,4.168751,3.2670932,1.0374719,0.38858038,0.30935526,1.6033657,6.8699503,3.7499893,5.96452,7.1340337,4.908185,0.9620194,2.6597006,2.2975287,2.293756,3.3727267,4.568649,7.303802,10.393582,11.876224,12.528888,15.871433,16.033657,16.26756,16.33924,16.4826,17.399347,16.7995,16.222288,15.354584,14.0983,12.566614,12.883514,11.92904,11.638548,12.1252165,11.676274,5.9682927,3.7348988,5.379763,7.7829256,4.3121104,5.485397,8.054554,11.3820095,15.803526,22.639523,19.67424,14.694374,9.303293,5.6325293,6.3342376,6.0211096,3.7009451,1.9768555,1.5316857,1.1091517,2.5917933,2.5993385,3.7198083,5.330719,3.5953116,2.6031113,3.1312788,3.3425457,2.5276587,1.1053791,3.712263,3.99521,3.2029586,2.4823873,2.8822856,3.1048703,3.2746384,3.7235808,4.4630156,5.2062225,4.9345937,5.0439997,5.194905,5.50426,6.5568223,6.688864,7.3075747,7.828197,8.0206,8.00551,9.446653,9.963503,10.050273,10.257768,11.174516,13.185325,12.759018,13.381501,15.16218,14.849052,13.649357,12.913695,12.064855,11.3820095,12.0082655,11.98563,12.67602,13.264549,13.196642,12.193124,11.080199,10.725573,10.672756,10.31813,8.929804,6.1531515,7.405663,8.503497,8.412953,9.246704,10.499215,11.7555,12.577931,13.008011,13.600313,15.569623,18.029375,20.040184,21.175745,21.503962,20.202406,17.53139,15.143317,13.641812,12.585477,14.037937,14.958458,13.562587,10.631257,9.5032425,9.982366,9.25425,8.379,7.6810646,6.7756343,7.194396,8.431817,10.495442,12.54775,12.917468,10.838752,9.669238,9.133525,8.959985,8.880759,8.710991,8.956212,9.310839,9.454198,9.031664,8.458225,8.254503,7.9828744,8.167733,10.310584,11.514051,12.789199,12.951422,11.864905,10.442626,10.891568,9.420244,8.262049,8.944894,12.321393,10.431308,8.36391,7.4509344,8.167733,10.140816,11.102836,11.921495,13.86817,15.943113,14.871688,11.717773,8.314865,7.2887115,8.480861,8.929804,6.1720147,3.832987,3.874486,6.3455553,9.371201,3.9159849,3.3274553,6.126743,9.133525,7.4509344,4.22534,6.1229706,7.6131573,7.0057645,6.4436436,8.14887,13.35132,15.445127,12.630749,7.911195,7.1264887,8.963757,8.68081,6.2889657,6.549277,6.8774953,6.790725,6.590776,6.3719635,6.017337,7.6886096,8.963757,9.884277,10.238904,9.563604,8.82417,8.394091,7.647111,6.771862,6.730363,6.7869525,6.0701537,5.311856,5.0138187,5.43258,5.6363015,5.975838,6.2889657,6.673774,7.496206,7.9036493,8.29223,8.209232,7.707473,7.33021,6.700182,6.405917,6.2436943,5.8966126,4.927048,5.6815734,6.349328,6.930312,7.3981175,7.7037,7.605612,6.9265394,6.8359966,7.4584794,7.9036493,7.5188417,7.3415284,7.001992,6.5832305,6.643593,6.5530496,6.8133607,6.832224,6.537959,6.4134626,5.5495315,5.9682927,6.7454534,7.2358947,7.0510364,6.7567716,6.439871,6.48137,6.7114997,6.398372,5.692891,5.5306683,5.9192486,6.515323,6.609639,6.5228686,6.1418333,5.904158,5.873977,5.753253,7.326438,8.107371,9.073163,10.170997,10.310584,9.442881,8.793989,9.039209,9.827688,9.759781,8.843033,7.6697464,7.020855,7.0472636,7.273621,6.6850915,6.1041074,5.832478,5.987156,6.470052,6.115425,5.745708,5.379763,4.9760923,4.4101987,3.259548,3.0822346,2.9954643,2.7087448,2.516341,3.0558262,3.380272,3.8292143,4.496969,5.2250857,6.066381,6.224831,6.156924,6.255012,6.8774953,7.062354,7.066127,7.2472124,7.858378,9.076936,9.922004,10.861387,11.46878,11.193378,9.35611,8.186596,7.2698483,6.530414,6.436098,7.9941926,7.6810646,7.4282985,7.2283497,7.111398,7.145352,8.329956,9.261794,9.371201,8.933576,9.0807085,9.737145,9.635284,9.612649,9.654147,8.899622,9.397609,9.952185,10.408672,10.887795,11.808316,12.340257,12.845788,13.853079,15.158407,15.818617,17.025856,19.97605,23.673222,26.944088,28.422956,28.60027,26.578144,25.933023,29.57738,39.763466,35.16841,18.776354,7.8432875,6.8737226,7.643338,8.22055,8.360137,7.352846,5.802297,5.6287565,4.7836885,4.6290107,4.7346444,4.9949555,5.643847,5.802297,5.726845,6.0739264,6.858632,7.432071,7.364164,6.94163,6.741681,6.911449,7.1793056,8.273367,9.378746,9.857869,9.42779,8.167733,8.66572,9.005256,9.1825695,9.220296,9.159933,8.790216,9.076936,9.235386,9.510788,11.200924,11.947904,10.469034,8.654402,7.564113,7.3905725,8.4544525,10.910432,12.113899,11.551778,10.834979,10.0276375,10.397354,11.555551,13.109872,14.683057,8.401636,10.7218,12.015811,12.853333,13.087236,11.838497,10.329447,10.091772,11.302785,12.955194,12.853333,12.781653,12.581704,12.762791,13.219278,13.241914,14.324657,15.007503,15.256495,15.350811,15.905387,15.433809,15.086727,14.871688,14.471789,13.2607765,13.615403,14.000212,13.951167,13.4644985,12.974057,13.917213,14.777372,15.309312,15.343266,14.7736,14.366156,14.007756,13.645585,13.381501,13.494679,13.5663595,12.89106,11.902632,11.234878,11.717773,12.0082655,11.378237,10.495442,9.88805,9.933322,10.457717,10.812344,11.068882,11.219787,11.18206,11.317875,11.729091,12.566614,13.177779,12.091263,10.974566,10.582213,10.26154,9.733373,9.06939,8.7751255,9.616421,10.834979,11.781908,11.891314,11.574413,10.982111,10.751981,11.042474,11.514051,13.238141,13.622949,13.268322,12.777881,12.728837,12.83447,13.12119,13.717264,14.392565,14.558559,13.396591,12.717519,12.51757,12.879742,13.9888935,13.751218,13.570132,13.400364,13.502225,14.4152,14.403882,14.667966,14.886778,14.875461,14.577423,13.890805,12.725064,11.646093,11.02361,11.004747,11.563096,12.411936,13.223051,13.702174,13.604086,14.064346,13.837989,13.377728,12.955194,12.672247,12.683565,11.861133,11.423509,11.634775,11.793225,11.887542,11.898859,11.974312,12.155397,12.393073,11.710228,11.476325,11.5857315,11.7555,11.506506,11.415963,10.570895,9.488152,8.612903,8.322411,7.9753294,7.911195,8.137552,8.586494,9.122208,9.250477,10.220041,11.16697,11.796998,12.385528,13.879487,15.743164,16.444872,16.03743,16.143063,15.588487,15.39231,14.7321005,13.536179,12.498707,12.540206,12.276122,12.15917,11.864905,10.310584,9.156161,9.035437,9.291975,9.669238,10.280403,10.801025,11.321648,12.049765,12.804289,13.000465,13.585222,13.70972,14.268067,15.460217,16.795727,16.961721,18.87067,18.802763,16.143063,13.36641,12.030901,11.732863,11.332966,10.514306,9.793735,8.612903,7.665974,7.224577,7.0774446,6.511551,6.043745,5.6778007,5.50426,5.409944,5.0854983,5.726845,5.9796104,6.2625575,6.598321,6.6134114,7.0585814,7.605612,8.262049,8.993938,9.748463,10.925522,11.732863,11.978085,11.634775,10.846297,9.865415,9.616421,10.023865,10.729345,11.076427,11.09529,10.684074,9.439108,7.956466,7.835742,6.5228686,6.760544,7.541477,8.409182,9.461743,10.914205,11.393328,11.09529,10.514306,10.453944,11.0613365,11.774363,12.649611,13.20796,12.453435,12.166716,10.065364,8.6581745,8.756263,9.465516,8.778898,9.639057,10.280403,10.167224,10.008774,10.178542,9.771099,9.574923,9.661693,9.386291,6.1003346,6.515323,9.110889,11.664956,11.25374,7.466025,7.3075747,8.639311,9.382519,7.5263867,8.213005,8.412953,8.016829,7.4094353,7.466025,4.6931453,3.482133,3.078462,3.0331905,3.2105038,1.690136,3.500996,4.9723196,7.567886,17.852062,6.4134626,4.9232755,4.6818275,2.5238862,0.814887,2.5540671,3.7952607,5.617439,7.665974,8.122461,11.299012,12.147853,12.261031,13.238141,16.682549,15.69412,15.192361,14.460471,14.117163,16.097792,16.018566,16.090246,15.30554,13.822898,12.970284,13.023102,12.423254,12.362892,11.902632,7.9451485,4.82896,4.738417,5.9720654,6.439871,3.6707642,5.8928404,9.582467,12.755245,15.973294,22.326395,20.594759,10.484125,3.6443558,2.9954643,2.7540162,1.3317367,4.4630156,5.111907,3.0030096,4.5988297,4.5950575,3.5802212,5.462761,9.159933,8.59404,3.9725742,2.6521554,3.5123138,4.1574326,0.90920264,3.199186,3.651901,3.1350515,2.463524,2.4031622,3.6896272,4.0593443,4.255521,4.636556,5.168496,5.458988,5.485397,5.523123,5.9003854,6.9944468,6.692637,6.590776,6.752999,7.1604424,7.7187905,8.76758,9.695646,10.212496,10.601076,11.717773,11.634775,12.027128,13.521088,15.313085,15.158407,14.094527,14.124708,13.562587,12.543978,13.030646,11.32542,12.706201,14.015302,13.9888935,13.234368,11.808316,11.140562,10.770844,10.514306,10.450171,8.677037,9.473062,10.33322,10.325675,10.084227,11.242422,11.853588,12.223305,12.709973,13.72481,15.939341,17.689838,19.278114,20.711712,21.719002,21.073883,19.17248,17.139036,15.641303,14.898096,13.675766,13.109872,11.98563,10.257768,9.073163,9.87296,9.22784,8.473316,7.9526935,7.0510364,7.4169807,9.216523,10.552032,10.842525,10.819888,10.121953,10.20495,10.612394,10.967021,10.985884,9.74469,9.510788,9.748463,9.854096,9.137298,8.080963,7.665974,7.3000293,7.405663,9.420244,10.95193,12.955194,13.777626,12.947649,11.200924,10.457717,9.590013,9.220296,9.476834,9.989911,11.042474,9.774872,8.843033,9.608876,12.14408,16.350557,17.938831,18.395319,19.168707,21.677504,13.298503,9.393836,10.11818,12.551523,10.676529,4.696918,7.533932,13.158916,16.263786,12.294985,4.06689,4.957229,7.4735703,7.6584287,5.0741806,3.9159849,6.6624556,7.7225633,6.0550632,5.13077,5.5306683,9.424017,13.8870325,16.203424,13.860624,8.688355,8.224322,7.5112963,5.292993,4.032936,6.537959,7.141579,6.8963585,6.549277,6.5530496,7.6320205,8.83926,9.669238,9.740918,8.797762,8.812852,8.703445,8.27714,7.647111,7.254758,6.79827,6.221059,5.7419353,5.492942,5.5306683,5.3458095,5.4665337,6.043745,6.9793563,7.9300575,8.13378,8.560086,8.122461,6.9944468,6.5756855,6.0286546,5.783434,5.2552667,4.5196047,4.3083377,5.6061206,5.8664317,6.2889657,7.001992,7.066127,7.201941,6.7643166,6.9491754,7.828197,8.333729,7.8734684,7.273621,6.760544,6.541732,6.79827,6.6850915,6.4247804,6.217286,6.1003346,5.9607477,5.2137675,5.7117543,6.1795597,6.228604,6.330465,6.820906,6.647365,6.560595,6.688864,6.511551,6.017337,5.4438977,5.455216,5.9682927,6.1418333,5.753253,5.4363527,5.323174,5.5382137,6.1908774,7.039718,8.171506,9.710737,10.978339,10.49167,9.922004,9.759781,10.336992,11.031156,10.27663,8.499724,8.726082,8.390318,7.2283497,7.284939,7.1076255,6.911449,6.439871,6.006019,6.466279,5.938112,5.402399,5.0477724,4.889322,4.7836885,3.62172,3.2029586,2.9954643,2.7351532,2.4522061,2.9049213,3.308592,3.8443048,4.534695,5.247721,5.7570257,5.873977,5.945657,6.2021956,6.722818,6.651138,6.5756855,6.790725,7.492433,8.76758,9.74469,10.627484,11.046246,10.714255,9.408927,7.9036493,6.903904,6.470052,6.628502,7.3792543,7.194396,7.17176,7.0284004,6.9755836,7.696155,9.159933,9.669238,9.612649,9.439108,9.669238,10.133271,10.336992,10.325675,9.854096,8.397863,9.137298,9.9257765,10.495442,10.93684,11.717773,12.2119875,12.283667,12.894833,14.007756,14.551015,16.048746,17.701157,19.010258,19.579924,19.112118,18.71222,16.444872,15.245177,16.509007,20.085455,17.139036,11.438599,7.466025,6.590776,7.069899,8.175279,8.179051,7.2358947,5.8966126,5.100589,4.6856003,4.6516466,4.745962,4.961002,5.5268955,5.406172,5.3986263,5.6589375,6.1342883,6.549277,6.9944468,6.930312,7.2396674,7.858378,7.7829256,7.888559,9.148616,9.827688,9.495697,9.039209,8.386545,8.66572,9.148616,9.491924,9.7296,9.159933,9.540969,9.95973,10.284176,11.170743,12.521342,11.925267,9.74469,7.405663,7.394345,8.09228,9.473062,10.7557535,11.442371,11.344283,10.484125,10.510533,11.000975,12.012038,14.109617,9.046755,11.442371,11.151879,10.751981,11.117926,11.434827,10.702937,10.978339,12.396846,13.9888935,13.671993,13.400364,13.117417,13.343775,13.928532,14.030393,15.218769,15.554533,15.46399,15.377219,15.724301,15.554533,15.452672,15.060319,14.068119,12.215759,12.857106,13.075918,13.215506,13.189097,12.449662,13.098554,14.226569,14.856597,14.671739,14.022847,13.860624,13.841762,13.487134,12.898605,12.781653,12.445889,11.962994,11.314102,10.759526,10.834979,11.487643,11.563096,11.219787,10.661438,10.159679,11.027383,11.321648,11.480098,11.631002,11.589504,10.906659,11.476325,12.3289385,12.491161,11.004747,9.88805,9.431562,9.220296,9.092027,9.159933,9.193887,10.057818,11.0613365,11.77059,12.0082655,12.196897,12.0233555,12.264804,12.996693,13.588995,14.864142,14.6302395,13.898351,13.434318,13.747445,13.234368,13.287186,13.928532,14.781145,15.0905,13.441863,13.117417,13.313594,13.739901,14.600059,14.11339,13.800262,13.687083,13.679539,13.585222,13.622949,13.502225,13.155144,12.736382,12.626976,12.883514,12.276122,11.3971,10.751981,10.759526,11.446144,12.106354,12.826925,13.336229,13.000465,13.396591,13.140053,12.868423,12.721292,12.340257,12.268577,12.019584,11.7555,11.551778,11.400873,11.306557,10.985884,11.212241,11.989402,12.5326605,11.751727,11.133017,11.072655,11.314102,10.974566,10.93684,10.087999,9.125979,8.303548,7.435844,6.937857,6.9567204,7.2962565,7.9300575,8.98262,9.167479,10.023865,10.7557535,11.170743,11.646093,12.291212,13.690856,14.354838,14.237886,14.728328,14.743419,14.690601,14.102073,12.992921,11.849815,11.6008215,11.514051,11.653639,11.574413,10.291721,9.22784,8.952439,8.918486,8.963757,9.303293,9.639057,10.133271,10.891568,11.7894535,12.494934,13.513543,13.837989,14.758509,16.422237,17.829426,17.527617,18.395319,17.550251,14.901869,13.12119,12.438345,12.091263,11.423509,10.427535,9.763554,8.650629,7.779153,7.2660756,6.8359966,5.828706,5.413717,5.406172,5.3609,5.0968165,4.6931453,5.3194013,5.6891184,5.994701,6.258785,6.3644185,7.032173,7.665974,8.179051,8.688355,9.533423,10.646348,11.465008,11.642321,11.295239,11.034928,10.072908,9.552286,9.548513,9.820143,9.786189,9.163706,9.359882,8.918486,7.7716074,7.250985,6.255012,6.647365,7.643338,8.793989,9.989911,10.895341,11.083972,11.072655,11.133017,11.32542,11.4838705,12.064855,12.453435,12.291212,11.465008,11.759273,10.453944,9.450426,9.597558,10.691619,9.6201935,10.091772,10.197406,9.608876,9.582467,9.81637,9.544742,9.49947,9.371201,7.854605,5.27413,6.511551,9.012801,10.725573,10.103089,7.492433,8.073418,8.726082,8.080963,6.560595,6.6020937,6.911449,7.0812173,6.587003,4.8025517,3.127506,2.1579416,1.8900851,3.9084394,11.3820095,4.8629136,5.243949,6.4210076,9.231613,21.4436,8.386545,5.5985756,4.2102494,1.780679,2.2786655,4.7535076,5.983383,8.461998,11.544232,11.449917,13.502225,12.804289,12.543978,13.766309,15.365902,14.592513,14.007756,13.038192,12.362892,13.894578,13.558814,14.04171,13.943622,13.068373,12.396846,11.864905,11.649866,11.442371,9.80128,4.172523,4.644101,5.243949,6.228604,6.643593,4.323428,7.594294,12.091263,14.260523,14.4152,16.761772,17.025856,8.7751255,2.9615107,2.7087448,3.3048196,2.5729303,5.836251,6.258785,4.1008434,6.741681,6.247467,4.538468,6.375736,10.782163,11.072655,5.66271,2.848332,3.059599,3.99521,0.59230214,3.1463692,3.92353,3.4783602,2.546522,2.052308,3.92353,4.7308717,4.8440504,4.768598,5.1345425,5.7570257,6.270103,6.417235,6.48137,7.281166,7.0812173,6.436098,6.273875,6.832224,7.6622014,8.194141,9.250477,10.054046,10.736891,12.359119,11.774363,12.717519,14.381247,15.845025,16.086473,15.958203,15.905387,15.260268,14.283158,14.173752,11.608367,12.898605,14.079436,13.766309,13.124963,12.257258,12.1101265,11.879996,11.431054,11.314102,10.917976,11.2650585,11.69891,11.898859,11.9064045,12.15917,12.294985,12.321393,12.400619,12.845788,14.852824,15.845025,16.965494,18.663176,20.68153,19.953413,18.58395,17.629477,17.346529,17.150352,14.260523,12.623203,11.415963,10.238904,9.122208,9.574923,9.0957985,8.601585,8.356364,7.9941926,8.284684,9.763554,10.238904,9.544742,9.540969,10.023865,11.076427,12.053536,12.649611,12.902377,11.227332,10.585986,10.427535,10.212496,9.397609,7.54525,7.0472636,6.94163,7.0585814,8.016829,9.759781,12.355347,13.86817,13.717264,12.706201,11.106608,10.3634,10.416218,10.291721,8.137552,10.850069,11.415963,11.370691,11.864905,13.675766,19.595015,24.21648,24.17498,21.047476,21.349285,17.984104,16.678776,18.99894,21.802,17.237123,7.7414265,10.819888,18.440592,22.213217,13.381501,4.327201,5.59103,6.937857,5.251494,4.5309224,4.930821,7.194396,8.329956,7.956466,8.262049,8.431817,8.963757,12.083718,16.690092,18.35382,9.797507,6.4021444,6.4021444,7.001992,4.402653,5.3986263,5.4250345,5.3609,5.5759397,5.9230213,7.914967,9.001483,9.42779,9.352338,8.854351,8.710991,8.420499,8.243186,8.099826,7.5716586,6.9944468,6.466279,5.9796104,5.6551647,5.7607985,5.643847,5.4967146,6.1041074,7.3377557,8.167733,7.884786,8.254503,7.9225125,6.858632,6.387054,5.7796617,5.4476705,5.010046,4.5120597,4.4177437,5.6061206,5.4891696,5.696664,6.3644185,6.1078796,6.6624556,6.651138,7.118943,8.065872,8.469543,8.031919,7.1981683,6.541732,6.387054,6.8171334,6.63982,6.1418333,5.7079816,5.534441,5.617439,4.979865,5.2326307,5.481624,5.485397,5.6325293,6.832224,6.964266,6.8850408,6.760544,6.066381,6.224831,5.4665337,5.0553174,5.3759904,5.9418845,5.8136153,5.66271,5.4288073,5.353355,5.983383,6.598321,8.197914,10.035183,11.227332,10.767072,10.657665,10.533169,11.00852,11.61214,10.77839,8.684583,7.9941926,8.039464,8.031919,7.0849895,7.152897,7.586749,7.3792543,6.670001,6.7341356,5.9494295,5.1647234,4.7044635,4.6327834,4.772371,3.9650288,3.4934506,3.180323,2.9124665,2.6408374,2.8822856,3.1463692,3.663219,4.436607,5.2326307,5.349582,5.704209,6.096562,6.4247804,6.6813188,6.356873,6.2625575,6.3908267,6.8699503,7.9753294,9.156161,10.012547,10.1294985,9.601331,9.031664,7.937603,6.673774,6.3229194,6.7944975,6.828451,7.1038527,7.039718,6.7152724,6.7077274,8.111144,9.1976595,9.556059,9.491924,9.378746,9.669238,9.774872,9.895596,9.87296,9.408927,8.050782,8.582722,9.14107,9.669238,10.201178,10.887795,11.114153,11.144334,11.649866,12.536433,12.96274,13.951167,14.377474,14.019074,13.034419,11.944131,10.929295,9.416472,8.624221,9.012801,10.310584,10.469034,9.073163,7.541477,6.7567716,7.0812173,7.91874,7.7301087,7.145352,6.296511,4.8365054,4.538468,4.5309224,4.6856003,4.8553686,4.9119577,4.715781,5.138315,5.59103,5.8400235,5.9796104,6.700182,6.8850408,7.466025,8.265821,7.9791017,8.062099,9.258021,9.710737,9.454198,10.423763,8.99771,8.986393,9.510788,9.971047,10.076681,9.839006,9.978593,10.291721,10.627484,10.899114,12.098808,12.393073,10.921749,8.643084,8.3525915,8.812852,9.261794,9.993684,10.782163,10.899114,10.336992,10.023865,9.88805,10.469034,12.936331,9.688101,11.581959,10.948157,10.533169,11.11038,11.491416,11.895086,12.472299,13.27964,13.951167,13.705947,13.430545,13.185325,13.313594,13.93985,14.992412,16.116653,15.961976,15.339493,14.852824,14.894323,15.611122,16.03743,15.441354,13.856852,12.095036,12.770335,12.555296,12.796744,13.45318,13.091009,13.083464,13.287186,13.268322,12.936331,12.540206,12.796744,13.249459,13.272095,12.777881,12.2119875,11.378237,10.985884,10.7218,10.321902,9.540969,9.831461,10.374719,10.808571,10.970794,10.884023,11.944131,11.853588,11.548005,11.344283,10.93684,10.114408,10.751981,11.480098,11.551778,10.853842,10.1294985,9.767326,9.631512,9.691874,10.023865,10.231359,10.653893,11.1631975,11.664956,12.098808,13.50977,14.162435,14.939595,15.935568,16.448645,15.882751,14.996184,14.626467,14.792462,14.7170105,13.441863,12.887287,13.098554,13.788944,14.335975,13.777626,14.279386,14.939595,15.154634,14.622695,13.902123,13.694629,13.687083,13.422999,12.298758,12.2119875,11.868678,11.514051,11.3669195,11.619685,12.468526,12.54775,12.4307995,12.193124,11.434827,11.657412,11.861133,12.15917,12.479843,12.577931,12.808062,12.687338,12.81938,13.057055,12.498707,12.925014,13.275867,12.96274,12.147853,11.744182,10.914205,10.933067,11.449917,12.064855,12.336484,12.853333,12.279895,11.7555,11.506506,10.853842,11.136789,10.148361,8.99771,8.047009,6.907676,6.126743,6.228604,6.6549106,7.2962565,8.503497,8.91094,9.627739,10.284176,10.665211,10.729345,11.00852,11.853588,12.453435,12.668475,13.034419,13.460726,13.562587,13.189097,12.449662,11.714001,11.216014,11.208468,11.404645,11.329193,10.310584,9.329701,8.8618965,8.66572,8.6581745,8.907167,9.092027,9.26934,9.540969,9.97482,10.612394,11.589504,12.687338,14.403882,16.463736,17.84829,17.482344,17.20317,16.033657,14.1926155,13.098554,12.728837,12.181807,11.517824,10.853842,10.336992,9.371201,8.563859,7.665974,6.677546,5.881522,5.613666,5.560849,5.409944,5.1458607,5.05909,5.4778514,5.7306175,5.945657,6.1720147,6.4134626,7.0548086,7.4773426,7.5603404,7.673519,8.6732645,9.661693,10.597303,11.133017,11.302785,11.502733,10.653893,9.971047,9.616421,9.544742,9.510788,8.111144,8.431817,9.167479,9.295748,8.084735,7.001992,6.8473144,7.8734684,9.488152,10.238904,11.23865,11.419736,11.706455,12.31762,12.740154,11.581959,11.065109,10.899114,10.797253,10.480352,11.034928,10.691619,10.231359,10.287949,11.363147,11.336739,11.091517,10.336992,9.473062,9.616421,9.748463,9.039209,8.778898,8.495952,5.945657,5.6098933,7.6508837,8.963757,8.835487,8.948667,7.937603,8.239413,7.303802,5.379763,5.515578,5.247721,5.9984736,6.398372,5.5457587,3.0143273,1.5958204,0.8262049,0.7922512,4.8100967,19.440336,7.6810646,4.1612053,3.5689032,5.73439,15.629986,7.5112963,7.0585814,6.1606965,3.5877664,4.961002,8.141325,8.145098,10.386037,14.260523,13.132507,14.302021,13.694629,13.573905,14.139798,13.521088,14.022847,13.917213,13.109872,12.076173,11.891314,10.314357,10.9594755,11.77059,11.691365,10.646348,9.793735,9.631512,8.695901,6.258785,2.3163917,4.7950063,4.779916,5.8136153,7.375482,4.859141,8.318638,13.505998,15.558306,13.404137,9.786189,9.578695,6.56814,4.29702,4.217795,5.6853456,4.13857,4.9232755,5.5759397,5.621211,6.541732,6.4926877,5.1458607,6.224831,9.559832,11.091517,7.5112963,4.0178456,2.474842,2.293756,0.4376245,3.4972234,4.485651,3.9650288,2.7804246,2.0485353,3.7273536,4.9987283,5.2175403,4.878004,5.6325293,5.8702044,6.971811,7.3113475,6.851087,7.1302614,7.5112963,6.952948,6.696409,7.0963078,7.6093845,8.024373,8.786444,9.4013815,10.106862,11.887542,12.96274,14.320885,15.735619,16.731592,16.580687,17.565342,16.7995,15.961976,15.596032,15.101818,12.864652,13.20796,13.441863,12.713746,12.019584,12.076173,12.943876,13.189097,12.521342,11.808316,11.823407,11.91395,12.257258,12.860879,13.562587,13.045737,13.12119,13.192869,12.940104,12.291212,13.430545,13.981348,14.811326,16.286423,18.263277,17.372938,16.542961,16.950403,18.248188,18.587723,16.233604,14.5132885,12.713746,10.774617,9.303293,9.397609,9.129752,8.907167,8.899622,9.06939,9.295748,9.914458,9.986138,9.5032425,9.4013815,9.865415,11.16697,12.261031,12.868423,13.456953,12.162943,11.2801485,10.61994,9.95973,9.046755,6.8737226,6.4511886,6.670001,6.7944975,6.439871,8.526133,11.472552,13.415455,14.0983,14.883006,13.219278,12.181807,11.785681,11.23865,8.975075,11.249968,13.177779,14.652876,15.584714,15.912932,23.129965,39.186256,44.864056,34.87792,17.852062,26.080156,27.253443,27.90988,28.773811,24.752193,17.53516,15.041456,17.674747,20.29295,12.200669,4.8742313,5.1798143,5.172269,3.5349495,5.5797124,6.0286546,7.424526,9.778644,12.626976,15.033911,15.222542,11.996947,9.899368,11.234878,16.056292,8.356364,5.541986,8.511042,13.000465,9.590013,4.9760923,3.7801702,4.395108,5.2099953,4.6252384,7.9036493,8.967529,9.046755,8.990166,9.25425,8.533678,7.8017883,7.5603404,7.6810646,7.4169807,7.194396,6.771862,6.1305156,5.613666,5.9305663,6.19465,6.0701537,6.4964604,7.4811153,8.122461,7.541477,7.61693,7.537705,7.1793056,7.1076255,6.356873,5.772116,5.715527,5.8890676,5.3269467,5.873977,5.723072,5.828706,6.092789,5.3458095,6.270103,6.7114997,7.3679366,8.156415,8.22055,7.9791017,7.33021,6.617184,6.2097406,6.507778,6.387054,6.1078796,5.6061206,5.1760416,5.4665337,4.606375,4.5837393,4.9119577,5.2250857,5.281675,6.670001,7.175533,7.333983,7.0170827,5.413717,6.066381,5.409944,4.821415,4.9760923,5.828706,6.439871,6.541732,6.1531515,5.594803,5.5004873,6.2927384,8.231868,10.042727,11.019837,11.012292,11.321648,10.899114,11.016065,11.574413,11.125471,9.084481,6.043745,6.56814,9.265567,6.7944975,7.032173,7.809334,8.265821,8.084735,7.4811153,6.304056,5.3759904,4.7836885,4.515832,4.4630156,4.0216184,3.832987,3.6443558,3.3350005,2.9464202,3.029418,3.059599,3.3764994,4.006528,4.67051,4.727099,5.564622,6.319147,6.643593,6.722818,6.307829,6.1305156,6.039973,6.1531515,6.8737226,8.171506,9.175024,9.171251,8.45068,8.296002,8.054554,6.6058664,6.0739264,6.6624556,6.6549106,7.394345,7.1604424,6.6020937,6.5568223,8.07719,8.458225,9.156161,9.393836,9.137298,9.122208,8.714764,8.488406,8.480861,8.514814,8.216777,8.348819,8.326183,8.533678,9.042982,9.590013,9.408927,9.740918,10.438853,11.133017,11.204697,11.544232,11.800771,11.295239,10.174769,9.431562,7.7225633,6.9680386,6.8699503,7.0548086,7.069899,7.9036493,7.752744,7.492433,7.466025,7.4999785,7.6508837,7.33021,7.069899,6.651138,5.1043615,4.402653,4.304565,4.508287,4.647874,4.2706113,4.0970707,4.8742313,5.6891184,6.1229706,6.2436943,6.802043,6.8850408,7.356619,8.009283,7.5792036,8.575176,9.567377,9.623966,9.514561,11.732863,10.555805,10.220041,10.34831,10.502988,10.201178,10.49167,10.352083,10.352083,10.646348,10.978339,11.246195,11.8045435,11.744182,10.997202,10.34831,10.408672,10.299266,10.167224,10.099318,10.163452,9.880505,9.623966,9.148616,9.046755,10.744436,10.604849,12.0082655,11.442371,10.638803,10.612394,11.6875925,12.238396,12.815607,13.381501,13.547497,12.559069,12.498707,13.004238,13.441863,13.70972,14.237886,14.5283785,14.445381,14.286931,14.2944765,14.649103,15.894069,16.131744,15.026365,13.377728,13.106099,12.728837,12.770335,13.102326,13.445636,13.396591,13.505998,13.04951,12.642066,12.393073,11.917723,12.1252165,12.396846,12.664702,12.600568,11.61214,10.7218,9.903141,9.329701,9.224068,9.857869,10.295494,10.287949,10.336992,10.868933,12.238396,12.370438,12.268577,11.491416,10.265312,9.461743,9.397609,9.650374,10.084227,10.729345,11.778135,11.34051,10.506761,10.091772,10.367173,11.0613365,10.574668,10.4049,10.948157,12.08749,13.200415,15.663939,16.463736,16.82968,17.21826,17.30503,17.399347,16.931541,16.150608,15.365902,14.939595,14.852824,14.747191,14.366156,13.981348,14.418973,14.079436,14.339747,14.071891,13.29473,13.185325,13.622949,13.853079,13.551269,12.762791,11.872451,12.457208,12.540206,12.551523,12.608112,12.498707,12.400619,11.7894535,11.197151,10.933067,11.091517,11.714001,11.962994,12.128989,12.189351,11.812089,12.370438,12.245941,12.294985,12.721292,13.060828,13.475817,13.332457,13.041965,12.54775,11.351829,10.729345,11.042474,11.664956,11.936585,11.155652,11.729091,11.879996,11.6008215,11.09529,10.804798,11.0613365,10.035183,8.601585,7.273621,6.224831,5.3948536,5.4250345,5.8664317,6.5040054,7.3717093,8.028146,8.314865,8.605357,8.971302,9.156161,9.57115,10.140816,10.770844,11.1782875,10.910432,11.434827,11.932813,11.944131,11.627231,11.747954,11.615912,11.434827,11.363147,11.204697,10.419991,9.665465,8.952439,8.801534,9.163706,9.446653,9.725827,9.58624,9.378746,9.273112,9.246704,10.453944,11.846043,13.513543,15.150862,16.052519,15.403628,14.886778,14.237886,13.392818,12.449662,12.415709,12.396846,12.261031,11.872451,11.091517,10.419991,8.816625,7.435844,6.809588,6.820906,5.96452,5.247721,4.9119577,4.98741,5.2779026,5.7079816,5.9796104,6.2851934,6.6549106,6.971811,7.1566696,7.303802,7.326438,7.4282985,8.088508,8.586494,9.397609,10.182315,10.891568,11.793225,11.465008,10.751981,9.97482,9.193887,8.194141,8.024373,8.446907,9.06939,9.74469,10.574668,7.9489207,7.273621,7.8017883,8.786444,9.507015,10.310584,11.106608,11.766817,12.325166,12.985375,11.970539,11.646093,11.204697,10.748209,11.261286,11.589504,12.095036,11.740409,10.838752,11.046246,12.121444,12.272349,11.570641,10.714255,11.031156,11.363147,9.65792,8.186596,7.066127,4.274384,7.1906233,9.639057,10.121953,8.98262,8.424272,8.99771,7.3905725,5.372218,3.9763467,3.5236318,3.561358,4.908185,4.561104,2.4522061,1.4637785,0.7205714,0.35839936,0.55080324,1.0299267,1.1317875,2.1051247,1.6071383,1.9127209,4.38379,9.476834,4.5950575,4.353609,4.3649273,4.2404304,7.598067,9.382519,9.680555,12.909923,16.74291,12.128989,14.962231,14.562332,13.592768,13.396591,14.007756,14.7170105,13.894578,12.355347,10.831206,9.963503,8.571404,9.533423,10.005001,9.26934,8.744945,8.473316,8.050782,6.156924,3.1576872,1.0827434,3.4745877,4.696918,5.2326307,5.0666356,3.663219,4.06689,9.714509,15.83748,17.621931,10.238904,10.653893,9.374973,8.062099,7.0170827,5.172269,3.5990841,5.6023483,9.435335,11.766817,7.6886096,6.017337,6.187105,6.187105,7.5263867,15.226315,10.480352,5.885295,3.3840446,2.5276587,0.48666862,2.9803739,3.7009451,3.8405323,3.572676,2.0598533,3.4745877,5.0213637,5.300538,5.010046,6.9265394,7.183078,8.209232,8.103599,6.8359966,6.224831,6.7756343,7.01331,7.3188925,7.673519,7.6584287,8.209232,8.246958,8.533678,9.397609,10.725573,12.925014,14.754736,16.26756,16.874952,15.335721,16.105335,16.11288,15.912932,16.018566,16.920223,14.664193,12.936331,11.9064045,11.446144,11.155652,11.385782,12.268577,12.706201,12.321393,11.427281,12.196897,12.306303,12.483616,12.902377,13.185325,13.27964,13.230596,13.849306,14.867915,14.954685,14.245432,14.298248,14.939595,15.456445,14.603831,14.784918,16.343012,18.312323,19.685556,19.395065,18.844261,17.708702,14.93205,11.219787,9.046755,9.756008,9.65792,9.537196,9.57115,9.337247,9.789962,10.212496,9.982366,9.0957985,8.179051,8.314865,9.49947,10.340765,10.661438,11.506506,10.650121,9.318384,8.356364,7.835742,7.0812173,5.8966126,5.342037,5.4891696,6.0739264,6.5002327,8.379,10.661438,12.2270775,13.551269,16.739138,15.347038,14.320885,14.203933,14.173752,12.038446,14.675511,16.97304,22.020813,27.974014,28.060785,40.269,85.61218,108.30452,86.56288,32.621887,32.59925,31.071339,29.181253,28.219234,29.64906,38.14124,28.400322,18.153872,13.434318,8.575176,5.0477724,5.1534057,4.776143,3.2105038,3.1727777,3.0407357,4.727099,9.092027,14.7170105,17.927513,15.841252,14.769827,10.291721,4.617693,6.609639,4.093298,9.092027,17.980331,24.423975,19.391293,9.005256,8.367682,10.095545,9.839006,6.2851934,6.40969,7.665974,8.507269,8.439363,8.009283,8.009283,7.752744,7.322665,6.9567204,7.066127,6.820906,6.319147,5.96452,5.915476,6.089017,5.8928404,6.221059,6.779407,7.4018903,8.024373,7.9526935,7.3490734,6.779407,6.741681,7.643338,7.118943,6.749226,6.730363,6.8435416,6.439871,6.6850915,7.2396674,7.654656,7.4697976,6.224831,6.7379084,7.232122,7.726336,7.964011,7.4169807,7.707473,7.635793,7.0548086,6.3229194,6.2851934,6.224831,6.1003346,5.5759397,4.9760923,5.292993,4.5120597,4.244203,4.5422406,5.1345425,5.4174895,6.307829,7.24344,7.8432875,7.6093845,5.9494295,5.5004873,5.093044,4.825187,4.8402777,5.342037,6.2927384,6.5040054,6.458734,6.379509,6.19465,6.8925858,8.582722,10.050273,10.691619,10.559577,11.144334,10.982111,10.967021,11.065109,10.284176,8.039464,7.605612,9.318384,10.921749,7.5527954,7.907422,7.6207023,8.194141,9.265567,8.605357,6.7643166,5.9984736,5.455216,4.768598,4.0593443,3.85185,3.9725742,4.217795,4.2517486,3.6179473,3.3463185,3.3727267,3.4444065,3.4029078,3.1576872,3.7198083,4.9119577,5.926794,6.477597,6.820906,6.6020937,6.0701537,5.832478,6.0286546,6.349328,7.1793056,8.171506,8.379,7.858378,7.673519,7.6395655,6.696409,5.915476,5.8513412,6.5455046,7.1076255,7.220804,7.1793056,7.3453007,8.16396,7.6282477,8.416726,9.325929,9.684328,9.352338,8.29223,8.182823,8.065872,7.7904706,8.009283,8.60913,8.66572,8.59404,8.552541,8.4544525,8.246958,9.035437,9.876732,10.069136,9.14107,9.774872,10.427535,10.427535,9.929549,9.918231,7.7338815,6.537959,6.6360474,7.6810646,8.68081,8.937348,8.854351,8.477088,7.816879,6.8661776,6.8774953,6.587003,6.2399216,5.8966126,5.43258,4.1272516,3.9273026,4.2027044,4.432834,4.2102494,3.7235808,4.123479,5.1232247,6.19465,6.560595,6.903904,6.971811,7.4207535,7.967784,7.3717093,8.503497,9.318384,9.688101,10.182315,12.098808,11.917723,11.59705,11.261286,10.997202,10.850069,10.774617,10.838752,11.133017,11.589504,11.993175,11.223559,11.299012,11.774363,12.264804,12.434572,11.947904,11.219787,10.152134,9.295748,9.857869,10.103089,10.740664,10.469034,9.25425,8.314865,9.846551,10.657665,11.291467,10.974566,10.529396,12.396846,12.838243,13.777626,13.909668,13.238141,13.057055,13.65313,14.162435,14.498198,14.675511,14.811326,14.056801,13.573905,13.151371,12.925014,13.36641,14.151116,14.607604,14.320885,13.615403,13.521088,13.8870325,14.320885,14.928277,15.448899,15.264041,14.769827,13.521088,12.404391,11.710228,11.136789,12.14408,12.81938,13.041965,12.759018,12.015811,10.480352,9.857869,9.827688,9.971047,9.797507,9.582467,10.038955,10.767072,11.4838705,12.030901,11.32542,11.004747,10.56335,10.084227,10.20495,10.103089,10.220041,10.570895,11.140562,11.876224,11.7026825,11.000975,10.593531,10.7557535,11.197151,11.031156,11.068882,11.849815,13.234368,14.381247,15.539442,15.90916,15.743164,15.62244,16.459963,16.550507,16.65614,16.45619,15.8676605,15.049001,15.596032,15.207452,14.743419,14.479335,14.079436,13.864397,13.694629,13.460726,13.287186,13.551269,13.920986,13.728582,13.128735,12.619431,13.057055,13.057055,12.879742,12.521342,12.068627,11.7026825,11.98563,11.389555,11.249968,11.763044,12.019584,12.185578,12.506252,12.411936,11.962994,11.846043,11.898859,11.751727,11.619685,11.653639,11.925267,12.117672,11.864905,11.491416,11.193378,11.0613365,10.544487,10.993429,11.449917,11.506506,11.314102,11.016065,10.86516,10.676529,10.472807,10.472807,10.408672,9.484379,8.179051,6.9982195,6.507778,5.9117036,5.8664317,6.047518,6.2927384,6.6020937,7.250985,8.0206,8.318638,8.243186,8.59404,9.058073,9.405154,9.869187,10.227587,9.8239155,9.654147,9.759781,9.797507,9.639057,9.367428,9.480607,9.805053,10.253995,10.502988,10.005001,9.386291,8.726082,8.303548,8.401636,9.2995205,10.11818,10.367173,10.265312,10.016319,9.797507,10.819888,12.136535,13.189097,13.622949,13.257004,12.845788,12.536433,12.340257,12.283667,12.438345,12.713746,12.611885,12.46098,12.019584,10.506761,9.650374,7.91874,6.930312,6.964266,6.9680386,5.987156,5.3458095,5.036454,5.0439997,5.3759904,5.5797124,5.832478,6.1229706,6.4474163,6.8133607,6.9189944,7.3188925,7.586749,7.7225633,8.14887,8.578949,9.446653,10.653893,11.955449,12.955194,12.664702,11.46878,10.340765,9.374973,7.779153,7.8508325,8.578949,9.42779,9.6201935,8.145098,6.8699503,6.5002327,6.9567204,7.91874,8.82417,10.076681,10.906659,11.227332,11.155652,10.982111,11.249968,11.374464,11.212241,11.068882,11.6875925,12.494934,13.551269,13.81158,13.306048,13.12119,13.377728,13.283413,12.37421,10.740664,9.065618,9.737145,8.786444,7.141579,5.624984,4.9685473,7.454707,8.620448,8.873214,8.631766,8.314865,8.98262,6.428553,3.7198083,2.1503963,1.2298758,1.1317875,2.252257,2.7615614,2.052308,0.7205714,0.482896,0.30181,0.5281675,1.2185578,2.1164427,4.8327327,5.304311,6.94163,8.956212,6.3644185,3.9122121,3.0633714,4.2291126,6.9680386,9.989911,10.502988,11.144334,12.725064,14.053028,11.947904,15.728074,14.064346,12.804289,13.483362,13.324911,12.868423,12.147853,10.834979,9.386291,9.035437,8.993938,9.382519,8.963757,8.035691,8.439363,8.09228,5.9796104,3.4179983,1.4260522,0.72811663,2.8785129,5.20245,7.1264887,7.986647,7.043491,3.2557755,3.199186,4.696918,6.537959,8.469543,8.816625,7.484888,8.786444,11.000975,6.356873,4.7044635,6.983129,12.283667,16.863634,14.136025,11.00852,9.031664,7.3981175,8.314865,17.022083,12.057309,7.0548086,4.1989317,3.0407357,0.47535074,2.4295704,3.7650797,4.0291634,3.3010468,2.2183034,3.1463692,4.2592936,5.0251365,5.4891696,6.2927384,6.3531003,7.375482,7.598067,6.7567716,6.066381,6.439871,7.2585306,8.616675,9.771099,9.125979,8.14887,8.130007,8.4544525,9.065618,10.446399,12.468526,14.136025,15.803526,16.848543,15.701665,16.060064,14.649103,15.373446,18.444365,20.353312,16.678776,14.177525,12.694883,11.7894535,10.763299,10.684074,11.053791,11.45369,11.7555,12.1252165,13.332457,13.604086,13.487134,13.283413,13.038192,12.811834,12.830698,13.521088,14.547242,14.807553,13.641812,13.841762,14.520834,14.966003,14.637785,15.07541,16.697638,18.044466,18.463226,18.101055,17.980331,16.776863,14.268067,11.136789,8.963757,9.046755,8.703445,8.533678,8.669493,8.790216,9.691874,10.167224,10.125726,9.812597,9.812597,9.529651,10.038955,10.242677,10.072908,10.518079,9.0957985,7.7904706,6.911449,6.375736,5.7381625,4.991183,4.8138695,5.062863,5.4174895,5.3646727,7.5565677,9.250477,10.672756,12.355347,15.150862,16.278877,15.094273,14.947141,15.939341,14.894323,17.953922,20.756983,27.559025,36.70387,40.65758,55.502857,95.892586,117.53613,97.348816,33.466957,27.404348,23.171463,20.904116,21.021067,24.227798,30.780848,25.872662,16.335466,8.3525915,7.4396167,3.3274553,3.8065786,4.2328854,3.270866,2.8822856,3.1576872,6.398372,7.937603,7.1000805,7.175533,10.702937,11.321648,8.296002,4.06689,4.2517486,2.6936543,8.880759,17.957695,24.537153,22.703657,12.604341,11.419736,13.272095,13.513543,8.703445,7.33021,7.673519,8.141325,8.058327,7.6697464,7.8244243,7.828197,7.496206,7.043491,7.0774446,7.224577,6.5568223,6.0512905,6.009792,6.0626082,5.8890676,5.7079816,5.8890676,6.3644185,6.647365,6.8359966,6.511551,6.198423,6.2135134,6.670001,6.368191,6.3116016,6.4738245,6.952948,7.9753294,7.567886,7.5565677,7.91874,8.126234,7.152897,6.749226,7.1604424,7.541477,7.4018903,6.609639,6.8246784,7.001992,6.9491754,6.6586833,6.3116016,5.994701,5.9230213,5.6815734,5.221313,4.8553686,5.138315,5.172269,5.0138187,5.05909,6.0512905,6.1720147,6.549277,6.828451,6.7379084,6.085244,5.4967146,5.304311,5.402399,5.4891696,5.070408,6.149379,6.5455046,6.349328,5.9532022,6.0739264,7.326438,8.914713,9.933322,10.11818,9.876732,10.344538,10.552032,10.570895,10.186088,8.903395,7.4697976,7.9413757,8.963757,9.495697,8.809079,8.578949,8.182823,8.465771,9.163706,8.873214,8.103599,7.032173,5.8966126,4.8930945,4.146115,3.9763467,4.085753,4.466788,4.878004,4.847823,4.247976,3.742444,3.4745877,3.3161373,2.867195,3.651901,4.90064,5.8890676,6.48137,7.1264887,6.9755836,6.3342376,5.9796104,6.149379,6.5568223,7.149124,7.7942433,8.311093,8.345046,7.383027,7.5301595,7.1906233,6.5945487,6.149379,6.4247804,6.730363,7.001992,7.118943,7.33021,8.235641,8.069645,8.741172,8.922258,8.639311,9.26934,8.009283,8.511042,8.710991,8.167733,8.047009,9.027891,9.099571,8.816625,8.348819,7.488661,8.677037,9.567377,10.38981,10.729345,9.5183325,9.997457,10.902886,11.087745,10.585986,10.612394,8.213005,6.934085,6.8850408,7.8810134,9.439108,9.4013815,8.43559,7.8244243,7.6584287,6.7944975,7.7037,7.0812173,6.3832817,6.0701537,5.6287565,4.06689,3.6443558,3.802806,4.1612053,4.52715,4.1272516,4.3875628,4.9987283,5.7079816,6.330465,6.8774953,7.250985,7.6395655,7.9791017,7.956466,8.858124,9.065618,9.748463,10.917976,11.427281,10.804798,10.902886,10.47658,9.6201935,9.786189,9.967276,9.654147,9.480607,9.793735,10.676529,9.857869,9.514561,9.906913,10.944386,12.178034,13.996439,13.004238,11.129244,9.880505,10.33322,10.401127,11.016065,10.642575,9.352338,8.83926,9.337247,10.582213,11.053791,11.125471,11.306557,12.234623,13.456953,13.88326,14.188843,14.600059,14.894323,15.55076,14.743419,13.830443,13.370183,13.12119,12.46098,12.1101265,12.030901,12.166716,12.423254,13.057055,14.068119,14.901869,15.245177,14.988639,15.260268,15.279131,15.335721,15.350811,14.852824,14.7321005,13.607859,12.830698,12.955194,13.732355,13.6833105,13.155144,12.464753,11.98563,12.151625,11.261286,11.442371,11.608367,11.276376,10.567122,10.834979,11.287694,11.672502,11.7894535,11.502733,10.608622,10.265312,10.155907,10.18986,10.49167,10.631257,10.499215,10.657665,11.185833,11.68382,12.057309,11.936585,11.868678,12.004493,12.128989,11.962994,12.310076,12.917468,13.588995,14.1926155,14.25675,14.490653,14.626467,14.562332,14.354838,15.516807,16.35433,16.42601,15.811071,15.131999,15.347038,14.924504,14.369928,14.124708,14.569878,15.17727,14.913187,14.418973,14.075664,14.000212,14.200161,13.86817,13.517315,13.449409,13.773854,13.728582,13.36641,12.728837,12.113899,12.083718,11.793225,11.25374,10.963248,11.02361,11.144334,11.457462,11.766817,11.751727,11.461235,11.314102,11.053791,10.940613,10.767072,10.627484,10.955703,10.812344,10.744436,10.518079,10.242677,10.38981,10.465261,10.989656,11.389555,11.431054,11.249968,10.944386,10.574668,10.250222,9.986138,9.7220545,9.371201,8.484633,7.462252,6.5643673,5.881522,5.6589375,5.5759397,5.5268955,5.6098933,6.126743,6.470052,6.6662283,6.802043,7.0510364,7.6395655,7.888559,8.43559,8.98262,9.303293,9.258021,9.246704,8.929804,8.661947,8.582722,8.616675,8.6581745,8.937348,9.337247,9.673011,9.703192,8.707218,8.14887,7.7640624,7.6093845,8.073418,8.643084,9.0543,9.408927,9.714509,9.876732,10.042727,10.631257,11.208468,11.378237,10.789707,10.355856,11.076427,11.978085,12.498707,12.498707,12.472299,12.47607,12.438345,11.917723,10.095545,8.948667,7.7338815,7.273621,7.4094353,7.020855,6.0814714,5.50426,5.27413,5.330719,5.5382137,5.5985756,5.7117543,5.847569,6.126743,6.858632,7.1679873,7.5112963,7.779153,8.062099,8.646856,9.224068,9.87296,10.702937,11.717773,12.83447,12.626976,11.261286,9.880505,8.707218,7.069899,6.700182,7.9526935,8.6732645,8.069645,6.7152724,6.0814714,5.9117036,6.4511886,7.6622014,9.239159,10.253995,10.914205,10.978339,10.627484,10.453944,10.801025,11.087745,11.487643,11.879996,11.868678,12.064855,13.332457,14.245432,14.611377,15.471535,15.396083,14.547242,13.245687,11.570641,9.363655,9.737145,9.035437,7.8206515,6.63982,6.013564,7.322665,7.8319697,7.707473,7.492433,8.084735,7.1906233,5.0439997,3.0935526,2.0258996,1.7731338,2.5238862,3.6368105,3.6292653,2.263575,0.52439487,0.27540162,0.25276586,0.4074435,1.6939086,6.0739264,3.531177,3.1652324,4.7610526,6.436098,4.6252384,3.7688525,3.289729,4.7836885,7.61693,8.933576,9.903141,11.25374,12.321393,12.698656,12.242168,13.943622,12.604341,12.306303,13.377728,12.393073,10.702937,10.208723,9.461743,8.669493,9.665465,9.831461,9.378746,8.529905,7.9300575,8.646856,6.911449,4.45547,2.1315331,0.6828451,0.73188925,2.263575,5.2137675,8.865668,11.921495,12.521342,6.579458,2.9086938,2.1843498,4.2404304,8.088508,7.145352,6.6549106,9.133525,12.7477,11.34051,6.6058664,7.375482,11.374464,15.214996,14.373701,12.223305,9.144843,7.424526,8.737399,14.166207,10.20495,6.013564,3.8782585,3.31991,1.0789708,2.1692593,3.6707642,4.3347464,3.783943,2.516341,2.7917426,3.4217708,3.9461658,4.5497856,6.0324273,6.2927384,7.0585814,7.3490734,7.062354,6.971811,7.1302614,7.6508837,8.412953,8.971302,8.537451,7.462252,7.8734684,8.563859,9.363655,11.144334,13.641812,15.32063,15.829934,15.596032,15.818617,16.056292,14.4152,14.690601,17.172989,18.636768,16.475054,14.769827,13.743673,13.075918,11.883769,11.393328,11.283921,11.351829,11.740409,12.921241,14.369928,14.381247,14.037937,13.660675,12.800517,12.472299,12.5326605,12.777881,12.894833,12.453435,11.7894535,12.174261,13.030646,13.981348,14.830189,15.260268,16.007248,16.746683,17.003222,16.146835,15.211224,14.11339,12.434572,10.457717,9.133525,9.318384,8.9788475,8.514814,8.156415,7.9753294,9.250477,9.8239155,9.673011,9.276885,9.6201935,9.593785,9.676784,9.454198,9.144843,9.582467,8.43559,7.3000293,6.688864,6.590776,6.462507,6.039973,6.1418333,6.273875,6.2399216,6.1342883,7.424526,8.801534,10.487898,12.404391,14.177525,15.663939,15.045229,14.7736,15.241405,14.796235,17.142809,20.187317,26.397057,34.870373,41.33665,51.92641,72.34763,78.791275,61.041073,22.469755,22.711203,21.545462,19.968504,17.972786,14.532151,21.228561,17.105082,10.95193,8.36391,11.725319,4.6818275,3.591539,4.4441524,4.5460134,2.5238862,3.4896781,5.455216,5.745708,4.255521,3.451952,8.054554,8.197914,5.956975,4.025391,5.7419353,4.429062,6.56814,10.733118,14.064346,12.287439,9.514561,9.64283,10.933067,11.461235,9.0807085,7.4999785,7.6395655,7.888559,7.6320205,7.24344,7.6508837,7.6622014,7.541477,7.326438,6.832224,6.907676,6.466279,6.096562,5.9607477,5.8098426,5.492942,5.2250857,5.492942,6.2361493,6.832224,6.3116016,5.9607477,6.1644692,6.5945487,6.205968,5.9305663,6.5228686,7.032173,7.326438,8.058327,7.707473,7.6282477,7.779153,7.8696957,7.375482,7.643338,7.7376537,7.54525,7.062354,6.398372,6.368191,6.2927384,6.198423,6.1531515,6.300284,5.9494295,6.0512905,6.3153744,6.221059,5.040227,4.919503,5.462761,5.5268955,5.2099953,5.855114,6.2625575,6.375736,6.217286,6.017337,6.2021956,5.9607477,5.80607,5.9984736,6.168242,5.3156285,6.3908267,7.1302614,7.213259,6.752999,6.3153744,7.745199,8.99771,9.676784,9.756008,9.574923,10.080454,10.416218,10.321902,9.665465,8.45068,7.665974,8.710991,9.26934,9.027891,9.684328,8.141325,8.582722,9.529651,9.808825,8.5563135,8.582722,7.594294,6.304056,5.292993,4.9987283,4.6931453,4.5950575,4.6327834,4.7572803,4.938366,4.745962,4.1310244,3.531177,3.2105038,3.2670932,3.9499383,5.138315,5.975838,6.3531003,6.9265394,6.7114997,6.4738245,6.33801,6.417235,6.79827,7.3792543,7.5716586,7.8206515,8.039464,7.6207023,7.835742,7.435844,6.6247296,5.8702044,5.8702044,6.417235,7.1000805,7.3792543,7.435844,8.182823,7.9828744,8.465771,8.756263,8.771353,9.22784,7.6282477,7.809334,8.118689,8.080963,8.386545,9.408927,9.386291,9.250477,9.050528,7.9338303,8.284684,9.0543,10.238904,11.083972,10.080454,9.42779,10.763299,11.506506,10.887795,9.9257765,8.14887,7.5829763,7.7640624,8.228095,8.52236,8.213005,7.0548086,6.9869013,7.745199,6.858632,7.605612,7.1264887,6.8171334,6.8397694,6.1078796,4.9157305,4.115934,3.772625,3.85185,4.2328854,4.0593443,4.353609,4.610148,4.851596,5.621211,6.417235,7.33021,7.7112455,7.586749,7.6810646,8.714764,8.83926,9.465516,10.518079,10.419991,9.876732,10.26154,9.910686,8.892077,9.016574,8.926031,8.907167,8.854351,8.873214,9.303293,9.725827,9.684328,10.03141,10.917976,11.8045435,13.721037,13.219278,11.574413,10.03141,9.793735,10.412445,10.608622,10.536942,10.529396,11.114153,9.654147,10.921749,11.159425,11.536687,12.272349,12.623203,13.962485,14.045483,14.520834,15.535669,15.739391,16.086473,14.698147,13.211733,12.313848,11.732863,11.438599,11.287694,11.480098,11.910177,12.14408,12.344029,13.400364,14.7170105,15.860115,16.546734,16.135517,14.973549,14.200161,13.951167,13.370183,13.29473,12.58925,12.751472,13.958713,15.067864,14.120935,12.728837,11.69891,11.442371,11.970539,12.717519,13.117417,12.668475,11.631002,11.019837,11.578186,11.910177,12.030901,11.879996,11.287694,10.484125,10.208723,10.416218,10.884023,11.234878,11.442371,11.234878,11.219787,11.495189,11.649866,12.362892,12.494934,12.50248,12.525115,12.415709,12.498707,13.094781,13.577678,13.630494,13.253232,13.155144,13.377728,13.781399,13.947394,13.170234,14.260523,14.9358225,15.116908,14.9358225,14.758509,14.720782,14.298248,13.898351,14.011529,15.222542,15.584714,15.026365,14.4114275,14.1058445,13.973803,14.003984,13.739901,13.5663595,13.528633,13.3626375,13.011784,12.981603,12.913695,12.811834,13.026875,12.347801,11.895086,11.46878,11.065109,10.887795,11.0613365,11.344283,11.317875,11.031156,11.004747,10.393582,10.220041,10.0465,9.906913,10.321902,9.895596,9.81637,9.608876,9.2844305,9.367428,9.74469,10.18986,10.585986,10.808571,10.7218,10.589758,10.397354,9.971047,9.374973,8.937348,8.480861,7.6282477,6.7680893,6.0814714,5.5570765,5.379763,5.3080835,5.194905,5.2099953,5.8513412,5.802297,5.666483,5.621211,5.7909794,6.255012,6.881268,7.7150183,8.303548,8.635539,9.118435,9.469289,9.122208,8.646856,8.394091,8.507269,8.4544525,8.537451,8.631766,8.756263,9.073163,8.231868,7.8696957,7.61693,7.333983,7.115171,7.3868,7.6395655,8.028146,8.5563135,9.092027,9.058073,9.042982,9.242931,9.484379,9.22784,9.159933,10.668983,12.083718,12.574159,12.147853,12.166716,12.438345,12.400619,11.574413,9.563604,8.428044,7.6697464,7.432071,7.375482,6.6813188,5.945657,5.6061206,5.6287565,5.8513412,5.9532022,5.8211603,5.8098426,5.828706,6.0211096,6.749226,7.303802,7.7037,8.080963,8.495952,8.937348,9.435335,9.9257765,10.472807,11.136789,11.989402,11.778135,10.702937,9.307066,7.9526935,6.832224,6.0776987,7.175533,7.6697464,7.01331,6.5568223,6.0550632,6.0211096,6.609639,7.816879,9.476834,10.076681,10.106862,9.831461,9.574923,9.710737,10.178542,10.653893,11.419736,12.291212,12.623203,12.366665,13.004238,13.736128,14.618922,16.58446,16.343012,14.905642,13.430545,12.189351,10.601076,10.801025,10.008774,9.246704,8.643084,7.432071,7.84706,6.862405,6.6247296,7.3905725,7.5527954,4.719554,3.3840446,2.5238862,1.8825399,1.961765,3.0671442,3.8103511,3.7688525,2.7238352,0.6828451,1.2147852,1.0148361,0.8639311,2.8181508,10.193633,4.5799665,3.561358,4.074435,4.247976,3.3953626,3.138824,3.9348478,5.2250857,6.700182,8.333729,9.891823,10.623712,10.997202,11.32542,11.759273,11.736636,11.46878,12.0233555,12.694883,10.978339,9.439108,9.152389,9.0543,9.314611,11.336739,10.499215,9.454198,8.563859,8.107371,8.29223,5.5985756,3.289729,1.4675511,0.543258,1.2261031,2.3880715,5.0025005,9.009028,13.2607765,15.524352,9.114662,4.2630663,2.7691069,4.659192,8.186596,10.63503,8.409182,8.729855,12.393073,13.773854,8.488406,9.039209,10.7218,11.480098,11.891314,12.208215,9.21275,7.4999785,8.858124,12.238396,9.118435,5.0477724,3.0822346,3.0369632,1.4939595,2.1994405,3.6556737,4.425289,3.942393,2.4974778,2.6974268,3.0105548,3.3463185,4.036709,5.8702044,6.436098,7.043491,7.466025,7.7112455,8.009283,8.065872,8.197914,8.209232,8.031919,7.707473,7.115171,7.7716074,8.699674,9.914458,12.427027,14.879233,16.188334,15.833707,14.894323,16.026112,15.943113,14.320885,13.788944,14.735873,15.294222,15.0376835,14.407655,13.834216,13.483362,13.287186,12.344029,12.083718,11.951676,12.012038,12.970284,14.652876,14.803781,14.781145,14.766054,13.739901,12.925014,12.811834,12.585477,11.951676,11.125471,11.087745,11.529142,12.298758,13.27964,14.381247,14.769827,15.271586,16.078928,16.750456,16.18456,13.9888935,12.555296,11.457462,10.540714,9.910686,9.914458,9.408927,8.726082,8.054554,7.454707,8.801534,9.476834,9.22784,8.586494,8.880759,8.560086,8.318638,8.137552,8.175279,8.7751255,8.314865,7.5075235,6.952948,6.802043,6.7454534,6.4549613,6.507778,6.4964604,6.3908267,6.56814,6.9793563,8.2507305,10.386037,12.559069,13.128735,13.619176,13.819125,13.879487,13.909668,13.966258,15.931795,19.134754,24.107073,30.245134,35.81353,38.8769,41.993088,38.34496,27.78161,16.82968,18.45568,18.87067,18.791445,16.739138,8.99771,14.64533,13.238141,9.646602,7.9941926,11.664956,7.1981683,5.885295,6.7379084,7.281166,3.5689032,3.7009451,4.244203,6.1116524,8.028146,6.5266414,7.1000805,5.66271,5.040227,6.4738245,9.58624,7.443389,7.466025,9.22784,10.140816,5.4703064,6.228604,7.6848373,8.937348,9.42779,8.903395,8.111144,7.756517,7.5188417,7.2057137,6.7756343,7.2623034,7.213259,7.2358947,7.2924843,6.7152724,6.673774,6.205968,5.956975,6.0248823,5.975838,5.696664,5.0213637,4.9232755,5.832478,7.624475,6.515323,6.1720147,6.6247296,7.183078,6.4436436,6.115425,6.549277,6.9944468,7.149124,7.1566696,7.3453007,7.5716586,7.541477,7.326438,7.364164,8.069645,7.84706,7.3490734,6.934085,6.673774,6.7341356,6.5832305,6.398372,6.40969,6.8850408,6.598321,6.4134626,6.771862,7.17176,6.156924,5.4363527,5.9230213,5.907931,5.240176,5.3269467,5.9682927,6.156924,5.8890676,5.5683947,5.9984736,6.270103,6.326692,6.571913,6.809588,6.2436943,6.9454026,7.624475,7.9036493,7.6584287,7.0170827,8.643084,9.590013,9.87296,9.673011,9.35611,9.680555,10.042727,9.940866,9.250477,8.243186,7.7301087,8.914713,9.35611,9.035437,10.340765,8.424272,9.280658,10.47658,10.419991,8.397863,8.235641,7.4811153,6.428553,5.5495315,5.523123,5.2628117,5.1835866,5.0175915,4.749735,4.6327834,4.6856003,4.3611546,3.8254418,3.361409,3.3764994,3.9574835,5.062863,5.824933,6.145606,6.7152724,6.5002327,6.5945487,6.730363,6.832224,7.0510364,7.699928,7.696155,7.6508837,7.798016,8.00551,8.054554,7.3868,6.3153744,5.3646727,5.247721,6.217286,7.3679366,7.7904706,7.726336,8.552541,7.9413757,8.122461,8.518587,8.756263,8.654402,7.677292,7.6697464,7.884786,8.047009,8.337502,8.98262,9.178797,9.465516,9.57115,8.386545,8.258276,8.582722,9.507015,10.431308,9.963503,8.892077,10.26154,11.302785,10.993429,10.042727,8.873214,8.782671,8.907167,8.748717,8.186596,7.5263867,6.4021444,6.3832817,7.213259,6.820906,7.1378064,6.8473144,6.8171334,6.94163,6.1305156,5.3458095,4.6327834,4.134797,3.9159849,3.9461658,3.8669407,4.0706625,4.142342,4.2630663,5.2288585,6.319147,7.54525,8.14887,8.039464,7.779153,8.548768,8.816625,9.325929,9.978593,9.827688,9.835234,10.208723,9.899368,9.103344,9.231613,8.548768,8.692128,8.835487,8.635539,8.239413,9.046755,9.273112,9.763554,10.63503,11.261286,13.117417,13.555041,12.540206,10.665211,9.122208,9.695646,9.910686,10.397354,11.423509,12.921241,10.653893,11.498961,11.9064045,12.427027,13.162688,13.762536,14.452927,14.698147,14.996184,15.32063,15.109364,15.113135,14.324657,13.332457,12.445889,11.69891,11.532914,11.498961,11.631002,11.898859,12.170488,12.0082655,12.630749,13.6833105,15.079182,16.995676,15.758255,13.615403,12.37421,12.257258,11.917723,11.495189,11.276376,12.294985,13.93985,13.95494,12.943876,11.672502,11.034928,11.129244,11.216014,13.385274,13.426772,12.234623,10.891568,10.687846,10.989656,11.272603,11.532914,11.646093,11.329193,10.770844,10.616167,10.970794,11.61214,12.0082655,12.061082,11.970539,11.864905,11.778135,11.668729,12.272349,12.294985,12.2119875,12.170488,11.974312,12.408164,12.958967,13.385274,13.340002,12.355347,12.664702,12.917468,13.287186,13.585222,13.257004,13.204187,13.151371,13.415455,13.93985,14.302021,14.139798,13.604086,13.539951,14.211478,15.316857,14.754736,13.894578,13.430545,13.528633,13.822898,13.600313,13.328684,12.992921,12.611885,12.264804,11.446144,11.910177,12.713746,13.306048,13.517315,13.143826,12.90615,12.67602,12.362892,11.921495,11.7026825,11.781908,11.3971,10.725573,10.86516,10.103089,9.782416,9.616421,9.57115,9.87296,9.242931,8.8769865,8.518587,8.213005,8.307321,8.601585,8.8618965,9.220296,9.6051035,9.737145,9.733373,9.944639,9.590013,8.771353,8.465771,8.039464,7.2170315,6.3455553,5.7607985,5.7872066,5.3646727,5.240176,5.1458607,5.13077,5.572167,5.3080835,5.402399,5.2854476,4.9534564,4.9723196,6.089017,6.964266,7.537705,8.031919,8.952439,9.533423,9.488152,9.035437,8.495952,8.280911,8.182823,8.145098,8.028146,7.937603,8.235641,8.050782,7.9262853,7.8621507,7.7225633,7.2358947,7.4584794,7.4697976,7.484888,7.6848373,8.201687,8.5563135,8.401636,8.495952,8.918486,9.0957985,9.623966,11.283921,12.423254,12.434572,11.751727,11.951676,12.276122,12.076173,11.02361,9.110889,8.197914,7.541477,7.2170315,6.952948,6.1606965,5.715527,5.7117543,6.013564,6.379509,6.4738245,6.1531515,6.0324273,6.058836,6.217286,6.5341864,7.220804,7.877241,8.480861,8.914713,8.959985,9.171251,9.673011,10.223814,10.676529,10.948157,10.767072,10.155907,8.929804,7.575431,7.232122,6.470052,6.752999,7.0246277,7.0170827,7.24344,6.820906,6.8774953,7.2887115,8.009283,9.058073,9.435335,9.039209,8.563859,8.382772,8.563859,9.224068,9.933322,10.729345,11.717773,13.091009,13.27964,13.336229,13.622949,14.592513,16.784409,16.229834,14.84528,13.634267,12.853333,11.993175,12.012038,10.801025,9.95973,9.563604,8.186596,8.29223,5.7381625,5.6325293,7.6923823,6.2361493,2.5540671,1.8636768,1.8787673,1.5580941,1.1204696,1.7165444,1.7731338,2.3993895,3.5651307,4.0970707,3.832987,2.4107075,2.5125682,5.7117543,12.449662,8.397863,6.771862,5.594803,4.164978,3.0633714,2.263575,4.2064767,5.613666,6.3945994,9.654147,10.56335,9.831461,9.457971,9.982366,10.518079,10.242677,10.785934,11.32542,11.099063,9.416472,9.386291,9.325929,9.74469,10.86516,12.626976,10.604849,9.450426,8.75249,8.126234,7.2283497,4.5422406,2.4597516,1.0525624,0.73188925,2.252257,3.2972744,4.8138695,7.696155,11.438599,14.158662,9.971047,5.9494295,4.142342,5.0779533,7.7602897,16.173243,10.985884,7.9489207,11.25374,13.513543,9.782416,10.868933,10.442626,7.9413757,8.578949,10.608622,8.590267,7.3000293,8.714764,11.981857,9.574923,5.0025005,2.463524,2.4597516,1.780679,2.335255,3.7537618,4.304565,3.5236318,2.2371666,2.757789,2.9615107,3.470815,4.459243,5.6287565,6.368191,7.0284004,7.7829256,8.488406,8.695901,8.907167,8.956212,8.6732645,8.156415,7.8017883,7.6282477,8.201687,8.986393,10.216269,12.879742,14.766054,15.505488,15.294222,14.966003,15.999702,15.411173,13.902123,13.034419,13.04951,12.883514,13.460726,13.479589,12.985375,12.649611,13.777626,12.740154,12.751472,12.736382,12.487389,12.664702,14.377474,14.890551,15.4074,15.992157,15.580941,14.068119,13.630494,13.143826,12.340257,11.808316,12.038446,12.283667,12.683565,13.20796,13.626721,13.913441,14.766054,15.848798,16.81459,17.30503,14.332202,12.310076,11.359374,11.076427,10.536942,10.253995,9.654147,9.042982,8.495952,7.8508325,8.827943,9.450426,9.250477,8.601585,8.710991,7.537705,6.8850408,6.900131,7.4811153,8.303548,8.45068,8.062099,7.432071,6.7680893,6.1720147,5.8626595,5.6815734,5.6815734,5.8928404,6.330465,6.247467,7.3981175,9.831461,12.294985,12.2270775,11.59705,12.245941,12.872196,13.0646,13.324911,15.196134,18.0671,21.651094,25.174726,27.366621,24.054256,20.1345,16.856089,15.524352,17.53139,14.679284,14.162435,15.588487,16.033657,10.03141,12.268577,14.464244,11.668729,6.1229706,7.24344,9.242931,9.325929,10.95193,12.604341,7.809334,4.6516466,4.236658,8.27714,13.558814,11.962994,7.3490734,4.112161,4.8968673,9.178797,13.272095,10.767072,12.200669,14.992412,15.264041,7.8734684,5.455216,7.069899,9.186342,9.7220545,8.039464,8.216777,7.54525,6.9189944,6.6624556,6.5040054,6.8661776,6.802043,6.722818,6.7077274,6.4926877,6.628502,5.9003854,5.6023483,6.006019,6.356873,6.273875,5.149633,4.640329,5.5495315,7.8508325,6.72659,6.7152724,7.1076255,7.3188925,6.900131,6.3153744,5.9418845,6.175787,6.617184,6.058836,6.7831798,7.4282985,7.4999785,7.2358947,7.5829763,7.748972,7.4169807,7.0963078,7.01331,7.1302614,7.5226145,7.643338,7.635793,7.677292,7.9338303,7.8923316,7.2283497,7.1566696,7.654656,7.466025,6.507778,6.3945994,6.0022464,5.2175403,4.938366,5.3986263,5.7570257,5.696664,5.3609,5.372218,6.149379,6.677546,7.066127,7.3679366,7.5603404,7.7338815,8.031919,8.345046,8.495952,8.273367,9.839006,10.374719,10.223814,9.74469,9.288202,9.14107,9.367428,9.348565,8.858124,8.07719,7.4584794,8.382772,8.7751255,8.707218,10.38981,9.933322,10.54826,11.050018,10.555805,8.495952,7.575431,6.8699503,6.1229706,5.455216,5.3646727,5.4438977,5.6400743,5.523123,5.028909,4.447925,4.29702,4.327201,4.244203,3.8895764,3.2670932,3.7273536,4.7572803,5.523123,5.915476,6.530414,6.3719635,6.5568223,6.888813,7.1868505,7.277394,7.9225125,8.028146,7.99042,8.080963,8.469543,8.122461,7.277394,6.1003346,5.0968165,5.089271,6.2927384,7.7112455,8.175279,7.99042,8.971302,7.884786,7.7640624,8.013056,8.137552,7.745199,7.8696957,7.9791017,8.050782,8.043237,7.8696957,7.960239,8.605357,9.2995205,9.435335,8.299775,8.68081,8.801534,9.050528,9.416472,9.495697,9.265567,10.197406,10.79348,10.725573,10.853842,10.235131,10.005001,9.710737,9.25425,8.892077,7.7904706,6.587003,5.9494295,6.006019,6.3945994,6.6247296,6.40969,6.349328,6.3832817,5.772116,5.13077,4.8327327,4.644101,4.395108,3.9499383,3.7273536,3.6858547,3.712263,4.006528,5.0741806,6.5341864,7.828197,8.778898,9.0957985,8.345046,8.533678,8.903395,9.2995205,9.6051035,9.767326,10.401127,10.638803,10.435081,10.072908,10.148361,9.061845,9.133525,9.2995205,8.9788475,8.088508,7.77538,7.858378,8.544995,9.646602,10.555805,12.792972,14.422746,14.400109,12.577931,9.7069645,9.137298,9.559832,10.461489,11.664956,13.313594,11.457462,12.864652,13.487134,13.792717,14.1058445,14.618922,15.230087,15.784663,15.501716,14.622695,14.388792,14.449154,14.264296,13.800262,13.162688,12.58925,12.113899,12.276122,12.193124,11.717773,11.476325,12.3289385,12.928786,13.694629,14.554788,14.909414,13.358865,12.310076,11.717773,11.491416,11.491416,11.52537,11.993175,12.864652,13.502225,12.649611,11.747954,10.917976,10.306811,9.884277,9.446653,10.676529,10.978339,10.740664,10.272858,9.797507,9.895596,10.246449,10.589758,10.789707,10.86516,10.853842,10.895341,10.925522,10.948157,11.031156,11.046246,11.046246,10.933067,10.812344,11.031156,11.129244,11.393328,11.838497,12.23085,12.083718,12.098808,12.0082655,12.027128,12.208215,12.449662,12.306303,12.626976,12.985375,13.158916,13.12119,13.257004,13.600313,14.034165,14.48688,14.939595,13.826671,13.008011,13.075918,13.792717,14.083209,14.449154,14.203933,14.007756,14.203933,14.800008,13.970031,13.132507,12.393073,11.936585,12.0082655,11.581959,11.548005,11.664956,11.830952,12.098808,12.638294,12.955194,13.290957,13.517315,13.151371,13.287186,12.551523,11.3669195,10.291721,10.008774,9.95973,9.639057,9.484379,9.480607,9.14107,8.284684,7.6508837,7.254758,7.232122,7.8432875,8.231868,8.394091,8.537451,8.66572,8.590267,8.858124,9.035437,8.952439,8.695901,8.635539,8.111144,7.2283497,6.4134626,5.9192486,5.8588867,5.455216,4.9723196,4.689373,4.719554,4.9760923,5.0213637,5.2099953,5.251494,5.093044,4.8968673,4.776143,5.1571784,5.8966126,6.8661776,7.964011,8.624221,8.631766,8.280911,7.8017883,7.4018903,7.1566696,7.115171,7.2585306,7.541477,7.858378,7.7112455,7.756517,8.069645,8.503497,8.710991,8.993938,9.246704,9.307066,9.205205,9.156161,8.959985,9.065618,9.703192,10.570895,10.86516,11.268831,12.702429,13.588995,13.373956,12.559069,11.642321,11.076427,10.714255,10.295494,9.416472,8.36391,7.5905213,7.273621,7.0887623,6.2097406,5.9909286,6.0626082,6.247467,6.436098,6.6058664,6.326692,6.009792,6.119198,6.5568223,6.6662283,7.326438,8.179051,8.782671,9.058073,9.276885,9.461743,9.982366,10.329447,10.336992,10.178542,10.446399,9.771099,8.654402,7.745199,7.8432875,7.3415284,7.1000805,7.092535,7.2924843,7.6584287,7.99042,8.073418,7.858378,7.6886096,8.299775,8.8618965,9.854096,9.914458,8.990166,8.329956,8.062099,8.793989,9.469289,9.891823,10.695392,12.479843,14.286931,15.894069,17.199398,18.248188,16.931541,16.490145,16.063837,15.082954,13.275867,12.091263,9.982366,8.009283,6.719045,6.1342883,6.1342883,4.908185,4.768598,5.2967653,3.3576362,1.539231,1.1846043,1.8674494,2.4522061,1.0827434,1.0827434,0.76207024,1.3543724,5.406172,16.769318,8.065872,3.2821836,5.881522,12.2270775,11.581959,9.446653,4.9647746,2.0296721,2.3088465,5.247721,2.6597006,3.6179473,6.888813,10.533169,11.902632,9.789962,9.42779,9.81637,10.152134,9.812597,9.6051035,9.533423,9.001483,8.303548,8.620448,9.940866,10.33322,10.985884,11.763044,11.200924,9.967276,9.137298,8.616675,7.937603,6.2399216,3.8367596,2.1088974,0.98465514,1.0940613,3.7537618,4.3385186,4.870459,6.620957,8.933576,9.201432,12.287439,9.948412,7.213259,6.1229706,5.723072,12.5326605,9.337247,7.8810134,11.793225,16.59955,10.155907,8.390318,6.741681,4.4894238,4.745962,4.1612053,3.308592,4.927048,8.307321,9.307066,8.892077,5.2628117,2.6898816,2.4522061,2.8521044,2.2069857,3.802806,4.304565,3.1048703,2.335255,2.505023,2.6106565,3.5538127,4.9685473,5.247721,5.836251,6.6322746,7.858378,9.035437,8.986393,9.756008,10.050273,9.623966,8.971302,9.337247,9.06939,9.623966,9.846551,9.654147,10.069136,12.034674,12.921241,13.664448,14.460471,14.754736,13.951167,13.317367,13.226823,13.422999,13.030646,12.981603,13.034419,12.464753,11.680047,12.193124,12.166716,12.709973,13.102326,13.238141,13.641812,14.592513,14.520834,14.6302395,15.388537,16.509007,15.045229,14.449154,13.894578,13.287186,13.275867,13.249459,12.958967,13.094781,13.675766,14.053028,13.8719425,14.079436,14.02662,13.962485,15.060319,12.826925,10.933067,10.163452,10.110635,9.171251,9.805053,10.091772,9.971047,9.695646,9.842778,9.97482,10.110635,10.072908,9.944639,10.054046,8.710991,7.2962565,6.802043,7.413208,8.499724,8.646856,8.60913,8.322411,7.6622014,6.4549613,6.1116524,5.9909286,6.356873,6.952948,6.9869013,6.2927384,6.9152217,9.050528,11.691365,12.619431,12.385528,12.37421,12.766563,13.140053,12.483616,12.992921,14.011529,15.358356,16.561823,16.82968,13.498452,10.367173,9.371201,10.008774,9.337247,11.487643,12.785426,14.381247,15.62244,14.022847,11.434827,10.001229,7.8508325,5.975838,8.209232,9.465516,9.81637,15.426264,22.518799,17.380484,8.371455,6.0550632,7.1340337,9.276885,11.106608,8.605357,4.1083884,2.4295704,5.6815734,13.2607765,14.3095665,16.712729,18.184053,17.286167,13.426772,6.126743,6.205968,9.608876,11.185833,4.7308717,4.7421894,5.8437963,6.119198,5.723072,6.881268,7.1378064,7.118943,6.507778,5.5985756,5.2967653,6.187105,5.6287565,5.119452,5.281675,5.904158,5.783434,5.4778514,6.2399216,7.352846,6.119198,5.3759904,6.25124,6.719045,6.375736,6.4247804,5.0062733,4.617693,5.624984,6.911449,5.873977,6.375736,7.1679873,7.9489207,8.461998,8.499724,7.462252,7.4018903,7.4509344,7.3113475,7.2623034,7.5301595,7.9451485,8.484633,8.8618965,8.544995,9.216523,8.99771,8.345046,7.635793,7.17176,6.19465,5.7419353,5.6551647,5.6098933,5.0968165,5.402399,5.485397,5.4703064,5.2250857,4.395108,5.6513925,6.752999,7.432071,7.8319697,8.514814,8.646856,9.001483,9.525878,10.03141,10.178542,10.495442,9.933322,9.548513,9.654147,9.812597,9.125979,8.782671,8.661947,8.567632,8.224322,7.322665,7.7640624,7.5075235,6.934085,8.850578,11.84227,12.468526,11.649866,10.095545,8.299775,7.605612,6.296511,5.342037,5.0213637,4.9119577,5.5004873,5.828706,5.643847,5.081726,4.6554193,4.2027044,3.9876647,4.3422914,4.7950063,4.074435,4.025391,4.957229,5.621211,5.7381625,5.9796104,5.726845,5.945657,6.458734,7.0472636,7.462252,7.8508325,8.114917,8.480861,8.944894,9.261794,8.420499,7.586749,6.511551,5.6400743,6.1041074,6.8850408,8.103599,8.337502,7.752744,8.118689,7.1302614,6.964266,7.1340337,7.3415284,7.4773426,7.122716,6.907676,7.0849895,7.5037513,7.6131573,7.515069,8.269594,8.8618965,8.7751255,7.9941926,8.533678,9.929549,10.469034,10.042727,10.178542,11.472552,11.91395,10.978339,9.559832,9.963503,10.574668,9.876732,9.333474,9.35611,9.307066,7.745199,6.1720147,5.142088,4.8666863,5.2326307,6.149379,6.039973,6.1078796,6.4210076,5.9192486,5.138315,4.696918,4.768598,4.938366,4.1800685,3.6669915,3.410453,3.3463185,3.5387223,4.195159,6.1720147,7.7112455,8.744945,9.065618,8.345046,8.552541,8.75249,8.843033,9.009028,9.703192,10.303039,10.827434,11.155652,11.125471,10.514306,10.023865,10.370946,10.38981,9.895596,9.673011,7.586749,7.1302614,7.635793,8.616675,9.752235,11.947904,14.958458,16.852316,16.471281,13.441863,10.940613,10.416218,10.978339,11.895086,12.604341,11.068882,12.355347,13.853079,14.015302,13.302276,14.166207,14.950912,16.218515,16.490145,15.79598,15.682802,14.728328,14.083209,13.717264,13.381501,12.611885,12.4307995,12.095036,11.717773,11.461235,11.548005,12.234623,12.566614,12.909923,13.162688,12.736382,12.113899,11.92904,11.710228,11.457462,11.61214,11.355601,11.529142,11.766817,11.838497,11.649866,11.185833,10.751981,10.646348,10.631257,9.910686,9.95973,10.072908,10.069136,9.861642,9.454198,9.895596,10.340765,10.684074,10.797253,10.559577,10.665211,10.770844,10.763299,10.702937,10.834979,11.053791,11.268831,11.314102,11.242422,11.32542,11.638548,11.638548,11.604594,11.747954,12.208215,11.966766,12.370438,12.611885,12.408164,12.00072,12.351574,13.008011,13.860624,14.351066,13.475817,13.649357,13.93985,13.913441,13.72481,14.109617,13.389046,13.12119,13.177779,13.234368,12.766563,12.54775,12.585477,12.826925,13.204187,13.615403,13.343775,12.90615,12.427027,11.902632,11.216014,10.533169,10.3634,10.729345,11.268831,11.234878,11.876224,12.411936,12.97783,13.588995,14.128481,14.166207,13.158916,11.849815,10.661438,9.669238,8.741172,8.503497,8.514814,8.484633,8.311093,7.7301087,7.1038527,6.752999,6.802043,7.2094865,7.5792036,7.786698,7.786698,7.7150183,7.907422,7.8810134,7.8998766,7.997965,8.09228,7.9526935,7.564113,7.0472636,6.4436436,5.828706,5.311856,4.957229,4.557331,4.398881,4.466788,4.447925,4.3422914,4.678055,5.010046,5.0968165,4.9119577,4.8666863,5.304311,5.8211603,6.3644185,7.220804,7.194396,7.4735703,7.5792036,7.4584794,7.484888,7.213259,7.1566696,7.2283497,7.4169807,7.7716074,7.673519,7.541477,7.6848373,8.111144,8.552541,9.978593,10.559577,10.552032,10.231359,9.899368,9.371201,9.661693,10.125726,10.7218,12.00072,12.37421,12.823153,13.000465,12.672247,11.729091,11.027383,10.616167,10.419991,10.125726,9.171251,8.296002,7.3679366,6.749226,6.4926877,6.356873,6.3342376,6.587003,6.7454534,6.6850915,6.5341864,6.3719635,6.2361493,6.48137,7.1038527,7.7414265,8.36391,8.52236,8.397863,8.348819,8.899622,9.288202,9.948412,10.216269,9.933322,9.431562,9.703192,8.801534,7.779153,7.2396674,7.3188925,7.3151197,7.3490734,7.2057137,7.0359454,7.3415284,7.575431,8.239413,8.744945,9.058073,9.718282,9.857869,10.93684,11.359374,10.699164,9.699419,8.560086,8.356364,8.379,8.446907,8.903395,10.997202,13.075918,14.664193,15.528125,15.660167,15.799753,16.807045,17.071129,16.120426,14.603831,13.068373,9.710737,7.7112455,7.3453007,5.938112,6.066381,5.323174,4.485651,3.5575855,1.780679,1.4071891,3.2746384,5.149633,5.5985756,3.9763467,3.1954134,6.6624556,8.59404,7.854605,7.9791017,6.1229706,4.7912335,4.8327327,5.87775,6.3342376,5.553304,3.5877664,2.3767538,2.5201135,3.2972744,4.8666863,9.865415,13.947394,14.634012,11.314102,9.507015,10.208723,10.763299,10.1294985,8.858124,9.910686,9.1825695,8.484633,8.465771,8.60913,9.820143,10.295494,10.47658,10.38981,9.661693,9.092027,8.707218,8.182823,7.3490734,6.1795597,3.4934506,1.7014539,0.8601585,1.2110126,3.169005,3.4594972,3.802806,4.0291634,4.3724723,5.4401255,6.2927384,7.4735703,11.536687,15.448899,10.604849,16.01102,9.95973,6.934085,11.974312,20.689075,11.676274,8.563859,7.0887623,5.1760416,2.9501927,3.742444,6.368191,8.013056,7.5527954,5.583485,6.2361493,4.323428,3.0935526,3.2746384,3.0746894,2.1051247,3.4745877,4.2404304,3.6254926,2.9803739,2.8219235,2.7200627,3.1425967,3.9461658,4.395108,5.66271,6.530414,7.541477,8.643084,9.171251,10.182315,9.906913,8.880759,8.09228,8.99771,9.948412,10.518079,10.178542,9.363655,9.446653,11.227332,11.970539,12.642066,13.245687,12.826925,13.505998,14.166207,15.135772,15.633758,13.788944,13.075918,13.679539,13.422999,12.347801,12.706201,12.027128,12.30253,12.815607,13.257004,13.739901,14.234114,14.558559,14.70192,14.864142,15.460217,14.883006,14.856597,14.381247,13.223051,11.872451,12.344029,12.294985,12.261031,12.562841,13.321139,13.468271,13.340002,12.679792,11.993175,12.5326605,11.41219,10.593531,10.3634,10.499215,10.291721,11.065109,11.729091,11.879996,11.400873,10.465261,9.884277,9.344792,9.25425,9.673011,10.310584,10.453944,9.371201,8.548768,8.552541,9.024119,8.329956,8.311093,8.650629,8.729855,7.6395655,7.2396674,7.232122,7.424526,7.5490227,7.2924843,6.247467,6.3644185,7.786698,10.242677,13.045737,13.664448,12.838243,11.955449,11.476325,10.944386,11.710228,12.796744,13.083464,12.90615,14.083209,12.762791,11.136789,9.684328,8.616675,7.8998766,10.035183,11.646093,12.687338,12.996693,12.276122,7.443389,6.217286,6.156924,6.587003,8.586494,9.159933,11.891314,13.604086,14.056801,15.939341,12.506252,8.420499,6.5568223,7.9753294,11.925267,14.249205,13.275867,11.570641,10.540714,10.47658,10.18986,10.838752,9.552286,7.8432875,11.619685,8.831716,8.7600355,8.190369,6.7077274,6.696409,7.432071,9.635284,9.088254,5.8588867,4.293247,6.1116524,6.79827,6.5756855,5.855114,5.247721,6.175787,5.7117543,5.956975,6.888813,6.368191,6.0512905,5.983383,6.7869525,7.7187905,6.692637,5.194905,4.5724216,4.6931453,5.119452,5.13077,4.2404304,4.640329,5.2288585,5.3382645,4.7535076,5.8664317,6.7643166,7.665974,8.529905,9.035437,8.537451,8.75249,8.36391,7.5226145,7.8244243,7.4584794,7.6697464,8.401636,9.193887,9.178797,9.997457,9.759781,9.265567,8.744945,7.8319697,6.63982,6.3719635,6.198423,5.5985756,4.3649273,4.327201,4.5988297,5.05909,5.413717,5.198677,6.2625575,7.4094353,7.9262853,7.745199,7.4509344,7.7338815,7.8961043,8.560086,9.7296,10.812344,11.080199,10.608622,9.669238,8.884532,9.250477,9.092027,8.793989,8.514814,8.333729,8.224322,7.24344,7.3377557,7.6320205,8.09228,9.522105,12.562841,13.275867,12.51757,10.93684,8.98262,7.8395147,6.4926877,5.5004873,4.870459,4.0480266,4.2517486,4.9534564,5.292993,5.028909,4.5309224,4.304565,3.9650288,4.1762958,4.7648253,4.708236,4.247976,4.889322,5.723072,6.168242,5.934339,5.1081343,5.2552667,5.8400235,6.56814,7.364164,7.8131065,7.7376537,7.91874,8.416726,8.578949,8.088508,7.254758,6.5040054,6.043745,5.8702044,6.8171334,7.9489207,8.439363,8.13378,7.54525,6.5341864,6.730363,7.001992,7.01331,7.24344,7.605612,7.2585306,7.0887623,7.3113475,7.4811153,6.8058157,7.564113,8.360137,8.707218,9.020347,8.299775,9.0807085,10.303039,11.208468,11.363147,11.921495,12.396846,12.162943,11.465008,11.378237,11.32542,10.352083,9.103344,8.182823,8.122461,7.5490227,6.7643166,5.772116,4.8553686,4.587512,4.9949555,4.859141,5.3344917,6.217286,5.9682927,5.353355,5.0477724,4.798779,4.5535583,4.4630156,4.183841,3.7348988,3.5538127,3.7877154,4.3196554,6.277648,7.677292,8.420499,8.718536,9.092027,9.748463,9.7296,9.205205,8.729855,9.22784,9.525878,9.952185,10.408672,10.597303,10.038955,9.861642,10.27663,10.450171,10.072908,9.35611,7.1906233,6.832224,7.360391,8.2507305,9.333474,10.967021,13.743673,15.784663,15.603577,12.08749,11.038701,10.921749,11.317875,11.69891,11.419736,10.386037,12.200669,13.223051,13.087236,12.611885,13.807808,14.049255,14.494425,15.218769,15.712983,14.890551,14.019074,13.215506,12.872196,12.826925,12.381755,12.411936,12.513797,12.47607,12.261031,12.015811,12.623203,12.385528,12.147853,12.076173,11.615912,11.947904,12.189351,12.147853,11.846043,11.506506,11.374464,11.744182,12.0724,12.019584,11.442371,11.099063,11.0613365,11.038701,10.819888,10.291721,10.016319,10.208723,10.453944,10.495442,10.227587,10.514306,10.657665,10.623712,10.555805,10.79348,11.155652,11.46878,11.623458,11.725319,12.106354,12.287439,12.66093,12.755245,12.574159,12.570387,12.694883,12.857106,12.947649,13.060828,13.4644985,13.604086,13.52486,13.306048,12.898605,12.132762,12.419481,13.343775,14.124708,14.0983,12.740154,13.370183,13.377728,13.04951,12.736382,12.838243,12.543978,12.581704,12.638294,12.366665,11.393328,11.34051,11.491416,11.830952,12.272349,12.66093,12.872196,12.562841,12.027128,11.472552,11.016065,10.461489,10.370946,10.665211,11.072655,11.155652,12.1252165,12.725064,13.072145,13.272095,13.411682,13.396591,12.2119875,10.804798,9.567377,8.329956,7.232122,7.066127,6.983129,6.730363,6.647365,6.3153744,5.987156,5.938112,6.1908774,6.5002327,6.470052,6.519096,6.488915,6.4549613,6.749226,6.7944975,6.771862,6.930312,7.2472124,7.3981175,7.0585814,6.5341864,5.9192486,5.300538,4.7610526,4.447925,4.22534,4.0404816,3.8858037,3.8254418,3.9688015,4.266839,4.666737,4.9949555,4.9232755,4.927048,5.198677,5.492942,5.7494807,6.119198,6.349328,6.7077274,6.930312,7.145352,7.8734684,7.6810646,7.7942433,7.8206515,7.6697464,7.5603404,7.194396,7.2962565,7.61693,8.028146,8.514814,9.540969,10.038955,10.220041,10.076681,9.337247,9.084481,9.016574,9.14107,9.661693,10.974566,11.774363,12.147853,12.181807,11.932813,11.438599,10.797253,10.514306,10.442626,10.121953,8.771353,7.99042,7.2396674,6.628502,6.2927384,6.3945994,6.2135134,6.398372,6.4738245,6.330465,6.258785,6.2851934,6.356873,6.5455046,6.8850408,7.3981175,7.605612,7.4471617,7.303802,7.5527954,8.575176,9.103344,9.480607,9.805053,9.891823,9.2844305,9.325929,8.590267,7.6320205,7.039718,7.435844,7.5565677,7.6282477,7.432071,7.043491,6.8133607,7.0887623,8.016829,8.8769865,9.522105,10.3634,10.751981,11.574413,11.706455,10.910432,9.839006,8.431817,7.84706,7.6584287,7.726336,8.216777,9.940866,12.079946,13.468271,13.747445,13.358865,14.562332,16.392056,17.753973,17.501207,14.445381,12.989148,10.182315,8.710991,8.412953,6.2663302,6.930312,6.326692,4.4441524,2.1692593,1.2713746,1.5505489,4.0782075,5.0515447,3.731126,2.4559789,2.2711203,3.682082,4.406426,4.036709,4.0517993,5.281675,5.1043615,4.6818275,5.8437963,11.072655,7.3792543,5.7683434,4.979865,4.9459114,6.790725,11.151879,13.826671,14.7321005,14.068119,12.321393,11.019837,10.612394,10.242677,9.6051035,8.967529,9.265567,8.469543,8.141325,8.575176,8.797762,9.967276,10.487898,10.265312,9.650374,9.461743,9.144843,8.816625,8.262049,7.375482,6.145606,3.5575855,1.8070874,0.80734175,0.87147635,2.727608,3.9499383,4.4177437,4.055572,4.3196554,8.190369,7.575431,7.8810134,10.099318,11.936585,7.835742,10.514306,10.438853,9.963503,11.423509,17.14658,10.616167,7.394345,5.6589375,4.568649,4.2592936,9.835234,15.78089,14.551015,7.5188417,4.983638,7.1604424,4.217795,2.41448,3.0822346,2.625747,1.8372684,3.2557755,4.187614,3.92353,3.7386713,3.983892,4.014073,3.9461658,3.9348478,4.191386,5.617439,5.9192486,6.149379,6.7869525,7.707473,8.488406,8.582722,8.333729,8.179051,8.646856,9.201432,9.5183325,9.303293,8.89585,9.291975,10.220041,10.676529,12.140307,14.075664,13.947394,14.434063,14.475562,14.924504,15.784663,16.218515,16.131744,16.712729,16.705183,15.686575,14.079436,12.721292,12.162943,12.095036,12.611885,14.203933,14.618922,14.517061,14.154889,13.902123,14.264296,14.275613,14.468017,14.169979,13.140053,11.593277,11.751727,11.944131,12.23085,12.73261,13.6682205,14.120935,13.849306,13.102326,12.245941,11.7555,11.102836,10.838752,11.004747,11.404645,11.6008215,12.272349,13.158916,13.494679,12.981603,11.800771,10.933067,10.106862,9.910686,10.450171,11.374464,12.774108,12.7477,12.166716,11.336739,9.997457,7.9753294,7.6886096,8.348819,9.110889,9.0957985,8.258276,7.84706,7.6320205,7.435844,7.115171,6.587003,6.436098,7.537705,9.850324,12.438345,13.819125,13.079691,12.049765,11.438599,10.842525,11.393328,12.577931,13.004238,12.830698,13.773854,12.792972,11.18206,9.473062,8.111144,7.435844,8.597813,9.261794,8.967529,9.009028,12.464753,9.631512,7.8923316,7.6207023,7.6282477,5.168496,9.971047,11.84227,10.616167,8.45068,9.80128,12.181807,9.759781,7.4999785,7.99042,11.442371,13.068373,14.086982,14.6151495,13.88326,10.227587,7.7376537,7.8131065,6.779407,5.7909794,10.812344,10.70671,9.046755,7.6508837,7.092535,6.6850915,13.539951,13.630494,10.978339,9.186342,11.472552,10.63503,7.3075747,5.5457587,5.915476,5.4703064,5.987156,5.745708,7.118943,9.239159,7.986647,7.77538,8.643084,8.586494,7.4697976,7.0284004,5.13077,4.1310244,4.2819295,4.881777,4.266839,3.904667,4.183841,4.5309224,4.7648253,5.1043615,5.624984,6.2436943,7.069899,8.080963,9.133525,9.646602,9.759781,9.0957985,8.213005,8.597813,7.756517,7.598067,8.296002,9.291975,9.303293,9.827688,9.193887,8.76758,8.733627,8.096053,7.3490734,7.122716,6.620957,5.5457587,4.115934,4.191386,4.4705606,5.0553174,5.6023483,5.3269467,6.187105,7.17176,7.7640624,7.77538,7.333983,7.4811153,7.726336,8.473316,9.718282,11.034928,11.102836,11.18206,10.374719,8.990166,8.533678,8.707218,8.903395,8.959985,8.643084,7.6584287,7.6093845,7.220804,7.0472636,7.635793,9.533423,11.642321,12.73261,12.472299,11.102836,9.465516,8.669493,7.492433,6.488915,5.6287565,4.29702,3.9386206,4.304565,4.727099,4.908185,4.930821,4.3422914,3.7801702,3.7386713,4.274384,4.9760923,4.4894238,5.010046,5.8966126,6.549277,6.4247804,5.5382137,5.50426,5.8966126,6.470052,7.1566696,7.6131573,7.748972,7.9338303,8.141325,7.9489207,7.8621507,6.7831798,6.0211096,5.934339,5.9418845,6.7680893,7.3905725,7.9451485,8.107371,7.115171,6.3229194,6.790725,7.0849895,6.8963585,7.0585814,7.594294,7.356619,7.2094865,7.4282985,7.6848373,6.8359966,7.2396674,7.564113,7.6131573,8.314865,8.669493,9.480607,10.54826,11.521597,11.91395,12.034674,11.714001,11.438599,11.389555,11.46878,10.529396,9.714509,8.571404,7.394345,7.213259,7.303802,7.0849895,6.228604,5.070408,4.5988297,4.610148,4.696918,5.3080835,6.0626082,5.7607985,5.643847,5.670255,5.4967146,5.138315,5.0062733,4.6856003,4.187614,4.115934,4.538468,4.979865,6.0022464,7.1981683,7.9791017,8.322411,8.756263,10.038955,10.774617,10.536942,9.601331,8.963757,8.82417,8.907167,9.276885,9.710737,9.688101,9.665465,9.703192,9.710737,9.461743,8.616675,7.3113475,7.118943,7.5301595,8.239413,9.129752,11.087745,13.6682205,14.464244,12.830698,9.880505,10.216269,11.838497,12.479843,11.710228,10.9594755,10.280403,12.076173,12.713746,12.6345215,12.566614,13.536179,13.328684,13.585222,14.743419,15.924251,14.962231,13.86817,12.970284,12.46098,12.268577,12.083718,12.151625,12.691111,13.117417,13.158916,12.868423,13.124963,12.626976,12.064855,11.627231,10.997202,11.559323,12.600568,12.932558,12.291212,11.351829,11.529142,12.079946,12.566614,12.562841,11.646093,11.155652,11.431054,11.4838705,11.068882,10.710483,11.11038,11.404645,11.619685,11.774363,11.883769,11.947904,11.883769,11.710228,11.581959,11.808316,11.9064045,12.528888,13.113645,13.449409,13.694629,13.909668,14.339747,14.385019,14.1058445,14.230342,14.27184,14.535924,14.796235,14.886778,14.720782,14.618922,14.392565,14.124708,13.79649,13.309821,13.996439,14.588741,14.543469,13.8719425,13.151371,13.50977,13.094781,12.559069,12.257258,12.257258,12.083718,12.223305,12.121444,11.570641,10.710483,10.842525,10.967021,11.140562,11.374464,11.604594,11.751727,11.7555,11.514051,11.129244,10.917976,10.736891,10.804798,11.072655,11.465008,11.868678,12.664702,13.053283,13.057055,12.743927,12.234623,11.955449,10.714255,9.273112,7.9791017,6.7944975,5.7796617,5.553304,5.304311,4.9459114,5.1345425,4.847823,4.779916,4.957229,5.300538,5.6325293,5.4967146,5.243949,5.081726,5.0854983,5.221313,5.4703064,5.5495315,5.73439,6.047518,6.270103,6.1908774,5.7192993,5.1458607,4.6214657,4.1574326,3.6443558,3.4481792,3.3764994,3.3689542,3.470815,3.8405323,4.006528,4.5309224,5.304311,5.5080323,5.3458095,5.111907,5.1081343,5.3382645,5.5193505,5.945657,6.1003346,6.2361493,6.628502,7.564113,7.7829256,8.024373,8.13378,7.9715567,7.405663,6.881268,6.9793563,7.2887115,7.7301087,8.533678,9.129752,9.367428,9.461743,9.333474,8.60913,8.371455,8.231868,8.107371,8.246958,9.235386,10.186088,11.227332,11.747954,11.604594,11.155652,10.20495,10.091772,10.216269,9.967276,8.733627,7.6584287,6.828451,6.258785,6.006019,6.149379,6.0286546,6.1342883,6.2097406,6.221059,6.375736,6.598321,6.436098,6.221059,6.187105,6.470052,6.6586833,6.6058664,6.8925858,7.779153,9.205205,9.6201935,9.58624,9.442881,9.2844305,8.959985,8.499724,8.20546,7.6093845,7.0170827,7.515069,8.047009,8.197914,8.054554,7.7187905,7.326438,7.533932,8.179051,8.873214,9.533423,10.382264,11.117926,11.59705,11.649866,11.083972,9.680555,8.265821,7.537705,7.2358947,7.3151197,7.9451485,9.446653,11.46878,12.921241,13.370183,12.996693,14.279386,16.531643,18.572634,18.621677,14.298248,13.158916,11.476325,10.186088,9.0807085,6.832224,7.1906233,5.9117036,3.519859,1.5052774,2.354118,1.9693103,3.4368613,4.055572,3.180323,2.2371666,2.2258487,1.8599042,2.3767538,3.8556228,5.2062225,5.670255,4.9119577,4.7912335,6.820906,12.178034,9.2995205,8.446907,8.412953,8.820397,10.121953,14.124708,14.554788,13.690856,12.853333,12.366665,11.570641,10.7218,10.103089,9.567377,8.537451,8.473316,7.6810646,7.8432875,9.005256,9.574923,10.386037,10.906659,10.714255,10.18986,10.49167,9.4013815,9.114662,8.60913,7.360391,5.342037,3.5236318,2.535204,1.4335974,0.6111652,1.8146327,4.3196554,4.67051,3.7990334,4.587512,11.891314,11.959221,10.70671,8.322411,5.5193505,3.5500402,4.247976,7.779153,9.940866,10.676529,14.079436,8.322411,5.4174895,4.014073,3.772625,5.342037,15.128226,22.688566,19.481836,9.073163,7.115171,7.5565677,3.7537618,1.7089992,2.4823873,2.1956677,2.2220762,3.2029586,3.9122121,4.085753,4.432834,4.3913355,4.8327327,4.745962,4.2027044,4.3422914,5.4212623,5.3571277,5.032682,5.160951,6.2889657,6.911449,7.3000293,7.7376537,8.182823,8.280911,8.537451,8.605357,8.790216,9.276885,10.170997,9.997457,9.967276,11.619685,14.1926155,14.66042,15.0376835,15.24895,15.39231,15.954432,17.818108,17.991648,18.346275,18.26705,17.444618,15.882751,14.011529,12.755245,12.193124,12.804289,15.460217,15.607349,14.392565,13.498452,13.472044,13.743673,13.517315,13.611631,13.547497,13.011784,11.857361,11.574413,12.106354,13.057055,14.045483,14.705692,15.490398,15.1395445,14.064346,12.668475,11.348056,10.982111,10.838752,10.95193,11.310329,11.891314,13.075918,14.302021,14.524607,13.309821,10.861387,10.442626,10.435081,10.601076,10.997202,11.978085,13.766309,14.2944765,13.962485,12.645839,9.710737,7.5188417,7.6018395,8.597813,9.7220545,10.751981,9.273112,8.514814,8.314865,8.111144,6.9189944,7.224577,7.3113475,8.024373,9.5032425,11.174516,12.242168,12.0233555,11.5857315,11.25374,10.623712,10.657665,11.7555,12.551523,13.109872,14.93205,12.860879,9.752235,7.7150183,7.224577,7.1264887,7.7640624,7.7376537,7.647111,8.231868,10.3634,10.970794,10.401127,10.125726,9.469289,5.6363015,8.024373,8.631766,7.201941,5.1345425,5.462761,8.231868,7.5037513,5.907931,5.6589375,8.544995,8.918486,9.989911,11.800771,13.27964,12.238396,6.8963585,6.1078796,6.1606965,6.379509,9.103344,10.940613,8.182823,6.0701537,6.006019,5.5306683,13.441863,16.22606,15.049001,13.053283,15.343266,15.516807,8.820397,4.870459,5.6778007,5.6363015,5.9117036,5.7872066,6.7379084,8.265821,7.877241,8.518587,9.4013815,8.526133,6.537959,6.7039547,5.402399,4.67051,4.727099,5.0175915,4.2064767,3.92353,3.802806,4.0593443,4.745962,5.7570257,5.7796617,6.3153744,7.0963078,8.050782,9.288202,10.242677,10.38981,9.714509,8.718536,8.431817,7.9451485,7.6810646,8.039464,8.733627,8.793989,9.382519,8.959985,8.880759,9.26934,8.993938,8.45068,8.122461,7.232122,5.723072,4.244203,4.4818783,5.1798143,5.764571,5.885295,5.3948536,6.092789,6.7944975,7.24344,7.383027,7.356619,7.3981175,7.6923823,8.511042,9.865415,11.517824,11.261286,11.355601,10.684074,9.258021,8.246958,8.29223,8.518587,8.820397,8.620448,6.858632,7.6395655,7.5565677,7.1793056,7.3075747,8.967529,10.272858,11.310329,11.287694,10.235131,9.020347,9.122208,8.612903,7.786698,6.7567716,5.451443,4.6629643,4.5196047,4.7120085,5.028909,5.3269467,4.6327834,3.9763467,3.712263,4.0706625,5.149633,5.0515447,5.3759904,6.096562,6.8397694,6.900131,6.4511886,6.2135134,6.228604,6.477597,6.8699503,7.5226145,7.828197,7.9338303,7.884786,7.6093845,7.707473,6.8850408,6.187105,5.9796104,5.9796104,6.5002327,6.9755836,7.54525,7.752744,6.541732,6.375736,7.1302614,7.598067,7.484888,7.435844,7.798016,7.7678347,7.647111,7.586749,7.5565677,7.281166,7.1302614,7.0812173,7.2358947,7.8508325,8.080963,9.144843,10.419991,11.348056,11.46878,11.517824,11.00852,10.812344,11.099063,11.351829,10.084227,9.4127,8.461998,7.232122,6.609639,7.069899,7.111398,6.5002327,5.4401255,4.5912848,4.285702,4.485651,5.089271,5.6363015,5.311856,5.406172,5.5080323,5.5382137,5.4967146,5.4665337,4.98741,4.67051,4.7308717,5.05909,5.2175403,5.243949,6.205968,7.1868505,7.7338815,7.8508325,8.869441,10.502988,11.155652,10.299266,8.488406,8.284684,8.461998,8.6732645,8.756263,8.729855,9.167479,9.329701,9.288202,9.06939,8.6732645,7.986647,7.7187905,7.654656,7.84706,8.612903,10.695392,12.770335,12.551523,10.303039,8.83926,10.26154,13.075918,13.951167,12.555296,11.551778,10.419991,11.917723,12.649611,12.774108,12.751472,13.340002,13.487134,14.1926155,15.188588,15.984612,15.8676605,14.400109,13.570132,12.970284,12.464753,12.181807,12.098808,12.506252,13.04951,13.502225,13.743673,13.347548,13.008011,12.510024,11.766817,10.819888,10.876478,12.423254,13.106099,12.366665,11.457462,11.751727,12.257258,12.645839,12.668475,12.151625,11.69891,12.196897,12.359119,11.921495,11.646093,12.913695,13.27964,13.328684,13.479589,13.943622,14.049255,13.985121,13.826671,13.543724,13.026875,12.649611,13.445636,14.385019,14.905642,14.924504,15.297995,15.856343,15.878979,15.497944,15.682802,15.671484,15.920478,16.218515,16.222288,15.445127,14.694374,14.769827,14.803781,14.543469,14.369928,15.467763,15.403628,14.569878,13.792717,14.286931,13.849306,13.189097,12.623203,12.347801,12.464753,12.249713,12.136535,11.589504,10.763299,10.518079,10.646348,10.714255,10.665211,10.567122,10.623712,10.514306,10.9594755,11.249968,11.155652,10.906659,11.034928,11.016065,11.249968,11.823407,12.487389,12.706201,12.842015,12.774108,12.393073,11.570641,10.789707,9.408927,7.858378,6.4549613,5.3948536,4.564876,4.217795,3.8895764,3.640583,4.08198,3.7198083,3.6971724,3.85185,4.0970707,4.436607,4.5497856,4.104616,3.7877154,3.772625,3.6971724,4.0291634,4.2630663,4.4705606,4.6554193,4.7346444,5.040227,4.7572803,4.304565,3.8782585,3.482133,2.746471,2.5314314,2.6823363,3.0369632,3.410453,3.8443048,3.9159849,4.564876,5.6815734,6.1342883,5.6476197,5.0213637,4.8402777,5.13077,5.3571277,5.624984,5.5495315,5.6287565,6.0362,6.6247296,7.4282985,7.756517,8.001738,8.058327,7.322665,6.9227667,6.700182,6.677546,7.032173,8.107371,8.7751255,8.967529,8.865668,8.571404,8.07719,7.3981175,7.432071,7.375482,7.2472124,7.907422,8.710991,10.431308,11.570641,11.559323,10.736891,9.405154,9.42779,9.669238,9.522105,8.888305,7.4018903,6.349328,5.8588867,5.8173876,5.8702044,5.8928404,5.9909286,6.19465,6.470052,6.719045,6.771862,6.247467,5.7683434,5.6551647,5.9117036,6.549277,6.730363,7.4282985,8.756263,9.97482,10.072908,9.710737,8.922258,8.167733,8.314865,7.61693,7.745199,7.677292,7.333983,7.5792036,8.526133,8.797762,8.835487,8.820397,8.66572,8.578949,8.582722,8.801534,9.26934,9.9257765,10.884023,11.2650585,11.623458,11.623458,10.061591,8.643084,7.752744,7.1793056,7.043491,7.7904706,9.533423,11.283921,12.804289,13.819125,14.000212,14.592513,16.84477,18.968758,19.029121,14.950912,13.773854,12.913695,11.438599,9.224068,6.94163,6.368191,4.093298,2.022127,1.6373192,4.0216184,2.6295197,2.3956168,3.8254418,5.5683947,4.432834,4.168751,4.093298,5.4288073,7.6131573,8.299775,6.5945487,5.1232247,5.59103,7.541477,8.360137,9.967276,10.514306,11.529142,12.6345215,11.521597,12.642066,13.158916,13.087236,12.487389,11.476325,10.899114,10.646348,10.518079,9.865415,7.594294,8.069645,7.4509344,8.00551,9.831461,10.880251,11.691365,12.276122,12.272349,11.974312,12.366665,9.88805,9.454198,8.809079,6.952948,4.1612053,3.108643,3.1840954,2.252257,0.5470306,0.6790725,4.044254,4.45547,3.0520537,3.6254926,12.604341,13.4644985,11.581959,7.032173,2.463524,3.0822346,2.3428001,4.2064767,7.488661,11.212241,14.600059,7.01331,4.266839,3.4594972,3.5123138,5.1647234,15.539442,22.130219,19.549744,11.09529,8.733627,5.723072,2.6106565,1.4109617,1.9994912,2.0900342,2.9539654,3.308592,3.7084904,4.327201,4.9421387,4.142342,5.0439997,5.458988,4.9345937,4.745962,5.1269975,5.0779533,4.719554,4.5988297,5.6778007,6.4021444,6.6247296,7.0284004,7.6093845,7.6886096,8.2507305,8.36391,8.843033,9.903141,11.170743,10.661438,10.355856,11.23865,12.947649,13.792717,14.505743,16.078928,16.795727,16.735365,17.757746,17.652113,17.829426,17.440845,16.697638,16.859861,15.101818,13.815352,13.087236,13.513543,16.195879,16.252468,14.2944765,13.317367,13.822898,13.822898,13.000465,12.921241,13.166461,13.272095,12.713746,12.189351,13.275867,14.954685,16.143063,15.686575,16.28265,15.935568,14.596286,12.706201,11.197151,11.106608,10.831206,10.695392,10.933067,11.676274,13.223051,14.460471,14.260523,12.113899,8.145098,8.465771,9.563604,10.27663,10.570895,11.555551,12.536433,12.774108,12.50248,11.317875,8.156415,6.964266,7.798016,9.031664,10.155907,11.778135,10.159679,9.49947,9.835234,9.937095,7.2924843,8.258276,8.816625,8.975075,9.0957985,9.918231,10.0276375,10.521852,10.963248,10.95193,10.121953,9.4127,10.186088,11.091517,12.321393,15.614895,12.947649,8.552541,6.1305156,6.349328,6.858632,7.6584287,7.8961043,9.133525,10.1294985,6.8171334,9.035437,10.887795,11.993175,11.857361,9.880505,5.05909,4.5799665,4.3875628,3.8707132,5.881522,3.7877154,3.5160866,3.4934506,3.5500402,4.8930945,5.945657,6.187105,7.605612,10.872705,15.354584,8.439363,5.723072,5.9230213,7.232122,7.284939,9.714509,7.9941926,4.9685473,3.3878171,5.915476,8.07719,15.260268,17.36162,13.487134,11.966766,15.739391,9.5183325,4.9044123,5.2854476,5.828706,6.187105,5.907931,5.221313,4.817642,5.8513412,7.284939,7.435844,6.485142,5.3684454,5.7909794,5.692891,5.5268955,5.451443,5.3571277,4.8930945,4.22534,3.9084394,4.13857,4.878004,5.8400235,5.934339,6.851087,7.6810646,8.265821,9.201432,10.084227,10.4049,9.989911,8.98262,7.8319697,8.179051,7.937603,7.726336,7.84706,8.265821,9.14107,9.5032425,9.861642,10.208723,10.023865,9.439108,8.975075,7.865923,6.1720147,4.7535076,4.9119577,6.009792,6.4926877,6.085244,5.772116,6.1908774,6.6058664,6.779407,6.862405,7.3717093,7.356619,7.484888,8.224322,9.688101,11.619685,11.404645,11.151879,10.502988,9.457971,8.371455,8.103599,7.752744,7.888559,7.956466,6.25124,7.0548086,7.8206515,7.937603,7.726336,8.424272,9.6051035,9.944639,9.608876,8.8618965,8.047009,8.68081,9.208978,8.941121,7.8923316,6.8058157,5.8400235,5.3986263,5.281675,5.3156285,5.3759904,4.9949555,4.587512,4.3724723,4.568649,5.406172,5.836251,5.9532022,6.462507,7.232122,7.277394,7.3679366,7.039718,6.72659,6.6020937,6.617184,7.5716586,7.809334,7.6395655,7.375482,7.326438,7.424526,7.3868,6.971811,6.3229194,5.9796104,6.19465,6.8058157,7.356619,7.3151197,6.096562,6.643593,7.567886,8.194141,8.303548,8.137552,8.386545,8.560086,8.29223,7.654656,7.1679873,7.858378,7.2924843,7.1264887,7.7187905,8.122461,7.1076255,8.20546,9.903141,10.997202,10.585986,10.695392,10.751981,10.917976,11.212241,11.54046,10.687846,9.963503,8.926031,7.5905213,6.4511886,7.043491,7.115171,6.790725,6.092789,4.9119577,4.1762958,4.1498876,4.61392,5.0854983,4.8138695,4.878004,4.8553686,5.036454,5.402399,5.6098933,5.062863,5.1647234,5.3080835,5.2250857,4.9723196,4.5912848,5.243949,6.2889657,7.1000805,7.062354,7.145352,9.163706,10.650121,10.235131,7.6810646,7.699928,8.420499,8.631766,8.111144,7.6395655,8.511042,9.239159,9.352338,9.024119,9.050528,8.718536,8.201687,7.5301595,7.175533,8.035691,9.808825,11.23865,11.016065,9.680555,9.654147,11.45369,14.109617,14.920732,13.675766,12.642066,9.246704,11.9064045,12.574159,12.121444,11.7894535,13.170234,15.131999,14.754736,13.773854,13.449409,14.57365,14.32843,14.139798,14.169979,14.158662,13.426772,13.060828,12.540206,12.4307995,12.940104,13.917213,12.902377,12.706201,12.5326605,12.079946,11.506506,11.102836,10.680302,10.838752,11.566868,12.238396,11.955449,12.242168,12.287439,12.2270775,13.151371,13.713491,14.422746,14.403882,13.830443,13.917213,14.50197,15.022593,15.384765,15.580941,15.701665,16.324148,16.214743,15.437581,14.249205,13.075918,13.283413,13.645585,14.117163,14.7321005,15.611122,16.060064,17.172989,17.463482,16.769318,16.218515,15.535669,15.99593,16.437326,16.31283,15.701665,15.614895,15.339493,14.781145,13.8719425,12.528888,12.113899,12.128989,12.321393,12.615658,13.091009,12.849561,12.67602,12.498707,12.381755,12.528888,12.759018,11.691365,10.295494,9.397609,9.688101,9.933322,10.103089,10.072908,10.012547,10.38981,11.012292,11.442371,11.638548,11.615912,11.442371,11.348056,10.480352,10.174769,10.691619,11.231105,11.400873,11.800771,12.423254,12.830698,12.14408,10.827434,8.7751255,6.7379084,5.1156793,3.9688015,3.6141748,3.3161373,3.1312788,3.078462,3.127506,2.9313297,2.6823363,2.5729303,2.6182017,2.655928,2.8256962,2.7313805,2.6219745,2.6332922,2.7917426,2.8521044,3.059599,3.2972744,3.5387223,3.8292143,4.134797,3.9650288,3.4745877,2.9464202,2.7615614,2.4559789,2.6182017,2.71629,2.7615614,3.3123648,3.8254418,3.9989824,4.376245,4.949684,5.1571784,4.4743333,4.606375,4.8327327,4.821415,4.640329,4.798779,5.0741806,5.4476705,5.855114,6.2097406,7.1981683,7.8319697,8.009283,7.7376537,7.141579,7.092535,6.722818,6.307829,6.092789,6.2851934,7.1038527,7.967784,8.469543,8.311093,7.3075747,6.2097406,5.7796617,6.2927384,7.333983,7.798016,8.835487,9.955957,10.804798,11.053791,10.4049,9.465516,9.359882,9.231613,8.805306,8.379,7.2283497,6.620957,6.519096,6.587003,6.2097406,5.6476197,5.7570257,6.1418333,6.4511886,6.379509,5.2175403,5.2779026,5.772116,6.2889657,6.790725,7.7414265,7.643338,8.0206,8.816625,8.379,8.216777,7.7112455,7.443389,7.5716586,7.828197,8.29223,8.345046,8.375228,8.4544525,8.345046,8.503497,8.635539,9.020347,9.431562,9.14107,8.567632,8.14887,8.197914,8.66572,9.156161,10.340765,11.314102,11.827179,11.879996,11.732863,10.159679,8.8769865,7.673519,6.971811,7.828197,10.099318,11.442371,12.042219,12.438345,13.551269,13.721037,15.282904,17.354074,18.440592,16.463736,13.902123,13.023102,11.879996,9.420244,5.4778514,5.040227,2.897376,1.7127718,2.3126192,3.6934,3.4594972,3.218049,5.2137675,7.828197,5.5683947,6.398372,6.149379,5.8211603,5.994701,6.8359966,6.5568223,6.8699503,8.601585,10.785934,10.665211,12.313848,12.815607,13.487134,14.132254,13.045737,11.827179,12.811834,12.951422,11.955449,12.283667,11.246195,10.555805,9.989911,9.220296,7.828197,8.341274,8.744945,9.556059,10.842525,12.223305,15.101818,16.060064,15.445127,14.305794,14.403882,11.389555,9.884277,8.262049,6.1003346,4.195159,2.2560298,2.2560298,1.7014539,0.39989826,0.47157812,3.572676,5.594803,4.3196554,2.5314314,8.028146,4.327201,2.2409391,2.4672968,5.3646727,10.955703,6.8774953,7.194396,10.887795,15.430037,16.784409,9.763554,6.6850915,5.0666356,4.1762958,5.0062733,10.20495,13.034419,13.298503,10.480352,3.7537618,2.3616633,1.3166461,1.3128735,2.04099,2.2107582,2.625747,3.500996,4.3800178,4.979865,5.1873593,5.028909,6.0776987,7.1604424,7.2472124,5.4778514,5.100589,4.9685473,4.938366,5.0779533,5.6778007,6.617184,6.477597,6.3417826,6.5040054,6.4549613,7.213259,7.9791017,8.296002,8.537451,9.903141,11.45369,11.940358,11.857361,11.793225,12.449662,12.89106,15.131999,16.867407,17.244669,16.890041,17.293713,17.45971,16.935314,15.848798,14.909414,14.652876,14.351066,13.472044,12.581704,13.35132,14.803781,14.460471,14.286931,14.483108,13.521088,13.215506,13.358865,14.030393,14.826416,14.86037,14.252977,16.260014,18.304777,18.470772,15.501716,14.245432,14.151116,14.000212,13.332457,12.464753,12.50248,12.091263,12.370438,13.200415,13.151371,12.577931,12.306303,11.544232,9.952185,7.643338,7.779153,7.9225125,8.265821,8.9788475,10.223814,9.186342,8.843033,8.635539,8.13378,7.0359454,6.349328,6.930312,7.748972,8.703445,10.61994,10.582213,10.646348,11.6008215,12.151625,8.941121,9.955957,10.446399,10.103089,9.405154,9.612649,9.967276,11.363147,12.47607,12.381755,10.574668,8.8769865,9.186342,9.9257765,10.816116,12.879742,13.758763,11.751727,9.205205,7.54525,7.2623034,7.9338303,9.273112,9.786189,9.050528,7.7225633,6.013564,8.265821,11.989402,13.909668,9.978593,8.428044,5.3759904,3.4745877,4.719554,10.484125,4.2706113,4.1083884,7.7640624,10.469034,4.927048,8.590267,9.616421,10.744436,13.373956,17.56157,14.011529,8.197914,6.2323766,8.333729,8.835487,8.186596,11.046246,9.318384,5.4401255,12.37421,8.967529,8.043237,6.752999,5.2175403,6.5455046,6.462507,5.560849,4.881777,5.1081343,6.560595,6.9755836,6.1908774,5.251494,4.666737,4.4101987,4.496969,5.1760416,5.3458095,4.927048,4.851596,5.1345425,5.6061206,6.0512905,6.224831,5.8588867,4.749735,4.7535076,4.889322,4.8025517,4.7912335,5.1571784,6.907676,7.7376537,7.4207535,7.798016,9.239159,9.359882,9.408927,9.567377,8.956212,9.273112,8.428044,7.647111,7.726336,9.031664,9.363655,10.057818,10.167224,9.6051035,9.156161,9.167479,8.748717,7.8508325,6.696409,5.7683434,5.4250345,5.4703064,5.553304,5.7570257,6.5756855,6.2361493,6.488915,6.903904,7.322665,7.8734684,7.605612,7.273621,7.4811153,8.326183,9.4013815,10.510533,10.899114,10.661438,9.812597,8.284684,8.311093,7.4471617,6.94163,6.911449,6.3644185,6.0814714,6.8171334,7.696155,8.375228,9.031664,10.7557535,10.03141,8.967529,8.439363,8.073418,7.277394,8.68081,9.559832,8.854351,7.17176,6.19465,5.915476,5.7117543,5.3382645,4.8968673,4.749735,5.1458607,5.6098933,5.8702044,5.8437963,6.3455553,6.617184,7.3113475,8.156415,7.9489207,7.914967,7.8017883,7.564113,7.164215,6.590776,7.567886,7.6923823,7.0849895,6.3153744,6.4247804,6.670001,7.224577,7.194396,6.5756855,6.270103,6.466279,6.560595,6.8925858,7.194396,6.620957,7.145352,7.752744,7.9791017,7.9036493,8.14887,9.001483,9.307066,8.695901,7.6207023,7.3377557,8.3525915,8.009283,7.54525,7.586749,8.14887,8.488406,8.922258,9.771099,10.710483,10.7557535,10.514306,10.763299,10.997202,11.212241,11.932813,11.857361,10.944386,9.510788,8.001738,6.9869013,7.564113,7.643338,7.54525,7.352846,6.911449,5.300538,4.61392,4.7120085,5.0477724,4.67051,5.1345425,5.342037,5.523123,5.6325293,5.342037,5.05909,5.723072,5.9796104,5.5193505,5.081726,5.3269467,5.4703064,6.013564,6.8435416,7.232122,7.2094865,8.631766,9.869187,9.58624,6.730363,6.5832305,7.635793,8.318638,8.224322,8.103599,8.273367,8.91094,9.088254,8.526133,7.598067,8.477088,7.9828744,7.24344,7.1679873,8.439363,10.072908,11.434827,12.14408,12.14408,11.717773,12.562841,13.970031,14.245432,13.328684,12.800517,9.967276,11.69891,11.121698,10.374719,10.725573,12.581704,12.966512,13.230596,13.336229,13.86817,16.026112,14.969776,14.373701,14.169979,13.985121,13.13628,12.943876,12.555296,12.3289385,12.3289385,12.3289385,12.381755,12.242168,12.166716,12.2119875,12.272349,11.208468,11.000975,11.302785,11.7555,12.019584,11.796998,11.849815,12.064855,12.626976,13.996439,14.664193,15.011275,15.16218,15.350811,15.894069,16.165699,16.807045,17.067356,16.795727,16.471281,16.029884,15.271586,14.403882,13.498452,12.50248,12.593022,12.898605,13.687083,14.822643,15.769572,16.131744,16.569368,16.437326,15.743164,15.147089,15.528125,15.543215,15.490398,15.343266,14.7736,14.611377,14.211478,13.781399,13.087236,11.442371,11.415963,11.099063,11.16697,11.506506,11.212241,11.272603,10.963248,11.1782875,11.774363,11.5857315,11.438599,10.401127,9.601331,9.473062,9.725827,9.7069645,10.303039,10.876478,11.193378,11.404645,12.045992,12.128989,11.872451,11.431054,10.906659,10.985884,10.895341,11.18206,11.819634,12.23085,12.694883,12.510024,11.910177,10.925522,9.363655,7.624475,5.9230213,4.8327327,4.191386,3.1010978,2.8558772,2.4559789,2.2296214,2.2220762,2.2107582,2.1843498,2.1956677,2.2786655,2.3993895,2.4484336,2.335255,2.2786655,2.2560298,2.233394,2.1579416,2.1013522,2.1315331,2.2975287,2.5314314,2.6597006,2.8558772,2.7011995,2.3616633,2.0447628,2.0183544,1.9957186,2.052308,2.033445,2.1353056,2.9086938,2.9124665,3.1048703,3.591539,4.1989317,4.4743333,4.5233774,4.5422406,4.564876,4.534695,4.3347464,4.5497856,4.7912335,4.8365054,4.851596,5.3910813,5.9532022,6.1531515,6.356873,6.6134114,6.688864,6.398372,6.039973,5.7909794,5.7494807,5.945657,5.934339,6.2436943,6.677546,6.851087,6.221059,6.217286,5.96452,6.258785,7.0548086,7.4811153,8.439363,9.673011,10.344538,10.220041,9.650374,8.76758,8.816625,8.880759,8.59404,8.107371,7.752744,7.394345,7.066127,6.802043,6.651138,6.3116016,6.0739264,5.8664317,5.6098933,5.2062225,5.119452,5.704209,6.4021444,7.0548086,7.877241,8.563859,9.371201,9.789962,9.7069645,9.416472,9.420244,8.76758,8.243186,8.024373,7.643338,8.088508,8.386545,8.597813,8.7600355,8.89585,8.126234,7.937603,8.0206,8.194141,8.409182,8.167733,8.269594,8.503497,8.756263,9.009028,9.352338,10.182315,10.850069,11.151879,11.317875,10.914205,10.272858,9.533423,9.0543,9.390063,10.431308,11.7026825,13.124963,14.392565,14.966003,15.086727,15.79598,15.912932,15.271586,14.7321005,13.015556,12.562841,12.4307995,11.4838705,8.371455,6.1342883,4.7308717,3.8367596,3.4972234,4.0970707,4.7308717,3.7914882,4.304565,6.149379,6.058836,6.19465,6.3116016,7.032173,8.360137,9.680555,8.186596,7.1000805,8.933576,12.491161,12.875969,11.057564,11.068882,12.030901,12.73261,11.604594,11.197151,12.310076,13.27964,13.245687,12.162943,11.69891,10.70671,10.702937,11.087745,9.159933,9.408927,9.993684,11.019837,12.657157,15.1395445,16.516552,16.207197,14.471789,12.068627,10.242677,11.932813,10.887795,8.111144,5.3646727,5.149633,3.108643,1.6146835,1.1883769,1.3996439,0.8262049,3.6141748,5.6589375,4.851596,2.323937,2.4484336,1.931584,1.9504471,2.8822856,5.1458607,9.224068,8.865668,11.204697,15.528125,18.904623,16.199652,10.095545,6.1041074,4.2592936,4.485651,6.56814,9.952185,9.507015,6.7756343,3.5839937,2.033445,1.0601076,0.65643674,1.0110635,1.81086,2.2371666,2.3880715,3.531177,4.557331,4.82896,4.187614,4.772371,6.40969,7.3000293,6.809588,5.4891696,5.6287565,5.2967653,4.9647746,5.0477724,5.907931,6.9152217,7.3415284,7.0510364,6.217286,5.3194013,5.753253,6.9680386,8.567632,10.057818,10.819888,11.781908,11.955449,11.52537,11.219787,12.3289385,12.936331,13.7700815,14.70192,15.380992,15.245177,16.407146,17.765291,18.534906,18.033148,15.675257,14.279386,13.317367,12.525115,11.978085,12.083718,13.973803,15.264041,15.878979,15.671484,14.422746,12.536433,11.84227,12.294985,13.347548,13.958713,16.999449,17.931286,17.852062,17.357847,16.52787,14.705692,14.520834,14.332202,13.890805,14.320885,15.011275,15.350811,15.347038,15.033911,14.445381,13.034419,12.340257,12.053536,11.627231,10.269085,10.238904,10.265312,10.540714,10.914205,10.917976,9.725827,8.809079,8.190369,7.8508325,7.7301087,7.2623034,7.696155,8.60913,9.986138,12.257258,13.204187,12.996693,11.947904,10.159679,7.5263867,9.133525,9.971047,9.997457,9.684328,10.0276375,9.952185,10.759526,11.551778,11.649866,10.574668,9.14107,9.273112,9.627739,9.6201935,9.435335,10.646348,10.812344,9.918231,8.458225,7.4471617,7.5603404,8.307321,9.058073,9.582467,10.0276375,9.265567,10.065364,12.555296,14.143571,9.525878,13.992666,9.250477,5.032682,7.907422,21.28515,14.1058445,9.337247,9.989911,12.879742,8.627994,7.9338303,7.9451485,9.235386,12.434572,18.221779,10.227587,6.700182,7.0246277,9.1976595,9.835234,6.8246784,6.741681,6.670001,6.511551,8.98262,9.491924,8.409182,7.066127,6.0512905,5.20245,4.9119577,4.5837393,4.908185,5.8664317,6.730363,6.3455553,6.0211096,5.5495315,4.9760923,4.5912848,4.5120597,5.0062733,5.221313,4.8968673,4.376245,4.636556,5.1269975,5.802297,6.319147,6.043745,5.0666356,5.028909,5.070408,4.8629136,4.606375,5.3458095,6.2135134,6.5756855,6.5530496,7.039718,8.179051,8.76758,9.363655,9.88805,9.627739,9.34102,8.477088,7.5490227,7.220804,8.314865,8.937348,9.982366,9.842778,8.722309,8.643084,8.235641,7.5792036,7.277394,7.3113475,7.0510364,6.326692,5.2326307,4.9044123,5.4174895,5.80607,5.621211,6.228604,6.688864,6.700182,6.617184,6.688864,6.2814207,5.4778514,4.696918,4.6742826,6.6850915,7.9791017,8.273367,7.7112455,6.8699503,7.284939,7.3113475,7.0849895,6.722818,6.2889657,5.9682927,6.862405,8.062099,8.831716,8.643084,10.450171,10.601076,9.839006,8.948667,8.718536,7.9828744,8.499724,8.986393,8.850578,8.22055,7.118943,6.477597,5.9230213,5.413717,5.2288585,4.6818275,5.040227,5.8400235,6.6058664,6.8435416,7.2283497,7.7187905,8.484633,9.163706,8.8769865,8.3525915,8.194141,8.27714,8.209232,7.322665,7.0887623,7.5112963,7.6207023,7.17176,6.6549106,6.2663302,6.477597,6.4964604,6.304056,6.673774,6.851087,6.7944975,7.111398,7.537705,6.9152217,7.605612,8.533678,8.907167,8.507269,7.696155,8.854351,10.574668,10.661438,9.016574,7.6320205,9.035437,10.008774,9.914458,8.907167,7.914967,8.590267,9.020347,9.544742,10.280403,11.099063,10.963248,11.23865,11.261286,11.174516,11.944131,12.438345,11.457462,9.906913,8.52236,7.8923316,8.213005,7.786698,7.4169807,7.3981175,7.533932,7.17176,6.5002327,6.1003346,5.9117036,5.2288585,5.587258,5.8928404,6.3116016,6.6247296,6.2436943,5.7683434,6.2135134,6.405917,5.983383,5.3986263,5.5268955,5.3684454,5.775889,6.741681,7.4169807,7.488661,8.254503,9.024119,9.092027,7.7301087,7.0170827,7.8131065,8.495952,8.59404,8.7751255,8.2507305,8.82417,9.310839,8.956212,7.4509344,8.0206,7.9300575,8.14887,9.099571,10.672756,10.559577,11.00852,11.18206,11.016065,11.193378,11.246195,11.578186,12.73261,14.245432,14.656648,9.81637,10.631257,10.54826,10.510533,11.174516,12.913695,12.796744,12.879742,13.200415,13.8719425,15.079182,14.750964,14.143571,13.630494,13.313594,13.008011,13.562587,13.513543,13.098554,12.653384,12.600568,11.717773,11.449917,11.815862,12.468526,12.706201,11.815862,11.646093,11.864905,12.098808,11.936585,11.581959,11.487643,11.781908,12.540206,13.804035,14.856597,15.347038,15.758255,16.218515,16.497688,15.603577,15.494171,15.47908,15.294222,15.124454,14.68683,14.2944765,13.932304,13.528633,12.936331,12.645839,12.728837,13.355092,14.317112,15.011275,15.565851,15.856343,15.603577,14.981093,14.611377,15.222542,15.23386,15.128226,14.9358225,14.249205,14.071891,13.622949,12.985375,12.027128,10.408672,10.253995,10.272858,10.242677,10.170997,10.321902,10.155907,10.1294985,10.303039,10.570895,10.638803,10.246449,9.944639,9.714509,9.627739,9.827688,9.9257765,10.412445,10.914205,11.291467,11.668729,11.721546,11.536687,11.102836,10.582213,10.325675,10.718028,11.257513,11.668729,12.027128,12.766563,13.302276,12.996693,12.049765,10.616167,8.812852,6.9265394,5.745708,4.7912335,3.7801702,2.6182017,2.2069857,2.04099,2.0183544,2.0372176,1.9844007,1.9579924,1.961765,1.9994912,2.0598533,2.093807,1.991946,2.0145817,2.0372176,1.9881734,1.8523588,1.7580433,1.7240896,1.7580433,1.8221779,1.8448136,1.9353566,1.7052265,1.4449154,1.3166461,1.3355093,1.5543215,1.5769572,1.6222287,1.841041,2.3126192,2.323937,2.6898816,3.2105038,3.6934,3.9725742,4.3649273,4.406426,4.496969,4.6252384,4.3686996,4.534695,4.678055,4.7120085,4.727099,4.9760923,5.149633,5.3080835,5.4665337,5.624984,5.7419353,5.4250345,5.2288585,5.149633,5.2326307,5.5759397,5.7306175,5.96452,6.115425,6.149379,6.1531515,6.3832817,6.519096,6.971811,7.605612,7.7225633,8.469543,8.967529,9.386291,9.6051035,9.239159,8.571404,8.771353,9.118435,9.133525,8.590267,8.197914,8.069645,7.907422,7.665974,7.54525,7.303802,6.7379084,6.432326,6.462507,6.4134626,6.9793563,7.8206515,8.182823,8.107371,8.439363,8.624221,9.0543,9.110889,8.873214,9.107117,9.039209,8.729855,8.431817,8.239413,8.084735,8.348819,8.122461,7.9413757,7.9828744,8.080963,8.326183,8.461998,8.52236,8.578949,8.737399,8.865668,9.25425,9.578695,9.684328,9.593785,9.201432,9.533423,9.918231,10.393582,11.69891,12.3289385,12.347801,11.91395,11.193378,10.374719,10.582213,11.16697,12.562841,14.237886,14.679284,13.879487,14.362384,13.773854,12.355347,12.943876,12.585477,12.928786,13.102326,12.14408,9.020347,6.760544,6.217286,5.9532022,5.353355,4.644101,5.2364035,4.8365054,5.040227,6.1305156,7.0963078,6.9944468,7.224577,7.809334,8.458225,8.578949,8.533678,8.529905,9.914458,12.015811,12.1101265,10.589758,10.427535,10.499215,10.359629,10.231359,10.197406,10.880251,11.578186,11.962994,12.076173,12.37421,11.419736,11.502733,12.08749,9.812597,9.835234,9.820143,10.861387,13.52486,17.863379,15.886524,15.007503,13.626721,11.45369,9.476834,11.721546,10.910432,8.122461,5.2854476,5.149633,4.0216184,2.3277097,1.3128735,1.1280149,0.80734175,1.9127209,3.4783602,3.5839937,2.1390784,0.8865669,2.082489,2.8596497,3.350091,4.346064,7.3075747,11.050018,15.350811,17.70493,16.625957,11.649866,8.458225,5.975838,5.0062733,5.8966126,8.52236,5.534441,3.9008942,2.335255,0.8526133,0.77716076,0.4376245,0.5093044,1.1016065,1.9730829,2.535204,2.9652832,3.6141748,4.214022,4.4818783,4.1197066,5.745708,7.4094353,7.303802,5.9117036,6.006019,5.915476,5.6476197,5.413717,5.4174895,5.855114,6.405917,7.462252,7.8131065,7.0548086,5.621211,6.0701537,7.4169807,9.322156,11.295239,12.706201,12.608112,11.978085,11.41219,11.25374,11.604594,12.66093,12.800517,13.083464,13.645585,13.705947,15.0905,17.101309,18.632996,18.614132,16.014793,14.053028,12.483616,11.732863,11.751727,12.019584,13.098554,13.894578,14.475562,14.875461,15.086727,12.642066,11.34051,11.864905,13.36641,13.456953,17.787928,18.417955,17.176762,15.958203,16.712729,15.143317,15.086727,14.924504,14.505743,15.150862,15.46399,15.871433,15.731846,14.984866,14.139798,12.619431,11.887542,11.638548,11.521597,11.144334,11.517824,12.178034,12.3289385,11.793225,11.019837,11.000975,10.842525,10.438853,10.0276375,10.155907,9.835234,9.835234,9.989911,10.661438,12.7477,13.9888935,13.573905,11.857361,9.540969,7.665974,9.26934,10.891568,11.61214,11.427281,11.249968,11.080199,10.601076,10.56335,10.997202,11.197151,10.861387,11.050018,11.076427,10.4049,8.646856,8.710991,9.322156,9.522105,9.009028,8.152642,8.390318,8.560086,9.26934,10.461489,11.41219,11.487643,12.50248,14.441608,16.180788,15.475307,15.505488,13.2607765,11.480098,17.05981,41.04239,41.053707,22.56407,9.552286,7.9715567,5.715527,7.4773426,6.960493,7.6207023,10.103089,12.234623,7.8810134,9.009028,9.280658,7.745199,8.850578,7.7187905,6.971811,7.1868505,8.213005,9.186342,8.529905,7.2358947,6.270103,5.783434,5.1232247,4.919503,4.606375,5.1156793,6.3945994,7.3717093,6.6020937,6.115425,5.6589375,5.304311,5.455216,4.847823,4.8553686,5.036454,4.9760923,4.266839,4.134797,4.7120085,5.4174895,5.7909794,5.511805,5.4665337,5.2967653,4.8930945,4.504514,4.7346444,5.4703064,5.704209,5.7796617,5.983383,6.549277,6.907676,7.3717093,8.031919,8.597813,8.412953,8.209232,8.341274,8.179051,7.6622014,7.3000293,8.473316,9.231613,8.741172,7.635793,8.0206,7.273621,6.8397694,6.971811,7.326438,6.9944468,6.851087,5.8664317,5.330719,5.4363527,5.2854476,5.3571277,5.511805,5.3910813,5.142088,5.406172,5.4174895,5.1345425,4.8742313,4.4177437,3.0181,3.7499893,4.98741,5.8098426,5.8588867,5.3269467,5.9984736,6.677546,7.020855,6.934085,6.5455046,6.398372,7.2585306,8.726082,9.940866,9.590013,9.989911,10.559577,10.272858,9.303293,9.027891,8.650629,8.458225,8.028146,7.4509344,7.303802,6.964266,6.692637,6.255012,5.7004366,5.3382645,4.9232755,4.851596,5.409944,6.4549613,7.3981175,8.028146,8.6581745,9.250477,9.522105,8.918486,8.254503,8.084735,8.239413,8.296002,7.5905213,7.2660756,7.699928,7.877241,7.5037513,7.0057645,6.598321,6.356873,6.1644692,6.119198,6.5455046,6.4738245,6.458734,6.9152217,7.575431,7.4811153,7.9941926,8.797762,8.933576,8.345046,7.8961043,8.703445,11.299012,12.340257,11.133017,9.627739,9.5032425,9.95973,10.382264,10.299266,9.348565,9.756008,10.023865,10.355856,10.887795,11.69891,11.974312,12.2119875,12.238396,12.313848,13.13628,13.611631,12.449662,10.880251,9.612649,8.850578,8.797762,8.688355,8.43559,8.254503,8.650629,8.89585,7.6923823,6.7077274,6.356873,5.828706,5.9984736,6.5568223,7.281166,7.654656,6.862405,6.198423,6.368191,6.560595,6.3531003,5.7079816,5.349582,5.1458607,5.5457587,6.4738245,7.3415284,8.084735,8.318638,8.511042,8.737399,8.684583,7.865923,8.299775,8.729855,8.873214,9.397609,9.114662,9.175024,9.276885,8.986393,7.7640624,7.665974,8.035691,9.148616,10.729345,11.955449,11.793225,11.668729,11.219787,10.582213,10.412445,10.359629,10.231359,11.16697,12.902377,13.739901,9.895596,9.839006,10.676529,10.982111,11.11038,13.185325,13.143826,13.057055,13.155144,13.505998,13.992666,14.32843,13.996439,13.385274,12.89106,12.921241,13.539951,13.626721,13.475817,13.275867,13.0646,11.257513,10.906659,11.502733,12.347801,12.551523,11.932813,11.793225,11.936585,12.136535,12.1252165,11.955449,11.729091,11.91395,12.66093,13.804035,15.015047,15.490398,15.829934,16.135517,16.003475,14.735873,14.151116,13.909668,13.879487,14.166207,13.909668,13.777626,13.604086,13.377728,13.223051,12.781653,13.0646,13.656902,14.25675,14.70192,15.060319,15.169725,15.015047,14.747191,14.7170105,14.999957,15.218769,15.218769,14.867915,14.060574,13.951167,13.894578,13.200415,11.812089,10.306811,10.03141,9.854096,9.703192,9.608876,9.703192,9.480607,9.457971,9.514561,9.529651,9.367428,9.393836,9.812597,9.922004,9.718282,9.876732,9.865415,10.197406,10.638803,11.053791,11.378237,11.449917,11.083972,10.631257,10.253995,9.95973,10.691619,11.461235,11.921495,12.276122,13.27964,13.536179,13.302276,12.355347,10.653893,8.345046,6.647365,5.462761,4.22534,2.886058,1.9278114,1.7240896,1.8749946,2.033445,2.0296721,1.8787673,1.9542197,1.9994912,2.0258996,2.0296721,1.9881734,2.0145817,2.0070364,1.9504471,1.8599042,1.81086,1.6486372,1.5505489,1.4977322,1.478869,1.4939595,1.5316857,1.2864652,1.0186088,0.84884065,0.7582976,0.9318384,1.0827434,1.2525115,1.4562333,1.6712729,1.931584,2.4182527,2.8558772,3.180323,3.5274043,4.0480266,4.183841,4.2819295,4.3611546,4.146115,4.395108,4.5233774,4.606375,4.6818275,4.7648253,4.6214657,4.7346444,4.8100967,4.8138695,4.961002,4.67051,4.6554193,4.7233267,4.8855495,5.3571277,5.666483,5.9796104,6.0626082,5.9909286,6.1531515,6.5756855,6.6662283,7.0472636,7.605612,7.5075235,8.069645,8.348819,8.699674,9.050528,8.869441,8.461998,8.741172,9.118435,9.231613,8.933576,8.560086,8.703445,8.786444,8.601585,8.322411,8.096053,7.4509344,7.2283497,7.4999785,7.54525,8.273367,9.084481,9.1825695,8.650629,8.439363,8.443134,8.386545,8.254503,8.254503,8.801534,8.605357,8.36391,8.401636,8.695901,8.846806,8.816625,8.307321,8.07719,8.288457,8.495952,9.231613,9.390063,9.261794,9.167479,9.431562,9.963503,10.978339,11.45369,11.197151,10.850069,10.152134,9.718282,9.797507,10.623712,12.415709,13.377728,13.472044,12.992921,12.012038,10.355856,10.050273,10.280403,11.283921,12.543978,12.762791,11.664956,11.868678,11.45369,10.495442,11.057564,11.947904,12.570387,12.728837,12.113899,10.325675,7.220804,6.858632,6.9189944,6.4210076,5.7192993,5.715527,6.224831,6.8133607,7.492433,8.729855,9.786189,9.242931,8.820397,8.933576,8.688355,9.446653,10.299266,10.7557535,10.552032,9.661693,10.378491,10.18986,9.631512,9.14107,9.076936,9.084481,9.250477,9.567377,10.201178,11.495189,12.442118,12.140307,12.068627,12.336484,11.680047,11.891314,10.540714,10.801025,13.6682205,17.980331,15.079182,14.124708,13.494679,12.287439,10.355856,11.234878,10.401127,8.337502,6.115425,5.3873086,4.5535583,2.957738,1.5241405,0.76584285,0.7696155,2.2598023,3.8254418,4.327201,3.6368105,2.625747,3.229367,3.0935526,2.987919,3.8556228,6.809588,13.460726,15.792209,14.822643,11.653639,7.4811153,6.4964604,6.6134114,7.122716,7.224577,6.017337,1.9051756,0.84884065,0.66775465,0.4376245,0.4979865,0.5470306,1.0186088,1.9127209,2.9049213,3.3463185,4.323428,4.164978,4.1272516,4.4818783,4.496969,6.6662283,8.288457,7.7904706,6.0701537,6.488915,6.1531515,6.006019,5.938112,5.9192486,6.009792,6.149379,7.194396,8.009283,7.9526935,6.8850408,7.032173,7.99042,9.4013815,11.034928,12.759018,12.555296,11.838497,11.570641,11.717773,11.2801485,11.570641,11.434827,11.61214,12.31762,13.230596,14.705692,16.927769,18.470772,18.651857,17.512526,15.516807,13.656902,12.736382,12.789199,13.053283,12.608112,12.2119875,12.359119,13.098554,14.015302,12.845788,12.034674,12.649611,14.007756,13.694629,17.999193,18.961214,17.157898,14.815099,15.833707,14.652876,14.634012,14.50197,14.154889,14.671739,15.011275,15.501716,15.629986,15.128226,13.985121,12.698656,12.193124,11.9064045,11.664956,11.664956,12.657157,12.808062,12.253486,11.3971,10.910432,12.034674,13.283413,13.306048,12.181807,11.41219,11.144334,11.099063,11.091517,11.431054,12.947649,13.377728,13.253232,12.351574,11.016065,10.193633,11.415963,13.045737,13.79649,13.211733,11.68382,12.362892,11.487643,11.034928,11.487643,11.84227,12.0082655,12.064855,11.974312,11.219787,8.820397,8.269594,8.537451,8.948667,9.076936,8.729855,8.8769865,9.020347,9.631512,10.767072,12.057309,12.147853,12.796744,15.569623,19.425245,20.730574,14.535924,14.622695,16.4411,21.636003,38.07333,37.564026,20.662666,9.129752,7.6207023,3.6896272,7.424526,7.496206,7.092535,7.6508837,8.854351,9.005256,13.128735,12.66093,8.084735,8.933576,8.948667,8.273367,8.382772,9.076936,8.465771,6.571913,5.775889,5.511805,5.3759904,5.1043615,5.0138187,4.7346444,5.2326307,6.541732,7.7678347,7.2660756,6.6586833,6.0512905,5.8173876,6.6020937,5.692891,5.2137675,5.168496,5.1043615,4.0782075,3.7348988,4.3800178,4.927048,4.98741,4.851596,5.2665844,5.221313,4.881777,4.640329,5.1156793,5.243949,5.643847,5.8098426,5.7494807,5.987156,6.175787,6.439871,6.670001,6.8397694,6.990674,6.628502,7.111398,7.798016,7.9753294,6.8435416,7.643338,7.752744,7.3679366,6.9982195,7.4697976,6.6020937,6.2361493,6.2361493,6.3832817,6.3832817,6.934085,6.1644692,5.523123,5.372218,4.991183,5.20245,4.425289,3.7462165,3.9348478,5.4401255,4.5535583,4.191386,4.768598,5.3458095,3.6330378,2.8445592,3.1161883,3.92353,4.5497856,4.063117,4.8930945,6.0324273,6.952948,7.405663,7.443389,7.537705,8.016829,9.265567,10.668983,10.61994,9.937095,10.431308,10.446399,9.691874,9.239159,8.865668,8.322411,7.352846,6.224831,5.753253,5.9909286,6.432326,6.590776,6.258785,5.485397,5.43258,5.300538,5.6513925,6.6058664,7.816879,8.733627,9.484379,9.778644,9.522105,8.782671,8.375228,8.262049,8.280911,8.235641,7.91874,7.8734684,8.069645,7.9338303,7.405663,6.937857,6.696409,6.33801,6.1418333,6.228604,6.5756855,6.417235,6.398372,6.7077274,7.281166,7.8131065,8.284684,8.831716,8.756263,8.175279,7.986647,8.375228,10.770844,12.076173,11.619685,11.140562,10.137043,9.49947,9.691874,10.419991,10.627484,10.801025,11.136789,11.52537,11.936585,12.423254,12.653384,12.638294,12.6345215,12.90615,13.70972,13.758763,12.751472,11.457462,10.329447,9.522105,9.250477,9.457971,9.408927,9.092027,9.231613,9.65792,8.390318,7.1793056,6.696409,6.519096,6.3116016,6.8473144,7.6923823,8.20546,7.5603404,6.779407,6.485142,6.349328,6.149379,5.7872066,5.2062225,4.8553686,5.1647234,6.1116524,7.2283497,8.231868,8.36391,8.3525915,8.499724,8.6732645,8.548768,8.922258,9.231613,9.476834,10.223814,10.435081,9.997457,9.5183325,9.129752,8.4544525,8.4544525,9.1825695,10.38981,11.642321,12.306303,12.068627,11.6875925,11.038701,10.26154,9.759781,9.903141,9.948412,10.502988,11.438599,11.891314,10.099318,9.612649,11.019837,11.295239,10.797253,13.29473,13.441863,13.272095,13.045737,13.091009,13.792717,13.992666,14.019074,13.619176,13.019329,12.928786,12.951422,13.026875,13.536179,14.0983,13.539951,11.823407,11.2801485,11.52537,12.049765,12.234623,11.668729,11.548005,11.710228,12.08749,12.73261,12.883514,12.657157,12.698656,13.283413,14.298248,15.147089,15.373446,15.433809,15.433809,15.128226,14.460471,13.981348,13.63804,13.592768,14.2077055,13.951167,13.675766,13.264549,12.89106,13.019329,12.792972,13.615403,14.392565,14.7321005,14.947141,14.815099,14.588741,14.626467,14.9358225,15.196134,14.84528,15.184815,15.147089,14.479335,13.754991,13.634267,14.083209,13.728582,12.355347,10.917976,10.695392,9.827688,9.537196,9.789962,9.307066,9.208978,8.854351,8.846806,8.9788475,8.231868,8.843033,9.457971,9.582467,9.363655,9.58624,9.137298,9.367428,9.827688,10.201178,10.27663,10.8576145,10.61994,10.408672,10.352083,9.839006,10.668983,11.261286,11.857361,12.638294,13.721037,13.70972,13.52486,12.540206,10.518079,7.598067,6.5228686,4.7912335,3.0331905,1.7014539,1.0902886,1.327964,1.629774,1.8259505,1.8334957,1.6486372,1.8863125,2.11267,2.2371666,2.2107582,2.0560806,2.173032,2.0296721,1.8485862,1.7618159,1.8221779,1.6373192,1.478869,1.418507,1.4562333,1.5505489,1.5807298,1.3770081,1.026154,0.6451189,0.362172,0.29426476,0.5696664,0.8111144,0.9318384,1.1242423,1.539231,1.9957186,2.2409391,2.4031622,3.0181,3.531177,3.8065786,3.8254418,3.6783094,3.591539,4.093298,4.247976,4.285702,4.353609,4.496969,4.2027044,4.1762958,4.2291126,4.3196554,4.5422406,4.3007927,4.4101987,4.5988297,4.8327327,5.3194013,5.511805,5.8098426,6.0814714,6.2097406,6.1078796,6.5530496,6.296511,6.360646,6.809588,6.7077274,7.2358947,7.9413757,8.390318,8.518587,8.661947,8.544995,8.7751255,8.884532,8.843033,9.0543,8.892077,9.152389,9.265567,9.042982,8.710991,8.661947,8.269594,8.141325,8.228095,7.809334,8.262049,8.899622,8.963757,8.443134,8.062099,8.386545,8.348819,8.288457,8.439363,8.929804,8.793989,8.59404,8.929804,9.673011,9.989911,9.808825,9.420244,9.390063,9.80128,10.269085,10.367173,9.997457,9.420244,9.107117,9.733373,10.419991,12.015811,12.687338,12.170488,11.785681,11.385782,10.574668,10.623712,11.725319,12.985375,13.604086,13.340002,12.691111,11.706455,9.989911,9.276885,9.639057,10.242677,10.582213,10.484125,9.895596,9.684328,9.650374,9.582467,9.25425,10.929295,11.299012,11.400873,11.69891,12.117672,7.8206515,6.911449,7.115171,7.3000293,7.488661,6.85486,7.575431,8.341274,9.058073,10.819888,13.849306,12.170488,10.412445,10.4049,11.193378,10.782163,11.004747,10.597303,9.25425,7.654656,10.559577,10.197406,9.631512,9.58624,8.461998,8.14887,8.035691,8.465771,9.476834,10.79348,11.676274,12.453435,12.464753,12.283667,13.721037,14.4152,12.091263,11.136789,12.702429,14.679284,14.02662,13.487134,13.483362,13.521088,12.223305,11.691365,10.284176,8.726082,7.3377557,6.006019,4.6252384,3.1350515,1.7844516,0.9242931,0.9997456,4.395108,6.33801,6.719045,5.9909286,5.194905,3.7952607,2.3578906,2.2447119,3.9084394,6.900131,14.600059,12.657157,9.771099,8.707218,6.2927384,5.3269467,7.4169807,8.89585,7.183078,0.7809334,1.116697,1.2298758,1.0525624,0.8337501,1.146878,1.267602,1.9994912,3.1539145,4.266839,4.6214657,5.5570765,4.8063245,4.5799665,5.172269,4.9987283,6.802043,8.254503,8.375228,7.488661,7.2472124,6.7756343,6.63982,6.643593,6.643593,6.5643673,6.700182,7.273621,8.031919,8.548768,8.22055,7.745199,8.09228,8.850578,9.820143,10.997202,11.61214,11.714001,12.019584,12.423254,12.0082655,10.782163,10.555805,11.016065,12.034674,13.634267,15.011275,16.735365,17.667202,17.980331,19.164934,18.116146,16.595778,15.116908,14.109617,13.917213,12.355347,11.348056,11.080199,11.415963,11.91395,12.96274,13.147598,13.656902,14.468017,14.324657,17.836971,19.074392,17.142809,14.000212,14.449154,13.604086,13.27964,13.174006,13.257004,13.800262,14.592513,15.143317,15.471535,15.294222,14.030393,13.336229,13.264549,13.204187,13.008011,12.974057,14.147344,13.264549,11.823407,10.827434,10.770844,12.162943,14.27184,14.705692,13.094781,11.087745,10.457717,10.714255,11.212241,11.785681,12.770335,12.321393,12.989148,13.521088,13.539951,13.505998,14.109617,14.84528,14.966003,13.902123,11.272603,12.958967,12.645839,12.457208,12.792972,12.325166,12.113899,11.895086,11.872451,11.54046,9.688101,9.159933,8.843033,8.639311,8.533678,8.586494,8.371455,8.98262,9.480607,9.929549,11.393328,11.32542,10.842525,14.947141,21.492645,21.156881,12.713746,13.234368,16.697638,19.240387,19.168707,9.718282,6.066381,9.314611,13.570132,5.9796104,8.654402,8.858124,7.2396674,6.2097406,9.940866,11.291467,15.169725,14.569878,10.106862,10.005001,9.175024,8.669493,8.801534,8.695901,6.307829,4.9534564,5.149633,5.4174895,5.1647234,4.7006907,4.749735,4.738417,5.2137675,6.270103,7.515069,7.7602897,7.3377557,6.620957,6.2814207,7.281166,6.4549613,5.7570257,5.43258,5.111907,3.8405323,3.4783602,3.9650288,4.221567,4.2102494,4.957229,4.7006907,4.8365054,4.859141,4.8365054,5.4363527,4.870459,5.907931,6.3832817,5.87775,5.7117543,5.9305663,6.1041074,5.904158,5.6363015,6.2361493,5.4665337,5.5004873,6.507778,7.647111,7.039718,6.617184,6.2851934,6.405917,6.820906,6.8774953,6.0362,5.553304,5.138315,5.0251365,5.994701,6.4021444,5.6023483,5.111907,5.142088,4.587512,4.4139714,2.9803739,2.3993895,3.4557245,5.6061206,3.85185,3.5424948,4.689373,6.4247804,7.001992,4.214022,3.1161883,3.4029078,4.13857,3.7462165,4.508287,5.847569,7.043491,7.84706,8.480861,8.835487,9.046755,9.767326,10.782163,10.989656,10.314357,10.559577,10.574668,10.035183,9.435335,8.790216,8.118689,7.0963078,5.783434,4.6290107,4.8402777,5.8928404,6.7114997,6.7454534,5.934339,6.0814714,6.3531003,6.7831798,7.3679366,8.043237,9.073163,9.978593,10.140816,9.590013,9.016574,9.024119,8.933576,8.707218,8.458225,8.420499,8.401636,8.171506,7.7187905,7.118943,6.530414,6.349328,6.1229706,6.126743,6.417235,6.7944975,6.952948,6.983129,6.960493,7.1000805,7.786698,8.303548,8.6581745,8.635539,8.2507305,7.7225633,7.8395147,9.382519,10.352083,10.480352,11.234878,10.770844,9.559832,8.926031,9.439108,10.887795,11.257513,11.910177,12.483616,12.811834,12.928786,12.789199,12.50248,12.494934,12.845788,13.317367,12.913695,12.393073,11.555551,10.555805,9.880505,9.756008,10.035183,10.050273,9.597558,8.933576,9.224068,8.552541,7.647111,7.0359454,7.0548086,6.507778,6.56814,7.2358947,8.054554,8.137552,7.4094353,6.7643166,6.1305156,5.6476197,5.6778007,5.2967653,4.708236,4.957229,6.126743,7.352846,7.937603,8.224322,8.405409,8.409182,7.8923316,8.843033,9.424017,9.793735,10.20495,11.02361,11.438599,10.661438,9.895596,9.57115,9.337247,9.835234,10.63503,11.423509,12.00072,12.279895,11.729091,11.336739,10.782163,10.057818,9.446653,9.793735,10.38981,10.853842,11.00852,10.899114,9.110889,9.367428,10.785934,12.030901,12.830698,13.977575,14.037937,13.192869,12.7477,13.20796,14.283158,13.660675,13.822898,13.879487,13.5663595,13.2607765,13.321139,13.7851715,14.705692,15.580941,15.335721,14.70192,13.324911,12.47607,12.50248,12.83447,12.245941,11.955449,12.14408,12.842015,13.917213,13.645585,13.8719425,14.109617,14.27184,14.664193,14.566105,14.796235,15.030138,15.101818,15.030138,14.626467,14.305794,13.936077,13.671993,13.977575,13.721037,13.400364,13.023102,12.725064,12.785426,12.932558,13.849306,14.652876,14.909414,14.618922,14.532151,14.109617,14.290704,15.064092,15.441354,14.354838,14.366156,13.81158,12.657157,12.498707,11.947904,11.974312,12.340257,12.370438,10.955703,10.770844,9.993684,9.556059,9.650374,9.733373,9.2844305,8.850578,8.741172,8.809079,8.4544525,8.318638,8.296002,8.09228,7.9262853,8.499724,7.6810646,7.594294,7.564113,7.443389,7.6131573,7.798016,8.401636,9.035437,9.495697,9.767326,10.008774,10.272858,11.034928,12.291212,13.551269,14.136025,13.841762,12.528888,10.4049,8.024373,8.122461,5.9607477,3.4330888,1.6260014,0.80734175,0.8337501,0.8299775,0.95824677,1.1959221,1.3430545,1.5015048,1.8787673,2.0749438,1.9730829,1.7391801,1.7882242,1.5618668,1.4600059,1.5430037,1.5430037,1.6373192,1.5165952,1.4675511,1.5882751,1.7693611,1.780679,1.5279131,1.0940613,0.6187105,0.29049212,0.19240387,0.1659955,0.32821837,0.6149379,0.80734175,0.87147635,1.1959221,1.1657411,1.1129243,2.335255,2.7011995,3.1312788,3.289729,3.1765501,3.127506,3.8858037,3.8820312,3.783943,3.8405323,3.874486,3.7650797,3.682082,3.953711,4.3686996,4.2102494,4.1762958,4.3309736,4.617693,4.9760923,5.3571277,5.6363015,5.643847,6.0211096,6.6662283,6.730363,5.983383,5.96452,6.0776987,6.085244,6.0739264,6.8171334,7.5263867,7.8734684,8.137552,9.186342,9.431562,9.473062,9.239159,9.065618,9.688101,9.310839,9.088254,8.741172,8.431817,8.7751255,9.446653,9.612649,9.540969,9.163706,8.103599,7.9791017,8.616675,8.575176,7.816879,7.7225633,8.646856,9.220296,9.092027,8.646856,9.001483,9.393836,10.499215,11.144334,11.268831,11.917723,12.196897,11.68382,10.955703,10.574668,11.0613365,10.623712,9.635284,8.60913,8.122461,8.820397,8.831716,9.623966,10.355856,10.627484,10.469034,11.004747,11.423509,11.891314,12.434572,12.925014,13.143826,13.008011,12.657157,12.064855,11.000975,9.646602,9.986138,10.412445,10.359629,10.299266,9.895596,9.669238,9.258021,8.605357,7.9338303,9.81637,10.27663,10.453944,10.812344,11.155652,8.858124,7.3868,8.424272,10.687846,9.918231,9.295748,8.243186,7.6584287,8.744945,13.030646,16.754227,15.275358,12.604341,11.461235,13.306048,10.412445,8.692128,8.526133,9.22784,9.031664,11.951676,10.819888,10.174769,10.623712,8.865668,7.7301087,7.7112455,8.967529,10.7218,11.246195,10.427535,12.098808,13.155144,12.683565,11.962994,12.804289,12.019584,10.740664,9.612649,8.7600355,10.725573,11.2801485,11.853588,13.223051,15.516807,15.067864,11.940358,9.190115,7.677292,6.1041074,4.515832,3.5689032,2.5804756,1.659955,1.7089992,3.9801195,5.5268955,6.205968,5.8664317,4.3649273,2.203213,1.9466745,2.886058,4.06689,4.2894745,11.442371,10.080454,10.9594755,14.128481,8.941121,5.534441,6.881268,7.069899,4.357382,1.1581959,2.3428001,2.173032,1.3355093,0.86770374,2.1353056,2.3088465,2.927557,3.8971217,5.0251365,6.0286546,4.878004,4.3724723,5.349582,6.719045,5.462761,5.975838,6.5530496,7.6886096,9.042982,9.446653,8.4544525,8.080963,8.088508,8.065872,7.432071,8.114917,8.82417,9.26934,9.186342,8.329956,7.5603404,7.8998766,8.914713,9.971047,10.238904,11.117926,12.106354,12.751472,13.181552,14.083209,13.034419,12.725064,13.13628,13.758763,13.611631,14.147344,14.034165,14.200161,15.23386,17.395575,19.191343,19.006485,16.376965,12.89106,12.208215,11.634775,11.69891,11.427281,10.985884,11.717773,13.355092,12.921241,13.011784,14.056801,14.313339,16.301512,16.535416,14.984866,13.12119,13.902123,13.619176,12.487389,12.438345,13.679539,14.679284,14.924504,14.747191,14.019074,13.057055,12.604341,13.275867,13.8719425,14.603831,15.414946,15.977067,15.939341,16.633503,15.46399,12.513797,10.574668,11.050018,11.717773,12.525115,12.796744,11.246195,9.26934,9.378746,9.763554,10.023865,11.170743,12.257258,13.781399,14.551015,14.275613,13.58145,13.358865,13.27964,13.124963,12.642066,11.506506,12.178034,11.921495,12.294985,13.192869,12.864652,12.291212,12.117672,12.147853,12.264804,12.434572,10.763299,9.748463,8.518587,7.24344,7.1566696,7.118943,8.054554,8.273367,7.7414265,8.073418,9.695646,9.186342,12.702429,18.229324,15.580941,11.744182,11.676274,12.208215,15.618668,29.630198,17.278622,6.7643166,8.590267,17.395575,11.962994,12.73261,8.83926,6.0701537,6.7944975,9.978593,8.088508,9.344792,10.155907,9.480607,8.835487,7.6131573,7.6848373,7.99042,7.699928,6.2097406,5.832478,6.3229194,6.047518,4.881777,4.2102494,4.7120085,5.040227,5.2779026,5.6476197,6.515323,7.394345,7.3113475,6.6586833,6.0626082,6.379509,5.7570257,5.353355,5.05909,4.708236,4.074435,3.3312278,3.1425967,3.0218725,3.6745367,7.0170827,4.919503,4.5497856,3.9386206,3.3236825,5.142088,5.0439997,5.9720654,6.4738245,6.3719635,6.7756343,5.323174,5.372218,5.7192993,5.904158,6.2097406,5.696664,5.881522,6.2851934,6.7114997,7.2472124,6.0512905,6.356873,6.7114997,6.477597,5.828706,4.889322,4.644101,4.466788,4.689373,6.590776,4.9685473,4.3347464,4.6742826,5.0138187,3.4029078,1.7542707,1.0940613,1.901403,3.1765501,2.4559789,2.04099,3.0105548,4.5912848,7.6886096,14.875461,7.224577,5.3194013,5.1798143,5.0251365,5.292993,5.5004873,6.560595,7.4169807,7.8206515,8.345046,9.0543,10.163452,10.842525,10.831206,10.453944,10.585986,11.114153,10.906659,9.986138,9.522105,9.178797,8.114917,6.8737226,5.7419353,4.715781,4.557331,5.5797124,6.2851934,6.4247804,6.971811,6.6813188,7.220804,7.8923316,8.152642,7.6131573,8.518587,9.639057,10.306811,10.321902,9.978593,10.076681,9.733373,9.318384,9.005256,8.7751255,8.043237,7.281166,7.001992,7.020855,6.470052,6.1041074,5.6476197,5.6023483,6.039973,6.5756855,7.5527954,8.088508,8.186596,7.967784,7.673519,7.7376537,8.054554,8.382772,8.333729,7.3717093,7.224577,8.624221,9.782416,10.114408,10.223814,10.687846,10.374719,9.529651,9.009028,10.253995,11.363147,12.257258,12.781653,12.894833,12.649611,12.868423,12.849561,13.185325,13.622949,13.060828,12.755245,12.58925,11.996947,11.004747,10.223814,10.759526,11.170743,10.985884,9.971047,8.103599,7.956466,7.9300575,7.7150183,7.2887115,6.8963585,6.6020937,5.798525,6.043745,7.281166,7.8432875,7.4773426,7.3113475,6.72659,5.873977,5.692891,5.643847,5.100589,5.726845,7.375482,8.073418,7.9753294,8.024373,8.345046,8.537451,7.6584287,8.892077,9.465516,9.797507,10.242677,11.106608,10.985884,9.891823,9.582467,10.167224,10.133271,9.680555,10.054046,11.219787,12.574159,12.940104,13.158916,12.894833,11.936585,10.559577,9.522105,9.88805,10.838752,11.491416,11.7894535,12.498707,9.548513,11.408418,13.124963,13.630494,13.35132,14.18507,15.143317,15.535669,15.226315,14.320885,13.158916,13.249459,13.313594,13.026875,12.67602,13.162688,13.087236,13.268322,13.6682205,14.200161,14.735873,13.947394,13.132507,12.81938,12.762791,11.92904,11.3820095,10.929295,11.099063,11.98563,13.245687,14.754736,15.414946,15.667711,15.558306,14.735873,14.015302,13.943622,14.139798,14.302021,14.200161,14.215251,14.0907545,13.65313,13.0646,12.804289,12.781653,12.842015,12.955194,13.117417,13.373956,13.804035,14.128481,14.1926155,14.139798,14.422746,13.985121,14.351066,14.875461,15.158407,15.0376835,14.588741,14.479335,13.864397,12.917468,12.826925,12.091263,11.465008,11.216014,11.140562,10.56335,9.7296,9.099571,8.933576,9.129752,9.235386,8.948667,8.416726,8.27714,8.4544525,8.14887,8.503497,8.3525915,7.986647,7.654656,7.533932,6.971811,7.0963078,7.432071,7.665974,7.6622014,8.443134,8.726082,8.922258,9.107117,9.046755,9.865415,10.695392,11.631002,12.755245,14.158662,16.014793,15.629986,13.717264,11.408418,10.246449,8.216777,5.6098933,3.169005,1.4222796,0.663982,0.6073926,0.482896,0.482896,0.633801,0.7809334,0.7922512,0.9393836,1.0336993,1.0186088,0.935611,0.8262049,0.7507524,0.91674787,1.1695137,1.0035182,1.267602,1.2902378,1.2562841,1.297783,1.4901869,1.6675003,1.5279131,1.2600567,0.95824677,0.6073926,0.31312788,0.211267,0.29803738,0.45648763,0.45648763,0.4979865,0.67152727,0.79602385,0.95447415,1.478869,1.6712729,2.033445,2.3126192,2.4823873,2.7879698,3.62172,3.6745367,3.6066296,3.6971724,3.85185,3.9386206,4.0480266,4.285702,4.5535583,4.5912848,4.5422406,4.82896,4.821415,4.5799665,4.8327327,5.6400743,5.643847,5.764571,5.96452,5.2628117,5.4288073,5.5683947,5.753253,6.0739264,6.647365,6.971811,7.062354,7.6584287,8.650629,9.076936,9.484379,9.525878,9.171251,8.926031,9.812597,9.473062,9.110889,8.888305,8.865668,9.042982,9.480607,9.733373,9.971047,10.227587,10.446399,10.012547,9.861642,9.601331,9.34102,9.673011,9.574923,9.869187,9.559832,8.778898,8.782671,9.7220545,10.250222,10.93684,11.872451,12.672247,11.774363,10.763299,10.378491,10.544487,10.367173,10.638803,10.27663,9.525878,8.801534,8.684583,8.43559,9.26934,10.280403,11.087745,11.846043,11.91395,11.763044,11.668729,11.827179,12.313848,12.974057,13.151371,12.958967,12.555296,12.136535,11.1631975,10.887795,10.748209,10.47658,10.103089,10.084227,9.771099,9.076936,8.235641,7.8508325,8.790216,9.597558,9.684328,9.22784,9.14107,8.065872,6.85486,7.394345,9.737145,12.102581,11.725319,10.057818,8.345046,7.84706,9.846551,12.377983,12.792972,11.778135,10.231359,9.25425,6.907676,6.741681,8.627994,10.714255,9.424017,10.533169,10.435081,10.593531,10.921749,9.782416,9.288202,8.707218,9.476834,11.200924,11.649866,10.340765,11.012292,11.812089,11.883769,11.389555,11.283921,11.812089,10.552032,7.8621507,6.8925858,9.129752,9.737145,10.623712,12.193124,13.343775,14.992412,12.90615,10.020092,7.8508325,6.470052,5.594803,4.293247,2.686109,1.4977322,2.0636258,2.6634734,4.1800685,4.6327834,3.5575855,1.9957186,2.637065,3.0445085,4.8930945,7.567886,8.156415,13.113645,14.200161,13.777626,12.091263,7.24344,4.768598,5.560849,4.749735,1.9844007,1.4524606,2.384299,2.2371666,2.1654868,2.535204,2.916239,3.772625,4.3196554,4.6327834,4.6931453,4.402653,4.504514,4.5837393,5.221313,6.1305156,6.1342883,5.6815734,6.205968,7.2585306,8.514814,9.786189,10.310584,10.174769,9.688101,9.050528,8.360137,8.650629,9.163706,9.224068,8.926031,9.125979,7.0963078,6.4738245,7.141579,8.386545,8.907167,9.971047,10.525623,10.567122,10.661438,11.936585,13.230596,15.022593,16.637276,17.30503,16.161926,15.313085,14.898096,14.656648,14.667966,15.343266,17.372938,19.247932,18.946123,16.109108,12.034674,11.442371,11.615912,11.423509,10.9594755,11.536687,11.45369,11.151879,11.653639,13.106099,14.78869,16.301512,16.01102,15.147089,14.750964,15.660167,16.022339,13.909668,12.442118,12.566614,13.019329,13.947394,13.426772,12.140307,11.0613365,11.46878,12.042219,12.498707,13.449409,14.784918,15.660167,14.558559,14.6151495,13.977575,12.038446,9.4013815,10.699164,12.510024,14.6302395,15.467763,12.049765,9.691874,9.171251,9.2844305,9.582467,10.38981,11.61214,12.913695,13.170234,12.570387,12.615658,13.109872,13.328684,12.604341,11.242422,10.518079,11.510279,11.608367,11.9064045,12.672247,13.340002,13.487134,12.800517,12.528888,12.917468,13.204187,11.729091,11.144334,9.57115,7.405663,7.3377557,6.94163,6.8925858,7.232122,7.375482,6.092789,7.7678347,8.718536,10.193633,12.136535,13.185325,12.528888,13.215506,14.27184,24.239115,61.161797,47.98779,20.689075,5.50426,7.8319697,12.23085,7.9526935,8.7600355,7.643338,5.13077,9.2844305,7.4396167,9.325929,10.438853,9.669238,9.288202,8.884532,8.137552,7.756517,7.677292,7.0284004,7.0887623,7.1038527,6.8397694,5.9796104,4.13857,4.112161,4.5460134,5.194905,5.8437963,6.319147,6.643593,6.56814,6.1720147,5.753253,5.8173876,5.643847,4.7006907,4.1574326,4.255521,4.293247,3.2557755,2.8521044,3.0709167,4.5799665,8.714764,7.6207023,5.915476,5.240176,5.5004873,4.847823,5.2288585,5.7419353,5.802297,5.6061206,6.126743,4.9685473,5.6400743,6.228604,5.945657,5.1345425,5.0251365,5.753253,6.2135134,6.33801,7.0887623,5.481624,5.553304,5.3759904,4.5724216,4.315883,4.3309736,4.436607,4.5233774,4.8742313,6.1644692,4.647874,4.2894745,3.4142256,2.2673476,2.9992368,5.4438977,5.111907,5.100589,5.938112,5.5683947,4.1272516,3.9310753,3.7462165,5.745708,15.513034,10.993429,7.375482,5.3873086,4.983638,5.3194013,5.4401255,6.9680386,8.246958,8.850578,9.578695,9.937095,10.502988,10.967021,11.151879,11.038701,10.978339,10.9594755,10.502988,9.703192,9.22784,9.491924,8.650629,7.5829763,6.7379084,6.1305156,5.3684454,6.228604,6.6549106,6.3229194,6.6549106,6.7039547,7.2057137,7.9791017,8.375228,7.273621,8.069645,8.975075,9.58624,9.906913,10.355856,10.269085,9.49947,8.646856,8.028146,7.699928,7.4735703,7.062354,6.647365,6.319147,6.043745,6.2021956,6.1041074,6.1116524,6.519096,7.5527954,7.5829763,7.4282985,7.5716586,7.960239,8.016829,8.262049,8.137552,7.9941926,7.888559,7.5792036,7.605612,8.428044,9.593785,10.63503,11.065109,10.729345,10.163452,9.431562,9.1825695,10.631257,11.714001,12.23085,12.800517,13.45318,13.63804,13.788944,13.996439,14.200161,14.539697,15.354584,14.173752,13.35132,12.947649,12.638294,11.747954,11.415963,11.544232,11.46878,10.668983,8.7751255,8.118689,7.7904706,7.54525,7.2623034,6.9227667,6.56814,5.5306683,5.281675,6.039973,6.7567716,6.3719635,6.3417826,6.4926877,6.598321,6.387054,6.0550632,5.80607,6.4134626,7.6395655,8.265821,7.3981175,7.6282477,8.107371,8.299775,7.9791017,9.042982,9.5032425,9.484379,9.42779,10.057818,10.56335,9.80128,9.129752,9.103344,9.484379,9.35611,9.484379,9.695646,10.167224,11.449917,12.283667,13.475817,14.011529,13.600313,12.657157,12.291212,12.344029,12.370438,12.291212,12.362892,10.582213,11.925267,13.505998,14.049255,13.626721,13.649357,13.649357,14.803781,15.026365,13.849306,12.419481,12.864652,12.83447,12.510024,12.325166,12.96274,13.124963,13.189097,13.400364,13.6682205,13.551269,12.781653,12.257258,12.264804,12.419481,11.676274,11.329193,10.582213,10.182315,10.521852,11.657412,13.649357,14.924504,15.316857,14.830189,13.656902,13.321139,13.45318,13.577678,13.521088,13.389046,13.656902,13.687083,13.3626375,12.774108,12.219532,12.525115,12.936331,13.373956,13.758763,14.003984,14.290704,14.626467,14.837734,14.898096,14.924504,14.596286,14.600059,14.667966,14.532151,13.920986,13.9888935,13.917213,13.547497,13.000465,12.717519,12.053536,11.631002,11.299012,10.876478,10.174769,9.510788,9.088254,8.801534,8.744945,9.22784,8.816625,8.548768,8.495952,8.533678,8.329956,8.239413,7.752744,7.3905725,7.2660756,7.073672,6.9982195,7.24344,7.567886,7.8131065,7.8961043,8.156415,8.390318,8.7751255,9.114662,8.865668,10.18986,10.9594755,12.140307,14.000212,16.15438,16.486372,15.614895,14.181297,12.649611,11.299012,7.673519,4.4177437,2.2786655,1.2751472,0.69793564,0.69039035,0.5357128,0.38858038,0.31312788,0.28294688,0.2678564,0.32067314,0.36971724,0.38480774,0.392353,0.34330887,0.35085413,0.47912338,0.6488915,0.63002837,0.8262049,0.97333723,1.0336993,1.0714256,1.2449663,1.5015048,1.4901869,1.1732863,0.7507524,0.63002837,0.32067314,0.241448,0.271629,0.29803738,0.2565385,0.30935526,0.392353,0.5885295,0.8601585,1.0827434,1.1695137,1.478869,1.8334957,2.1541688,2.425798,3.1840954,3.1576872,3.127506,3.4142256,3.8820312,4.112161,4.2027044,4.429062,4.7648253,4.8968673,4.7308717,4.9345937,4.8138695,4.402653,4.4630156,4.7572803,4.6742826,4.7120085,4.949684,5.0175915,5.27413,5.342037,5.6325293,6.2927384,7.175533,7.254758,7.6131573,8.394091,9.273112,9.469289,9.714509,9.420244,9.012801,8.937348,9.650374,10.103089,9.718282,9.578695,9.884277,9.952185,9.940866,10.303039,10.423763,10.412445,11.087745,10.785934,10.386037,10.072908,9.929549,9.940866,10.386037,10.370946,9.793735,9.133525,9.450426,9.97482,10.423763,11.053791,11.774363,12.147853,11.408418,10.612394,10.137043,10.03141,10.0276375,10.529396,10.518079,10.065364,9.495697,9.382519,9.390063,9.940866,11.144334,12.706201,13.913441,14.332202,14.8339615,14.358611,13.215506,13.094781,13.038192,13.189097,13.290957,13.268322,13.253232,12.411936,11.480098,10.850069,10.502988,10.001229,9.933322,9.574923,9.084481,8.631766,8.394091,8.7751255,9.273112,9.220296,8.710991,8.616675,7.635793,6.5002327,6.828451,8.6581745,10.453944,10.933067,10.608622,9.522105,8.296002,8.141325,9.665465,10.63503,11.121698,10.929295,9.593785,7.4282985,7.224577,8.703445,10.370946,9.548513,10.250222,10.329447,10.8576145,11.438599,10.227587,9.737145,9.563604,10.167224,11.249968,11.759273,11.053791,11.359374,11.608367,11.532914,11.657412,11.404645,12.438345,11.548005,8.469543,5.855114,8.111144,9.144843,10.223814,11.223559,10.631257,11.932813,12.47607,11.200924,8.461998,6.013564,6.2814207,4.568649,3.4896781,4.1762958,6.270103,4.5950575,4.4516973,3.802806,2.3126192,1.3656902,3.6330378,3.7462165,5.7570257,9.582467,10.982111,12.694883,12.223305,10.77839,8.488406,4.38379,4.2328854,3.5802212,2.3578906,1.3958713,2.3880715,3.0633714,2.7426984,2.6672459,3.1840954,3.7462165,4.9534564,5.05909,5.040227,5.040227,4.3649273,4.0970707,4.376245,4.7836885,5.093044,5.2590394,4.8930945,5.7079816,6.9227667,8.080963,9.046755,10.506761,10.940613,10.47658,9.582467,9.065618,9.107117,9.239159,9.175024,9.035437,9.367428,7.24344,6.149379,6.398372,7.6131573,8.703445,8.8618965,8.9788475,8.959985,9.107117,10.106862,11.593277,12.842015,13.86817,14.475562,14.25675,15.154634,15.954432,16.376965,16.275105,15.63753,15.931795,18.376457,19.515789,17.663431,12.928786,12.08749,11.3971,10.533169,9.918231,10.710483,10.412445,10.155907,10.56335,11.763044,13.396591,15.339493,15.569623,15.045229,14.566105,14.781145,15.47908,14.317112,12.826925,11.819634,11.41219,12.789199,12.709973,11.955449,11.287694,11.476325,11.902632,12.362892,13.132507,14.154889,15.049001,13.694629,12.875969,12.310076,11.476325,9.623966,11.351829,13.147598,14.132254,13.721037,11.604594,9.669238,8.763808,8.722309,9.280658,10.084227,10.650121,11.921495,13.072145,13.8870325,14.728328,15.267814,14.136025,11.891314,9.688101,9.273112,10.725573,10.902886,11.140562,11.898859,12.770335,12.955194,12.596795,12.313848,12.351574,12.608112,11.502733,11.559323,10.495442,8.382772,7.643338,7.5716586,7.152897,7.4282985,7.8395147,6.258785,7.322665,8.646856,9.650374,10.137043,10.336992,12.038446,16.739138,17.516298,22.337713,54.061718,51.205837,23.273323,4.8365054,6.1418333,13.102326,6.462507,9.171251,9.590013,6.224831,7.7187905,8.567632,9.714509,10.216269,9.839006,9.061845,9.159933,8.409182,7.854605,7.726336,7.435844,7.9036493,7.748972,7.575431,7.062354,4.961002,4.1008434,4.395108,5.240176,6.066381,6.326692,6.039973,6.2135134,5.9607477,5.311856,5.2099953,5.5004873,4.515832,3.9348478,4.1800685,4.432834,3.0709167,2.6144292,2.8936033,4.0706625,6.63982,6.319147,4.8968673,4.5912848,5.3344917,4.776143,4.8138695,5.032682,5.1043615,5.0968165,5.4703064,5.270357,6.0248823,6.5945487,6.4134626,5.481624,5.409944,5.8890676,5.9796104,5.8211603,6.620957,5.240176,5.270357,5.168496,4.7044635,4.927048,4.353609,4.568649,5.0741806,5.4401255,5.3080835,4.346064,4.7912335,3.9763467,3.078462,7.1302614,9.431562,14.883006,16.463736,12.321393,5.772116,5.5457587,4.5309224,4.025391,5.696664,11.570641,16.580687,9.895596,4.90064,5.3873086,5.572167,5.2175403,6.6360474,8.22055,9.49947,11.151879,11.155652,11.374464,11.664956,11.978085,12.37421,12.061082,11.140562,10.106862,9.405154,9.420244,9.0807085,8.646856,7.9715567,7.24344,6.960493,6.043745,6.6624556,7.183078,7.039718,6.7152724,6.7077274,6.9567204,7.5905213,8.073418,7.194396,7.9300575,8.499724,8.797762,9.125979,10.197406,10.001229,9.118435,8.27714,7.7376537,7.273621,7.0548086,6.952948,6.688864,6.3531003,6.428553,6.48137,6.7756343,7.1793056,7.8395147,9.159933,8.337502,7.413208,7.194396,7.594294,7.61693,8.084735,8.111144,7.9715567,7.756517,7.3905725,7.2660756,7.707473,8.552541,9.57115,10.469034,10.518079,10.272858,10.001229,10.050273,10.86516,12.136535,12.751472,13.283413,13.924759,14.479335,15.07541,15.173498,14.890551,14.875461,16.305285,15.494171,14.362384,13.849306,13.856852,13.257004,13.087236,12.574159,11.751727,10.691619,9.480607,8.262049,7.4584794,6.8171334,6.221059,5.7117543,5.7381625,5.413717,5.4740787,6.047518,6.651138,6.3116016,5.824933,6.126743,7.0774446,7.484888,7.164215,6.888813,6.907676,7.3151197,8.050782,7.4282985,7.5226145,7.8017883,8.028146,8.2507305,9.34102,10.18986,10.265312,9.756008,9.574923,10.310584,10.291721,9.955957,9.7296,10.054046,9.846551,9.767326,9.616421,9.64283,10.529396,11.423509,13.109872,14.358611,14.667966,14.268067,14.954685,14.93205,14.317112,13.340002,12.336484,12.268577,12.921241,14.003984,14.445381,14.04171,13.430545,12.721292,13.747445,14.173752,13.385274,12.464753,12.472299,12.498707,12.604341,12.894833,13.505998,13.804035,13.649357,13.419228,13.079691,12.162943,11.608367,11.3971,11.627231,11.978085,11.69891,11.461235,10.672756,10.208723,10.397354,11.02361,12.132762,13.234368,13.807808,13.713491,13.192869,13.045737,13.343775,13.58145,13.536179,13.264549,13.275867,13.298503,13.200415,12.955194,12.626976,12.823153,13.147598,13.517315,13.834216,13.992666,14.196388,14.611377,15.045229,15.335721,15.331948,15.16218,14.671739,14.313339,13.95494,12.898605,13.162688,13.249459,13.147598,12.868423,12.442118,11.996947,11.747954,11.302785,10.54826,9.673011,9.424017,9.110889,8.778898,8.616675,8.959985,8.786444,8.729855,8.737399,8.763808,8.744945,8.382772,7.7338815,7.3075747,7.2170315,7.183078,7.277394,7.515069,7.6282477,7.6395655,7.865923,7.7942433,8.058327,8.443134,8.733627,8.737399,10.069136,10.733118,12.411936,15.188588,17.512526,16.4826,15.9695215,15.79598,15.388537,13.781399,7.967784,3.7084904,1.5241405,0.97710985,0.65643674,0.5998474,0.6073926,0.45648763,0.17354076,0.056589376,0.03772625,0.049044125,0.071679875,0.094315626,0.11317875,0.12826926,0.15467763,0.23013012,0.33576363,0.41121614,0.6375736,0.7884786,0.98842776,1.20724,1.2713746,1.2185578,1.1732863,0.9016574,0.543258,0.5885295,0.331991,0.35462674,0.3734899,0.31312788,0.32444575,0.38103512,0.41121614,0.51684964,0.70170826,0.87147635,1.0223814,1.1996948,1.5165952,1.9429018,2.2975287,2.9011486,2.7502437,2.727608,3.138824,3.712263,4.0706625,4.3007927,4.5761943,4.908185,5.149633,4.927048,4.9760923,4.825187,4.4818783,4.425289,4.357382,4.112161,4.055572,4.315883,4.768598,4.8968673,4.98741,5.2250857,5.828706,7.0170827,7.4471617,8.152642,8.831716,9.2995205,9.495697,9.752235,9.393836,8.959985,8.801534,9.0807085,10.314357,9.922004,9.7296,10.208723,10.484125,10.684074,11.151879,11.3669195,11.442371,12.136535,11.993175,11.449917,10.891568,10.370946,9.623966,10.272858,10.355856,10.012547,9.7069645,10.220041,10.370946,10.740664,11.23865,11.68382,11.808316,11.706455,11.268831,10.736891,10.329447,10.265312,10.450171,10.751981,10.744436,10.487898,10.514306,10.687846,11.087745,12.400619,14.3095665,15.467763,16.260014,17.14658,16.622187,15.150862,15.17727,14.6302395,14.675511,14.837734,14.803781,14.418973,13.558814,12.359119,11.400873,10.740664,9.940866,9.654147,9.1976595,8.907167,8.801534,8.590267,8.6581745,8.907167,8.831716,8.529905,8.722309,7.8432875,6.937857,7.2698483,8.499724,8.695901,9.001483,9.529651,9.442881,8.703445,8.088508,9.250477,9.540969,10.035183,10.763299,10.718028,9.337247,8.035691,8.314865,9.835234,10.427535,10.842525,10.257768,10.242677,10.695392,9.827688,9.601331,9.691874,10.295494,11.136789,11.491416,11.46878,11.887542,11.695138,11.197151,12.049765,10.985884,11.857361,11.763044,9.627739,6.2361493,7.8131065,8.944894,10.272858,11.32542,10.533169,10.54826,11.517824,10.997202,8.8769865,7.4018903,6.587003,5.2967653,5.4174895,7.2660756,9.608876,6.307829,5.0213637,3.904667,2.5012503,1.7316349,3.3538637,3.8556228,6.688864,10.827434,10.733118,10.016319,8.986393,7.17176,4.659192,2.0975795,2.8445592,2.0296721,1.6184561,2.4220252,4.08198,4.3083377,4.044254,4.0782075,4.6026025,5.1798143,6.1418333,5.975838,5.6325293,5.323174,4.504514,3.8669407,4.1574326,4.3007927,4.1197066,4.3347464,4.4630156,5.8437963,7.250985,8.088508,8.394091,9.929549,10.665211,10.408672,9.593785,9.261794,9.397609,9.092027,8.959985,9.190115,9.552286,7.8734684,6.8058157,6.6662283,7.533932,9.239159,8.684583,8.616675,8.89585,9.378746,9.929549,10.529396,10.650121,10.797253,11.208468,11.830952,13.306048,15.007503,16.343012,16.810818,15.98084,16.331694,18.202915,19.395065,18.433046,14.569878,13.102326,11.962994,10.684074,9.691874,10.295494,10.11818,9.857869,10.167224,11.227332,12.770335,14.924504,15.475307,14.562332,13.045737,12.510024,13.321139,13.377728,12.698656,11.555551,10.472807,11.714001,12.181807,12.083718,11.717773,11.506506,11.272603,11.676274,12.219532,12.7477,13.449409,12.717519,11.212241,10.397354,10.442626,10.250222,12.449662,13.645585,13.132507,11.487643,10.578441,9.574923,8.6581745,8.492179,9.050528,9.601331,9.861642,11.510279,13.547497,15.328176,16.58446,17.150352,14.78869,11.608367,9.314611,9.205205,9.88805,9.9257765,10.54826,11.77059,12.415709,12.136535,11.876224,11.25374,10.774617,11.834724,11.140562,11.638548,11.642321,10.472807,8.439363,8.179051,7.8395147,7.9338303,8.118689,7.1793056,7.6131573,8.386545,9.363655,10.152134,10.11818,11.3820095,17.05981,16.569368,14.132254,28.762493,31.090202,15.456445,6.19465,9.548513,13.671993,8.186596,10.26154,10.521852,7.745199,8.827943,12.132762,11.038701,9.665465,9.322156,8.503497,8.846806,8.586494,8.3525915,8.265821,7.9225125,8.284684,8.073418,8.00551,7.8621507,6.4926877,5.353355,5.13077,5.560849,6.187105,6.349328,5.723072,6.085244,6.043745,5.3194013,4.727099,5.1156793,4.534695,4.0517993,4.0291634,4.0970707,3.048281,2.625747,2.8256962,3.6179473,4.938366,4.738417,3.8292143,3.9159849,4.776143,4.2706113,4.346064,4.8025517,4.851596,4.4894238,4.4705606,5.13077,5.824933,6.2814207,6.417235,6.3531003,6.2135134,6.217286,5.956975,5.594803,5.885295,5.0477724,5.062863,5.292993,5.5193505,5.938112,4.478106,5.1269975,6.1531515,6.1795597,4.183841,5.2062225,5.726845,4.52715,4.1498876,10.86516,13.060828,18.685812,18.504726,11.830952,6.5341864,6.7341356,4.817642,4.376245,6.224831,8.424272,16.863634,9.64283,4.538468,6.19465,6.1229706,5.934339,6.6549106,7.986647,9.797507,12.1101265,11.729091,11.619685,11.876224,12.506252,13.468271,13.151371,11.578186,10.087999,9.367428,9.469289,8.82417,8.741172,8.228095,7.3717093,7.3151197,7.0284004,7.5112963,8.13378,8.27714,7.322665,7.383027,7.2396674,7.484888,7.8319697,7.1340337,7.707473,8.16396,8.235641,8.314865,9.439108,9.295748,8.529905,7.858378,7.5188417,7.2623034,6.888813,6.7869525,6.7114997,6.72659,7.1793056,7.213259,7.6508837,8.171506,8.7600355,9.703192,8.782671,7.828197,7.462252,7.567886,7.281166,7.61693,7.7829256,7.8131065,7.696155,7.3717093,7.092535,7.3000293,7.8998766,8.835487,10.099318,10.257768,10.382264,10.552032,10.748209,10.86516,12.034674,12.970284,13.864397,14.705692,15.256495,15.539442,15.109364,14.460471,14.339747,15.754482,15.596032,14.407655,13.5663595,13.317367,12.774108,13.475817,13.317367,12.536433,11.45369,10.484125,8.926031,7.7338815,6.6662283,5.715527,5.1345425,5.2892203,5.6476197,6.25124,6.903904,7.1566696,6.719045,5.828706,5.938112,7.043491,7.6923823,7.7942433,7.5829763,7.092535,6.749226,7.3679366,7.484888,7.5037513,7.677292,8.043237,8.420499,9.631512,11.234878,11.759273,10.982111,9.895596,10.552032,11.057564,11.02361,10.642575,10.665211,10.054046,9.880505,9.906913,10.231359,11.272603,12.649611,14.4152,15.207452,14.796235,14.034165,15.475307,15.645076,14.981093,13.8719425,12.657157,14.071891,14.532151,15.098045,15.173498,14.622695,13.728582,13.3626375,13.826671,14.124708,13.807808,12.992921,12.223305,12.377983,12.985375,13.739901,14.471789,14.766054,14.268067,13.449409,12.510024,11.408418,11.363147,11.400873,11.649866,11.951676,11.876224,11.378237,10.831206,10.8576145,11.363147,11.54046,11.491416,11.781908,12.37421,13.094781,13.622949,13.245687,13.441863,13.815352,14.019074,13.743673,13.287186,13.211733,13.377728,13.607859,13.656902,13.306048,13.204187,13.257004,13.370183,13.43809,13.679539,14.037937,14.403882,14.724555,14.988639,14.9358225,14.373701,13.951167,13.543724,12.291212,12.306303,12.66093,12.774108,12.491161,12.106354,11.940358,11.551778,10.861387,9.978593,9.21275,9.314611,8.907167,8.661947,8.688355,8.544995,8.914713,8.986393,9.046755,9.190115,9.2995205,9.031664,8.333729,7.745199,7.5188417,7.6093845,7.496206,7.643338,7.594294,7.3981175,7.605612,7.696155,7.8961043,7.907422,7.9413757,8.722309,9.563604,10.34831,12.702429,15.90916,16.939087,16.493916,16.867407,17.938831,18.65563,17.063583,9.35611,4.025391,1.3166461,0.62625575,0.5017591,0.29426476,0.47912338,0.482896,0.2263575,0.120724,0.06413463,0.026408374,0.026408374,0.0452715,0.02263575,0.049044125,0.06413463,0.15467763,0.30181,0.34330887,0.694163,0.7092535,0.9507015,1.3619176,1.2600567,0.84884065,0.7394345,0.62248313,0.49421388,0.6790725,0.5093044,0.6111652,0.58475685,0.43385187,0.5696664,0.58475685,0.5998474,0.5583485,0.5281675,0.7054809,1.0186088,1.0412445,1.267602,1.7467253,2.1013522,2.6823363,2.6408374,2.7087448,3.1161883,3.5689032,3.953711,4.3724723,4.6856003,4.908185,5.194905,5.0213637,4.961002,4.881777,4.749735,4.659192,4.636556,4.285702,4.123479,4.2291126,4.2630663,4.349837,4.610148,4.6931453,4.9459114,6.4021444,7.33021,8.058327,8.495952,8.733627,9.046755,9.439108,9.21275,8.726082,8.288457,8.186596,9.556059,9.231613,9.020347,9.578695,10.401127,11.200924,11.955449,12.694883,13.400364,13.996439,13.9888935,13.2607765,12.419481,11.510279,9.986138,9.993684,10.321902,10.529396,10.570895,10.804798,10.774617,10.917976,11.234878,11.6008215,11.744182,12.030901,11.879996,11.615912,11.332966,10.872705,10.506761,11.057564,11.517824,11.574413,11.623458,11.800771,12.253486,13.517315,15.184815,15.920478,16.878725,17.542706,17.293713,16.678776,17.4333,17.105082,17.093763,17.097536,16.72782,15.494171,14.667966,13.645585,12.596795,11.521597,10.250222,9.661693,8.941121,8.541223,8.465771,8.280911,8.273367,8.499724,8.499724,8.3525915,8.6732645,8.235641,7.816879,8.239413,9.167479,9.125979,8.643084,8.650629,8.586494,8.439363,8.7600355,10.269085,9.669238,9.027891,9.420244,10.963248,10.725573,8.541223,8.028146,9.756008,11.234878,11.2650585,10.054046,9.224068,9.190115,9.175024,9.574923,9.623966,10.091772,10.850069,10.868933,11.261286,11.872451,11.465008,10.653893,11.895086,9.857869,10.155907,10.789707,10.367173,8.111144,8.439363,9.084481,10.487898,12.140307,12.608112,11.2650585,10.834979,10.091772,9.378746,10.608622,6.9491754,6.2135134,7.1302614,8.612903,9.771099,6.7680893,5.772116,4.979865,3.7990334,2.8219235,2.3088465,4.123479,8.420499,12.136535,9.027891,7.141579,7.0359454,5.2288585,1.9429018,1.0789708,1.3958713,1.8599042,2.7879698,4.2328854,5.975838,5.80607,5.8211603,6.300284,6.9944468,7.1302614,6.9491754,6.7152724,6.0362,5.070408,4.52715,4.1612053,4.304565,4.146115,3.8254418,4.4139714,5.3269467,7.111398,8.243186,8.337502,8.137552,9.4127,10.20495,10.174769,9.559832,9.159933,9.597558,8.993938,8.7751255,9.265567,9.669238,8.273367,7.7338815,7.515069,7.805561,9.533423,9.012801,9.009028,9.597558,10.378491,10.484125,10.291721,10.005001,9.835234,10.023865,10.846297,11.193378,12.781653,14.302021,15.147089,15.396083,17.870924,18.72731,19.346022,19.349794,16.588232,14.0907545,12.955194,11.751727,10.480352,10.574668,10.163452,9.952185,10.367173,11.532914,13.27964,14.875461,14.924504,13.272095,10.982111,10.355856,11.019837,11.54046,11.736636,11.427281,10.442626,11.117926,11.623458,11.751727,11.536687,11.23865,10.038955,10.246449,10.631257,10.79348,11.151879,11.529142,10.167224,9.21275,9.58624,10.970794,13.460726,14.045483,12.706201,10.495442,9.533423,9.42779,8.941121,8.850578,9.26934,9.635284,9.978593,11.910177,14.037937,15.743164,17.172989,17.693611,14.905642,11.887542,10.253995,10.174769,8.918486,8.677037,9.922004,11.834724,12.306303,11.676274,11.106608,9.81637,8.850578,11.0613365,10.77839,11.476325,12.574159,12.638294,9.367428,8.582722,8.175279,7.964011,7.8508325,7.7942433,8.043237,8.137552,8.793989,10.238904,12.208215,11.668729,14.188843,12.468526,7.5527954,8.816625,8.0206,6.964266,8.654402,12.264804,13.132507,11.306557,11.604594,10.269085,8.213005,11.016065,15.207452,12.291212,9.144843,8.318638,8.00551,8.416726,8.567632,8.726082,8.805306,8.375228,8.480861,8.420499,8.367682,8.27714,7.8961043,7.364164,6.5568223,6.175787,6.319147,6.458734,5.798525,6.1041074,6.2399216,5.674028,4.4705606,4.5950575,4.6290107,4.29702,3.6971724,3.3048196,3.1010978,2.795515,2.897376,3.5500402,4.5460134,3.9801195,3.4368613,3.731126,4.3422914,3.4255435,4.2781568,5.0666356,4.851596,4.08198,4.587512,4.7836885,5.160951,5.6589375,6.2889657,7.1264887,6.990674,6.677546,6.273875,5.80607,5.2665844,5.1873593,5.1835866,5.66271,6.4436436,6.7341356,4.8025517,6.089017,7.405663,6.7831798,3.4557245,8.793989,8.5563135,5.4363527,4.191386,11.634775,15.199906,15.731846,11.329193,6.7114997,13.215506,9.884277,5.764571,4.4818783,6.466279,8.941121,11.046246,6.5530496,4.647874,6.802043,6.749226,7.1981683,6.8774953,7.598067,9.748463,12.264804,11.638548,11.151879,11.355601,12.393073,13.985121,13.456953,11.864905,10.401127,9.616421,9.431562,9.016574,9.084481,8.507269,7.432071,7.2660756,8.201687,8.986393,9.646602,9.7220545,8.265821,8.367682,8.031919,7.865923,7.7678347,6.9189944,7.273621,7.8621507,7.956466,7.752744,8.360137,8.605357,8.118689,7.537705,7.281166,7.5565677,7.1679873,6.881268,6.9265394,7.3377557,7.9828744,8.228095,8.631766,8.944894,9.114662,9.242931,8.827943,8.329956,8.009283,7.7942433,7.273621,7.149124,7.1679873,7.2472124,7.3490734,7.466025,7.356619,7.61693,8.296002,9.35611,10.665211,10.518079,10.748209,11.038701,11.125471,10.770844,11.472552,12.66093,14.196388,15.543215,15.773345,15.23386,14.128481,13.283413,13.241914,14.252977,14.558559,13.441863,12.381755,11.808316,11.087745,12.193124,13.015556,13.290957,12.913695,11.951676,10.103089,8.601585,7.1566696,5.9192486,5.481624,5.553304,6.1078796,7.043491,7.8810134,7.779153,7.175533,6.2361493,6.0248823,6.5756855,6.911449,7.4509344,7.5188417,7.009537,6.3945994,6.722818,7.4735703,7.4999785,7.647111,8.114917,8.465771,9.786189,11.766817,12.751472,12.238396,10.872705,11.25374,11.864905,11.887542,11.283921,10.789707,9.929549,9.839006,10.27663,11.200924,12.774108,14.8339615,16.437326,16.188334,14.3095665,12.638294,13.920986,14.275613,14.351066,14.245432,13.536179,14.875461,15.0376835,15.671484,15.769572,15.0376835,13.902123,14.400109,15.230087,15.769572,15.297995,13.015556,12.453435,12.498707,12.709973,13.151371,14.373701,14.909414,14.173752,13.419228,13.041965,12.604341,13.505998,13.283413,12.985375,12.853333,12.3289385,10.899114,10.56335,10.646348,10.955703,11.747954,12.479843,12.593022,12.725064,13.147598,13.732355,13.4644985,13.377728,13.396591,13.547497,13.962485,13.792717,13.7851715,14.162435,14.584969,14.143571,13.3626375,13.094781,13.124963,13.241914,13.230596,13.264549,13.558814,13.63804,13.45318,13.36641,13.622949,13.487134,13.192869,12.755245,11.962994,11.204697,11.970539,12.3289385,11.861133,11.642321,11.740409,11.234878,10.536942,9.861642,9.201432,9.567377,8.809079,8.405409,8.714764,8.971302,9.4127,9.876732,10.159679,10.18986,10.054046,9.556059,8.386545,7.6886096,7.707473,7.7678347,7.4999785,7.605612,7.77538,7.8131065,7.6282477,7.6886096,7.5792036,7.2924843,7.4773426,9.431562,9.673011,10.823661,13.649357,16.203424,13.822898,16.58446,16.486372,17.486116,19.274342,17.271078,10.853842,5.1534057,1.7165444,0.6111652,0.42630664,0.16976812,0.08677038,0.28294688,0.5357128,0.29049212,0.1659955,0.056589376,0.0,0.0,0.0,0.02263575,0.06790725,0.16976812,0.3169005,0.42630664,0.67152727,0.4376245,0.3772625,0.5394854,0.38103512,0.5281675,0.7469798,0.6149379,0.3961256,1.0676528,1.056335,1.0450171,0.7394345,0.3734899,0.7167987,0.59607476,0.6451189,0.66020936,0.59607476,0.59607476,0.935611,0.9393836,1.2336484,1.599593,0.97710985,2.0258996,2.7841973,3.2821836,3.6669915,4.1800685,4.2404304,4.3309736,4.5120597,4.7044635,4.67051,4.5837393,4.5988297,4.798779,5.0251365,4.8666863,4.610148,4.4630156,4.3724723,4.3007927,4.22534,4.3724723,4.7120085,4.8629136,5.119452,6.439871,6.6850915,7.092535,7.673519,8.314865,8.790216,8.850578,8.171506,7.533932,7.2698483,7.232122,7.647111,7.6584287,7.9036493,8.741172,10.253995,10.646348,12.2270775,13.751218,14.7170105,15.365902,15.803526,14.988639,14.483108,14.2077055,12.449662,11.853588,11.619685,11.729091,11.864905,11.41219,10.729345,10.650121,10.77839,10.838752,10.680302,10.510533,10.70671,11.174516,11.555551,11.216014,10.751981,11.212241,11.766817,12.064855,12.223305,12.672247,13.098554,13.9888935,15.067864,15.275358,16.55428,17.195625,17.354074,17.357847,17.701157,17.882242,17.863379,17.863379,17.569115,16.127972,15.712983,14.969776,14.162435,13.204187,11.642321,10.604849,9.310839,8.382772,8.047009,8.13378,8.401636,8.469543,8.420499,8.231868,7.7829256,7.647111,7.8244243,8.22055,9.408927,12.619431,13.215506,12.00072,9.654147,7.624475,8.14887,10.370946,10.597303,9.699419,9.06939,10.61994,10.412445,9.590013,9.420244,9.808825,9.307066,9.699419,9.676784,9.469289,9.397609,9.87296,10.544487,11.004747,10.759526,10.087999,10.023865,10.868933,11.125471,10.582213,9.895596,10.589758,9.869187,9.525878,9.812597,10.540714,11.076427,10.272858,10.005001,10.661438,11.925267,12.815607,10.291721,11.170743,11.608367,11.18206,12.879742,8.2507305,5.8702044,5.5193505,6.3531003,6.8661776,7.3792543,7.809334,6.911449,5.1798143,4.8365054,3.3350005,6.247467,11.189606,14.483108,11.140562,8.345046,6.620957,4.2894745,1.6524098,0.9922004,2.5917933,3.8895764,4.67051,5.3156285,6.8058157,6.9755836,7.1000805,7.888559,8.959985,8.850578,6.2851934,5.726845,4.9949555,4.0970707,5.2326307,5.4665337,5.149633,4.798779,4.9421387,6.089017,8.492179,9.699419,9.314611,8.054554,7.7376537,9.752235,10.978339,11.1782875,10.499215,9.476834,9.963503,9.446653,9.163706,9.352338,9.231613,7.1679873,7.6131573,8.07719,7.8508325,7.9941926,8.080963,8.137552,8.567632,9.0543,8.590267,8.956212,9.544742,9.812597,10.0276375,11.261286,12.019584,12.940104,12.785426,12.306303,14.237886,17.667202,18.13878,19.58747,21.424738,18.55377,14.709465,12.721292,11.54046,10.842525,11.0613365,9.831461,9.869187,10.529396,11.544232,13.045737,13.313594,12.0724,10.442626,9.461743,10.084227,10.182315,10.042727,10.167224,10.650121,11.200924,11.555551,11.012292,10.804798,11.129244,11.155652,9.540969,9.480607,9.654147,9.552286,9.431562,10.589758,11.027383,10.774617,10.627484,12.128989,13.875714,14.422746,12.932558,10.253995,8.91094,8.8618965,9.261794,9.891823,10.782163,12.223305,11.989402,12.838243,14.151116,15.731846,17.80679,17.440845,14.622695,12.362892,11.457462,10.469034,7.598067,7.0284004,8.299775,10.291721,11.231105,11.41219,10.846297,9.159933,7.6923823,9.476834,9.669238,10.627484,12.0724,12.528888,9.291975,9.231613,7.605612,6.85486,7.3415284,7.356619,8.160188,8.892077,8.563859,8.60913,12.894833,14.003984,13.328684,12.645839,14.237886,20.889025,18.617905,16.32792,10.770844,5.4778514,10.789707,12.253486,12.178034,9.876732,7.001992,7.537705,11.261286,10.929295,9.193887,7.8810134,7.9791017,8.371455,8.058327,7.8432875,7.960239,8.058327,8.98262,9.665465,9.390063,8.360137,7.673519,8.443134,7.7112455,6.960493,6.802043,6.971811,6.349328,6.270103,6.145606,5.6061206,4.4705606,4.3611546,4.82896,4.5535583,3.4142256,2.4861598,2.7804246,2.7615614,2.8294687,3.0558262,3.187868,2.516341,2.8256962,3.1425967,3.1350515,3.097325,4.9534564,4.8968673,4.2404304,4.8440504,9.076936,5.80607,4.9534564,6.009792,7.5905213,7.432071,7.4811153,7.2094865,6.8171334,6.304056,5.462761,6.488915,6.560595,6.907676,7.6508837,7.798016,5.9909286,7.322665,8.080963,6.79827,4.2706113,17.101309,16.32792,9.246704,3.9348478,9.231613,14.260523,16.177015,12.642066,11.959221,33.063286,18.953669,9.303293,4.7912335,6.013564,13.456953,4.644101,3.742444,5.089271,6.043745,6.9567204,7.1038527,5.9494295,6.537959,9.322156,12.193124,11.838497,10.944386,10.676529,11.714001,14.268067,12.057309,11.23865,10.612394,9.955957,10.038955,9.393836,9.352338,8.937348,7.9262853,6.851087,8.888305,10.834979,11.721546,11.072655,8.91094,8.265821,8.52236,8.401636,7.5301595,6.4549613,6.771862,7.4811153,7.805561,7.643338,7.567886,8.83926,8.726082,7.986647,7.4811153,8.179051,8.141325,8.069645,8.137552,8.375228,8.66572,8.922258,9.510788,9.869187,9.831461,9.597558,9.318384,8.45068,7.7301087,7.4169807,7.3075747,6.8435416,6.4926877,6.2361493,6.270103,6.9869013,7.7225633,8.635539,9.812597,11.068882,11.947904,12.242168,12.204442,12.049765,11.736636,10.955703,11.189606,12.242168,13.958713,15.539442,15.565851,15.467763,14.177525,12.932558,12.472299,13.045737,13.679539,12.604341,12.0233555,12.257258,11.732863,10.770844,11.106608,12.283667,13.573905,13.977575,11.242422,9.239159,7.2887115,5.6287565,5.43258,6.0286546,6.379509,7.0774446,7.914967,7.888559,7.413208,6.7643166,6.255012,6.0701537,6.2399216,6.2889657,6.7152724,6.8774953,6.809588,7.1868505,7.7716074,7.5527954,7.277394,7.466025,8.394091,9.673011,10.33322,11.155652,12.045992,12.0082655,12.0082655,12.577931,12.691111,11.947904,10.544487,10.457717,10.684074,11.234878,11.872451,12.113899,13.630494,14.649103,14.305794,12.868423,11.732863,12.81938,13.385274,14.750964,16.248695,15.196134,15.743164,15.803526,15.558306,15.286676,15.120681,15.049001,15.928022,16.32792,16.478827,16.03743,14.064346,13.211733,12.864652,13.011784,13.698401,15.045229,14.958458,14.7321005,14.603831,14.611377,14.581196,13.920986,13.543724,13.072145,12.272349,11.02361,10.521852,10.993429,11.099063,10.63503,10.540714,11.419736,11.932813,12.238396,12.536433,13.072145,12.940104,12.672247,12.762791,13.257004,13.728582,13.970031,13.977575,13.985121,13.951167,13.570132,13.072145,12.883514,13.124963,13.472044,13.155144,12.694883,12.694883,12.838243,12.898605,12.743927,13.019329,13.253232,13.166461,12.81938,12.623203,12.4307995,12.434572,12.034674,11.329193,11.117926,10.736891,10.47658,10.084227,9.556059,9.152389,9.167479,9.152389,8.941121,8.669493,8.790216,9.5032425,10.087999,10.257768,9.940866,9.2995205,8.89585,8.416726,8.009283,7.8319697,8.047009,7.624475,7.454707,7.356619,7.250985,7.164215,7.1378064,6.673774,6.56814,7.3679366,9.382519,10.035183,11.729091,15.256495,18.368912,15.7657995,18.806536,17.40312,16.505234,17.127718,16.346785,9.876732,4.7308717,1.6788181,0.55080324,0.23013012,0.14335975,0.23390275,0.35085413,0.36971724,0.20372175,0.16976812,0.07922512,0.0150905,0.0,0.0,0.003772625,0.049044125,0.15845025,0.271629,0.24522063,0.34330887,0.4678055,0.7205714,0.91674787,0.6149379,0.6526641,0.875249,0.73188925,0.35839936,0.58098423,0.7054809,0.72811663,0.56589377,0.452715,0.9016574,0.83752275,1.026154,1.1921495,1.1996948,1.0827434,1.3770081,1.4034165,1.5467763,1.8070874,1.8184053,2.3126192,2.6068838,2.8558772,3.2746384,4.168751,4.123479,4.104616,4.1612053,4.2404304,4.2064767,4.3347464,4.636556,5.093044,5.4174895,5.0741806,4.644101,4.5196047,4.4743333,4.398881,4.2894745,4.3083377,4.7006907,5.010046,5.3458095,6.3908267,7.0548086,7.443389,7.7225633,8.024373,8.458225,8.345046,7.6207023,7.0963078,7.0170827,7.0359454,6.7869525,6.8963585,7.5527954,8.424272,8.68081,9.733373,10.785934,11.521597,11.92904,12.30253,12.51757,13.000465,12.875969,12.08749,11.41219,11.185833,11.457462,11.6008215,11.355601,10.827434,11.072655,11.106608,10.967021,10.608622,9.910686,9.537196,9.929549,10.344538,10.555805,10.850069,11.204697,12.106354,12.928786,13.385274,13.517315,13.615403,13.434318,13.313594,13.411682,13.687083,15.369675,16.007248,15.803526,15.362129,15.675257,16.452417,18.16519,19.357338,19.342249,18.214233,17.067356,16.177015,15.147089,14.011529,13.230596,11.955449,10.567122,9.424017,8.854351,9.144843,9.473062,9.144843,8.812852,8.635539,8.269594,8.096053,8.431817,9.042982,10.095545,12.14408,15.222542,15.520579,12.800517,8.8769865,7.624475,10.11818,11.393328,10.834979,9.220296,8.729855,8.590267,8.7600355,9.0807085,9.020347,7.6584287,8.880759,10.544487,10.917976,10.125726,10.152134,10.295494,10.412445,10.114408,9.676784,10.038955,10.284176,10.005001,10.03141,10.419991,10.442626,10.18986,10.125726,9.933322,9.831461,10.56335,11.310329,10.872705,10.604849,10.93684,11.34051,12.47607,14.034165,14.396337,12.970284,10.193633,8.182823,6.138061,4.798779,4.659192,5.96452,8.16396,6.673774,6.058836,7.273621,7.643338,9.031664,10.733118,12.830698,12.955194,6.2814207,6.7944975,4.7874613,2.6332922,1.8334957,2.969056,4.6252384,6.296511,7.1679873,7.0774446,6.5228686,5.9230213,6.8661776,8.118689,8.820397,8.495952,6.2361493,4.991183,4.610148,5.040227,6.330465,5.9984736,5.8966126,6.092789,6.5266414,7.039718,8.643084,9.861642,10.11818,9.574923,9.14107,9.220296,9.635284,9.5032425,8.888305,8.778898,8.624221,8.235641,7.8395147,7.7414265,8.3525915,7.4811153,7.99042,8.571404,8.560086,7.9338303,7.7187905,7.515069,7.798016,8.401636,8.541223,9.092027,10.325675,11.385782,11.891314,11.932813,12.913695,13.951167,14.143571,13.928532,15.067864,18.0671,18.961214,20.157135,20.907888,17.297485,15.852571,14.290704,12.811834,11.378237,9.733373,9.242931,9.5183325,10.265312,11.174516,11.921495,11.966766,10.763299,9.95973,10.238904,11.332966,12.31762,12.449662,11.91395,11.208468,11.151879,11.027383,10.657665,10.34831,10.26154,10.435081,10.306811,10.416218,10.680302,11.076427,11.627231,12.925014,13.166461,12.1252165,10.933067,12.095036,13.079691,11.98563,10.227587,8.790216,8.228095,8.412953,9.7069645,11.0613365,12.279895,14.003984,13.890805,14.136025,14.8339615,15.961976,17.391802,16.731592,14.234114,12.336484,11.532914,10.355856,8.446907,7.835742,7.8696957,8.526133,10.423763,10.872705,10.816116,9.854096,8.854351,9.963503,9.552286,9.582467,11.068882,13.407909,14.369928,13.343775,10.638803,8.088508,6.900131,7.6848373,7.1604424,8.265821,8.280911,7.6508837,9.963503,13.026875,13.162688,11.676274,10.099318,10.220041,13.389046,10.521852,6.752999,6.40969,13.008011,13.174006,10.280403,9.857869,11.050018,6.587003,7.914967,8.677037,8.6732645,7.9941926,7.0170827,7.9338303,8.126234,8.296002,8.82417,9.740918,10.650121,11.1631975,10.729345,9.488152,8.284684,8.175279,8.360137,8.114917,7.541477,7.533932,6.8133607,6.2889657,5.564622,4.689373,4.1762958,4.214022,4.689373,4.5309224,3.5839937,2.6106565,2.8256962,2.9237845,3.2859564,3.6179473,2.969056,2.4333432,2.8143783,3.1199608,3.3727267,4.587512,4.636556,3.7801702,3.059599,4.745962,12.351574,9.480607,6.6813188,6.168242,7.466025,7.405663,7.515069,7.6320205,7.3679366,6.881268,6.8774953,7.443389,8.062099,9.261794,10.370946,9.529651,8.054554,9.031664,9.608876,8.499724,5.994701,13.20796,18.983849,20.270313,18.881989,21.473782,35.13823,43.268234,35.821075,23.593996,38.20537,34.561016,20.82489,8.888305,3.863168,4.085753,2.6898816,3.8707132,4.8930945,5.3986263,7.3981175,5.3571277,3.9574835,4.659192,7.284939,10.005001,10.091772,10.370946,10.702937,11.351829,12.985375,10.823661,10.253995,9.906913,9.363655,9.137298,9.107117,9.092027,9.25425,9.125979,7.6320205,9.593785,10.993429,11.076427,9.850324,8.080963,7.6886096,8.016829,7.7301087,6.741681,6.221059,6.8925858,7.3453007,7.5490227,7.5263867,7.3868,8.790216,9.4013815,9.461743,9.333474,9.473062,8.66572,8.52236,8.892077,9.491924,9.910686,10.216269,10.699164,10.993429,10.985884,10.782163,10.265312,9.480607,9.224068,9.288202,8.4544525,7.3188925,6.651138,6.7114997,7.5226145,8.869441,9.8239155,10.47658,11.102836,11.563096,11.287694,11.631002,12.1101265,12.15917,11.815862,11.747954,12.351574,13.162688,14.634012,16.014793,15.343266,15.618668,14.78869,14.279386,14.358611,14.132254,14.143571,13.758763,13.226823,12.853333,12.992921,13.109872,12.5326605,12.287439,12.717519,13.45318,12.1252165,10.612394,8.809079,7.1264887,6.48137,6.6813188,6.7341356,6.7643166,6.8737226,7.1302614,6.273875,5.6891184,5.43258,5.492942,5.7909794,6.356873,6.888813,7.4735703,8.016829,8.246958,7.7301087,7.073672,6.7944975,6.971811,7.24344,7.9225125,8.488406,9.552286,11.031156,12.166716,11.8045435,11.940358,12.242168,12.581704,13.034419,12.276122,12.223305,13.460726,15.369675,16.131744,15.124454,14.4152,14.11339,14.120935,14.124708,14.996184,15.120681,15.554533,16.124199,15.418718,15.475307,15.554533,14.969776,14.758509,15.343266,16.505234,17.139036,17.28994,16.87118,15.901614,14.494425,14.128481,13.920986,14.045483,14.5283785,15.241405,14.807553,15.094273,15.528125,15.62244,14.984866,14.124708,13.736128,13.038192,11.834724,10.533169,10.453944,11.148107,11.053791,10.103089,9.725827,10.642575,11.634775,12.491161,13.13628,13.622949,13.166461,12.864652,13.030646,13.539951,13.800262,14.347293,14.592513,14.543469,14.18507,13.483362,13.20796,13.264549,13.58145,13.853079,13.513543,12.743927,12.555296,12.585477,12.683565,12.898605,12.506252,12.604341,12.857106,13.038192,13.034419,12.992921,12.562841,11.932813,11.23865,10.54826,10.250222,10.012547,9.718282,9.473062,9.57115,9.703192,9.774872,9.710737,9.669238,10.023865,10.453944,10.665211,10.438853,9.835234,9.1825695,8.722309,8.458225,8.303548,8.262049,8.428044,7.745199,7.394345,7.2472124,7.183078,7.0849895,6.9793563,6.3908267,6.247467,6.8699503,7.9489207,8.9788475,11.751727,15.022593,17.56157,18.172735,20.1345,20.281631,20.77962,21.364376,19.346022,11.185833,4.9685473,1.720317,0.97333723,0.7507524,0.5772116,0.6488915,0.6413463,0.482896,0.32067314,0.241448,0.15845025,0.090543,0.0452715,0.0,0.0,0.018863125,0.07922512,0.150905,0.124496624,0.3470815,0.5696664,0.72811663,0.73188925,0.47912338,0.41876137,0.49044126,0.41498876,0.23013012,0.30181,0.56212115,0.68661773,0.7205714,0.77716076,1.0110635,1.3732355,1.6825907,1.7467253,1.6486372,1.780679,2.2258487,2.263575,2.2560298,2.3277097,2.3956168,2.757789,3.0331905,3.410453,3.821669,3.9461658,4.055572,3.8858037,3.8895764,4.0895257,4.0895257,4.2517486,4.52715,4.859141,5.0175915,4.606375,4.406426,4.3347464,4.2592936,4.168751,4.183841,4.429062,4.817642,5.0854983,5.4476705,6.617184,7.5226145,7.8017883,7.858378,7.9526935,8.167733,8.269594,7.937603,7.7716074,7.8206515,7.564113,7.375482,7.673519,8.29223,8.888305,8.937348,9.65792,10.567122,11.329193,11.751727,11.800771,12.019584,12.73261,12.770335,11.853588,10.578441,10.955703,11.272603,11.581959,11.751727,11.457462,11.408418,11.314102,11.031156,10.589758,10.178542,9.646602,10.076681,10.461489,10.570895,10.948157,11.883769,13.0646,14.04171,14.641558,14.984866,14.818871,14.675511,14.02662,13.094781,12.868423,14.173752,15.052773,15.316857,15.211224,15.369675,16.316603,17.91997,19.934551,21.35683,20.432537,17.569115,16.452417,15.460217,14.27184,13.845533,12.940104,11.853588,10.819888,10.069136,9.812597,9.910686,10.001229,9.982366,9.691874,8.89585,9.190115,9.495697,9.850324,10.604849,12.434572,14.735873,16.305285,15.218769,11.955449,9.386291,10.427535,10.170997,9.35611,8.83926,9.608876,8.484633,8.254503,8.337502,8.186596,7.284939,8.118689,9.382519,10.080454,10.310584,11.257513,11.6008215,11.480098,10.695392,9.646602,9.371201,9.661693,9.563604,9.808825,10.299266,10.095545,10.27663,10.253995,10.125726,10.005001,10.023865,10.714255,10.38981,10.329447,10.891568,11.529142,13.140053,15.475307,15.362129,12.898605,11.434827,9.318384,7.213259,5.149633,4.142342,6.187105,7.3075747,5.5382137,6.2097406,9.910686,12.510024,13.204187,11.774363,10.446399,10.076681,10.163452,7.4999785,3.9310753,2.2447119,2.795515,3.4745877,5.59103,6.8397694,7.2283497,6.8737226,6.013564,6.013564,6.858632,7.997965,8.688355,7.986647,6.300284,5.402399,5.1043615,5.4250345,6.6247296,6.187105,5.8588867,6.19465,7.1000805,7.828197,8.243186,9.039209,9.797507,10.121953,9.665465,9.416472,9.608876,9.397609,8.993938,9.695646,8.646856,7.7225633,7.1906233,7.2094865,7.8508325,7.884786,7.99042,8.065872,7.964011,7.488661,7.3151197,7.5565677,7.986647,8.563859,9.435335,10.050273,11.038701,11.978085,12.623203,12.925014,13.573905,13.856852,13.93985,13.8870325,13.664448,14.958458,16.859861,19.063074,20.398582,18.814081,18.12369,17.037174,15.362129,13.238141,11.148107,10.042727,10.110635,10.514306,10.95193,11.623458,11.766817,10.978339,10.831206,11.7026825,12.785426,13.555041,13.604086,13.13628,12.574159,12.54775,11.808316,11.59705,11.996947,12.608112,12.551523,11.895086,11.102836,10.668983,10.86516,11.7555,13.52486,13.396591,12.287439,11.223559,11.363147,11.978085,11.374464,10.54826,9.778644,8.650629,7.7904706,8.624221,9.7220545,10.397354,10.695392,11.52537,12.37421,13.487134,14.943368,16.667458,17.354074,16.192106,14.268067,12.242168,10.340765,9.039209,8.190369,7.665974,7.8508325,9.627739,10.469034,10.023865,9.0957985,8.322411,8.16396,9.21275,9.378746,10.340765,12.411936,14.543469,15.335721,13.245687,10.382264,8.243186,7.665974,6.900131,7.24344,7.5527954,7.828197,9.21275,10.782163,11.25374,11.276376,10.702937,8.597813,9.714509,9.382519,8.537451,7.986647,8.412953,10.736891,9.024119,7.884786,8.296002,7.5829763,7.303802,8.07719,8.254503,7.5792036,7.1793056,7.877241,8.269594,8.6732645,9.322156,10.3634,11.736636,12.419481,12.076173,10.797253,9.114662,8.171506,8.548768,8.748717,8.345046,7.9941926,7.032173,6.4511886,5.783434,4.9534564,4.2706113,4.3347464,4.610148,4.4931965,3.8707132,3.1237335,3.1463692,2.9916916,3.218049,3.62172,3.2255943,2.8785129,2.7389257,2.9652832,3.7499893,5.2892203,4.1762958,3.482133,3.9801195,7.5301595,17.105082,11.959221,7.5527954,6.33801,7.6395655,7.6395655,7.3075747,7.454707,7.3679366,7.2887115,8.439363,8.213005,9.167479,10.227587,10.578441,9.699419,9.971047,10.642575,10.521852,9.371201,7.907422,9.87296,14.396337,19.938324,25.001186,28.132465,39.2768,48.670635,43.6455,31.671186,40.36709,38.062016,19.957186,5.907931,2.2711203,1.8863125,2.2975287,4.0970707,5.4401255,6.277648,8.311093,5.4174895,3.9876647,4.327201,6.2927384,9.314611,8.865668,9.669238,10.382264,10.699164,11.355601,10.035183,9.733373,9.529651,9.024119,8.326183,9.163706,9.307066,9.665465,10.054046,9.163706,11.125471,11.853588,11.019837,9.186342,7.8017883,7.1264887,7.164215,7.1340337,6.888813,6.8963585,7.435844,7.4509344,7.333983,7.201941,6.9265394,8.544995,9.5032425,9.740918,9.608876,9.876732,9.235386,9.0957985,9.363655,9.884277,10.453944,11.034928,11.41219,11.491416,11.249968,10.748209,10.182315,9.846551,9.937095,10.035183,9.118435,7.907422,7.5527954,8.111144,9.171251,9.850324,10.306811,11.080199,11.778135,12.012038,11.408418,11.563096,11.502733,11.54046,11.8045435,12.257258,12.751472,13.151371,14.313339,15.758255,15.690348,15.75071,15.271586,15.301767,16.109108,17.195625,18.229324,18.097282,17.191853,16.075155,15.501716,13.404137,12.645839,12.479843,12.649611,13.404137,12.706201,11.32542,9.774872,8.458225,7.6886096,7.164215,6.809588,6.541732,6.4210076,6.651138,5.8588867,5.3910813,5.27413,5.3194013,5.1345425,6.006019,6.8737226,7.7829256,8.563859,8.82417,8.054554,7.375482,7.284939,7.7037,7.9753294,8.571404,9.205205,10.137043,11.234878,11.959221,11.544232,11.25374,11.472552,12.3893,13.977575,13.626721,12.804289,13.490907,15.652621,17.244669,14.958458,13.86817,14.924504,17.063583,17.195625,19.80251,22.643295,23.303505,20.764528,15.418718,15.211224,15.62244,15.62244,15.701665,16.173243,17.191853,17.63325,17.357847,16.51278,15.445127,14.683057,14.690601,14.683057,14.909414,15.32063,15.588487,15.260268,15.418718,15.603577,15.433809,14.600059,13.981348,13.411682,12.777881,11.962994,10.861387,10.744436,11.193378,11.117926,10.423763,10.038955,10.910432,12.034674,13.128735,13.970031,14.385019,13.958713,13.687083,13.815352,14.177525,14.166207,14.611377,14.841507,14.871688,14.543469,13.532406,13.355092,13.204187,13.230596,13.400364,13.502225,13.004238,12.740154,12.811834,13.091009,13.234368,12.261031,12.219532,12.626976,13.015556,12.943876,12.608112,12.083718,11.570641,11.019837,10.133271,10.050273,9.831461,9.718282,9.81637,10.087999,10.280403,10.359629,10.34831,10.419991,10.872705,11.151879,11.159425,10.661438,9.835234,9.273112,8.571404,8.197914,8.114917,8.197914,8.231868,7.5112963,7.1604424,7.020855,6.934085,6.7567716,6.590776,6.2135134,6.1229706,6.4021444,6.7152724,7.858378,11.2650585,14.532151,16.908905,19.300749,19.48938,20.832436,23.480818,25.733074,24.008986,15.282904,7.2887115,2.4823873,1.0072908,0.70170826,0.663982,0.8111144,0.77716076,0.5281675,0.35085413,0.24899325,0.25276586,0.21881226,0.116951376,0.02263575,0.033953626,0.02263575,0.026408374,0.0754525,0.17354076,0.3961256,0.4640329,0.43385187,0.35462674,0.25276586,0.17354076,0.150905,0.13958712,0.15467763,0.30181,0.8111144,0.91297525,0.9393836,1.1053791,1.5165952,1.8523588,2.1315331,2.203213,2.1994405,2.5087957,2.897376,2.867195,2.795515,2.8181508,2.8219235,3.2557755,3.519859,3.9461658,4.3800178,4.1612053,4.123479,3.85185,3.821669,4.06689,4.1498876,4.3007927,4.436607,4.538468,4.508287,4.164978,4.1272516,4.1498876,4.044254,3.9197574,4.1762958,4.82896,5.2665844,5.572167,6.0776987,7.3981175,8.348819,8.529905,8.412953,8.22055,7.9526935,8.186596,8.518587,8.952439,9.1825695,8.60913,8.650629,8.922258,9.314611,9.639057,9.650374,10.080454,10.748209,11.415963,11.898859,12.064855,12.1101265,12.54775,12.642066,12.038446,10.748209,11.521597,11.827179,11.887542,11.84227,11.732863,11.32542,11.11038,11.004747,10.955703,10.940613,10.570895,10.684074,10.770844,10.729345,10.887795,11.774363,12.759018,13.600313,14.369928,15.47908,15.924251,15.584714,14.252977,12.6345215,12.321393,12.751472,13.837989,14.652876,14.969776,15.23386,16.120426,17.04472,18.953669,20.99843,20.515535,17.942604,17.297485,16.33924,14.713238,13.932304,13.411682,12.611885,11.962994,11.3669195,10.182315,10.042727,10.465261,10.7557535,10.442626,9.250477,9.967276,10.435081,10.993429,11.887542,13.290957,13.951167,15.528125,16.301512,15.494171,13.287186,11.921495,9.763554,8.416726,8.612903,10.246449,8.080963,7.598067,7.745199,7.7904706,7.3377557,7.726336,7.8810134,8.518587,9.831461,11.465008,12.298758,13.083464,12.423254,10.540714,9.280658,9.582467,9.544742,9.684328,9.933322,9.631512,10.0465,9.937095,9.993684,10.216269,9.910686,9.74469,9.537196,9.997457,10.989656,11.548005,12.645839,14.237886,14.683057,13.705947,12.404391,9.854096,8.2507305,6.6624556,5.847569,8.273367,8.069645,7.6697464,9.103344,11.895086,13.087236,10.378491,7.9753294,6.349328,6.3455553,9.1825695,5.956975,3.3463185,2.8143783,3.8141239,3.7914882,6.356873,6.888813,6.651138,6.3455553,6.1003346,6.3945994,7.01331,7.786698,8.167733,7.1981683,6.0814714,5.66271,5.330719,5.1345425,5.772116,5.794752,5.624984,6.1795597,7.405663,8.254503,7.888559,8.379,9.25425,9.8239155,9.144843,9.337247,9.567377,9.337247,9.0807085,10.140816,8.152642,7.0774446,6.7680893,6.9793563,7.3490734,7.5792036,7.4811153,7.3717093,7.326438,7.164215,7.1981683,8.047009,8.624221,8.880759,9.80128,10.216269,10.899114,11.649866,12.355347,12.996693,13.573905,13.238141,12.985375,12.90615,12.215759,12.106354,13.807808,16.320375,18.53868,19.25925,17.961468,17.127718,15.746937,13.936077,12.928786,11.642321,11.148107,11.038701,11.125471,11.434827,11.3971,10.989656,11.400873,12.668475,13.660675,13.441863,13.257004,13.158916,13.355092,14.215251,13.038192,13.124963,14.064346,15.079182,15.049001,13.306048,11.449917,10.484125,10.661438,11.480098,13.555041,13.343775,12.419481,11.589504,10.884023,11.136789,11.52537,12.038446,11.98563,9.982366,8.118689,8.246958,8.586494,8.216777,7.0510364,8.443134,10.242677,12.2119875,13.913441,14.68683,16.4411,16.592005,15.328176,13.298503,11.627231,10.601076,9.322156,8.028146,7.424526,8.677037,9.895596,9.522105,8.763808,7.9753294,6.643593,8.431817,9.088254,9.752235,10.895341,12.313848,13.694629,13.943622,12.083718,8.99771,7.4094353,7.224577,7.0057645,7.250985,8.160188,9.627739,9.97482,10.023865,10.7218,11.442371,9.989911,8.563859,9.242931,9.171251,7.3717093,4.7610526,10.729345,10.280403,7.5527954,5.9418845,8.122461,7.2660756,7.9036493,7.8961043,7.141579,7.594294,7.986647,8.194141,8.52236,9.0957985,9.820143,11.329193,12.045992,12.121444,11.517824,10.03141,8.484633,8.624221,8.865668,8.631766,8.326183,7.24344,6.730363,6.273875,5.6023483,4.666737,4.7308717,4.8666863,4.776143,4.3649273,3.7047176,3.3915899,3.0181,3.1124156,3.5953116,3.8065786,3.7613072,3.0633714,3.0709167,4.0517993,5.172269,3.9122121,3.8820312,4.8666863,7.537705,13.475817,10.061591,7.2170315,6.6134114,7.6697464,7.541477,7.356619,7.364164,7.466025,7.907422,9.295748,8.560086,9.774872,10.518079,10.1294985,9.748463,10.484125,10.751981,10.804798,10.284176,8.20546,9.80128,11.548005,16.807045,24.09953,27.09122,32.13522,37.488575,34.84019,28.619133,36.01725,29.716967,13.306048,3.1048703,2.4522061,1.659955,2.8747404,4.7610526,6.2814207,7.2924843,8.537451,7.073672,7.1906233,6.1531515,4.851596,7.7942433,8.047009,9.190115,10.061591,10.238904,10.023865,9.186342,9.122208,9.295748,9.1825695,8.258276,8.956212,9.325929,9.850324,10.299266,9.737145,11.291467,11.861133,10.880251,8.914713,7.654656,6.5341864,6.330465,6.647365,7.1340337,7.4773426,7.745199,7.4509344,7.2057137,7.0963078,6.6850915,8.186596,9.295748,9.533423,9.208978,9.390063,9.446653,9.601331,9.87296,10.265312,10.744436,11.321648,11.45369,11.2650585,10.876478,10.419991,10.321902,10.34831,10.133271,9.590013,8.903395,8.296002,8.548768,9.446653,10.340765,10.186088,10.3634,11.359374,11.9064045,11.646093,11.114153,11.299012,11.1631975,11.419736,12.185578,12.974057,13.019329,12.706201,13.298503,14.652876,15.252723,15.573396,15.807299,16.31283,17.501207,19.851553,23.126192,23.58645,22.171717,20.741892,22.081175,16.218515,13.211733,12.464753,12.909923,13.011784,12.691111,11.370691,10.008774,9.0543,8.461998,7.484888,6.8699503,6.515323,6.428553,6.730363,6.149379,5.8626595,5.8098426,5.7570257,5.270357,5.8400235,6.7152724,7.6093845,8.314865,8.695901,8.507269,8.047009,8.246958,9.118435,9.767326,10.231359,10.642575,11.102836,11.487643,11.434827,11.000975,10.834979,11.400873,12.600568,13.807808,14.068119,13.317367,13.698401,15.335721,16.335466,14.007756,13.592768,15.878979,19.447882,20.689075,27.600525,37.76775,43.038105,38.080875,20.360857,15.347038,16.177015,17.199398,17.595524,17.335213,17.176762,17.501207,16.735365,15.829934,15.267814,15.033911,15.056546,15.158407,15.486626,15.928022,16.075155,16.248695,15.705438,14.950912,14.324657,14.000212,13.585222,12.736382,12.366665,12.340257,11.476325,11.114153,11.291467,11.589504,11.695138,11.378237,12.049765,12.830698,13.713491,14.494425,14.781145,14.7170105,14.618922,14.698147,14.879233,14.796235,14.8339615,14.803781,14.849052,14.649103,13.419228,13.20796,12.626976,12.272349,12.423254,13.060828,13.151371,13.030646,13.283413,13.70972,13.336229,12.219532,12.102581,12.283667,12.347801,12.140307,11.661184,11.306557,10.989656,10.597303,9.978593,10.061591,9.918231,10.035183,10.374719,10.393582,10.506761,10.718028,10.729345,10.646348,11.000975,11.11038,11.136789,10.559577,9.533423,8.918486,8.047009,7.54525,7.3868,7.3981175,7.273621,6.790725,6.6020937,6.458734,6.258785,6.0211096,5.8588867,5.8211603,5.832478,5.9117036,6.198423,7.0812173,10.303039,13.751218,16.392056,18.293459,17.395575,18.53868,21.798227,25.51049,26.268787,19.021576,10.506761,3.92353,0.6451189,0.181086,0.422534,0.8337501,0.8299775,0.5696664,0.97333723,0.31312788,0.30935526,0.32067314,0.15467763,0.056589376,0.071679875,0.0452715,0.02263575,0.06413463,0.2565385,0.3055826,0.1659955,0.060362,0.060362,0.094315626,0.06413463,0.0754525,0.1358145,0.31312788,0.7092535,1.2223305,1.1129243,1.1091517,1.5203679,2.2409391,2.123988,2.3767538,2.6106565,2.795515,3.2520027,3.2746384,3.1463692,3.1199608,3.2142766,3.218049,3.4934506,3.6745367,4.044254,4.5120597,4.610148,4.1574326,3.8895764,3.8367596,3.9650288,4.1762958,4.3083377,4.3347464,4.266839,4.134797,3.9650288,3.9159849,4.074435,4.0291634,3.9122121,4.38379,5.2967653,5.885295,6.4247804,7.1981683,8.488406,9.424017,9.601331,9.374973,8.884532,8.065872,8.254503,9.027891,9.9257765,10.393582,9.805053,9.793735,9.756008,9.903141,10.144588,10.087999,10.47658,10.748209,10.974566,11.242422,11.642321,11.487643,11.589504,11.695138,11.5857315,11.09529,11.917723,12.257258,11.849815,11.102836,11.129244,10.819888,10.695392,11.00852,11.581959,11.8045435,11.653639,11.1782875,10.751981,10.555805,10.559577,11.012292,11.472552,11.944131,12.7477,14.505743,15.607349,14.84528,13.174006,11.744182,11.910177,11.615912,12.581704,13.5663595,14.147344,14.70192,15.671484,16.252468,17.542706,19.134754,19.123436,18.561316,18.795218,17.674747,15.124454,13.13628,13.170234,12.845788,12.728837,12.419481,10.525623,10.170997,10.56335,10.933067,10.70671,9.495697,10.250222,11.099063,12.264804,13.479589,13.985121,13.434318,14.139798,16.143063,18.289686,18.23687,14.822643,11.129244,8.75249,8.22055,8.990166,6.828451,6.6549106,7.2623034,7.7678347,7.6207023,8.065872,7.3679366,7.61693,9.118435,10.393582,11.302785,13.298503,13.543724,11.717773,10.016319,9.955957,9.533423,9.473062,9.680555,9.246704,9.786189,9.608876,9.820143,10.469034,10.518079,9.64283,9.627739,10.336992,11.129244,10.834979,11.287694,11.61214,13.313594,14.913187,11.955449,9.488152,8.567632,8.114917,8.345046,10.748209,10.661438,11.136789,11.34051,10.552032,8.156415,3.0181,2.0749438,2.5201135,2.7540162,2.3880715,2.8936033,3.308592,4.0178456,4.768598,4.67051,7.1906233,7.1566696,6.5643673,6.488915,7.066127,6.983129,7.4396167,7.748972,7.4999785,6.5568223,6.039973,5.80607,5.43258,4.8553686,4.38379,5.070408,5.5306683,6.432326,7.6697464,8.390318,7.9338303,8.303548,8.89585,9.076936,8.171506,8.809079,9.107117,8.82417,8.461998,9.276885,6.8473144,6.3342376,6.5756855,6.8774953,7.0170827,6.730363,6.63982,6.7869525,7.043491,7.1000805,7.3151197,8.469543,9.088254,8.986393,9.288202,9.514561,10.148361,10.906659,11.581959,12.027128,12.777881,12.438345,12.0082655,11.830952,11.570641,10.974566,11.502733,13.147598,15.343266,17.006994,15.01882,14.456699,13.973803,13.430545,13.902123,13.328684,12.393073,11.830952,11.710228,11.419736,11.034928,10.710483,11.442371,13.072145,14.27184,13.143826,12.619431,12.585477,13.177779,14.758509,13.536179,13.777626,14.577423,15.328176,15.712983,13.694629,11.54046,10.7218,11.272603,11.796998,13.951167,13.909668,12.989148,11.98563,11.18206,11.080199,11.962994,13.29473,13.826671,11.619685,9.650374,9.525878,8.986393,7.352846,5.5004873,6.8473144,9.171251,11.631002,13.079691,12.068627,13.615403,14.494425,14.671739,14.34352,13.951167,12.989148,11.548005,9.371201,7.4018903,7.7829256,9.092027,9.4013815,9.205205,8.397863,6.300284,7.3188925,8.420499,9.258021,9.771099,10.167224,10.325675,12.894833,12.494934,8.956212,7.3377557,8.016829,7.9451485,7.877241,8.348819,9.684328,10.220041,9.733373,9.910686,10.902886,11.310329,9.382519,8.68081,7.352846,5.4438977,4.90064,11.249968,11.5857315,8.843033,6.387054,8.016829,6.990674,7.699928,7.7829256,7.1076255,7.7716074,8.00551,7.8923316,8.088508,8.650629,9.031664,10.061591,10.423763,10.955703,11.502733,10.902886,9.137298,8.76758,8.620448,8.356364,8.473316,7.5565677,7.164215,6.8246784,6.25124,5.342037,5.383536,5.406172,5.2854476,4.9119577,4.1800685,3.5085413,3.0520537,3.1463692,3.7613072,4.52715,4.749735,3.9008942,3.6707642,4.323428,4.689373,4.123479,4.5988297,4.8440504,4.6856003,5.0251365,6.719045,6.530414,6.6586833,7.3717093,7.020855,7.752744,7.7376537,7.9225125,8.567632,9.258021,8.586494,9.665465,10.193633,9.87296,10.38981,9.789962,9.7296,10.838752,11.332966,7.001992,13.200415,13.664448,15.656394,19.817598,20.16468,21.262514,20.655123,18.142553,17.20317,24.99364,16.407146,9.710737,6.0211096,4.2630663,1.1657411,4.323428,6.2399216,7.062354,7.2924843,7.7904706,8.6581745,10.891568,8.318638,3.029418,5.3646727,7.303802,8.741172,9.654147,9.929549,9.352338,8.258276,8.280911,8.944894,9.495697,8.89585,8.627994,9.133525,9.80128,10.008774,9.144843,9.80128,10.589758,10.201178,8.669493,7.3679366,6.1418333,5.8928404,6.3531003,7.115171,7.6395655,7.6320205,7.149124,6.9793563,7.141579,6.8661776,7.8810134,8.892077,9.175024,8.801534,8.639311,9.224068,9.7069645,10.220041,10.725573,11.00852,11.295239,11.189606,10.868933,10.521852,10.352083,10.7557535,10.7557535,9.839006,8.495952,8.231868,8.514814,9.235386,10.140816,10.744436,10.321902,10.47658,11.581959,11.717773,10.714255,10.155907,10.612394,11.11038,11.84227,12.781653,13.694629,13.475817,12.50248,12.23085,12.985375,13.95494,14.988639,15.943113,16.833452,18.168962,20.95316,26.15561,27.453392,25.933023,25.10682,30.92798,21.345512,14.622695,12.464753,13.264549,12.098808,11.989402,10.86516,9.646602,8.816625,8.424272,7.4811153,6.937857,6.771862,6.9265394,7.3000293,6.7643166,6.6624556,6.670001,6.5568223,6.1795597,5.987156,6.379509,6.9680386,7.5716586,8.239413,8.914713,8.710991,9.208978,10.61994,11.819634,11.759273,11.6875925,11.563096,11.336739,10.970794,10.668983,11.02361,12.042219,13.109872,12.996693,13.494679,13.762536,14.600059,15.565851,14.966003,13.230596,13.626721,16.150608,19.828917,22.730066,33.840446,51.662327,64.040306,59.93192,29.36234,15.516807,16.252468,17.320122,17.882242,17.810562,17.701157,17.335213,16.58446,16.094019,16.01102,15.961976,16.0827,16.324148,16.463736,16.376965,16.03743,16.818363,15.79598,14.392565,13.513543,13.551269,13.268322,12.521342,12.064855,11.902632,11.291467,10.963248,11.5857315,12.468526,13.038192,12.815607,12.96274,13.091009,13.713491,14.57365,14.649103,14.4152,14.898096,15.230087,15.275358,15.641303,15.467763,15.418718,15.211224,14.505743,12.894833,12.577931,12.423254,12.400619,12.525115,12.879742,12.940104,13.373956,13.607859,13.422999,12.970284,12.079946,11.555551,11.076427,10.627484,10.469034,11.200924,11.091517,10.729345,10.4049,10.103089,10.370946,10.246449,10.306811,10.518079,10.223814,10.49167,10.789707,10.9594755,11.099063,11.551778,10.47658,10.182315,9.461743,8.171506,7.232122,6.8435416,6.6360474,6.4436436,6.187105,5.8437963,5.6853456,5.66271,5.564622,5.3609,5.20245,5.168496,5.0741806,4.8553686,4.8553686,5.8437963,6.1003346,8.582722,11.02361,12.849561,15.165953,16.01102,16.686321,16.94286,17.538933,20.247679,15.62244,10.812344,5.323174,0.72811663,0.65643674,0.694163,1.478869,1.358145,1.0827434,3.8292143,0.8262049,0.24899325,0.23767537,0.041498873,0.030181,0.018863125,0.00754525,0.00754525,0.011317875,0.0,0.0,0.00754525,0.0150905,0.02263575,0.0452715,0.0452715,0.12826926,0.392353,0.90543,1.7240896,1.1506506,0.7130261,1.2826926,2.4107075,2.3503454,2.203213,2.916239,3.1614597,3.059599,4.1800685,3.7047176,3.640583,3.7009451,3.7273536,3.6934,2.9237845,3.2633207,3.8669407,4.244203,4.255521,3.7462165,3.6179473,3.5500402,3.5424948,3.9197574,3.9461658,3.9801195,3.8707132,3.682082,3.7084904,3.7688525,4.104616,4.2706113,4.3121104,4.776143,5.3382645,6.126743,7.066127,8.088508,9.125979,10.284176,10.582213,10.423763,9.933322,8.956212,9.261794,9.393836,9.869187,10.54826,10.63503,9.952185,9.450426,9.420244,9.797507,10.163452,10.148361,10.238904,10.152134,9.835234,9.446653,9.737145,9.782416,9.869187,9.850324,9.156161,9.839006,10.072908,9.903141,9.703192,10.178542,10.287949,10.63503,11.276376,12.034674,12.513797,11.853588,10.853842,10.121953,9.95973,10.374719,10.887795,11.099063,11.2650585,11.589504,12.223305,11.589504,11.11038,11.016065,11.336739,11.887542,12.019584,12.193124,12.800517,13.698401,14.173752,15.958203,17.071129,18.58395,20.115637,19.821371,19.444109,19.613878,18.02183,14.354838,10.314357,11.962994,13.117417,13.494679,12.917468,11.306557,10.56335,10.914205,11.276376,11.091517,10.359629,10.627484,11.759273,12.894833,13.487134,13.290957,12.14408,12.853333,15.546988,19.312067,22.21699,18.968758,13.358865,8.695901,6.319147,5.583485,5.6589375,5.6476197,6.2663302,7.484888,8.560086,9.559832,8.812852,8.567632,9.159933,9.001483,8.563859,9.424017,10.627484,11.332966,10.834979,9.989911,8.967529,9.050528,9.846551,9.246704,10.137043,10.114408,10.570895,11.6008215,11.993175,11.638548,12.3289385,12.6345215,11.872451,10.103089,9.295748,11.438599,13.008011,12.808062,11.978085,9.416472,7.6093845,6.971811,7.7225633,9.918231,12.272349,8.82417,4.376245,1.7240896,1.6637276,1.5052774,0.94315624,0.5998474,0.7922512,1.50905,4.2706113,5.05909,5.50426,6.1229706,6.330465,7.748972,7.707473,7.4169807,7.624475,8.650629,8.443134,8.428044,8.141325,7.54525,7.020855,7.4697976,7.2094865,6.8246784,6.1041074,4.0291634,4.7346444,5.66271,6.63982,7.594294,8.560086,8.473316,8.526133,8.612903,8.552541,8.088508,8.477088,8.76758,8.3525915,7.5301595,7.5075235,5.994701,6.3832817,7.0548086,7.3453007,7.5527954,6.466279,5.956975,6.085244,6.6247296,7.066127,7.1981683,7.9941926,8.639311,8.809079,8.650629,9.408927,10.065364,10.70671,11.159425,11.000975,11.344283,11.529142,11.657412,11.646093,11.231105,10.729345,11.363147,11.955449,12.196897,12.649611,12.174261,12.657157,13.487134,14.124708,14.0983,14.305794,13.8719425,13.140053,12.506252,12.419481,12.347801,11.706455,12.151625,13.966258,16.06761,15.445127,14.335975,13.298503,12.672247,12.574159,11.793225,11.321648,11.291467,11.732863,12.58925,12.355347,11.631002,11.710228,12.604341,13.030646,15.448899,15.282904,13.751218,12.242168,12.3289385,12.31762,12.826925,13.343775,13.404137,12.574159,11.7555,12.136535,10.868933,7.9300575,6.149379,7.6018395,9.329701,10.853842,11.619685,10.970794,10.982111,11.921495,13.434318,14.924504,15.546988,14.694374,14.279386,12.185578,8.903395,7.537705,8.269594,8.7751255,9.201432,8.888305,6.349328,6.3116016,7.7225633,8.892077,9.495697,10.544487,10.555805,11.9064045,11.9064045,10.084227,8.179051,9.190115,9.665465,9.540969,8.778898,7.3415284,8.024373,8.488406,9.408927,10.884023,12.419481,10.054046,8.518587,7.4509344,6.779407,6.7454534,2.6936543,6.119198,8.126234,7.224577,9.322156,7.0284004,7.7640624,8.348819,7.858378,7.6131573,7.6131573,7.6584287,8.299775,9.363655,9.948412,10.106862,9.680555,10.076681,11.234878,11.61214,10.099318,9.024119,8.311093,8.0206,8.360137,7.9338303,7.84706,7.541477,6.9189944,6.330465,6.247467,5.87775,5.492942,5.119452,4.5460134,3.7160356,3.1048703,3.199186,4.0291634,5.1873593,5.27413,5.0213637,4.8440504,4.8365054,4.776143,5.0213637,4.9723196,4.304565,4.4894238,8.7751255,10.982111,7.5263867,5.6778007,6.8246784,6.470052,8.179051,8.643084,8.586494,8.537451,8.820397,8.722309,8.495952,8.68081,9.646602,11.61214,9.525878,9.718282,11.389555,11.808316,6.3153744,17.7917,18.225552,17.463482,17.625704,13.106099,16.305285,14.928277,12.30253,10.536942,10.514306,11.638548,20.255224,18.485863,6.221059,1.1280149,7.062354,8.937348,7.5301595,5.349582,6.670001,7.0472636,8.578949,6.541732,2.4710693,4.1800685,6.0626082,7.594294,8.650629,9.216523,9.397609,7.6886096,7.466025,8.130007,9.042982,9.507015,9.092027,9.371201,9.846551,9.876732,8.66572,8.288457,8.714764,8.710991,7.9036493,6.8058157,6.439871,6.2361493,6.3908267,6.930312,7.7376537,7.3717093,6.5002327,6.2361493,6.779407,7.4169807,7.854605,8.258276,8.601585,8.835487,8.89585,8.846806,8.937348,9.650374,10.740664,11.216014,11.434827,11.555551,11.510279,11.25374,10.740664,10.3634,9.80128,8.831716,7.937603,8.314865,8.963757,9.435335,10.035183,10.676529,10.895341,10.393582,11.404645,11.619685,10.484125,9.216523,9.789962,10.612394,11.653639,12.740154,13.536179,14.109617,13.392818,12.102581,11.427281,13.015556,14.079436,14.600059,15.588487,17.572887,20.598532,24.774828,26.212198,25.767029,26.883726,35.61358,23.797718,15.943113,13.358865,13.72481,11.125471,10.710483,10.0465,9.129752,8.13378,7.4018903,6.828451,6.7944975,7.3868,8.118689,7.9338303,6.971811,6.911449,7.0510364,7.0359454,6.851087,6.1305156,5.775889,6.1003346,7.092535,8.424272,9.156161,9.027891,9.748463,11.574413,13.321139,12.283667,11.970539,11.555551,11.042474,11.276376,11.778135,12.178034,12.427027,12.434572,12.068627,12.166716,13.272095,14.852824,15.992157,15.380992,13.634267,13.426772,14.958458,17.591751,19.836462,29.052984,44.852737,59.811195,62.10118,35.477764,16.090246,16.052519,16.4826,16.912678,17.101309,17.040947,17.682293,16.588232,15.603577,15.328176,15.143317,15.656394,15.935568,15.935568,15.777118,15.754482,15.55076,15.335721,15.184815,15.071637,14.905642,14.339747,13.747445,12.826925,11.861133,11.717773,11.9064045,12.344029,12.770335,13.04951,13.170234,13.600313,13.853079,14.347293,15.079182,15.599804,16.305285,17.037174,17.123945,16.622187,16.335466,16.097792,15.829934,15.505488,14.969776,13.943622,14.075664,14.739646,15.188588,15.033911,14.245432,14.249205,13.841762,13.430545,13.109872,12.691111,11.623458,11.41219,11.091517,10.552032,10.540714,11.106608,11.219787,11.087745,10.850069,10.552032,10.54826,10.4049,10.382264,10.419991,10.125726,10.257768,10.269085,10.70671,11.299012,10.989656,10.18986,9.397609,8.329956,7.141579,6.428553,5.6551647,5.142088,4.8063245,4.538468,4.195159,4.183841,4.134797,4.104616,4.0517993,3.8367596,3.6254926,3.7084904,3.7914882,4.063117,5.198677,5.455216,9.024119,11.246195,11.92904,15.362129,15.414946,17.093763,16.893814,14.754736,14.083209,9.125979,5.73439,2.6974268,0.271629,0.181086,0.14713238,0.38480774,0.38480774,0.271629,0.80356914,0.211267,0.7582976,0.9205205,0.38103512,0.018863125,0.00754525,0.0,0.0,0.003772625,0.011317875,0.003772625,0.08299775,0.116951376,0.071679875,0.00754525,0.5470306,0.7922512,0.97710985,1.1016065,0.94315624,0.62248313,1.297783,2.1956677,2.7615614,2.6295197,2.9237845,3.229367,3.5047686,3.6934,3.7047176,3.1614597,2.9841464,2.7879698,2.474842,2.252257,2.4408884,3.31991,3.8292143,3.802806,3.953711,3.712263,3.8065786,3.7348988,3.4632697,3.4217708,2.9954643,3.270866,3.6028569,3.640583,3.3048196,3.3350005,3.6934,4.2102494,4.7912335,5.409944,6.058836,6.6020937,7.1038527,7.647111,8.329956,9.548513,10.223814,10.457717,10.284176,9.639057,9.778644,9.937095,10.269085,10.597303,10.378491,10.0276375,9.857869,9.424017,9.009028,9.650374,9.461743,9.329701,9.416472,9.612649,9.540969,9.307066,9.771099,10.170997,10.114408,9.593785,9.027891,8.797762,8.669493,8.616675,8.809079,9.261794,9.608876,10.242677,11.125471,11.766817,11.3820095,10.789707,10.397354,10.303039,10.27663,10.148361,10.465261,10.914205,11.461235,12.370438,12.513797,12.355347,11.883769,11.544232,12.242168,12.921241,13.558814,14.249205,15.143317,16.45619,17.067356,16.7995,17.139036,18.421728,19.794964,18.704676,16.048746,12.457208,9.246704,8.397863,12.08749,13.875714,14.302021,13.864397,13.004238,11.898859,11.774363,11.744182,11.487643,11.2650585,11.902632,12.570387,12.887287,12.800517,12.543978,12.951422,13.917213,15.984612,18.16519,17.946377,20.730574,17.904879,12.887287,8.669493,7.8319697,7.356619,6.304056,5.9720654,6.5530496,7.118943,8.646856,9.337247,10.416218,11.747954,11.834724,11.083972,10.401127,9.967276,10.03141,10.906659,9.899368,9.016574,8.929804,9.348565,9.016574,9.593785,9.906913,10.570895,11.415963,11.506506,11.133017,12.095036,12.872196,12.37421,9.929549,8.695901,10.416218,10.299266,7.7904706,6.571913,5.6778007,4.5460134,4.214022,4.938366,6.205968,6.307829,4.4177437,2.6295197,1.9202662,2.1503963,1.3694628,1.418507,1.7655885,2.5012503,4.353609,6.156924,6.9567204,7.7829256,8.390318,7.2585306,8.492179,8.59404,8.013056,7.3717093,7.4811153,7.066127,7.1340337,6.964266,6.571913,6.700182,7.0170827,7.3717093,7.220804,6.360646,4.919503,4.9723196,6.0512905,6.8246784,7.2358947,8.511042,8.612903,8.299775,7.9828744,7.748972,7.356619,7.707473,7.7376537,7.322665,6.6850915,6.398372,5.9682927,6.436098,6.930312,7.2283497,7.798016,7.0510364,6.187105,5.6513925,5.5570765,5.6853456,6.2021956,6.971811,7.537705,7.7301087,7.6886096,8.024373,8.386545,9.205205,10.201178,10.355856,10.246449,10.359629,10.54826,10.574668,10.084227,9.669238,10.27663,11.042474,11.649866,12.306303,13.63804,15.99593,17.172989,16.395828,14.332202,14.539697,14.434063,14.094527,13.528633,12.702429,13.739901,14.762281,15.388537,15.648849,15.9695215,15.716756,14.864142,14.279386,13.966258,13.04951,11.68382,11.227332,11.106608,11.272603,12.185578,12.736382,12.5326605,12.513797,12.838243,12.883514,14.694374,14.637785,13.441863,12.249713,12.596795,12.381755,11.936585,11.46878,11.2801485,11.766817,11.231105,10.917976,10.099318,8.827943,7.8961043,8.333729,9.408927,11.019837,12.506252,12.679792,11.8045435,11.257513,11.465008,11.959221,11.3971,11.676274,13.140053,13.59654,12.117672,9.050528,7.986647,7.9828744,8.805306,9.250477,7.141579,6.6549106,7.424526,8.069645,8.635539,10.604849,10.79348,11.498961,11.498961,10.899114,11.133017,10.827434,8.933576,7.8810134,8.047009,7.779153,7.956466,8.963757,9.695646,10.582213,13.604086,12.427027,11.5857315,10.159679,8.329956,7.352846,5.1760416,7.9451485,9.273112,8.156415,8.956212,7.677292,7.911195,8.235641,8.160188,8.152642,7.877241,7.7904706,7.726336,7.8696957,8.729855,10.0276375,10.31813,10.159679,10.050273,10.438853,9.601331,8.612903,7.9489207,7.914967,8.66572,8.054554,8.103599,8.07719,7.677292,7.0510364,6.6360474,6.058836,5.6476197,5.3759904,4.8402777,4.398881,4.1310244,4.217795,4.610148,5.0175915,5.0553174,5.119452,5.323174,5.6061206,5.7419353,6.149379,5.0062733,3.6066296,3.663219,7.322665,9.952185,7.0887623,5.621211,7.0548086,7.5188417,8.2507305,8.375228,8.122461,7.6886096,7.2585306,8.29223,9.031664,9.337247,9.491924,10.197406,9.0957985,10.597303,11.027383,9.861642,9.710737,16.87118,18.274595,15.660167,11.864905,10.823661,15.75071,15.603577,15.848798,17.093763,15.067864,13.094781,29.181253,36.266243,24.506971,1.2751472,4.006528,5.492942,4.8327327,3.7198083,6.4247804,6.273875,7.484888,5.983383,2.9539654,4.82896,5.7419353,7.0887623,8.356364,9.084481,8.888305,8.084735,8.073418,8.484633,9.186342,10.27663,10.170997,9.850324,9.993684,10.265312,9.288202,8.518587,8.944894,8.975075,8.031919,6.571913,6.149379,6.519096,7.020855,7.364164,7.6131573,7.1679873,6.6247296,6.6020937,7.0849895,7.4282985,8.122461,8.571404,8.710991,8.703445,8.967529,9.537196,10.050273,10.597303,11.18206,11.714001,12.012038,12.166716,12.095036,11.853588,11.646093,10.416218,8.692128,7.443389,7.1566696,7.828197,8.661947,9.393836,10.069136,10.604849,10.785934,10.438853,10.419991,10.18986,9.661693,9.190115,9.288202,10.178542,11.23865,12.151625,12.925014,13.283413,12.491161,11.498961,11.065109,11.732863,11.751727,12.479843,13.664448,14.947141,15.875206,17.599297,18.806536,18.980076,19.21398,22.213217,16.418465,13.792717,13.109872,12.774108,10.819888,10.774617,10.336992,9.171251,7.6584287,6.8774953,6.537959,6.428553,6.8359966,7.5716586,7.9941926,7.273621,7.322665,7.696155,7.937603,7.5603404,6.477597,6.0701537,6.1041074,6.5756855,7.6886096,9.850324,10.238904,10.314357,10.7557535,11.465008,11.932813,12.559069,12.510024,11.910177,11.849815,12.525115,12.566614,11.879996,11.11038,11.642321,12.483616,13.068373,13.947394,14.777372,14.332202,13.189097,12.898605,13.675766,15.158407,16.418465,19.240387,23.692085,27.159128,26.449873,17.814335,16.70141,15.739391,15.863888,16.199652,16.452417,16.931541,17.301258,17.37671,17.18808,16.58446,15.267814,14.539697,14.049255,13.717264,13.664448,14.1926155,14.517061,14.490653,14.441608,14.584969,15.022593,14.815099,13.905896,12.917468,12.362892,12.67602,12.453435,12.464753,12.789199,13.396591,14.18507,14.1926155,14.373701,14.811326,15.467763,16.16947,17.297485,18.018057,17.799244,16.905132,16.41092,15.931795,15.618668,15.475307,15.347038,14.901869,15.430037,16.090246,16.331694,15.935568,14.999957,14.124708,13.324911,12.913695,12.687338,11.9064045,11.6008215,11.548005,11.114153,10.47658,10.642575,10.997202,11.2650585,11.348056,11.174516,10.7218,10.770844,10.567122,10.423763,10.336992,10.001229,9.805053,10.005001,10.34831,10.438853,9.733373,8.888305,7.9413757,6.858632,5.828706,5.27413,4.5912848,3.9574835,3.4368613,3.0671442,2.8407867,2.8294687,2.8106055,2.8596497,2.9313297,2.8521044,2.6408374,2.7426984,3.0105548,3.5085413,4.5120597,5.1156793,8.541223,10.280403,10.733118,15.192361,13.604086,14.003984,14.120935,12.792972,9.95973,6.25124,3.8178966,1.8561316,0.35462674,0.07922512,0.02263575,0.049044125,0.056589376,0.026408374,0.018863125,0.02263575,0.46026024,0.5470306,0.20372175,0.02263575,0.018863125,0.02263575,0.018863125,0.011317875,0.0150905,0.003772625,0.28294688,0.4376245,0.52439487,1.0601076,1.2336484,1.056335,1.0714256,1.3468271,1.478869,1.6184561,2.191895,2.9011486,3.3727267,3.1765501,3.440634,3.3010468,3.2482302,3.3236825,3.1010978,2.6710186,2.4295704,2.1353056,1.8636768,1.9844007,2.3088465,2.8445592,3.180323,3.2218218,3.2067313,3.2255943,3.2633207,3.3727267,3.470815,3.3689542,2.8822856,2.9200118,3.1840954,3.3915899,3.2784111,3.4557245,3.6745367,4.06689,4.7572803,5.8626595,6.7454534,7.3075747,7.605612,7.8734684,8.499724,9.5183325,10.012547,9.986138,9.684328,9.582467,10.450171,10.552032,10.661438,10.819888,10.314357,10.038955,9.601331,9.042982,8.597813,8.669493,9.242931,9.408927,9.5183325,9.650374,9.6051035,9.348565,9.612649,9.865415,9.710737,8.888305,8.341274,8.314865,8.397863,8.439363,8.560086,8.937348,9.295748,9.774872,10.367173,10.914205,10.536942,10.035183,9.597558,9.307066,9.175024,9.114662,9.393836,9.993684,10.785934,11.52537,12.00072,11.68382,11.16697,10.989656,11.642321,12.366665,13.7700815,15.603577,17.448391,18.731083,17.89356,17.18808,16.859861,17.172989,18.417955,18.765038,15.894069,11.336739,7.699928,8.631766,12.596795,14.664193,15.467763,15.460217,14.894323,13.521088,13.019329,12.849561,12.585477,11.902632,10.797253,11.034928,11.672502,12.283667,12.936331,13.313594,13.592768,14.634012,16.120426,16.546734,19.153618,18.229324,14.475562,10.114408,8.903395,7.6508837,6.5455046,6.273875,6.7114997,6.952948,8.428044,9.582467,10.642575,11.578186,12.121444,12.543978,11.52537,10.038955,9.092027,9.733373,9.2844305,8.692128,8.345046,8.356364,8.563859,9.325929,9.661693,10.110635,10.876478,11.793225,11.7026825,11.649866,11.895086,11.657412,9.144843,9.186342,9.461743,8.552541,6.466279,4.640329,3.2444575,4.4403796,5.8702044,6.7114997,7.696155,3.5651307,2.3390274,2.263575,2.546522,3.3727267,2.6672459,2.4295704,2.8521044,4.123479,6.4210076,7.2660756,8.235641,9.333474,9.914458,8.68081,8.605357,8.699674,8.382772,7.6886096,7.2962565,7.175533,7.122716,6.79827,6.330465,6.2927384,6.258785,6.7831798,7.2358947,7.2660756,6.790725,6.300284,6.673774,7.454707,8.269594,8.809079,7.5565677,7.1302614,7.069899,7.069899,6.960493,7.1264887,6.930312,6.417235,5.8173876,5.515578,5.926794,6.7077274,7.3075747,7.4811153,7.3000293,6.617184,5.956975,5.4665337,5.2099953,5.149633,5.832478,6.507778,7.1076255,7.5112963,7.5188417,7.1566696,7.201941,7.914967,8.907167,9.129752,9.393836,9.948412,10.340765,10.34831,9.952185,9.525878,9.793735,10.408672,11.1631975,12.012038,13.588995,14.988639,15.724301,15.55076,14.490653,14.57365,13.675766,13.030646,12.894833,12.525115,13.389046,14.777372,15.720529,15.807299,15.184815,13.951167,13.302276,13.555041,14.3095665,14.460471,12.483616,11.133017,10.3634,10.265312,11.02361,12.1252165,12.574159,12.796744,13.0646,13.498452,14.3095665,13.920986,13.072145,12.411936,12.491161,12.310076,11.581959,10.668983,10.038955,10.246449,10.012547,9.597558,9.4013815,9.431562,9.318384,9.378746,10.352083,11.498961,12.200669,11.925267,11.646093,10.974566,10.714255,10.79348,10.26154,10.49167,12.162943,13.981348,14.600059,12.615658,9.540969,8.167733,8.518587,9.261794,7.707473,6.9982195,7.3981175,7.643338,7.8395147,9.457971,10.069136,10.427535,10.061591,9.408927,9.820143,9.148616,7.6018395,7.1604424,7.835742,7.6697464,7.673519,8.737399,9.424017,10.095545,12.940104,11.766817,11.2801485,10.3634,8.858124,7.564113,9.420244,12.6345215,12.842015,10.238904,9.590013,8.035691,7.3717093,7.4207535,7.8131065,8.001738,7.8206515,8.031919,7.9413757,7.6923823,8.231868,9.684328,9.857869,9.224068,8.537451,8.846806,8.578949,8.062099,7.6508837,7.752744,8.82417,8.333729,8.265821,8.329956,8.29223,8.001738,7.3113475,6.5228686,5.9720654,5.6325293,5.149633,5.191132,4.983638,4.889322,4.938366,4.8365054,4.817642,4.817642,5.0138187,5.481624,6.1908774,6.571913,5.4288073,3.7914882,5.010046,14.728328,14.102073,9.258021,6.515323,7.394345,8.616675,7.7187905,8.001738,8.171506,7.6923823,6.7643166,7.6093845,8.299775,8.809079,9.303293,10.125726,9.899368,10.880251,10.63503,9.608876,11.136789,13.20796,12.845788,10.797253,8.805306,9.58624,10.872705,9.778644,11.45369,16.071383,18.821627,13.140053,21.96045,26.438557,18.48209,0.7432071,2.916239,3.9084394,3.6066296,3.0030096,4.2027044,6.066381,6.4926877,6.330465,5.794752,4.466788,5.323174,7.073672,8.612903,9.333474,9.0957985,8.43559,8.635539,8.963757,9.318384,10.220041,9.97482,9.65792,9.97482,10.672756,10.533169,9.87296,9.673011,9.21275,8.239413,6.971811,6.511551,6.7869525,7.24344,7.4999785,7.356619,6.8963585,6.771862,6.9567204,7.24344,7.2094865,8.246958,8.99771,9.216523,9.039209,9.005256,9.952185,10.804798,11.32542,11.653639,12.298758,12.864652,13.140053,12.702429,11.672502,10.691619,9.967276,8.314865,7.115171,7.0246277,7.99042,8.537451,9.405154,10.235131,10.725573,10.638803,10.370946,9.918231,9.57115,9.239159,8.480861,8.258276,8.922258,9.929549,10.974566,11.993175,12.438345,12.068627,11.510279,11.0613365,10.680302,10.672756,11.661184,12.668475,13.340002,13.936077,14.517061,15.290449,15.456445,15.17727,15.592259,14.4114275,13.826671,13.456953,12.826925,11.348056,10.902886,10.310584,9.231613,7.8319697,6.790725,6.7454534,6.7379084,7.0849895,7.7225633,8.194141,7.865923,7.865923,8.00551,7.914967,7.0510364,6.2889657,6.228604,6.3342376,6.677546,7.937603,9.748463,10.284176,10.231359,10.152134,10.480352,11.306557,12.366665,13.041965,13.158916,12.981603,13.158916,13.004238,12.525115,12.132762,12.6345215,13.204187,13.27964,13.392818,13.739901,14.188843,13.000465,12.611885,13.079691,13.88326,13.943622,14.667966,15.671484,16.078928,15.264041,12.883514,16.177015,15.060319,15.188588,15.535669,15.82239,16.524097,16.991903,17.542706,17.53516,16.720274,15.226315,14.211478,13.430545,12.872196,12.751472,13.50977,14.796235,14.977322,14.498198,14.049255,14.577423,14.694374,13.875714,13.226823,13.177779,13.494679,12.713746,12.483616,12.898605,13.860624,15.113135,15.071637,15.124454,15.260268,15.592259,16.346785,17.267305,17.870924,17.72002,17.010767,16.603323,15.82239,15.4074,15.252723,15.252723,15.309312,16.309057,16.859861,16.833452,16.21097,15.098045,13.630494,12.868423,12.528888,12.2119875,11.41219,11.204697,11.242422,10.963248,10.521852,10.79348,11.140562,11.291467,11.246195,10.978339,10.47658,10.702937,10.536942,10.370946,10.227587,9.763554,9.416472,9.454198,9.408927,9.001483,8.156415,7.3490734,6.48137,5.485397,4.496969,3.863168,3.1916409,2.584248,2.123988,1.8485862,1.7542707,1.780679,1.7882242,1.8334957,1.8938577,1.871222,1.7957695,1.8146327,2.022127,2.463524,3.127506,4.1762958,7.443389,9.156161,9.612649,13.200415,11.461235,11.004747,11.763044,12.223305,9.431562,8.688355,7.062354,4.134797,0.97333723,0.1358145,0.049044125,0.026408374,0.02263575,0.0150905,0.00754525,0.0150905,0.124496624,0.150905,0.10186087,0.1659955,0.30935526,0.3470815,0.392353,0.44894236,0.4074435,0.46026024,0.935611,1.1544232,1.1581959,1.690136,1.3468271,1.3392819,1.7580433,2.2862108,2.2069857,2.5691576,2.7200627,3.0822346,3.4255435,2.8407867,3.1539145,2.9803739,2.886058,2.9916916,2.9766011,2.493705,2.3692086,2.1994405,2.0447628,2.4295704,2.5767028,2.6106565,2.7728794,2.938875,2.6031113,2.9992368,2.9124665,3.199186,3.8254418,3.85185,3.2255943,2.848332,2.9200118,3.2784111,3.4255435,3.5877664,3.7084904,3.8405323,4.3196554,5.772116,6.6020937,7.3490734,7.956466,8.567632,9.5183325,9.978593,9.944639,9.654147,9.450426,9.797507,10.529396,10.457717,10.431308,10.495442,9.869187,9.676784,9.276885,8.820397,8.397863,8.028146,8.907167,9.318384,9.533423,9.623966,9.450426,9.129752,9.167479,9.171251,8.8769865,8.175279,8.062099,8.356364,8.582722,8.601585,8.650629,9.167479,9.703192,10.246449,10.687846,10.804798,10.325675,9.759781,9.291975,8.990166,8.7751255,8.812852,9.107117,9.665465,10.310584,10.672756,11.1782875,10.808571,10.427535,10.453944,10.834979,11.461235,13.038192,15.562078,18.30855,19.828917,19.183798,18.591496,17.50498,16.4411,16.954176,18.082191,16.780636,13.196642,9.590013,10.31813,12.917468,14.351066,14.962231,15.079182,15.052773,14.43029,14.079436,13.807808,13.181552,11.510279,9.88805,10.201178,11.208468,12.166716,12.857106,13.290957,13.147598,13.498452,14.584969,15.833707,16.271332,16.135517,14.305794,11.461235,10.084227,8.329956,7.224577,6.9944468,7.3151197,7.3188925,8.620448,10.020092,10.834979,11.11038,11.627231,12.89106,12.483616,11.012292,9.4013815,8.91094,8.707218,8.243186,7.677292,7.3792543,7.9338303,8.873214,9.148616,9.529651,10.352083,11.532914,11.721546,10.612394,10.370946,10.808571,9.348565,11.02361,9.367428,7.484888,5.994701,3.0105548,3.5085413,5.674028,7.54525,8.179051,7.635793,2.886058,1.9655377,2.5540671,3.4481792,4.5799665,4.285702,4.0480266,4.459243,5.7570257,7.8319697,8.069645,9.088254,10.310584,10.861387,9.590013,8.299775,8.065872,8.058327,7.964011,7.9941926,7.9451485,7.201941,6.56814,6.300284,6.0776987,5.723072,6.187105,6.9793563,7.5792036,7.443389,6.673774,6.628502,7.424526,8.345046,7.835742,6.19465,6.1833324,6.5266414,6.6813188,6.832224,6.9189944,6.5832305,6.0211096,5.5683947,5.6551647,6.1305156,6.7680893,7.432071,7.745199,7.073672,6.187105,5.481624,5.1043615,5.036454,5.081726,5.802297,6.470052,7.152897,7.7376537,7.8961043,7.232122,6.9755836,7.375482,8.182823,8.631766,9.137298,9.771099,10.137043,10.076681,9.646602,9.239159,9.314611,9.793735,10.514306,11.25374,12.472299,12.796744,13.336229,14.203933,14.532151,15.17727,13.721037,12.551523,12.427027,12.457208,12.898605,14.068119,15.203679,15.79598,15.607349,13.158916,12.30253,12.766563,13.966258,15.00373,13.355092,11.593277,10.38981,10.008774,10.310584,11.02361,11.868678,12.513797,13.038192,13.962485,13.943622,13.434318,12.875969,12.453435,12.08749,11.800771,11.314102,10.589758,9.80128,9.337247,9.012801,8.91094,9.261794,9.955957,10.578441,10.61994,11.423509,11.793225,11.480098,11.18206,11.793225,11.068882,10.495442,10.453944,10.231359,10.397354,11.661184,13.532406,15.026365,14.66042,11.385782,8.922258,8.345046,9.005256,8.548768,7.809334,7.707473,7.726336,7.8508325,8.537451,9.246704,9.6051035,9.442881,8.986393,8.850578,8.07719,7.032173,7.0510364,7.8621507,7.6018395,7.6207023,8.669493,9.310839,9.81637,12.151625,11.091517,10.642575,10.506761,10.33322,9.710737,11.740409,14.154889,13.743673,10.842525,9.318384,7.854605,6.5945487,6.379509,7.115171,7.786698,7.7942433,8.160188,8.29223,8.197914,8.492179,9.416472,9.382519,8.571404,7.6395655,7.7301087,7.7640624,7.8131065,7.7112455,7.756517,8.703445,8.484633,8.360137,8.480861,8.786444,8.990166,8.201687,7.352846,6.752999,6.3531003,5.7494807,5.772116,5.455216,5.2062225,5.0666356,4.689373,4.7233267,4.610148,4.696918,5.2250857,6.326692,5.987156,5.624984,4.3083377,5.6891184,18.010511,17.323895,11.974312,7.91874,7.4018903,8.952439,7.352846,7.7338815,8.265821,8.035691,7.069899,7.6282477,8.137552,8.726082,9.439108,10.212496,9.963503,10.382264,10.435081,10.208723,10.917976,10.238904,9.114662,8.582722,8.582722,7.937603,6.5643673,5.6589375,7.3113475,11.706455,17.13149,12.404391,14.683057,14.441608,8.616675,0.6111652,3.5236318,4.093298,3.7084904,4.4139714,8.907167,12.313848,10.49167,8.986393,8.627994,5.511805,5.4740787,7.454707,9.208978,9.771099,9.495697,8.850578,8.937348,9.103344,9.26934,9.922004,9.250477,9.265567,9.737145,10.386037,10.876478,10.469034,9.695646,8.846806,8.099826,7.5112963,7.213259,7.3679366,7.635793,7.6810646,7.17176,6.7379084,6.673774,6.858632,7.175533,7.4811153,8.578949,9.231613,9.333474,9.125979,9.190115,10.253995,11.400873,12.012038,12.219532,12.894833,13.20796,13.0646,12.381755,11.216014,9.74469,9.616421,8.329956,7.3188925,7.3151197,8.360137,8.722309,9.699419,10.665211,11.042474,10.303039,9.805053,9.405154,9.084481,8.529905,7.1076255,7.254758,8.001738,9.129752,10.355856,11.321648,11.506506,11.374464,11.291467,11.1782875,10.510533,10.763299,12.136535,13.072145,13.234368,13.505998,13.958713,14.498198,14.64533,14.11339,12.796744,13.174006,13.038192,12.974057,12.909923,12.1101265,10.978339,9.997457,8.98262,7.865923,6.6813188,6.688864,7.0510364,7.605612,8.126234,8.329956,8.371455,8.314865,8.118689,7.665974,6.779407,6.6247296,6.587003,6.5341864,6.8058157,8.20546,9.5032425,10.26154,10.223814,9.839006,10.235131,11.287694,12.223305,13.004238,13.528633,13.645585,13.996439,13.65313,12.951422,12.423254,12.792972,13.460726,13.758763,13.70972,13.747445,14.70192,13.558814,12.626976,12.574159,12.981603,12.344029,12.611885,13.52486,14.18507,14.037937,12.883514,14.901869,14.332202,14.807553,15.282904,15.430037,15.629986,16.569368,16.520325,15.988385,15.331948,14.762281,14.6151495,14.215251,13.687083,13.385274,13.917213,15.939341,16.592005,15.792209,14.396337,14.2077055,14.086982,13.600313,13.487134,13.822898,14.011529,13.124963,13.008011,13.52486,14.490653,15.675257,16.007248,15.826162,15.509261,15.501716,16.305285,17.056038,17.56157,17.610613,17.237123,16.735365,15.829934,15.369675,15.131999,15.060319,15.290449,16.486372,16.991903,16.897587,16.135517,14.483108,13.174006,12.736382,12.366665,11.781908,11.242422,10.472807,10.559577,10.661438,10.593531,10.834979,11.268831,11.121698,10.748209,10.374719,10.099318,10.419991,10.336992,10.212496,10.03141,9.371201,8.873214,8.3525915,7.8621507,7.3377557,6.620957,6.017337,5.27413,4.3083377,3.2331395,2.3654358,1.6260014,1.1695137,0.97333723,0.94692886,0.935611,1.0072908,1.0072908,0.9997456,0.97710985,0.8903395,0.97333723,0.9205205,0.935611,1.1091517,1.4260522,2.71629,6.1078796,8.265821,8.756263,10.054046,9.774872,9.5032425,10.487898,11.887542,10.785934,13.015556,11.472552,6.7680893,1.4826416,0.16976812,0.0754525,0.056589376,0.060362,0.05281675,0.02263575,0.05281675,0.071679875,0.10186087,0.18485862,0.36594462,0.8903395,0.91674787,0.995973,1.1808317,1.0450171,1.1355602,1.750498,1.9730829,1.7467253,1.8636768,1.3770081,2.082489,2.927557,3.1916409,2.4672968,2.7841973,2.655928,2.757789,2.8596497,1.8297231,2.4220252,2.5012503,2.6446102,2.9803739,3.187868,2.6031113,2.7087448,2.7502437,2.655928,3.0218725,3.0746894,2.9313297,3.0558262,3.2255943,2.5540671,3.1954134,2.9916916,3.350091,4.2894745,4.425289,3.6934,3.0558262,3.0030096,3.4179983,3.5839937,3.5123138,3.5424948,3.5085413,3.7763977,5.251494,5.983383,6.832224,7.8810134,9.125979,10.484125,10.386037,9.903141,9.676784,9.839006,10.042727,9.918231,9.797507,9.914458,10.035183,9.454198,9.201432,9.1825695,8.922258,8.386545,7.9791017,8.511042,8.933576,9.4127,9.710737,9.1976595,8.684583,8.763808,8.66572,8.311093,8.269594,8.548768,8.8769865,8.944894,8.82417,8.944894,9.891823,10.79348,11.563096,11.910177,11.363147,10.767072,10.186088,9.857869,9.7069645,9.363655,9.393836,9.831461,10.20495,10.314357,10.231359,10.552032,10.450171,10.386037,10.487898,10.533169,11.016065,12.012038,14.102073,16.893814,19.029121,19.94964,19.655376,17.96524,15.924251,15.811071,16.478827,17.105082,15.739391,13.060828,12.404391,12.804289,12.928786,12.894833,12.97783,13.588995,14.177525,14.362384,13.977575,12.777881,10.469034,10.076681,10.797253,11.744182,12.306303,12.151625,12.940104,13.019329,13.287186,14.019074,14.864142,13.875714,13.6682205,13.449409,12.785426,11.619685,9.699419,8.186596,7.6018395,7.8131065,8.0206,8.873214,10.412445,11.34051,11.385782,11.329193,12.54775,13.038192,12.351574,10.804798,9.484379,8.831716,8.013056,7.2283497,6.85486,7.413208,8.182823,8.360137,8.846806,9.680555,10.0465,10.382264,9.1976595,9.035437,9.967276,9.608876,12.257258,8.990166,6.043745,4.715781,1.3656902,4.67051,5.772116,6.5341864,6.832224,4.5724216,3.127506,2.5276587,3.0331905,4.2894745,5.300538,5.462761,5.715527,6.1342883,6.934085,8.443134,8.443134,9.280658,10.374719,10.872705,9.669238,8.062099,7.3490734,7.394345,8.0206,9.027891,8.578949,7.1378064,6.270103,6.270103,6.145606,5.7570257,6.0626082,6.730363,7.232122,6.8435416,6.066381,6.096562,6.628502,6.9189944,5.7872066,5.247721,5.881522,6.4511886,6.587003,6.7944975,6.9189944,6.519096,6.0362,5.8890676,6.477597,6.3945994,6.537959,7.1264887,7.726336,7.254758,6.349328,5.353355,4.8968673,5.070408,5.406172,5.9984736,6.7567716,7.537705,8.182823,8.537451,8.273367,7.805561,7.7150183,8.141325,8.778898,9.152389,9.439108,9.710737,9.831461,9.495697,9.148616,9.193887,9.416472,9.752235,10.287949,11.208468,11.249968,11.872451,13.196642,14.02662,15.577168,14.634012,13.430545,12.913695,12.743927,12.996693,13.860624,14.898096,15.829934,16.509007,13.50977,12.46098,12.709973,13.5663595,14.302021,13.532406,12.3289385,11.317875,10.740664,10.453944,10.065364,10.785934,11.672502,12.487389,13.72481,13.332457,13.015556,12.67602,12.208215,11.472552,10.842525,10.518079,10.208723,9.774872,9.216523,8.616675,8.89585,9.593785,10.412445,11.223559,11.227332,11.631002,11.415963,10.789707,11.197151,12.204442,11.140562,10.227587,10.170997,10.148361,10.604849,11.408418,12.385528,13.27964,13.781399,12.283667,10.1294985,8.733627,8.631766,9.457971,8.914713,8.29223,8.243186,8.635539,8.578949,8.956212,9.476834,9.986138,10.167224,9.544742,8.582722,7.213259,6.937857,7.6131573,7.466025,7.907422,9.382519,10.140816,10.208723,11.393328,10.948157,10.552032,10.917976,11.947904,12.751472,11.92904,11.962994,11.219787,9.457971,7.8319697,7.009537,5.7004366,5.2665844,6.0550632,7.4207535,7.8017883,8.167733,8.499724,8.793989,9.050528,9.288202,9.26934,8.631766,7.6810646,7.3981175,7.4735703,7.960239,8.141325,8.073418,8.578949,8.586494,8.469543,8.560086,8.967529,9.58624,8.99771,8.314865,7.798016,7.364164,6.579458,6.168242,5.674028,5.3609,5.1873593,4.8100967,4.9421387,4.8365054,4.908185,5.3986263,6.3719635,4.7912335,5.3269467,4.881777,5.27413,13.245687,17.244669,14.403882,9.7296,6.9265394,8.412953,7.586749,7.9526935,8.394091,8.386545,8.00551,8.458225,8.922258,9.156161,9.337247,10.080454,9.393836,9.590013,10.069136,10.114408,8.899622,8.963757,8.382772,8.367682,8.228095,5.3986263,4.429062,5.4250345,6.72659,8.14887,11.000975,10.884023,14.094527,12.830698,6.5832305,2.1315331,4.817642,4.938366,4.315883,6.8850408,18.678267,25.759483,20.534397,13.630494,9.665465,7.2585306,5.674028,7.364164,9.208978,9.797507,9.424017,9.076936,8.843033,8.76758,8.929804,9.461743,8.590267,8.963757,9.295748,9.378746,10.069136,9.906913,8.892077,8.050782,7.798016,7.914967,7.9489207,8.07719,8.069645,7.7829256,7.145352,6.8397694,6.5530496,6.587003,7.118943,8.171506,9.099571,9.378746,9.26934,9.163706,9.6201935,10.438853,11.796998,12.581704,12.687338,13.038192,12.73261,11.785681,11.031156,10.484125,9.344792,9.544742,8.714764,7.9451485,7.828197,8.431817,8.854351,9.948412,11.053791,11.3669195,9.955957,8.967529,8.669493,8.360137,7.5263867,5.824933,6.670001,7.805561,9.193887,10.499215,11.057564,10.967021,10.853842,11.042474,11.393328,11.2801485,11.785681,13.445636,14.524607,14.505743,14.109617,14.988639,15.535669,15.671484,14.883006,12.242168,11.879996,11.23865,11.634775,12.789199,12.838243,11.216014,9.884277,8.726082,7.677292,6.719045,6.4926877,7.194396,7.997965,8.439363,8.424272,8.627994,8.461998,7.964011,7.3377557,6.9793563,7.496206,7.3717093,7.009537,7.020855,8.201687,9.42779,10.559577,10.521852,9.759781,10.253995,11.785681,12.449662,12.7477,13.026875,13.490907,14.551015,14.219024,12.974057,11.77059,12.0233555,13.456953,14.7170105,14.962231,14.569878,15.116908,14.728328,13.27964,12.453435,12.332711,11.3669195,11.427281,12.615658,13.800262,14.169979,13.234368,14.815099,14.4152,15.712983,16.38451,15.739391,14.724555,14.894323,14.607604,14.5283785,14.68683,14.479335,14.139798,13.8870325,13.679539,13.562587,13.671993,15.965749,17.21826,16.882498,15.46399,14.509516,13.192869,12.076173,12.264804,13.585222,14.57365,14.437836,14.7170105,15.154634,15.611122,16.052519,16.199652,15.467763,15.064092,15.46399,16.403374,18.500954,18.99894,18.45568,17.271078,15.686575,15.260268,15.23386,15.569623,15.897841,15.531898,15.863888,15.98084,15.920478,15.252723,13.091009,12.506252,12.396846,12.147853,11.521597,10.680302,10.291721,10.34831,10.416218,10.370946,10.4049,10.578441,10.325675,10.0465,9.989911,10.269085,10.416218,10.212496,9.993684,9.688101,8.835487,7.466025,6.6850915,6.126743,5.666483,5.4476705,5.032682,4.1612053,3.059599,1.9504471,1.0223814,0.694163,0.5017591,0.42630664,0.422534,0.3961256,0.27540162,0.271629,0.31312788,0.34330887,0.3055826,0.36594462,0.42630664,0.482896,0.58475685,0.83752275,1.780679,4.9421387,7.3792543,8.186596,8.514814,9.224068,8.729855,8.518587,8.903395,9.065618,10.699164,7.043491,2.8822856,0.573439,0.060362,0.071679875,0.056589376,0.0754525,0.10940613,0.060362,0.10940613,0.1659955,0.124496624,0.08677038,0.36594462,1.5241405,1.3656902,1.2638294,1.4939595,1.2525115,1.0676528,1.8297231,2.1466236,2.0598533,3.0369632,3.097325,3.7537618,3.2972744,1.9881734,2.0749438,2.4408884,2.2409391,2.2598023,2.4031622,1.6939086,2.5616124,2.4672968,2.4786146,2.806833,2.806833,2.686109,2.837014,2.8747404,2.8143783,3.0822346,3.399135,3.6896272,4.055572,4.1762958,3.3123648,3.4330888,3.078462,3.3425457,4.1197066,4.1197066,4.0216184,3.6330378,3.5085413,3.682082,3.6481283,3.3312278,3.0218725,3.0407357,3.6179473,4.8968673,6.4134626,6.85486,7.4282985,8.52236,9.703192,9.88805,9.669238,9.812597,10.005001,8.835487,9.14107,9.639057,10.393582,10.978339,10.469034,9.442881,9.295748,9.148616,8.699674,8.224322,8.786444,9.163706,9.963503,10.589758,9.246704,8.782671,9.178797,9.314611,9.137298,9.673011,10.235131,10.054046,9.450426,9.0807085,9.933322,11.106608,12.494934,13.162688,12.770335,11.59705,10.899114,10.627484,10.442626,10.167224,9.767326,10.167224,10.808571,10.993429,10.597303,10.069136,9.97482,10.352083,10.944386,11.423509,11.3971,11.521597,11.796998,12.498707,13.856852,16.052519,17.41821,17.338985,16.26756,14.969776,14.543469,15.1395445,16.022339,15.826162,14.539697,13.502225,12.381755,11.476325,11.532914,12.321393,12.649611,12.857106,13.249459,12.849561,11.589504,10.284176,10.578441,11.227332,11.830952,12.151625,12.113899,12.298758,12.774108,13.404137,13.924759,13.962485,13.50977,13.12119,13.215506,13.45318,12.755245,10.570895,8.296002,7.2094865,7.726336,9.397609,8.7751255,9.839006,11.272603,12.049765,11.41219,12.427027,13.038192,12.830698,12.121444,11.962994,10.461489,8.446907,7.220804,7.118943,7.5226145,7.6093845,7.4811153,7.7640624,8.130007,7.322665,7.6923823,8.2507305,8.646856,8.314865,6.470052,8.729855,5.247721,2.384299,2.161714,2.2598023,1.7354075,1.4109617,1.7957695,2.5201135,2.3503454,3.1425967,3.0860074,3.4934506,4.557331,5.3269467,5.802297,6.2323766,6.3832817,6.6134114,7.858378,7.6508837,8.137552,8.695901,9.046755,9.276885,8.66572,7.84706,7.5527954,8.111144,9.431562,8.307321,7.677292,6.9869013,6.3153744,6.379509,6.5228686,6.598321,6.937857,7.356619,7.1264887,6.4549613,6.349328,5.983383,5.2364035,4.7006907,5.2854476,5.9003854,6.375736,6.6134114,6.5756855,6.6020937,6.1418333,5.8702044,6.0512905,6.515323,6.089017,6.2927384,6.79827,7.2170315,7.0963078,7.2660756,6.5228686,5.9305663,5.9305663,6.330465,6.466279,7.2887115,8.186596,8.816625,9.110889,9.903141,9.442881,8.643084,8.107371,8.13378,8.424272,8.710991,9.495697,10.642575,11.336739,10.970794,10.733118,9.963503,9.190115,10.11818,11.204697,10.861387,10.842525,11.570641,12.147853,13.45318,14.4114275,14.622695,14.109617,13.306048,13.551269,14.305794,14.894323,14.973549,14.558559,12.298758,12.321393,13.321139,14.071891,13.411682,12.336484,12.215759,12.095036,11.623458,11.0613365,10.050273,9.933322,10.306811,11.099063,12.58925,12.294985,12.030901,11.883769,11.631002,10.725573,9.737145,8.394091,7.8244243,8.239413,8.91094,8.643084,8.89585,9.752235,10.612394,10.223814,9.650374,9.688101,9.903141,10.231359,11.000975,11.551778,10.4049,9.454198,9.367428,9.612649,10.272858,10.638803,10.601076,10.423763,10.740664,11.302785,11.955449,10.608622,8.360137,9.507015,9.480607,8.98262,8.918486,9.382519,9.627739,9.6051035,10.054046,10.54826,10.657665,9.948412,8.692128,6.7379084,5.915476,6.3455553,6.4549613,8.311093,11.272603,12.743927,11.808316,9.231613,9.4013815,9.710737,9.778644,10.137043,12.238396,13.264549,11.019837,8.83926,7.7338815,6.379509,5.485397,4.478106,3.9159849,4.304565,6.089017,7.515069,8.265821,8.68081,8.918486,8.941121,9.099571,9.186342,8.948667,8.348819,7.567886,7.605612,8.228095,8.646856,8.7600355,9.14107,9.0807085,8.771353,8.439363,8.412953,9.110889,9.159933,8.869441,8.405409,7.8621507,7.2623034,6.7152724,6.126743,5.7570257,5.6400743,5.613666,5.6400743,5.6815734,5.945657,6.360646,6.590776,4.063117,4.606375,5.5457587,5.7494807,5.617439,15.271586,16.969267,12.193124,6.1078796,7.5829763,8.537451,9.175024,9.012801,8.590267,9.507015,9.322156,9.578695,8.620448,7.541477,10.178542,10.408672,9.669238,8.571404,7.069899,4.45547,7.9489207,6.0626082,3.1237335,1.6637276,2.4559789,2.7879698,5.2137675,8.073418,9.439108,7.0963078,7.9262853,17.599297,21.292696,15.241405,6.7454534,5.0477724,4.3196554,3.92353,7.0849895,20.889025,41.98177,33.81781,18.184053,7.7225633,5.904158,4.2328854,5.1232247,6.971811,8.375228,8.118689,8.484633,8.280911,8.141325,8.265821,8.439363,8.412953,8.83926,8.729855,8.333729,9.14107,9.261794,8.22055,7.7376537,8.099826,8.14887,8.416726,8.228095,7.726336,7.2283497,7.2170315,7.3151197,7.111398,7.141579,7.624475,8.4544525,9.416472,9.989911,10.238904,10.291721,10.314357,10.352083,11.714001,12.698656,12.623203,11.84227,11.5857315,10.386037,9.397609,8.9788475,8.695901,9.5032425,9.767326,9.322156,8.394091,7.6131573,8.114917,9.303293,10.646348,11.299012,10.103089,8.684583,7.809334,7.3151197,6.900131,6.119198,6.730363,7.9451485,9.42779,10.653893,10.910432,11.838497,12.151625,12.0233555,11.891314,12.449662,13.317367,14.66042,15.852571,16.418465,16.052519,17.320122,17.803017,17.327667,15.901614,13.717264,13.472044,11.068882,10.823661,12.958967,13.59654,12.166716,10.914205,9.374973,7.914967,7.7225633,7.17176,7.492433,8.016829,8.424272,8.744945,8.669493,8.137552,7.273621,6.515323,6.6360474,7.858378,8.677037,8.60913,8.058327,8.299775,9.484379,10.880251,10.853842,9.718282,9.703192,11.744182,12.864652,13.151371,12.943876,12.83447,13.539951,13.95494,13.645585,12.830698,12.3893,14.479335,16.720274,16.758,14.909414,14.1926155,15.7657995,15.169725,13.88326,12.464753,10.574668,10.525623,10.970794,11.989402,12.966512,12.58925,13.170234,14.102073,14.520834,14.286931,13.645585,13.249459,12.928786,12.638294,12.894833,13.588995,13.966258,14.1058445,14.143571,13.905896,13.551269,13.573905,15.147089,16.70141,16.678776,15.0905,13.536179,13.106099,13.264549,13.483362,13.615403,13.902123,14.547242,14.626467,14.879233,15.535669,16.29774,15.592259,15.365902,15.516807,15.943113,16.550507,17.067356,16.950403,16.463736,15.754482,14.830189,15.516807,15.705438,15.973294,16.248695,15.814844,14.826416,14.298248,13.622949,12.73261,12.102581,12.132762,11.940358,11.589504,11.019837,10.069136,9.2995205,9.431562,9.507015,9.322156,9.416472,9.639057,9.808825,10.125726,10.457717,10.367173,10.182315,10.072908,9.805053,9.114662,7.7225633,6.8246784,6.5266414,6.307829,5.885295,5.2288585,4.459243,3.229367,2.0145817,1.0827434,0.4979865,0.31312788,0.20372175,0.14713238,0.13958712,0.150905,0.116951376,0.1659955,0.21881226,0.24899325,0.27917424,0.29426476,0.32067314,0.29803738,0.28294688,0.46026024,1.177059,3.187868,4.825187,5.7079816,6.719045,7.4094353,6.6322746,6.1908774,6.628502,7.2585306,5.564622,3.059599,1.116697,0.25276586,0.120724,0.0754525,0.05281675,0.0452715,0.041498873,0.011317875,0.060362,0.19240387,0.16976812,0.094315626,0.40367088,1.1053791,0.8526133,1.177059,2.0372176,1.81086,2.0183544,2.3428001,2.4031622,2.3767538,3.0105548,1.6675003,1.6335466,1.9278114,2.142851,2.4408884,2.4069347,2.493705,2.7087448,2.8709676,2.6219745,2.776652,2.2899833,1.9504471,1.8938577,1.6109109,1.8297231,2.463524,2.7615614,2.746471,3.240685,3.2444575,3.6254926,3.983892,4.187614,4.38379,3.470815,3.3274553,3.92353,4.666737,4.4139714,4.7836885,4.0706625,3.651901,3.8707132,4.036709,3.5236318,3.2859564,3.4783602,4.032936,4.6290107,5.7909794,6.205968,7.3000293,8.956212,9.495697,8.216777,8.084735,8.420499,8.601585,8.054554,8.367682,9.322156,10.280403,10.680302,10.038955,9.639057,9.020347,8.7600355,8.918486,9.031664,9.084481,8.918486,9.367428,10.170997,9.978593,9.623966,10.295494,10.521852,10.435081,11.763044,12.449662,11.883769,11.480098,11.59705,11.544232,11.672502,12.170488,12.630749,12.713746,12.15917,11.834724,11.898859,11.936585,11.778135,11.521597,11.065109,10.974566,10.729345,10.257768,9.88805,9.563604,9.9257765,10.7557535,11.649866,11.996947,12.498707,13.158916,13.845533,14.720782,16.222288,18.274595,17.882242,16.923996,16.248695,15.675257,15.716756,16.188334,16.063837,15.358356,15.150862,14.086982,13.343775,13.985121,15.169725,14.151116,13.185325,13.249459,13.000465,12.053536,10.944386,11.012292,10.733118,10.506761,10.344538,9.857869,10.653893,10.940613,11.295239,11.793225,11.98563,12.54775,12.487389,12.004493,11.185833,10.008774,8.382772,7.854605,8.288457,9.295748,10.253995,9.016574,9.835234,11.54046,12.668475,11.487643,12.638294,13.377728,12.67602,11.18206,11.219787,9.952185,9.012801,8.13378,7.4094353,7.3151197,8.043237,7.5301595,7.5037513,8.028146,7.496206,5.7607985,8.469543,8.52236,5.2062225,4.1762958,3.0445085,1.9542197,1.2562841,1.1091517,1.4524606,0.8903395,2.4522061,3.4142256,3.3840446,4.315883,4.8930945,4.5988297,4.7648253,5.6513925,6.458734,7.2396674,7.4169807,6.7567716,6.013564,6.9189944,7.7376537,8.333729,8.571404,8.529905,8.507269,7.858378,7.2623034,7.2170315,7.8621507,8.967529,7.364164,6.930312,6.72659,6.3531003,5.975838,6.7454534,7.194396,7.6584287,7.877241,6.990674,6.1644692,6.5341864,6.4474163,5.7004366,5.553304,6.3153744,6.8774953,7.0963078,6.9680386,6.6360474,6.934085,6.771862,6.990674,7.635793,7.9451485,7.1340337,7.17176,7.492433,7.7414265,7.752744,7.33021,6.63982,6.224831,6.3945994,7.2472124,7.4697976,8.107371,8.922258,9.359882,8.560086,8.601585,8.620448,8.27714,7.8810134,8.36391,9.261794,10.065364,10.79348,11.446144,11.98563,11.295239,10.544487,10.174769,10.140816,9.895596,10.552032,10.691619,10.514306,10.480352,11.2801485,12.223305,12.966512,14.007756,14.856597,14.049255,13.619176,13.981348,14.064346,13.588995,13.057055,12.427027,12.117672,11.838497,11.476325,11.080199,10.269085,10.842525,11.234878,10.876478,10.208723,10.287949,10.050273,9.963503,10.401127,11.634775,11.966766,11.653639,11.057564,10.216269,8.835487,7.9338303,6.8661776,6.2889657,6.4926877,7.3981175,8.13378,8.405409,8.511042,8.631766,8.809079,9.688101,9.771099,9.616421,9.627739,10.038955,11.2801485,10.974566,10.646348,10.49167,9.367428,8.2507305,9.088254,9.748463,9.982366,11.41219,11.653639,12.966512,12.664702,10.533169,8.809079,8.873214,8.60913,8.616675,9.122208,9.971047,9.680555,10.31813,10.567122,9.869187,8.409182,6.858632,6.4021444,6.651138,7.115171,7.1868505,7.696155,8.718536,10.18986,11.672502,12.366665,10.038955,10.910432,11.329193,10.861387,12.287439,12.559069,10.970794,8.865668,6.9454026,5.2665844,4.191386,4.014073,4.1612053,4.5761943,5.723072,6.8850408,7.360391,7.816879,8.382772,8.612903,9.307066,9.639057,9.314611,8.605357,8.299775,7.9941926,8.224322,8.311093,8.182823,8.394091,8.627994,8.503497,8.299775,8.262049,8.597813,8.869441,8.835487,8.420499,7.7037,6.9227667,6.549277,6.387054,6.089017,5.794752,6.1531515,5.8136153,5.723072,5.9682927,6.515323,7.2283497,5.5306683,4.447925,4.821415,6.017337,5.934339,13.04951,15.667711,13.083464,8.156415,7.277394,8.473316,8.7751255,9.7069645,11.310329,12.117672,8.827943,8.59404,8.160188,7.462252,9.639057,11.465008,9.695646,9.495697,9.850324,3.5764484,5.485397,6.760544,7.020855,6.722818,7.145352,3.6141748,3.6141748,5.8702044,8.107371,7.020855,5.168496,10.77839,16.03743,16.818363,12.67602,8.050782,5.353355,3.942393,4.349837,8.29223,14.154889,14.6302395,13.12119,10.650121,5.8437963,6.066381,5.1534057,5.621211,7.3490734,7.5792036,8.122461,7.8998766,7.7640624,7.9715567,8.182823,7.9413757,8.431817,8.6581745,8.560086,9.005256,8.590267,8.039464,8.103599,8.76758,9.235386,8.544995,7.816879,7.3151197,7.118943,7.1076255,7.1566696,7.224577,7.462252,7.7112455,7.5263867,8.031919,9.22784,10.103089,10.408672,10.657665,10.63503,11.272603,12.064855,12.272349,10.914205,11.329193,10.850069,10.442626,10.284176,9.759781,10.253995,10.54826,9.850324,8.52236,8.103599,8.552541,9.246704,10.001229,10.31813,9.344792,8.337502,7.858378,7.5490227,7.2698483,7.0812173,7.360391,8.001738,8.786444,9.484379,9.846551,11.321648,12.015811,12.253486,12.543978,13.573905,14.373701,14.841507,15.060319,14.93205,14.18507,15.784663,17.961468,18.693357,17.421982,15.071637,11.578186,10.710483,11.389555,12.672247,13.766309,13.04951,11.917723,10.163452,8.29223,7.4999785,7.4584794,7.937603,8.465771,8.778898,8.793989,8.552541,7.5037513,6.3455553,5.715527,6.198423,7.8395147,8.858124,9.129752,8.756263,8.043237,8.699674,9.854096,10.31813,10.310584,11.461235,12.113899,12.208215,12.245941,12.479843,12.917468,13.13628,13.43809,14.04171,14.6151495,14.283158,14.962231,16.290195,16.086473,14.48688,13.920986,13.555041,13.306048,13.264549,12.951422,11.344283,11.510279,12.038446,12.608112,12.96274,12.917468,11.649866,12.611885,13.3626375,13.057055,11.974312,11.532914,11.604594,12.0082655,12.427027,12.789199,13.253232,13.370183,13.472044,13.551269,13.649357,13.860624,14.219024,14.807553,14.713238,13.773854,12.54775,12.58925,13.011784,13.521088,13.721037,13.083464,13.879487,14.18507,14.584969,15.211224,15.724301,15.705438,15.62244,15.331948,14.988639,15.067864,15.724301,16.044973,15.920478,15.486626,15.1395445,15.049001,14.652876,14.64533,14.988639,14.943368,14.603831,13.736128,12.808062,12.136535,11.846043,11.672502,11.393328,10.955703,10.325675,9.488152,9.156161,9.344792,9.529651,9.58624,9.793735,9.548513,9.846551,10.34831,10.710483,10.56335,10.144588,9.9257765,9.265567,8.122461,7.0812173,6.3417826,5.8513412,5.3382645,4.7006907,4.0291634,3.0860074,2.04099,1.1695137,0.5998474,0.28294688,0.1659955,0.094315626,0.056589376,0.041498873,0.0452715,0.041498873,0.071679875,0.094315626,0.10186087,0.12826926,0.1659955,0.1659955,0.15845025,0.17354076,0.23767537,0.8601585,2.516341,3.8707132,4.4630156,4.7346444,5.292993,5.3609,5.0854983,4.851596,5.2967653,3.229367,1.5354583,0.55457586,0.22258487,0.08299775,0.041498873,0.041498873,0.041498873,0.033953626,0.018863125,0.060362,0.150905,0.150905,0.18485862,0.6488915,1.0072908,1.0110635,1.478869,2.173032,1.8070874,1.6561824,1.7089992,1.629774,1.478869,1.7052265,1.0714256,1.3392819,1.5769572,1.5543215,1.7542707,2.1994405,2.4484336,2.7540162,2.9841464,2.6144292,2.7653341,2.282438,2.0636258,2.2786655,2.354118,2.4710693,2.8181508,2.848332,2.7125173,3.2972744,3.180323,3.7877154,4.13857,4.146115,4.606375,3.8480775,3.682082,4.221567,5.119452,5.594803,5.13077,4.285702,3.9801195,4.2404304,4.191386,4.2894745,4.093298,3.9914372,4.2102494,4.82896,5.4778514,6.058836,7.17176,8.586494,9.235386,8.575176,8.646856,8.948667,9.046755,8.582722,8.963757,9.303293,9.578695,9.65792,9.291975,9.107117,8.884532,8.82417,9.035437,9.525878,9.699419,9.74469,10.193633,10.895341,11.012292,11.174516,11.408418,11.766817,12.3893,13.483362,13.483362,12.90615,12.664702,12.838243,12.687338,11.925267,11.834724,12.181807,12.664702,12.913695,12.826925,12.940104,13.004238,12.879742,12.513797,11.555551,10.695392,10.080454,9.831461,10.042727,9.789962,9.752235,10.152134,11.02361,12.200669,13.3626375,13.8719425,14.562332,15.7657995,17.335213,18.980076,19.289433,19.191343,18.742401,17.112627,15.901614,15.894069,15.845025,15.414946,15.181043,14.750964,14.920732,15.728074,16.376965,15.211224,13.4644985,12.898605,12.800517,12.604341,11.895086,11.54046,10.989656,10.457717,9.944639,9.239159,9.5032425,9.81637,10.005001,10.137043,10.502988,11.559323,11.2650585,10.280403,9.276885,8.918486,7.7376537,7.4471617,8.322411,9.903141,11.00852,10.487898,10.152134,10.744436,11.793225,11.623458,11.400873,12.3289385,12.513797,11.672502,11.114153,9.955957,9.344792,8.793989,8.096053,7.326438,8.122461,7.515069,7.1793056,8.043237,10.310584,8.412953,7.707473,5.9796104,3.399135,2.5389767,1.8561316,1.5015048,1.086516,0.70170826,0.875249,1.0487897,3.3312278,4.5196047,4.478106,6.1342883,6.4247804,6.5455046,7.001992,7.665974,7.752744,8.394091,8.443134,7.726336,6.8473144,7.1679873,8.103599,8.254503,8.375228,8.537451,8.152642,7.7187905,7.4018903,7.3188925,7.6282477,8.492179,6.851087,6.1418333,6.1833324,6.488915,6.2399216,6.9567204,7.488661,7.7942433,7.7150183,7.001992,6.7756343,6.9869013,6.858632,6.3531003,6.1720147,6.7114997,7.2623034,7.492433,7.284939,6.7341356,6.9567204,7.0849895,7.326438,7.7414265,8.246958,7.884786,7.707473,7.6207023,7.4697976,7.01331,6.8699503,6.375736,5.8664317,5.704209,6.2851934,7.0963078,7.937603,8.907167,9.484379,8.552541,8.2507305,7.8734684,7.488661,7.5075235,8.661947,9.507015,10.408672,11.087745,11.434827,11.487643,11.200924,10.650121,10.401127,10.484125,10.408672,10.672756,10.435081,10.057818,9.940866,10.521852,11.559323,12.049765,12.887287,13.917213,13.917213,13.860624,13.928532,13.837989,13.290957,11.974312,11.778135,11.751727,11.25374,10.367173,9.922004,9.835234,10.997202,11.691365,11.2801485,10.20495,10.280403,10.065364,9.861642,10.016319,10.902886,11.099063,10.759526,10.31813,9.57115,7.665974,6.9265394,6.379509,6.058836,6.1041074,6.790725,7.484888,7.8017883,7.6207023,7.5075235,8.718536,10.38981,10.925522,10.668983,10.023865,9.484379,10.7557535,11.476325,11.646093,11.019837,9.0807085,7.273621,8.937348,10.121953,10.065364,11.197151,11.355601,11.751727,11.668729,10.812344,9.295748,8.684583,8.122461,8.069645,8.6732645,9.763554,9.144843,9.337247,9.95973,10.453944,10.095545,8.45068,6.677546,6.1041074,6.828451,7.7187905,8.394091,8.084735,8.284684,9.465516,11.076427,10.582213,11.087745,11.129244,10.49167,10.201178,9.74469,8.914713,7.9791017,7.001992,5.8702044,4.7610526,4.1498876,4.06689,4.496969,5.383536,6.175787,6.6360474,7.2924843,8.130007,8.601585,9.405154,9.793735,9.393836,8.514814,8.126234,7.488661,7.7150183,7.9941926,8.054554,8.182823,8.495952,8.2507305,8.0206,8.084735,8.469543,8.75249,8.631766,8.288457,7.786698,7.073672,6.7077274,6.677546,6.587003,6.511551,7.001992,5.8702044,5.8928404,6.1795597,6.375736,6.670001,6.515323,4.9157305,4.979865,6.598321,6.4134626,8.386545,11.223559,12.215759,10.31813,6.149379,7.4282985,7.9262853,10.423763,14.234114,15.207452,8.409182,7.726336,8.3525915,8.639311,10.110635,11.827179,9.669238,8.190369,7.8696957,5.0968165,4.727099,4.7950063,9.231613,18.078419,27.476028,18.757492,9.601331,6.771862,10.072908,12.321393,6.1908774,9.590013,13.034419,12.615658,10.005001,9.971047,5.8588867,3.1727777,3.482133,4.436607,9.265567,10.733118,10.231359,8.495952,5.6098933,6.039973,5.1534057,5.1835866,6.485142,7.5565677,8.918486,8.76758,8.103599,7.7602897,8.409182,8.269594,9.005256,9.537196,9.616421,9.831461,9.129752,8.714764,8.695901,9.065618,9.699419,8.880759,7.7414265,7.043491,6.9265394,6.907676,6.9793563,7.175533,7.533932,7.8244243,7.5226145,7.7225633,8.6581745,9.623966,10.272858,10.623712,10.672756,11.000975,11.747954,12.31762,11.348056,11.438599,11.506506,11.589504,11.498961,10.804798,10.616167,10.718028,9.967276,8.499724,7.7301087,7.7678347,8.239413,9.224068,10.159679,9.850324,8.99771,8.6732645,8.477088,8.273367,8.186596,8.262049,8.68081,8.929804,9.073163,9.767326,11.355601,12.0724,12.596795,13.200415,13.728582,14.611377,14.43029,13.996439,13.758763,13.807808,14.2944765,15.939341,16.893814,16.044973,13.023102,11.151879,10.895341,11.344283,12.030901,12.940104,13.245687,12.694883,11.261286,9.337247,7.7678347,7.4697976,7.9526935,8.922258,9.763554,9.525878,9.076936,7.5490227,6.175787,5.6853456,6.326692,8.099826,8.903395,8.865668,8.371455,8.035691,8.443134,9.337247,10.170997,10.834979,11.646093,11.868678,11.781908,11.800771,12.128989,12.7477,12.58925,12.596795,13.140053,13.943622,14.124708,14.928277,16.373192,16.546734,15.497944,15.226315,14.34352,13.864397,13.875714,13.875714,12.751472,12.336484,12.30253,12.400619,12.453435,12.351574,11.00852,11.710228,12.664702,12.664702,11.672502,10.804798,11.385782,12.019584,12.491161,12.740154,12.875969,12.468526,12.279895,12.551523,13.098554,13.313594,13.128735,13.106099,12.996693,12.672247,12.132762,12.166716,12.543978,13.166461,13.483362,12.510024,13.302276,13.555041,13.902123,14.535924,15.211224,16.01102,15.928022,15.16218,14.298248,14.302021,14.981093,15.603577,15.75071,15.414946,15.01882,14.286931,13.758763,13.747445,14.079436,14.068119,14.053028,13.147598,12.298758,11.84227,11.498961,11.185833,10.970794,10.540714,9.944639,9.556059,9.590013,9.58624,9.627739,9.733373,9.842778,9.533423,9.937095,10.47658,10.850069,11.012292,10.208723,9.563604,8.469543,7.069899,6.2361493,5.3684454,4.7120085,4.0782075,3.4217708,2.8521044,1.9730829,1.2298758,0.70170826,0.38858038,0.21503963,0.12826926,0.071679875,0.049044125,0.0452715,0.0150905,0.011317875,0.026408374,0.033953626,0.026408374,0.018863125,0.060362,0.05281675,0.06790725,0.1056335,0.10940613,0.6413463,1.9429018,2.9803739,3.3048196,3.059599,3.4557245,4.074435,4.134797,3.6292653,3.3048196,1.9466745,0.98465514,0.44139713,0.22258487,0.08677038,0.060362,0.041498873,0.056589376,0.08677038,0.056589376,0.056589376,0.116951376,0.13204187,0.19994913,0.6375736,0.8224323,1.0827434,1.4109617,1.6071383,1.2751472,1.2110126,1.1921495,1.0714256,0.87902164,0.8639311,0.8941121,1.3392819,1.3732355,1.1129243,1.6146835,1.8749946,2.0108092,2.233394,2.4823873,2.4182527,2.8709676,2.8407867,2.795515,2.9049213,3.059599,2.8407867,3.029418,3.108643,3.0633714,3.3651814,3.2482302,3.7235808,4.134797,4.2404304,4.2102494,4.074435,4.2630663,4.768598,5.4665337,6.138061,5.3759904,4.610148,4.353609,4.4931965,4.274384,4.82896,4.5988297,4.3083377,4.429062,5.1873593,5.783434,6.6624556,7.515069,8.213005,8.809079,8.89585,9.201432,9.710737,10.148361,9.97482,9.922004,9.465516,9.295748,9.484379,9.476834,9.484379,9.397609,9.273112,9.408927,10.355856,10.940613,11.355601,11.853588,12.268577,12.027128,12.404391,12.37421,12.562841,13.132507,13.788944,13.615403,13.264549,13.196642,13.313594,12.96274,11.84227,11.695138,12.147853,12.815607,13.290957,12.83447,12.408164,12.174261,12.162943,12.249713,11.8045435,10.861387,10.231359,10.235131,10.702937,10.831206,10.729345,10.804798,11.400873,12.800517,14.068119,14.241659,14.724555,15.99593,17.637022,18.565088,19.24416,20.126955,20.36463,17.799244,16.177015,15.78089,15.531898,15.211224,15.467763,15.878979,16.618414,16.867407,16.293968,15.067864,13.324911,12.362892,12.208215,12.393073,11.955449,12.027128,11.604594,10.872705,10.0276375,9.280658,9.035437,9.397609,9.58624,9.514561,9.774872,10.804798,10.484125,9.424017,8.390318,8.322411,7.6923823,7.5829763,8.390318,9.854096,11.046246,11.3971,10.419991,9.971047,10.54826,11.306557,10.152134,10.427535,11.310329,11.993175,11.6875925,10.423763,10.306811,10.159679,9.220296,7.118943,7.8131065,7.647111,7.8998766,9.344792,12.234623,9.5183325,6.326692,3.7575345,2.2786655,1.7278622,2.2484846,2.1503963,1.6335466,1.1544232,1.418507,2.5993385,3.832987,4.7950063,5.7494807,7.5490227,8.650629,9.201432,9.4127,9.261794,8.503497,8.926031,8.990166,8.477088,7.673519,7.383027,7.8923316,8.013056,8.190369,8.375228,8.024373,7.8508325,7.7037,7.5226145,7.488661,7.9941926,6.7944975,6.0626082,6.205968,6.85486,6.858632,7.2094865,7.8508325,8.145098,7.964011,7.6584287,7.884786,7.7112455,7.2396674,6.7341356,6.628502,6.72659,7.4509344,7.8734684,7.624475,6.900131,6.9189944,6.9982195,7.0170827,7.141579,7.854605,8.273367,7.911195,7.3792543,6.903904,6.330465,6.3116016,6.0626082,5.6363015,5.2288585,5.1835866,6.0211096,6.7756343,7.786698,8.646856,8.179051,7.858378,7.624475,7.5112963,7.7602897,8.809079,9.559832,10.280403,10.925522,11.32542,11.200924,11.457462,11.461235,11.299012,11.117926,11.11038,11.291467,11.004747,10.484125,10.121953,10.453944,11.276376,11.646093,12.034674,12.608112,13.219278,13.800262,13.626721,13.407909,13.0646,11.736636,11.532914,11.69891,11.442371,10.70671,10.148361,10.197406,11.389555,12.166716,11.680047,9.752235,9.627739,9.318384,9.114662,9.220296,9.733373,9.914458,9.5183325,9.250477,8.975075,7.7150183,6.7454534,6.33801,6.228604,6.375736,6.94163,7.141579,7.484888,7.6320205,7.967784,9.627739,11.672502,11.978085,11.076427,9.699419,8.763808,9.842778,11.314102,11.92904,11.174516,9.2995205,8.00551,9.4013815,10.159679,9.57115,9.5183325,10.416218,10.423763,10.220041,10.008774,9.522105,8.929804,8.307321,8.039464,8.322411,9.144843,8.714764,8.345046,8.778898,9.81637,10.295494,9.363655,7.647111,6.930312,7.432071,7.798016,8.20546,7.699928,7.4169807,7.91874,9.224068,10.257768,10.518079,10.608622,10.087999,7.484888,9.06939,8.001738,6.937857,6.7077274,6.3342376,5.7419353,5.2665844,5.2062225,5.5495315,5.9796104,6.651138,7.1038527,7.6508837,8.3525915,9.024119,9.344792,9.556059,9.408927,8.91094,8.314865,7.2698483,7.364164,7.654656,7.828197,8.224322,8.635539,8.394091,8.073418,8.080963,8.66572,8.801534,8.605357,8.333729,8.043237,7.575431,7.1340337,7.073672,7.069899,7.111398,7.515069,5.885295,5.96452,6.2323766,6.0324273,5.560849,6.72659,5.379763,5.3684454,7.0284004,7.2094865,7.0887623,9.371201,12.053536,12.555296,7.7414265,7.3377557,6.752999,9.016574,13.177779,14.317112,8.45068,7.6848373,9.216523,10.985884,11.7026825,12.012038,9.590013,7.5565677,6.990674,6.952948,4.2404304,2.9011486,7.647111,19.149845,34.06303,22.601797,10.431308,5.798525,8.929804,12.012038,7.394345,11.087745,12.494934,9.156161,6.7454534,9.205205,5.96452,3.500996,4.002755,5.3571277,15.335721,17.372938,13.272095,6.858632,3.9914372,4.949684,5.036454,5.383536,6.277648,7.164215,9.216523,9.476834,8.60913,7.7602897,8.567632,8.669493,9.7220545,10.453944,10.521852,10.533169,9.869187,9.616421,9.465516,9.435335,9.861642,9.035437,7.809334,6.8435416,6.3531003,6.1116524,6.4210076,7.194396,7.7904706,7.937603,7.7602897,7.7037,8.235641,9.107117,9.955957,10.31813,10.680302,10.891568,11.491416,12.193124,11.876224,12.162943,12.645839,12.751472,12.215759,11.09529,10.423763,10.084227,9.378746,8.303548,7.5527954,7.3113475,7.533932,8.484633,9.740918,10.212496,9.7069645,9.495697,9.552286,9.688101,9.57115,9.5032425,9.552286,9.318384,9.208978,10.442626,12.15917,12.849561,13.336229,13.792717,13.721037,14.298248,14.045483,13.456953,13.132507,13.754991,13.739901,13.992666,14.079436,13.306048,10.7218,10.789707,10.77839,10.880251,11.310329,12.306303,13.411682,13.343775,12.140307,10.212496,8.36391,7.8244243,8.3525915,9.64283,10.834979,10.480352,9.374973,7.6395655,6.2097406,5.696664,6.379509,8.084735,8.563859,8.167733,7.54525,7.6697464,8.047009,9.0543,10.235131,11.076427,10.997202,11.170743,11.446144,11.710228,11.849815,11.77059,11.623458,11.54046,12.045992,13.132507,14.226569,15.705438,16.776863,16.403374,15.105591,14.947141,14.641558,14.222796,13.966258,13.804035,13.328684,12.513797,11.891314,11.487643,11.299012,11.287694,11.200924,11.864905,12.5326605,12.698656,12.174261,11.065109,12.064855,12.50248,13.023102,13.521088,13.158916,12.027128,11.378237,11.548005,12.196897,12.30253,12.276122,12.404391,12.400619,12.264804,12.283667,11.974312,12.30253,12.811834,13.015556,12.415709,12.985375,12.808062,12.894833,13.604086,14.637785,15.482853,15.433809,14.807553,14.215251,14.577423,14.735873,15.192361,15.362129,14.984866,14.124708,13.634267,13.490907,13.687083,13.879487,13.377728,12.823153,12.174261,11.59705,11.148107,10.774617,10.518079,10.423763,10.167224,9.884277,10.186088,10.012547,9.6201935,9.322156,9.22784,9.216523,9.510788,9.997457,10.412445,10.770844,11.332966,10.054046,8.948667,7.6886096,6.3116016,5.20245,4.2064767,3.6254926,3.1765501,2.7087448,2.2183034,1.5656394,1.0035182,0.5885295,0.33576363,0.19994913,0.124496624,0.071679875,0.060362,0.071679875,0.011317875,0.003772625,0.02263575,0.03772625,0.030181,0.0,0.011317875,0.018863125,0.02263575,0.026408374,0.03772625,0.41876137,1.1317875,1.6939086,1.9089483,1.8863125,2.1390784,2.5880208,2.9011486,2.7389257,1.7693611,1.1242423,0.84884065,0.55080324,0.20372175,0.17731337,0.124496624,0.056589376,0.071679875,0.1358145,0.071679875,0.041498873,0.10940613,0.120724,0.10940613,0.31312788,0.43007925,0.79602385,0.9280658,0.76584285,0.68661773,1.1959221,1.20724,1.1129243,1.0714256,1.0299267,0.94692886,1.1506506,1.0902886,1.026154,1.9881734,1.5580941,1.539231,1.6184561,1.8146327,2.4786146,2.9728284,3.3425457,3.3840446,3.1840954,3.1048703,2.727608,2.9916916,3.3651814,3.5538127,3.4783602,3.3123648,3.4029078,3.8707132,4.3007927,3.7613072,4.13857,4.8402777,5.4212623,5.723072,5.8702044,5.643847,5.142088,4.82896,4.7346444,4.4705606,5.0062733,4.776143,4.5988297,4.8930945,5.692891,6.439871,7.5527954,8.216777,8.322411,8.473316,8.692128,9.107117,9.944639,10.895341,11.148107,10.540714,9.771099,9.703192,10.291721,10.593531,10.917976,10.744436,10.370946,10.336992,11.408418,12.513797,13.253232,13.698401,13.721037,13.000465,13.075918,13.091009,12.845788,12.585477,13.004238,13.13628,13.011784,13.053283,13.075918,12.283667,11.408418,11.593277,12.340257,13.102326,13.29473,12.083718,10.948157,10.314357,10.355856,10.978339,11.548005,11.272603,11.038701,11.204697,11.59705,12.181807,12.487389,12.694883,13.094781,14.079436,14.886778,14.728328,14.747191,15.456445,16.765545,17.425755,18.044466,19.470518,20.428764,17.542706,17.191853,16.84477,16.13929,15.573396,16.497688,17.482344,18.214233,17.701157,16.060064,14.483108,13.472044,12.37421,11.830952,11.751727,11.332966,12.559069,12.510024,11.59705,10.393582,9.639057,9.2844305,9.488152,9.601331,9.439108,9.310839,10.076681,10.080454,9.405154,8.416726,7.779153,7.8017883,8.262049,8.8769865,9.552286,10.38981,11.136789,10.54826,9.850324,9.812597,10.729345,9.903141,9.042982,9.556059,11.257513,12.385528,11.302785,11.785681,11.868678,10.355856,6.828451,7.541477,8.348819,9.903141,11.615912,11.657412,7.594294,4.8855495,3.1124156,2.0900342,1.901403,2.746471,2.746471,2.3163917,2.0447628,2.686109,4.266839,4.036709,4.6931453,6.673774,8.145098,10.585986,11.593277,11.227332,9.952185,8.627994,8.793989,8.926031,8.6581745,8.013056,7.3717093,7.2623034,7.7037,7.956466,7.865923,7.854605,7.865923,7.745199,7.5829763,7.4735703,7.5112963,7.009537,6.5945487,6.6850915,7.1679873,7.4018903,7.4697976,8.224322,8.699674,8.688355,8.744945,9.001483,8.492179,7.6320205,6.903904,6.881268,6.470052,7.2283497,7.8131065,7.6886096,7.122716,7.1000805,6.820906,6.530414,6.560595,7.3415284,8.254503,7.8131065,7.0472636,6.5002327,6.2436943,6.039973,6.039973,5.9003854,5.50426,4.9232755,5.0062733,5.1835866,5.956975,7.0359454,7.3490734,7.039718,7.575431,8.099826,8.337502,8.575176,9.393836,9.820143,10.38981,11.072655,11.299012,11.887542,12.498707,12.604341,12.23085,11.966766,12.095036,12.061082,11.491416,10.767072,10.997202,11.227332,11.559323,11.747954,11.895086,12.457208,13.415455,13.057055,12.66093,12.585477,12.272349,12.015811,12.030901,12.0233555,11.793225,11.216014,10.714255,11.148107,11.646093,11.23865,8.892077,8.714764,8.167733,7.9338303,8.141325,8.386545,8.907167,8.567632,8.341274,8.465771,8.424272,7.1378064,6.511551,6.4436436,6.8359966,7.586749,7.454707,7.8810134,8.6581745,9.627739,10.672756,12.23085,11.672502,10.11818,8.646856,8.273367,9.190115,10.808571,11.480098,10.785934,9.548513,9.691874,9.910686,9.574923,8.5563135,7.232122,9.159933,9.646602,9.424017,9.076936,9.031664,8.963757,8.869441,8.518587,8.122461,8.314865,8.533678,7.937603,7.61693,7.8810134,8.2507305,8.348819,8.431817,8.744945,8.831716,7.5301595,6.7152724,6.903904,7.4999785,8.126234,8.643084,9.1976595,9.725827,10.340765,9.88805,5.9532022,10.838752,8.805306,6.4926877,6.2927384,6.349328,6.63982,6.9567204,7.2962565,7.533932,7.4018903,7.9451485,8.318638,8.597813,8.9788475,9.786189,9.49947,9.408927,9.64283,9.865415,9.314611,7.937603,7.624475,7.61693,7.786698,8.643084,9.050528,8.903395,8.563859,8.420499,8.884532,8.926031,8.869441,8.714764,8.499724,8.265821,7.665974,7.533932,7.4094353,7.2358947,7.356619,5.9230213,5.9909286,6.1720147,5.753253,4.7044635,6.3153744,5.523123,5.572167,7.0963078,8.096053,8.975075,11.170743,14.045483,15.445127,11.706455,8.201687,6.277648,6.907676,9.1825695,10.310584,8.741172,7.9753294,10.152134,13.837989,14.030393,12.574159,9.454198,7.6584287,8.280911,10.487898,6.6813188,4.353609,4.8666863,10.33322,23.597769,13.970031,8.20546,7.677292,9.740918,7.7376537,7.4999785,12.872196,13.924759,9.473062,7.0812173,7.1378064,6.405917,5.617439,5.553304,7.009537,21.4851,26.212198,19.206434,6.428553,1.81086,3.8254418,4.821415,5.783434,6.677546,6.4738245,8.507269,9.322156,8.8618965,7.9791017,8.443134,8.850578,10.072908,10.79348,10.710483,10.544487,10.242677,10.26154,10.170997,9.891823,9.688101,8.76758,7.6886096,6.571913,5.5985756,5.040227,5.583485,7.122716,8.050782,7.9941926,7.809334,7.4169807,7.7640624,8.567632,9.450426,9.944639,10.748209,10.940613,11.249968,11.740409,11.8045435,13.143826,13.962485,13.543724,12.042219,10.469034,9.827688,9.039209,8.367682,7.9300575,7.7112455,7.6131573,7.6207023,8.047009,8.873214,9.752235,9.857869,9.967276,10.495442,11.133017,10.853842,10.510533,10.001229,9.533423,9.654147,11.216014,13.132507,13.913441,14.139798,14.132254,13.932304,13.856852,13.902123,13.622949,13.226823,13.585222,13.947394,12.996693,11.846043,10.876478,9.7220545,10.34831,10.495442,10.453944,10.804798,12.415709,13.86817,13.913441,12.6345215,10.642575,9.065618,8.518587,9.042982,10.235131,11.2801485,10.93684,8.990166,7.3868,6.2814207,5.8928404,6.5341864,7.884786,8.145098,7.643338,7.020855,7.2585306,7.61693,8.846806,10.140816,10.725573,9.876732,10.057818,10.891568,11.54046,11.548005,10.831206,10.970794,10.801025,11.359374,12.913695,14.950912,16.905132,16.818363,15.188588,13.253232,13.000465,13.58145,13.6682205,13.370183,13.004238,13.087236,12.404391,11.314102,10.401127,10.005001,10.246449,11.3820095,12.2270775,12.766563,12.381755,11.3971,11.076427,12.751472,13.788944,14.505743,14.807553,14.222796,12.770335,12.00072,11.898859,12.276122,12.800517,12.521342,12.725064,12.683565,12.355347,12.404391,11.781908,11.940358,12.47607,12.955194,12.894833,12.419481,11.895086,12.061082,12.7477,12.894833,12.577931,12.770335,13.215506,13.72481,14.173752,14.286931,14.634012,14.652876,14.158662,13.36641,13.4644985,13.113645,13.094781,13.170234,12.083718,11.363147,11.219787,10.899114,10.287949,9.933322,9.273112,9.035437,9.163706,9.661693,10.589758,9.514561,8.899622,8.52236,8.424272,8.91094,10.095545,10.355856,10.220041,10.170997,10.63503,9.133525,8.228095,7.352846,6.1908774,4.6554193,4.104616,3.572676,3.059599,2.584248,2.1805773,1.7052265,1.1204696,0.6375736,0.34330887,0.19994913,0.124496624,0.071679875,0.05281675,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.03772625,0.0,0.0,0.1961765,0.41876137,0.6073926,0.7884786,1.0676528,1.2638294,1.3770081,1.5430037,1.6863633,1.5241405,1.3166461,1.5128226,1.1355602,0.31312788,0.27540162,0.1659955,0.071679875,0.049044125,0.060362,0.0,0.03772625,0.10186087,0.10186087,0.041498873,0.030181,0.041498873,0.40367088,0.69039035,0.79602385,0.9318384,1.4298248,1.3091009,1.2864652,1.50905,1.5580941,1.2864652,1.3392819,1.1506506,0.84129536,1.2223305,1.4524606,1.8485862,2.033445,2.161714,2.9313297,2.516341,2.1466236,2.3390274,2.9728284,3.2670932,3.4745877,3.3689542,3.2670932,3.3312278,3.6028569,3.0520537,3.2255943,3.5387223,3.783943,4.1498876,4.478106,4.817642,5.3571277,5.9192486,5.9796104,5.8588867,5.7381625,5.6589375,5.4967146,4.957229,5.349582,5.4212623,5.451443,5.7419353,6.6058664,6.5832305,7.5565677,8.582722,9.084481,8.865668,9.073163,9.25425,9.789962,10.453944,10.38981,10.427535,10.253995,10.321902,10.763299,11.3971,12.057309,12.762791,12.706201,12.030901,11.812089,13.532406,14.739646,15.033911,14.600059,14.222796,13.7700815,13.490907,12.966512,12.442118,12.83447,12.370438,12.1252165,11.989402,11.710228,10.880251,10.612394,11.019837,12.038446,13.174006,13.502225,12.08749,11.185833,10.627484,10.208723,9.65792,10.072908,10.653893,11.019837,11.2801485,12.0233555,12.657157,13.385274,14.1058445,14.86037,15.82239,16.395828,15.954432,15.380992,15.241405,15.777118,17.316349,18.587723,19.625195,19.640285,17.029629,19.7761,20.443855,19.338476,17.63325,17.365393,18.097282,18.829172,18.738628,17.595524,15.777118,15.705438,14.249205,12.913695,12.196897,11.61214,13.456953,13.970031,13.140053,11.589504,10.589758,10.087999,9.680555,9.107117,8.394091,7.858378,8.710991,8.8618965,8.7751255,8.488406,7.5829763,8.13378,8.975075,9.461743,9.537196,9.718282,10.280403,10.70671,10.56335,10.216269,10.804798,11.268831,10.386037,9.280658,9.310839,12.068627,12.559069,12.717519,12.223305,10.589758,7.17176,8.186596,10.269085,12.528888,13.04951,8.91094,5.775889,4.1574326,3.802806,3.9273026,3.218049,3.3538637,2.7200627,2.2069857,2.282438,2.9916916,3.138824,4.3196554,5.458988,6.2889657,7.3377557,9.329701,11.491416,11.747954,10.103089,8.650629,8.262049,8.280911,8.397863,8.360137,7.9791017,7.394345,7.3868,7.435844,7.356619,7.2924843,7.3905725,7.24344,7.3377557,7.5603404,7.1566696,7.0963078,6.8058157,6.590776,6.7077274,7.356619,7.586749,8.14887,8.624221,8.941121,9.367428,9.514561,8.892077,8.099826,7.405663,6.760544,5.9305663,5.7683434,6.145606,6.8058157,7.352846,7.7716074,7.24344,6.692637,6.6850915,7.4169807,7.7716074,7.454707,7.0170827,6.6850915,6.379509,6.439871,6.6549106,6.6058664,6.217286,5.753253,4.8968673,4.3007927,4.5497856,5.6023483,6.7756343,6.006019,6.6850915,7.5075235,7.8432875,7.7225633,8.537451,8.7600355,9.110889,9.846551,10.774617,11.370691,12.427027,13.128735,13.309821,13.441863,12.721292,12.019584,11.45369,11.18206,11.41219,11.291467,11.378237,11.830952,12.370438,12.298758,13.128735,12.694883,12.178034,12.234623,13.015556,12.672247,12.423254,12.344029,12.276122,11.827179,10.933067,9.81637,9.35611,9.454198,9.001483,8.695901,7.9791017,7.6093845,7.7640624,8.058327,8.850578,9.012801,8.986393,8.827943,8.194141,7.5603404,7.0510364,6.888813,7.2585306,8.329956,8.695901,9.431562,10.3634,10.989656,10.453944,9.49947,8.695901,8.333729,8.567632,9.382519,10.201178,11.174516,10.819888,9.280658,8.314865,10.159679,10.144588,9.363655,8.258276,6.620957,8.258276,8.650629,8.903395,9.114662,8.345046,7.466025,8.439363,8.748717,7.9225125,7.5075235,8.167733,8.084735,7.5829763,7.092535,7.141579,6.9944468,7.2057137,8.137552,8.907167,7.3717093,5.3080835,6.0550632,8.001738,9.544742,9.0957985,8.458225,9.473062,10.0276375,9.2995205,7.7376537,11.3971,9.310839,7.394345,7.4509344,7.1566696,7.914967,8.047009,8.243186,8.575176,8.514814,8.050782,8.394091,9.001483,9.688101,10.604849,10.627484,10.4049,10.435081,10.718028,10.740664,9.484379,8.729855,8.590267,9.046755,9.948412,9.789962,9.348565,9.21275,9.250477,8.590267,8.944894,9.318384,9.439108,9.26934,8.986393,8.035691,7.888559,7.533932,6.832224,6.515323,6.0286546,6.3153744,6.439871,5.983383,5.081726,5.873977,5.323174,5.451443,6.8133607,8.499724,7.865923,13.015556,18.648085,20.19109,13.792717,8.09228,8.4544525,9.110889,8.529905,9.382519,8.458225,6.8774953,9.955957,15.9695215,16.188334,14.0907545,9.224068,5.753253,7.997965,20.462717,18.814081,12.936331,8.20546,9.031664,18.859352,16.150608,19.885506,26.853544,29.07562,13.792717,7.567886,13.106099,16.120426,13.109872,11.351829,8.130007,8.52236,9.016574,7.8998766,5.2628117,17.912424,25.32186,18.191597,2.9803739,1.9089483,3.9348478,4.67051,5.7796617,7.069899,6.485142,7.435844,8.314865,8.571404,8.284684,8.16396,8.967529,9.865415,10.250222,10.069136,9.812597,10.103089,10.325675,10.38981,10.03141,8.7751255,7.967784,6.907676,5.9984736,5.3571277,4.821415,5.040227,6.405917,7.5603404,7.8810134,7.492433,6.5530496,6.903904,7.745199,8.699674,9.812597,10.850069,11.136789,11.197151,11.219787,11.046246,13.392818,14.535924,13.309821,10.593531,9.322156,9.322156,8.537451,7.7678347,7.405663,7.432071,7.956466,8.216777,8.2507305,8.2507305,8.544995,9.205205,10.1294985,11.306557,12.076173,11.125471,10.084227,9.239159,9.2844305,10.140816,10.970794,12.838243,13.864397,14.079436,13.932304,14.298248,13.88326,13.834216,14.04171,14.158662,13.59654,13.656902,12.415709,11.23865,10.578441,9.978593,10.955703,11.155652,10.782163,10.853842,13.200415,14.588741,14.407655,12.928786,10.910432,9.567377,8.933576,9.031664,9.646602,10.242677,9.948412,7.8734684,6.651138,6.5832305,7.303802,7.7678347,8.265821,8.492179,8.145098,7.624475,8.024373,8.013056,8.661947,9.314611,9.363655,8.239413,8.473316,9.639057,10.540714,11.0613365,12.162943,12.370438,11.359374,11.151879,12.46098,14.694374,16.403374,15.32063,13.690856,12.683565,12.3893,12.951422,13.385274,13.513543,13.441863,13.5663595,13.223051,11.472552,10.091772,9.7220545,9.857869,12.434572,12.83447,12.89106,12.536433,11.947904,11.555551,12.593022,13.313594,13.932304,14.286931,13.819125,13.65313,12.830698,12.506252,12.849561,13.023102,12.408164,12.377983,12.147853,11.695138,11.732863,11.434827,11.551778,12.498707,13.751218,13.845533,12.4307995,12.0724,11.966766,11.876224,12.098808,12.377983,12.453435,12.725064,13.117417,13.053283,13.317367,13.4644985,13.290957,12.992921,13.147598,12.823153,12.506252,12.313848,12.162943,11.778135,10.748209,9.948412,9.495697,9.446653,9.786189,9.265567,9.250477,9.175024,9.159933,10.0276375,9.861642,9.193887,8.956212,9.21275,9.156161,9.4013815,9.639057,9.65792,9.57115,9.831461,8.329956,7.5603404,6.7869525,5.828706,5.081726,4.881777,3.9122121,3.4444065,3.712263,3.9159849,2.354118,1.3241913,0.69793564,0.35839936,0.17354076,0.090543,0.071679875,0.0452715,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.049044125,0.271629,0.63002837,0.95447415,0.9205205,0.98842776,1.2751472,1.3091009,1.1242423,1.2562841,1.3996439,1.7278622,1.3732355,0.47912338,0.18863125,0.26408374,0.18485862,0.120724,0.10186087,0.0,0.00754525,0.026408374,0.033953626,0.02263575,0.018863125,0.07922512,0.4678055,0.90543,1.2185578,1.3317367,1.7542707,1.7919968,1.418507,1.0487897,1.50905,1.1431054,1.20724,1.3317367,1.297783,0.9997456,1.3204187,1.6939086,1.7429527,1.5958204,1.9051756,2.0447628,1.9542197,1.8033148,1.6712729,1.5430037,1.9089483,2.173032,2.282438,2.323937,2.516341,2.9615107,3.2746384,3.5764484,3.9876647,4.640329,4.6931453,5.406172,6.013564,6.3531003,6.8359966,6.9491754,7.118943,6.9944468,6.360646,5.13077,4.9459114,4.8553686,5.3156285,6.2851934,7.2283497,7.0284004,7.6207023,8.424272,8.963757,8.903395,9.020347,9.74469,10.408672,10.702937,10.661438,11.378237,11.099063,11.3820095,12.064855,11.2650585,11.423509,11.551778,11.517824,11.446144,11.725319,12.362892,13.570132,14.34352,14.407655,14.245432,14.075664,13.373956,13.223051,13.747445,14.079436,13.068373,12.96274,13.275867,13.2607765,11.940358,11.544232,11.763044,12.204442,12.536433,12.464753,11.664956,11.034928,10.306811,9.635284,9.58624,9.552286,10.291721,11.216014,12.042219,12.770335,13.600313,13.970031,14.50197,15.354584,16.248695,17.274849,16.795727,16.433554,16.920223,18.119919,19.413929,20.598532,21.451145,20.53817,15.222542,19.7761,22.149082,23.065828,22.609343,20.232588,18.357594,18.263277,18.787672,19.146072,18.938578,17.165443,15.505488,14.320885,13.739901,13.664448,14.332202,14.9358225,14.864142,13.88326,12.140307,10.944386,9.937095,8.778898,7.6810646,7.4169807,7.8810134,7.8017883,7.7338815,7.7414265,7.424526,7.7678347,8.480861,9.352338,10.272858,11.208468,10.79348,10.974566,10.970794,10.536942,9.95973,9.654147,9.684328,9.774872,9.952185,10.544487,13.113645,13.079691,12.132762,10.601076,7.4773426,10.627484,13.151371,12.958967,9.861642,5.5683947,4.353609,4.357382,4.870459,5.5457587,6.428553,6.700182,4.5196047,2.384299,1.6033657,2.2711203,3.500996,4.0517993,5.458988,7.273621,7.0849895,7.586749,8.692128,9.310839,9.084481,8.394091,8.726082,8.782671,8.971302,9.137298,8.552541,8.360137,7.745199,7.6018395,7.964011,7.99042,7.2170315,6.4134626,6.3719635,6.903904,6.8133607,6.6247296,6.779407,6.9680386,7.183078,7.7338815,8.443134,8.605357,8.850578,9.276885,9.442881,8.786444,8.477088,8.337502,8.179051,7.798016,7.496206,7.3415284,7.220804,7.3151197,8.099826,7.9791017,8.054554,7.726336,7.118943,7.111398,7.141579,7.2472124,7.3075747,7.152897,6.5228686,6.4210076,6.5568223,6.688864,6.6662283,6.4474163,5.6325293,5.198677,5.247721,5.5797124,5.6891184,4.957229,5.036454,5.5985756,6.2814207,6.7077274,7.594294,8.084735,8.318638,8.669493,9.733373,11.106608,11.883769,12.404391,12.879742,13.392818,12.4307995,11.506506,11.11038,11.431054,12.366665,11.834724,11.446144,11.449917,11.883769,12.593022,13.705947,14.25675,13.641812,12.400619,12.234623,12.770335,12.242168,11.917723,12.030901,11.763044,11.529142,10.570895,9.333474,8.52236,9.125979,9.276885,8.959985,8.224322,7.4697976,7.4584794,8.458225,9.4013815,9.616421,8.835487,7.2057137,6.688864,7.073672,7.4018903,7.5905213,8.428044,8.812852,8.4544525,8.60913,9.4127,9.842778,8.597813,7.9526935,7.779153,8.156415,9.382519,9.352338,9.95973,10.016319,9.027891,7.194396,8.782671,10.042727,10.374719,9.6051035,7.99042,7.888559,7.748972,8.031919,8.495952,8.175279,7.405663,7.492433,7.673519,7.8017883,8.375228,7.61693,7.2396674,6.971811,6.6813188,6.360646,6.047518,6.0701537,5.9117036,5.564622,5.5495315,6.2135134,6.3455553,6.3945994,6.8058157,8.031919,7.6886096,8.688355,9.940866,9.831461,6.2097406,11.329193,9.559832,7.5263867,7.5829763,7.828197,8.6732645,8.710991,8.627994,8.60913,8.345046,7.7414265,7.816879,8.499724,9.333474,9.469289,10.510533,11.185833,11.219787,10.801025,10.570895,10.133271,9.416472,9.0957985,9.34102,9.812597,10.152134,9.944639,9.639057,9.446653,9.322156,9.258021,9.64283,9.567377,9.020347,8.8769865,7.9828744,7.756517,7.6131573,7.2698483,6.749226,7.0585814,7.0887623,7.1000805,7.01331,6.4134626,6.326692,6.3229194,6.379509,6.722818,7.8508325,8.175279,9.344792,12.344029,15.116908,12.596795,7.4735703,7.854605,7.8319697,7.752744,14.181297,10.087999,6.4021444,10.880251,17.625704,7.0963078,21.058792,15.32063,8.246958,7.8432875,11.732863,21.609596,23.548725,20.289177,19.63274,34.459156,38.446823,56.99682,70.13687,61.546604,18.542452,6.379509,7.564113,10.831206,12.370438,15.807299,8.865668,8.643084,10.623712,11.25374,7.9753294,10.435081,11.936585,8.843033,3.138824,2.4559789,3.270866,4.3649273,6.3116016,7.956466,6.4247804,7.356619,7.9526935,8.258276,8.394091,8.567632,9.125979,10.110635,10.431308,10.174769,10.593531,10.47658,10.103089,9.933322,9.854096,9.152389,8.024373,6.458734,5.3194013,4.90064,4.919503,5.13077,5.8400235,6.507778,6.8359966,6.749226,6.432326,6.881268,7.816879,8.741172,8.944894,9.073163,9.405154,10.133271,10.812344,10.340765,12.253486,13.626721,12.577931,9.691874,8.043237,7.884786,7.7602897,7.594294,7.3981175,7.2962565,8.00551,8.488406,8.646856,8.605357,8.692128,8.812852,9.480607,10.397354,10.933067,10.099318,9.58624,9.371201,9.5032425,9.929549,10.506761,12.042219,13.298503,13.430545,12.826925,13.124963,12.868423,12.902377,13.117417,13.241914,12.826925,12.672247,12.0082655,11.193378,10.714255,11.200924,11.3669195,10.989656,10.733118,10.993429,11.879996,13.087236,13.230596,12.325166,10.782163,9.420244,9.001483,8.567632,8.52236,8.654402,8.118689,7.3905725,6.5832305,6.579458,7.2170315,7.2924843,7.2924843,7.1906233,7.1604424,7.432071,8.280911,8.379,8.326183,8.390318,8.714764,9.352338,9.612649,9.371201,9.190115,9.661693,11.404645,12.128989,10.933067,10.137043,10.850069,12.985375,14.109617,14.34352,14.169979,13.649357,12.438345,12.5326605,12.600568,12.483616,12.457208,13.223051,12.196897,11.016065,10.412445,10.480352,10.661438,12.464753,12.121444,12.042219,11.895086,11.634775,11.498961,12.487389,13.113645,13.385274,13.445636,13.562587,13.853079,12.853333,12.151625,12.23085,12.464753,11.849815,11.887542,11.744182,11.415963,11.721546,11.883769,11.921495,12.381755,13.023102,12.81938,12.204442,12.004493,11.861133,11.664956,11.563096,12.113899,12.457208,12.593022,12.653384,12.879742,12.936331,12.838243,12.770335,12.679792,12.294985,11.766817,11.631002,11.559323,11.268831,10.514306,10.272858,9.665465,9.201432,9.152389,9.540969,9.242931,9.646602,9.861642,9.680555,9.574923,9.220296,9.125979,9.06939,9.005256,9.0957985,8.986393,9.06939,9.250477,9.239159,8.567632,8.126234,7.598067,6.72659,5.8702044,5.994701,4.961002,5.111907,6.066381,6.670001,4.979865,2.5691576,1.3091009,0.6413463,0.271629,0.13958712,0.06790725,0.03772625,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.15845025,0.35462674,0.56589377,0.86770374,0.94692886,1.0638802,0.98465514,0.8262049,1.0336993,1.2449663,1.2713746,1.0827434,0.7394345,0.3772625,0.32444575,0.211267,0.116951376,0.060362,0.0,0.0,0.003772625,0.033953626,0.08299775,0.1056335,0.07922512,0.43007925,0.90543,1.2411937,1.1581959,1.6373192,1.7919968,1.4600059,0.9808825,1.2223305,1.056335,0.91297525,0.97333723,1.1355602,1.0110635,1.1242423,1.5807298,1.7919968,1.750498,2.04099,2.425798,2.3578906,2.233394,2.214531,2.2409391,2.3428001,2.1202152,2.0598533,2.2673476,2.4522061,2.5276587,3.0030096,3.712263,4.4215164,4.8440504,4.961002,5.2326307,5.330719,5.4438977,6.2814207,6.8397694,7.3075747,7.039718,6.1078796,5.292993,5.168496,4.745962,5.2137675,6.439871,6.971811,7.3377557,7.7112455,7.9791017,8.262049,8.918486,8.4544525,8.771353,9.367428,9.993684,10.646348,11.785681,11.774363,12.057309,12.411936,10.963248,11.000975,11.148107,11.2801485,11.415963,11.721546,11.98563,12.4307995,12.894833,13.234368,13.343775,13.966258,13.788944,13.81158,14.124708,13.920986,13.355092,13.332457,13.619176,13.781399,13.204187,12.7477,12.102581,11.781908,11.623458,10.770844,10.736891,10.367173,9.952185,9.827688,10.3634,10.223814,10.970794,12.162943,13.385274,14.245432,15.147089,15.094273,15.120681,15.62244,16.376965,17.863379,18.052011,17.670975,17.584206,18.791445,18.68204,19.440336,20.492899,20.432537,17.033401,19.794964,22.115128,23.348776,22.884743,20.16468,17.172989,17.67852,18.648085,18.749947,18.365139,16.724047,16.135517,15.807299,15.475307,15.39231,15.245177,14.901869,14.735873,14.603831,13.853079,12.200669,10.7218,9.295748,7.986647,7.043491,7.5263867,7.533932,7.273621,7.043491,7.2396674,8.284684,9.092027,9.835234,10.676529,11.7555,11.3820095,11.276376,11.102836,10.748209,10.336992,8.801534,8.401636,9.288202,10.668983,10.812344,13.8719425,14.758509,14.102073,12.215759,9.092027,11.891314,13.728582,12.37421,8.280911,4.5460134,4.5460134,4.9760923,5.1081343,5.349582,7.2698483,7.1076255,5.5382137,3.8178966,2.6672459,2.3013012,3.3764994,3.3576362,4.142342,5.798525,6.541732,8.016829,8.809079,9.133525,8.937348,7.865923,8.669493,8.511042,8.2507305,8.246958,8.367682,8.477088,8.118689,8.07719,8.3525915,8.152642,7.1076255,6.1342883,5.798525,6.089017,6.3908267,6.436098,6.651138,6.8737226,7.1302614,7.61693,8.401636,8.507269,8.688355,8.990166,8.7751255,7.9715567,7.7338815,7.865923,7.997965,7.598067,7.092535,7.326438,7.654656,7.937603,8.560086,8.428044,8.763808,8.809079,8.431817,8.141325,7.696155,7.4697976,7.5112963,7.484888,6.688864,6.375736,6.983129,7.7338815,7.9941926,7.3075747,6.3644185,6.19465,6.145606,5.9532022,5.7381625,4.9949555,4.606375,4.7308717,5.20245,5.5193505,6.48137,7.0472636,7.4018903,7.8923316,9.035437,10.714255,11.419736,11.996947,12.566614,12.513797,11.676274,11.427281,11.729091,12.494934,13.592768,13.200415,12.472299,12.038446,12.147853,12.691111,13.585222,14.071891,13.7851715,13.019329,12.762791,13.81158,12.875969,11.921495,11.661184,11.521597,11.155652,10.774617,9.778644,8.484633,8.122461,8.14887,8.348819,7.91874,7.092535,7.152897,8.216777,9.039209,9.031664,8.047009,6.379509,6.1720147,6.7869525,7.405663,7.726336,7.960239,8.013056,7.6886096,7.91874,8.729855,9.231613,8.654402,8.941121,9.1976595,9.314611,9.978593,9.903141,10.329447,10.657665,9.982366,7.0963078,7.586749,9.26934,10.137043,9.273112,6.8133607,7.9300575,8.213005,7.9036493,7.4094353,7.326438,8.039464,8.379,8.062099,7.605612,8.296002,7.1000805,6.590776,6.5002327,6.304056,5.2326307,5.7909794,6.300284,6.156924,5.383536,4.5912848,5.832478,6.039973,5.7079816,5.723072,7.356619,6.937857,8.107371,9.1976595,8.933576,6.405917,8.511042,7.84706,8.265821,9.771099,8.507269,8.82417,8.82417,8.688355,8.526133,8.394091,7.6395655,7.809334,8.571404,9.378746,9.488152,9.654147,10.382264,10.789707,10.601076,10.163452,9.797507,9.646602,9.74469,9.895596,9.654147,10.26154,10.386037,10.163452,9.808825,9.616421,9.378746,9.548513,9.25425,8.511042,8.209232,8.171506,7.888559,7.7301087,7.7037,7.435844,7.77538,7.7301087,7.7301087,7.726336,7.201941,7.213259,7.066127,6.828451,6.832224,7.6810646,9.046755,9.442881,9.906913,10.646348,11.046246,8.231868,7.9225125,7.8923316,9.163706,16.022339,14.705692,11.306557,11.148107,12.506252,6.6247296,20.300495,15.818617,8.597813,6.598321,10.329447,14.890551,16.22606,16.316603,18.448135,27.200626,30.501673,53.239285,72.67962,66.730194,13.936077,5.089271,4.4101987,6.930312,10.495442,15.758255,9.710737,11.563096,13.539951,12.555296,10.216269,9.099571,8.213005,6.1644692,3.6179473,3.289729,3.5160866,4.7535076,6.8850408,8.3525915,6.1342883,7.2962565,7.567886,7.699928,8.07719,8.703445,8.537451,9.623966,10.193633,9.989911,10.238904,9.918231,9.963503,9.87296,9.416472,8.631766,7.462252,6.1606965,5.2364035,4.878004,4.9723196,4.8138695,5.251494,5.9192486,6.511551,6.771862,6.628502,6.934085,7.5565677,8.29223,8.884532,8.567632,8.858124,9.903141,11.004747,10.646348,11.664956,12.66093,11.925267,9.789962,8.646856,8.507269,8.194141,7.828197,7.496206,7.2358947,8.578949,9.129752,9.454198,9.58624,9.031664,8.627994,9.159933,9.839006,10.103089,9.6051035,9.835234,9.65792,9.291975,9.42779,11.242422,12.498707,12.966512,12.883514,12.604341,12.611885,12.766563,12.970284,12.97783,12.702429,12.223305,11.962994,12.1252165,12.113899,11.879996,11.891314,11.170743,10.423763,10.412445,10.993429,11.129244,11.966766,12.359119,11.993175,10.974566,9.842778,9.21275,8.511042,7.8734684,7.3075747,6.7152724,6.911449,6.692637,6.7756343,7.1378064,6.9869013,6.9982195,6.862405,6.8397694,7.0774446,7.586749,8.088508,8.639311,9.242931,9.906913,10.642575,10.642575,10.416218,9.940866,9.737145,10.850069,11.336739,10.510533,10.080454,10.910432,13.015556,13.962485,13.837989,13.12119,12.291212,11.838497,11.827179,11.487643,11.18206,11.2801485,12.147853,11.25374,10.797253,10.49167,10.193633,9.910686,12.242168,11.54046,11.193378,11.087745,11.1631975,11.427281,12.174261,12.811834,13.079691,13.102326,13.392818,13.226823,12.083718,11.302785,11.2650585,11.389555,11.295239,11.400873,11.321648,11.065109,11.000975,11.133017,11.261286,11.449917,11.551778,11.219787,11.299012,11.336739,11.234878,11.000975,10.740664,11.106608,11.389555,11.6008215,11.793225,12.083718,12.049765,12.162943,12.347801,12.351574,11.747954,11.491416,11.174516,10.940613,10.601076,9.635284,9.967276,9.612649,9.246704,9.1976595,9.484379,9.578695,10.084227,10.20495,9.782416,9.2844305,8.907167,9.333474,9.378746,9.039209,9.495697,9.280658,9.220296,9.322156,9.201432,8.088508,8.179051,7.564113,6.7152724,6.2625575,6.9869013,5.934339,7.492433,9.476834,9.446653,4.6742826,2.1843498,1.1280149,0.7130261,0.44894236,0.1358145,0.06413463,0.026408374,0.018863125,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.13204187,0.2565385,0.8224323,0.7809334,0.7432071,0.66775465,0.6149379,0.754525,0.8337501,0.7054809,0.633801,0.5998474,0.33576363,0.23013012,0.14335975,0.071679875,0.018863125,0.0,0.0,0.0,0.03772625,0.1056335,0.1659955,0.09808825,0.331991,0.7130261,1.0374719,1.0450171,1.3770081,1.448688,1.2562841,0.94315624,0.7809334,0.784706,0.784706,0.8601585,0.9997456,1.1091517,1.0110635,1.4750963,1.7769064,1.841041,2.2258487,2.686109,2.655928,2.6031113,2.686109,2.757789,2.886058,2.4107075,2.1956677,2.5012503,2.9916916,2.8898308,3.5047686,4.134797,4.5535583,5.040227,5.481624,5.3344917,5.1043615,5.1647234,5.7872066,6.4474163,7.0548086,6.937857,6.221059,5.828706,5.523123,5.342037,5.80607,6.730363,7.194396,7.956466,8.20546,8.07719,8.00551,8.707218,8.156415,8.20546,8.533678,9.125979,10.272858,11.3669195,11.563096,11.808316,12.004493,11.019837,10.876478,10.853842,10.963248,11.114153,11.106608,11.627231,11.98563,12.0724,12.068627,12.442118,13.302276,13.702174,13.902123,13.996439,13.8870325,13.215506,12.770335,12.853333,13.317367,13.570132,13.306048,12.204442,11.306557,10.79348,9.971047,10.152134,10.054046,9.97482,10.201178,10.997202,11.415963,12.287439,13.404137,14.584969,15.675257,16.58446,16.686321,16.542961,16.52787,16.810818,18.014284,18.421728,18.070873,17.682293,18.666948,18.285913,18.75372,19.942095,21.009748,20.406128,21.553007,22.50748,22.53389,21.292696,18.832945,17.429527,18.700903,19.470518,18.76881,17.833199,17.048492,16.97304,17.033401,16.840998,16.192106,16.16947,15.513034,14.852824,14.483108,14.381247,12.894833,11.299012,9.793735,8.379,6.8925858,7.1340337,7.33021,7.224577,7.01331,7.3490734,8.873214,9.842778,10.514306,11.065109,11.608367,11.415963,11.261286,10.872705,10.321902,10.001229,8.688355,8.114917,9.21275,11.336739,12.283667,15.584714,16.580687,14.396337,10.63503,9.367428,10.329447,10.891568,9.480607,6.6134114,4.878004,4.9459114,5.481624,5.5080323,5.462761,7.1906233,5.873977,5.160951,4.666737,4.0291634,2.9124665,2.8407867,2.5012503,2.9803739,4.4139714,5.994701,8.537451,9.789962,9.805053,8.918486,7.752744,8.612903,8.458225,8.141325,8.13378,8.495952,8.66572,8.484633,8.326183,8.194141,7.7376537,7.009537,6.398372,5.9607477,5.764571,5.926794,6.1720147,6.4134626,6.7379084,7.1679873,7.6584287,8.428044,8.537451,8.66572,8.831716,8.409182,7.6395655,7.322665,7.443389,7.6810646,7.4094353,6.7756343,6.9189944,7.220804,7.5075235,8.065872,8.118689,8.465771,8.782671,8.850578,8.567632,8.160188,7.696155,7.4697976,7.352846,6.79827,6.5832305,7.5490227,8.582722,8.827943,7.7187905,6.9567204,6.964266,6.952948,6.6586833,6.300284,5.6778007,5.20245,5.0666356,5.221313,5.3873086,6.0550632,6.436098,6.85486,7.5188417,8.529905,9.895596,10.533169,11.083972,11.593277,11.487643,11.257513,11.9064045,12.838243,13.641812,14.068119,13.483362,12.706201,12.106354,11.830952,11.819634,12.679792,12.679792,12.73261,13.091009,13.347548,14.136025,13.547497,12.698656,12.057309,11.491416,10.993429,10.767072,10.050273,8.831716,7.84706,7.360391,7.5075235,7.2887115,6.741681,6.937857,7.805561,8.224322,7.9036493,7.043491,6.326692,6.7379084,7.1981683,7.5263867,7.575431,7.2283497,7.1076255,7.2358947,7.8395147,8.699674,9.152389,8.718536,9.318384,9.793735,9.895596,10.26154,10.287949,10.072908,10.167224,10.057818,8.16396,7.598067,8.805306,9.544742,8.635539,5.9984736,7.3415284,7.8696957,7.5226145,6.771862,6.6322746,7.7640624,8.66572,8.60913,7.9526935,8.107371,7.1038527,6.4926877,6.326692,6.217286,5.3344917,5.7117543,5.8173876,5.8173876,5.515578,4.398881,4.8025517,5.2590394,5.2590394,5.292993,6.8435416,6.4511886,7.443389,8.296002,8.182823,6.9982195,6.730363,7.2660756,9.107117,10.853842,9.208978,8.718536,8.458225,8.311093,8.126234,7.7376537,7.322665,7.647111,8.216777,8.843033,9.635284,9.386291,9.582467,9.857869,9.88805,9.382519,9.144843,9.371201,9.850324,10.186088,9.786189,10.601076,10.79348,10.555805,10.193633,10.1294985,9.473062,9.186342,8.627994,7.888559,7.786698,8.22055,8.00551,7.745199,7.696155,7.7602897,7.8395147,7.9753294,8.194141,8.333729,8.0206,8.235641,7.9300575,7.4509344,7.2094865,7.6584287,9.465516,10.687846,10.457717,9.616421,10.7218,10.133271,8.959985,8.492179,10.084227,15.16218,17.16167,15.271586,13.973803,13.641812,10.544487,22.10381,29.44911,21.74541,6.4436436,9.273112,10.110635,9.767326,12.193124,16.822134,18.576405,23.262005,38.824085,52.179176,47.923656,8.367682,8.29223,6.368191,7.6697464,12.611885,16.97304,10.582213,14.358611,16.090246,12.792972,10.70671,10.216269,8.288457,5.7117543,3.6669915,3.7462165,4.4630156,5.723072,7.3453007,8.22055,6.3116016,7.488661,7.699928,7.5527954,7.6093845,8.394091,7.99042,9.171251,10.008774,9.933322,9.718282,9.348565,9.635284,9.691874,9.0957985,7.865923,6.7567716,5.975838,5.5080323,5.2552667,5.0439997,4.768598,4.8629136,5.304311,6.0324273,6.9567204,7.039718,7.4811153,7.865923,8.213005,8.975075,8.707218,9.118435,10.223814,11.329193,11.012292,11.151879,11.676274,11.16697,9.786189,9.273112,9.650374,9.21275,8.537451,7.9225125,7.3717093,8.899622,9.635284,9.982366,9.884277,8.83926,8.778898,9.34102,9.789962,9.839006,9.665465,10.159679,10.310584,9.955957,9.854096,11.69891,12.642066,12.551523,12.562841,12.770335,12.2270775,12.445889,12.785426,12.73261,12.215759,11.5857315,11.502733,12.294985,12.823153,12.66093,12.083718,11.102836,10.397354,10.408672,10.884023,10.880251,11.393328,11.781908,11.551778,10.70671,9.737145,9.042982,8.3525915,7.5565677,6.72659,6.0814714,6.4926877,6.7379084,6.9793563,7.115171,6.8133607,6.8359966,6.79827,6.8661776,7.118943,7.5490227,8.186596,8.98262,9.8239155,10.502988,10.748209,10.552032,10.782163,10.70671,10.435081,10.899114,10.540714,10.20495,10.469034,11.536687,13.234368,13.79649,13.083464,12.00072,11.208468,11.125471,10.884023,10.627484,10.601076,10.850069,11.197151,10.61994,10.63503,10.570895,10.18986,9.703192,12.166716,11.559323,10.872705,10.54826,10.740664,11.314102,11.619685,12.310076,12.89106,13.140053,13.102326,11.910177,10.789707,10.344538,10.49167,10.461489,11.046246,11.117926,10.9594755,10.608622,9.846551,9.548513,9.842778,10.193633,10.325675,10.238904,10.238904,10.397354,10.336992,10.061591,9.944639,10.069136,10.016319,10.378491,10.967021,10.831206,10.948157,11.480098,11.796998,11.717773,11.510279,11.714001,10.978339,10.378491,10.152134,9.665465,9.861642,9.488152,9.224068,9.322156,9.58624,10.061591,10.235131,9.891823,9.310839,9.2844305,9.2995205,9.759781,9.797507,9.556059,10.220041,9.899368,9.7296,9.563604,9.1825695,8.299775,8.024373,7.2094865,6.7944975,7.145352,8.050782,8.420499,11.050018,12.562841,10.49167,3.2444575,1.4071891,0.8601585,0.8186596,0.7167987,0.20372175,0.08299775,0.041498873,0.041498873,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.08299775,0.20749438,0.6488915,0.44894236,0.39989826,0.4074435,0.42630664,0.4376245,0.36971724,0.34330887,0.271629,0.15845025,0.071679875,0.05281675,0.033953626,0.018863125,0.011317875,0.0,0.0,0.0,0.0150905,0.060362,0.150905,0.14713238,0.23013012,0.41876137,0.7054809,1.0751982,1.1242423,0.95824677,0.8639311,0.83752275,0.5772116,0.62248313,0.95447415,1.1393328,1.1129243,1.1732863,1.0714256,1.5354583,1.7580433,1.7014539,2.1164427,2.5767028,2.6446102,2.6936543,2.7653341,2.5767028,2.867195,2.7087448,2.5125682,2.6898816,3.6481283,3.802806,4.3649273,4.4630156,4.3083377,5.1798143,5.934339,5.670255,5.5268955,5.7909794,5.885295,6.398372,6.862405,7.0170827,6.8699503,6.7039547,6.115425,6.5756855,7.0548086,7.3377557,8.001738,8.552541,8.605357,8.495952,8.43559,8.465771,8.473316,8.710991,8.82417,9.024119,10.091772,10.608622,10.887795,11.136789,11.344283,11.287694,10.985884,10.631257,10.555805,10.665211,10.435081,11.193378,12.042219,12.027128,11.427281,11.766817,12.106354,12.713746,13.140053,13.389046,13.894578,12.838243,11.917723,11.691365,12.147853,12.67602,12.921241,12.136535,11.106608,10.401127,10.359629,10.303039,10.284176,10.291721,10.465261,11.125471,12.336484,13.52486,14.50197,15.422491,16.776863,17.738882,18.414183,18.459454,18.033148,17.787928,18.187824,18.35382,18.119919,17.855835,18.43682,19.04421,19.523335,20.711712,22.465982,23.650587,24.623924,23.933533,22.352802,20.368402,18.146326,19.557287,20.790936,20.77962,19.568605,18.342503,18.399092,18.150099,17.897333,17.482344,16.28265,17.08999,16.946632,15.845025,14.452927,14.128481,13.298503,11.895086,10.340765,8.801534,7.17176,6.79827,7.183078,7.5829763,7.7678347,7.997965,9.318384,10.242677,10.921749,11.283921,11.019837,10.963248,10.876478,10.321902,9.390063,8.733627,9.027891,9.118435,10.035183,11.846043,13.630494,17.89356,17.584206,12.47607,6.5568223,7.9941926,6.7114997,6.047518,5.2326307,4.5912848,5.5495315,4.9949555,5.5268955,6.255012,6.6850915,6.730363,4.22534,3.640583,4.5535583,5.383536,3.3878171,2.8106055,2.4408884,2.848332,4.0895257,5.692891,8.461998,10.49167,10.427535,8.782671,7.911195,8.692128,8.926031,9.1976595,9.559832,9.548513,9.559832,9.024119,8.337502,7.6810646,7.0359454,6.730363,6.752999,6.56814,6.1305156,5.8664317,6.096562,6.368191,6.8435416,7.462252,7.937603,8.537451,8.563859,8.586494,8.643084,8.231868,7.537705,7.141579,7.152897,7.3981175,7.4471617,7.118943,6.888813,6.6134114,6.488915,7.066127,7.213259,7.4773426,7.9413757,8.356364,8.126234,8.096053,7.8017883,7.3151197,6.8359966,6.6850915,6.8246784,7.6923823,8.469543,8.575176,7.6697464,7.3490734,7.394345,7.4735703,7.352846,6.907676,6.5341864,6.330465,6.205968,6.1342883,6.1305156,6.221059,6.2851934,6.6058664,7.24344,8.00551,8.854351,9.454198,9.910686,10.321902,10.785934,11.555551,12.898605,13.958713,14.226569,13.551269,12.540206,11.955449,11.529142,11.087745,10.574668,11.415963,11.272603,11.706455,12.81938,13.234368,13.068373,13.355092,13.370183,12.777881,11.61214,11.295239,10.684074,9.884277,9.050528,8.360137,7.432071,7.152897,6.888813,6.5945487,6.8397694,7.2887115,7.375482,7.0246277,6.643593,7.149124,8.114917,8.209232,7.816879,7.2057137,6.5002327,6.5643673,7.175533,8.096053,9.076936,9.876732,8.873214,8.858124,9.118435,9.333474,9.574923,9.639057,8.771353,8.507269,9.099571,9.495697,8.575176,8.778898,8.89585,8.235641,6.6360474,6.7114997,6.7152724,6.696409,6.673774,6.628502,6.8246784,7.835742,8.492179,8.473316,8.296002,7.7640624,7.0585814,6.4926877,6.2021956,6.1305156,5.621211,4.6742826,4.478106,4.930821,4.640329,3.7198083,4.323428,4.8327327,5.081726,6.3531003,6.4210076,6.790725,7.352846,7.6886096,7.073672,6.700182,7.5075235,9.163706,10.484125,9.408927,8.488406,8.001738,7.907422,7.8017883,6.9152217,6.888813,7.4169807,7.7150183,7.937603,9.175024,9.507015,9.371201,9.291975,9.242931,8.635539,8.763808,8.971302,9.476834,10.099318,10.287949,11.227332,11.208468,10.850069,10.642575,10.948157,9.6201935,8.778898,7.956466,7.3453007,7.786698,8.009283,7.8131065,7.4169807,7.1340337,7.3717093,7.2698483,7.677292,8.243186,8.661947,8.684583,8.892077,8.677037,8.197914,7.752744,7.77538,9.310839,11.559323,12.223305,11.355601,11.393328,11.879996,10.574668,9.597558,10.295494,13.223051,15.83748,16.784409,18.97253,20.62494,15.294222,26.729048,47.301174,39.329617,9.224068,7.4999785,9.952185,9.812597,12.494934,17.003222,15.916705,23.778856,27.528845,26.449873,20.104319,8.326183,14.977322,12.472299,13.751218,20.530624,23.292187,15.377219,18.670721,19.123436,13.698401,10.355856,11.517824,8.869441,5.560849,3.591539,3.7877154,5.6098933,6.749226,7.4735703,7.7112455,7.039718,7.779153,8.126234,7.752744,7.152897,7.6584287,7.6810646,8.827943,9.684328,9.737145,9.367428,9.092027,9.110889,9.125979,8.729855,7.4207535,6.571913,6.1078796,5.9720654,5.87775,5.292993,5.1835866,4.859141,4.7120085,5.1835866,6.771862,7.4584794,8.341274,8.729855,8.695901,9.065618,8.956212,9.567377,10.555805,11.287694,10.884023,10.393582,10.695392,10.419991,9.548513,9.442881,10.419991,9.997457,9.144843,8.360137,7.6584287,8.695901,9.58624,9.835234,9.303293,8.182823,9.073163,9.789962,10.11818,10.144588,10.253995,10.250222,10.850069,11.057564,10.876478,11.299012,11.812089,11.812089,12.128989,12.51757,11.668729,11.691365,12.132762,12.223305,11.747954,11.050018,11.461235,12.453435,12.96274,12.645839,11.891314,11.091517,10.725573,10.612394,10.631257,10.7218,11.027383,11.1631975,10.748209,9.842778,8.937348,8.465771,7.9941926,7.462252,6.858632,6.187105,6.2851934,6.832224,7.2358947,7.175533,6.6247296,6.515323,6.670001,7.039718,7.537705,8.043237,8.45068,8.733627,9.125979,9.544742,9.593785,9.522105,10.020092,10.510533,10.759526,10.884023,9.789962,9.933322,10.808571,11.932813,12.83447,12.792972,11.947904,11.276376,10.985884,10.514306,9.955957,10.186088,10.725573,11.076427,10.733118,10.299266,10.431308,10.63503,10.61994,10.303039,12.313848,11.668729,11.140562,10.521852,10.095545,10.61994,11.02361,11.774363,12.336484,12.491161,12.344029,10.295494,9.514561,9.612649,10.167224,10.740664,11.231105,11.299012,10.948157,10.419991,10.178542,9.846551,10.012547,10.299266,10.555805,10.850069,10.506761,10.220041,10.170997,10.310584,10.359629,11.129244,11.268831,11.408418,11.551778,11.0613365,11.306557,11.46878,11.3971,11.083972,10.680302,10.668983,10.023865,9.627739,9.797507,10.299266,10.020092,9.435335,9.099571,9.1825695,9.476834,9.903141,9.590013,9.303293,9.393836,9.797507,9.820143,9.669238,9.627739,9.831461,10.269085,9.646602,9.288202,9.016574,8.59404,7.752744,7.092535,6.8359966,7.5263867,8.831716,9.552286,12.042219,15.448899,14.551015,8.710991,1.8787673,0.8526133,0.62248313,0.513077,0.33953625,0.41121614,0.15467763,0.056589376,0.030181,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06790725,0.16222288,0.1358145,0.211267,0.19240387,0.23390275,0.3169005,0.24522063,0.29426476,0.21503963,0.1358145,0.1056335,0.1056335,0.071679875,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.090543,0.150905,0.20372175,0.19240387,0.2678564,0.7922512,0.8563859,0.58475685,0.5319401,0.845068,1.297783,1.4298248,1.3468271,1.297783,1.297783,1.1129243,1.3204187,2.1164427,2.2484846,1.7995421,2.1654868,2.5578396,2.5993385,3.0897799,3.7462165,3.2331395,2.8332415,3.1161883,3.0407357,2.8181508,3.904667,3.6481283,3.6669915,3.7763977,4.06689,4.8968673,5.5080323,5.1043615,5.168496,5.9003854,6.1795597,7.0359454,6.983129,6.79827,6.9227667,7.462252,7.643338,8.047009,8.20546,8.122461,8.269594,8.001738,7.5301595,7.9791017,9.001483,8.820397,9.295748,9.725827,10.18986,10.714255,11.276376,10.740664,11.310329,11.570641,11.204697,10.970794,11.117926,11.106608,11.046246,11.106608,11.521597,11.2650585,11.574413,11.691365,11.363147,10.86516,10.559577,11.068882,11.623458,11.955449,12.283667,12.626976,12.491161,11.710228,10.785934,10.895341,11.921495,11.864905,11.283921,10.774617,10.970794,11.117926,10.54826,10.310584,10.646348,11.000975,12.08749,13.6682205,15.041456,16.192106,17.7917,18.987621,19.68933,19.647831,19.180025,19.180025,19.47429,20.051502,19.844007,18.934805,18.568861,19.425245,20.096773,21.4436,23.492136,25.419947,26.434784,25.450129,23.933533,22.356575,20.232588,21.526598,21.247423,20.447628,19.50447,18.112373,18.636768,19.097027,18.542452,17.244669,16.708956,17.96524,17.912424,16.893814,15.645076,15.290449,14.9358225,13.664448,11.936585,10.054046,8.14887,7.2094865,7.786698,8.526133,8.926031,9.352338,10.001229,10.26154,10.514306,10.676529,10.238904,10.789707,10.386037,9.597558,8.771353,8.024373,9.307066,10.435081,11.336739,12.064855,12.785426,19.304522,16.98813,10.997202,6.1644692,7.020855,4.2102494,3.1161883,2.848332,3.3764994,5.523123,5.010046,4.9760923,6.72659,8.511042,5.5080323,3.2972744,2.0975795,4.538468,7.575431,2.4710693,5.05909,4.82896,4.063117,4.214022,5.873977,8.499724,10.665211,10.653893,8.763808,7.322665,8.643084,9.540969,10.597303,11.623458,11.672502,11.476325,10.103089,8.635539,7.5490227,6.6850915,5.926794,6.270103,6.72659,6.9152217,7.0510364,7.0849895,7.1038527,7.33021,7.7187905,7.9489207,7.828197,7.6508837,7.515069,7.3679366,6.9869013,6.587003,6.330465,6.379509,6.6662283,6.8963585,7.213259,7.5792036,7.435844,6.9793563,7.1264887,7.039718,7.3490734,8.062099,8.688355,8.224322,7.9300575,7.986647,7.454707,6.4436436,6.089017,6.3945994,6.670001,7.01331,7.413208,7.7678347,7.533932,7.594294,7.594294,7.432071,7.2472124,7.0510364,7.1679873,7.1868505,6.8737226,6.1795597,5.9494295,5.8702044,6.0248823,6.4549613,7.1868505,8.311093,9.129752,9.778644,10.295494,10.650121,12.543978,14.203933,14.596286,13.70972,12.574159,11.962994,11.589504,11.555551,11.563096,10.940613,10.710483,11.695138,13.019329,13.600313,12.162943,10.940613,11.23865,11.857361,12.015811,11.3669195,11.393328,10.453944,9.424017,8.639311,7.91874,7.333983,7.360391,7.2283497,6.900131,7.0963078,7.145352,7.0359454,7.3000293,7.9451485,8.469543,9.042982,8.590267,7.7414265,6.85486,6.013564,6.477597,7.5603404,8.586494,9.608876,11.427281,10.220041,9.480607,9.088254,8.661947,7.537705,7.805561,7.809334,8.182823,8.873214,9.156161,9.031664,8.424272,7.914967,7.7716074,7.9791017,8.262049,6.930312,6.0286546,6.3719635,7.567886,7.3377557,7.277394,7.364164,7.798016,9.016574,8.835487,8.167733,6.934085,5.5570765,4.961002,5.6778007,5.0175915,4.398881,4.4101987,4.776143,3.138824,3.7575345,4.696918,5.2288585,5.828706,6.9869013,6.590776,6.1078796,6.085244,6.1342883,6.0739264,4.8402777,7.17176,11.117926,8.043237,8.07719,8.152642,8.390318,8.526133,7.9036493,6.937857,8.024373,8.612903,8.065872,7.673519,8.296002,9.34102,10.099318,10.054046,8.880759,9.175024,9.25425,9.42779,9.933322,10.970794,11.763044,11.570641,11.314102,11.378237,11.59705,9.839006,8.601585,7.6207023,7.1038527,7.752744,7.677292,7.001992,6.4134626,6.2361493,6.40969,6.4210076,6.8359966,7.5188417,8.160188,8.269594,8.477088,8.473316,8.329956,8.201687,8.360137,9.397609,11.627231,12.513797,11.69891,11.000975,11.099063,11.672502,11.921495,12.038446,13.200415,12.649611,19.138527,22.137764,19.606333,18.006739,24.39002,32.787884,29.645287,16.471281,9.857869,8.345046,8.816625,10.465261,12.14408,12.37421,15.158407,16.659912,13.445636,9.9257765,18.372684,18.516043,18.040693,23.322369,32.72752,36.63596,31.972998,30.716713,26.019794,17.716248,12.283667,12.147853,9.205205,6.3417826,4.7648253,3.983892,6.168242,6.907676,7.009537,7.1378064,7.798016,7.6395655,7.854605,7.5188417,6.752999,6.730363,7.194396,7.960239,8.360137,8.428044,8.880759,8.854351,8.639311,8.122461,7.605612,7.8131065,7.7640624,7.001992,6.549277,6.4926877,5.96452,5.745708,5.3910813,4.7535076,4.4403796,5.783434,7.5527954,8.729855,9.208978,9.261794,9.507015,8.846806,9.367428,10.069136,10.374719,10.11818,9.21275,9.7296,10.103089,9.940866,10.038955,10.589758,9.49947,8.390318,7.9413757,7.9036493,8.209232,8.643084,8.922258,8.76758,7.888559,9.024119,9.876732,10.401127,10.7557535,11.291467,10.144588,10.076681,10.393582,10.593531,10.359629,10.227587,10.585986,10.774617,10.70671,10.86516,11.219787,11.827179,11.98563,11.574413,11.0613365,12.185578,12.932558,13.008011,12.419481,11.491416,10.269085,10.11818,10.212496,10.133271,9.903141,10.023865,9.827688,9.442881,8.914713,8.194141,7.937603,7.7716074,7.4999785,7.0812173,6.651138,6.541732,7.4207535,7.8508325,7.3075747,6.2097406,6.0022464,6.537959,7.3075747,7.7376537,7.1868505,7.432071,7.254758,7.1868505,7.54525,8.424272,8.937348,9.239159,9.488152,9.563604,9.065618,8.624221,9.393836,10.627484,11.627231,11.747954,11.480098,10.910432,10.435081,10.159679,9.903141,9.49947,9.929549,10.529396,10.842525,10.63503,10.084227,10.186088,10.419991,10.450171,10.133271,13.936077,13.536179,12.494934,11.876224,11.921495,12.083718,12.117672,11.472552,11.148107,11.219787,10.819888,9.58624,9.0807085,9.0807085,9.420244,9.97482,10.695392,10.77839,10.733118,10.676529,10.336992,10.661438,10.4049,9.846551,9.371201,9.469289,9.673011,9.899368,9.982366,10.167224,11.091517,12.3893,12.600568,12.510024,12.434572,12.208215,12.23085,11.574413,11.148107,11.012292,10.3634,9.552286,9.129752,8.858124,8.544995,8.088508,8.111144,8.375228,8.926031,9.420244,9.110889,9.476834,9.559832,9.488152,9.386291,9.367428,9.4013815,8.941121,8.605357,8.7600355,9.510788,9.81637,10.001229,9.699419,9.144843,9.129752,8.186596,7.9262853,8.827943,10.612394,12.261031,18.991394,18.312323,12.049765,4.346064,1.6825907,1.2034674,0.7884786,0.5017591,0.3734899,0.39989826,0.11317875,0.02263575,0.0150905,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.06790725,0.094315626,0.08677038,0.150905,0.14713238,0.150905,0.1961765,0.2678564,0.2867195,0.20749438,0.124496624,0.0754525,0.0452715,0.07922512,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.07922512,0.211267,0.271629,0.26031113,0.3169005,0.8941121,0.91674787,0.88279426,1.0072908,1.237421,1.2223305,1.116697,1.146878,1.2600567,1.1242423,1.4600059,1.6561824,1.9655377,2.2560298,1.9957186,1.9466745,2.7426984,3.199186,3.0331905,2.8936033,3.8782585,4.0178456,3.572676,3.138824,3.6481283,4.1762958,3.832987,3.5349495,3.6858547,4.164978,6.2097406,6.466279,6.571913,6.9944468,7.009537,7.0057645,7.149124,7.2396674,7.2283497,7.2283497,7.277394,7.020855,7.3453007,7.967784,7.4396167,7.5829763,8.650629,9.424017,9.5032425,9.318384,9.514561,9.929549,10.238904,10.38981,10.627484,10.725573,11.038701,10.914205,10.49167,10.691619,11.1782875,11.461235,11.5857315,11.604594,11.581959,10.808571,10.763299,10.831206,10.748209,10.608622,10.20495,9.944639,9.850324,9.989911,10.47658,10.47658,10.93684,11.261286,11.227332,11.004747,11.249968,11.268831,11.106608,10.933067,11.068882,11.517824,11.449917,11.415963,11.604594,11.830952,12.770335,14.139798,15.596032,16.784409,17.338985,18.350048,18.346275,17.912424,17.557796,17.70493,18.787672,19.787418,19.960958,19.56106,19.840235,20.832436,22.062311,23.318596,24.152346,23.895807,23.892035,23.431774,23.205416,22.771564,20.53817,20.534397,19.270569,18.738628,19.312067,19.749691,21.043703,21.571869,20.832436,19.312067,18.489635,17.471025,17.335213,16.999449,16.41092,16.535416,16.316603,15.301767,13.7700815,11.887542,9.699419,8.544995,8.028146,8.318638,9.186342,10.012547,10.631257,10.642575,10.638803,10.650121,10.152134,10.242677,9.918231,9.42779,9.178797,9.7220545,9.922004,10.284176,10.751981,11.359374,12.238396,18.033148,15.829934,10.167224,6.145606,9.4127,4.7308717,2.916239,2.5238862,2.8747404,4.0480266,6.356873,5.73439,5.945657,6.9680386,5.0213637,3.4368613,1.8485862,2.6823363,4.7044635,3.0105548,5.2854476,4.908185,4.7912335,5.926794,7.4018903,9.782416,11.45369,11.796998,10.884023,9.473062,10.567122,10.812344,11.68382,12.992921,12.894833,12.015811,10.687846,9.14107,7.677292,6.6850915,5.7683434,5.764571,6.2851934,6.8359966,6.8058157,6.937857,6.858632,6.7454534,6.6850915,6.643593,6.9793563,7.122716,7.0585814,6.8397694,6.598321,6.5266414,6.477597,6.590776,6.900131,7.3490734,7.3453007,7.7942433,7.91874,7.5565677,7.175533,7.5301595,7.220804,7.01331,7.254758,7.8810134,9.042982,8.262049,7.6093845,7.4094353,6.2361493,6.168242,6.368191,6.428553,6.4247804,6.937857,8.099826,8.729855,8.511042,7.8131065,7.6886096,7.149124,7.2170315,7.322665,7.0887623,6.3153744,5.907931,5.8437963,6.0248823,6.5002327,7.466025,8.111144,8.616675,9.480607,10.616167,11.321648,12.189351,13.324911,14.0907545,14.011529,12.770335,12.196897,12.004493,12.00072,11.959221,11.61214,11.740409,12.268577,13.117417,13.905896,13.917213,12.619431,11.947904,11.634775,11.219787,10.038955,10.834979,11.144334,10.193633,8.409182,7.394345,6.9755836,7.322665,7.364164,6.9793563,7.009537,7.1679873,7.183078,7.6886096,8.60913,9.163706,9.650374,8.75249,7.7602897,7.0170827,5.8890676,6.6549106,8.397863,9.465516,9.578695,9.805053,10.091772,9.831461,9.310839,8.654402,7.854605,7.8508325,8.122461,8.903395,9.552286,8.533678,8.314865,7.858378,7.8319697,8.284684,8.627994,9.220296,8.201687,7.0849895,6.8661776,8.043237,7.745199,7.383027,7.0246277,6.903904,7.432071,7.677292,7.726336,7.3075747,6.221059,4.323428,4.9459114,5.0213637,4.564876,3.893349,3.6028569,3.561358,4.6252384,5.458988,5.59103,5.4401255,5.847569,6.2851934,5.983383,5.342037,5.938112,6.198423,7.492433,10.412445,12.691111,9.21275,9.280658,8.254503,7.7112455,8.167733,9.088254,7.1868505,6.820906,7.5075235,8.526133,8.944894,8.367682,8.737399,9.507015,10.020092,9.491924,9.092027,9.374973,9.793735,10.178542,10.740664,11.736636,11.672502,11.249968,10.989656,11.219787,10.016319,9.110889,8.356364,7.858378,7.960239,7.964011,7.6131573,7.149124,6.6813188,6.175787,6.3455553,6.579458,7.1906233,7.858378,7.635793,7.598067,8.031919,8.167733,7.960239,8.080963,8.60913,9.986138,10.789707,10.653893,10.280403,9.635284,9.49947,9.782416,10.544487,11.966766,11.476325,11.778135,13.226823,14.637785,13.29473,17.297485,24.491882,25.695349,19.836462,13.920986,9.733373,8.394091,8.446907,8.722309,8.360137,10.008774,10.672756,10.0276375,12.649611,28.000423,27.574116,19.768555,18.414183,26.574371,36.5756,41.10275,35.402313,27.155355,20.485353,15.9695215,11.578186,8.20546,6.300284,5.624984,5.2628117,5.975838,6.7680893,7.122716,6.964266,6.6850915,6.9869013,7.356619,7.394345,6.964266,6.1795597,6.907676,7.3075747,7.303802,7.1076255,7.2094865,7.6508837,8.446907,8.590267,8.062099,7.8017883,8.141325,7.647111,7.284939,7.0849895,6.1116524,5.4740787,5.3986263,5.251494,5.1458607,5.9418845,7.0170827,7.911195,8.439363,8.646856,8.7751255,8.624221,9.088254,9.4127,9.420244,9.507015,8.884532,9.318384,9.842778,10.137043,10.529396,10.393582,8.9788475,7.6018395,7.0812173,7.756517,7.575431,8.084735,8.959985,9.408927,8.167733,8.631766,9.416472,9.993684,10.336992,10.914205,9.6201935,9.118435,9.250477,9.839006,10.691619,10.759526,10.827434,10.585986,10.314357,10.86516,11.363147,11.7555,11.876224,11.781908,11.759273,12.577931,12.766563,12.570387,12.030901,10.963248,9.469289,9.092027,8.975075,8.793989,8.76758,9.397609,9.544742,9.303293,8.801534,8.216777,8.235641,8.080963,7.677292,7.1076255,6.6058664,6.964266,7.564113,7.5263867,6.7831798,6.0776987,5.4476705,6.096562,7.2585306,7.877241,6.6247296,5.9909286,5.8928404,6.4134626,7.454707,8.75249,9.148616,9.216523,9.099571,8.956212,8.952439,9.510788,9.805053,10.1294985,10.585986,11.076427,10.661438,10.246449,9.6201935,9.156161,9.81637,10.536942,11.212241,11.566868,11.427281,10.733118,9.695646,9.242931,9.039209,8.975075,9.156161,14.618922,14.211478,13.890805,13.751218,13.573905,12.83447,11.514051,10.665211,10.212496,10.0465,10.054046,9.782416,9.9257765,10.1294985,10.054046,9.397609,9.363655,9.567377,9.759781,9.857869,9.899368,10.291721,9.955957,9.393836,9.129752,9.684328,9.042982,8.918486,8.959985,9.231613,10.186088,11.4838705,11.661184,11.895086,12.23085,11.608367,11.185833,10.631257,10.502988,10.589758,9.963503,9.476834,9.473062,9.190115,8.605357,8.416726,8.412953,8.963757,9.839006,10.480352,10.016319,9.835234,9.673011,9.574923,9.522105,9.435335,9.876732,9.733373,9.57115,9.691874,10.110635,10.0465,9.774872,9.771099,10.091772,10.382264,8.6581745,9.144843,9.767326,11.050018,16.143063,23.205416,19.017803,10.197406,2.5917933,1.237421,0.9393836,0.6111652,0.3734899,0.24899325,0.15845025,0.041498873,0.003772625,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.120724,0.23013012,0.06790725,0.0754525,0.116951376,0.14713238,0.1659955,0.211267,0.20749438,0.14335975,0.094315626,0.07922512,0.056589376,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.29426476,0.5357128,0.5998474,0.4640329,1.0035182,1.1053791,1.1732863,1.3505998,1.5128226,0.97333723,1.20724,1.3015556,1.0940613,1.146878,1.2562841,1.4977322,1.841041,2.0485353,1.6788181,1.6222287,1.8599042,2.1503963,2.2183034,1.7467253,2.8709676,3.1765501,3.2670932,3.3123648,3.0558262,3.6443558,4.183841,4.2630663,4.074435,4.4139714,5.541986,6.5040054,7.2396674,7.4584794,6.63982,6.802043,7.001992,7.2283497,7.375482,7.2283497,6.647365,6.7114997,7.3717093,8.039464,7.6093845,8.416726,9.118435,9.408927,9.348565,9.363655,9.359882,9.540969,9.405154,9.314611,10.469034,10.834979,10.853842,10.623712,10.321902,10.208723,11.02361,11.532914,11.793225,11.812089,11.532914,10.386037,9.963503,10.087999,10.329447,10.005001,9.6051035,9.623966,9.646602,9.669238,10.099318,9.8239155,10.170997,10.702937,11.136789,11.344283,11.774363,11.589504,11.68382,12.091263,12.00072,12.408164,12.453435,12.453435,12.585477,12.89106,13.449409,14.634012,16.275105,17.77661,18.116146,18.157644,17.991648,17.618158,17.14658,16.795727,18.184053,18.8254,19.010258,19.066847,19.36111,20.598532,22.424482,23.348776,23.145054,22.873425,22.432028,22.266033,22.545206,22.797974,21.934042,21.375692,19.08571,17.814335,18.417955,19.828917,21.571869,21.964222,20.821117,19.059301,18.689585,16.422237,15.580941,15.286676,15.230087,15.663939,15.863888,15.109364,13.788944,12.347801,11.302785,10.27663,8.733627,7.9489207,8.303548,9.2995205,10.401127,11.144334,11.374464,11.046246,10.242677,10.005001,9.752235,9.476834,9.488152,10.412445,10.801025,10.804798,10.736891,11.072655,12.457208,16.58446,15.060319,10.18986,6.1305156,8.858124,6.530414,5.372218,4.3347464,3.259548,2.8521044,5.2665844,5.2854476,4.991183,4.979865,4.357382,2.4672968,1.5015048,2.233394,3.712263,3.2821836,5.3986263,5.6363015,6.1833324,7.541477,8.514814,10.555805,11.766817,12.193124,11.902632,10.989656,11.793225,11.725319,12.272349,13.358865,13.373956,12.600568,11.208468,9.563604,8.0206,6.8925858,6.0362,5.772116,6.0362,6.5228686,6.651138,7.0812173,7.273621,7.118943,6.719045,6.3908267,6.9755836,7.4169807,7.4207535,7.020855,6.571913,6.7680893,6.9454026,7.001992,7.0284004,7.2887115,7.3868,7.9262853,8.179051,7.8923316,7.3075747,7.77538,7.8621507,8.047009,8.152642,7.3113475,8.367682,8.412953,8.062099,7.537705,6.6549106,6.3945994,6.515323,6.5756855,6.549277,6.8133607,8.054554,8.858124,8.782671,8.047009,7.5037513,7.432071,7.435844,7.7225633,7.967784,7.3377557,6.417235,5.983383,5.8966126,6.228604,7.254758,7.756517,8.050782,8.827943,10.140816,11.378237,11.815862,12.668475,13.6682205,14.290704,13.7700815,12.966512,12.393073,11.947904,11.548005,11.121698,11.932813,12.377983,12.713746,13.060828,13.389046,12.875969,12.2119875,12.079946,12.204442,11.32542,11.3971,11.868678,10.812344,8.499724,7.383027,7.194396,7.1566696,6.9454026,6.6360474,6.696409,7.5075235,7.6886096,8.194141,8.956212,8.873214,8.933576,8.590267,7.914967,7.01331,6.043745,7.250985,9.329701,10.423763,10.103089,9.363655,9.239159,9.382519,9.1825695,8.631766,8.337502,8.307321,7.997965,8.401636,9.163706,8.597813,8.126234,7.4471617,7.5263867,8.265821,8.495952,8.326183,7.914967,7.6697464,7.9300575,8.9788475,7.9941926,7.484888,7.009537,6.4926877,6.2021956,6.6134114,6.228604,5.836251,5.304311,3.5802212,3.7613072,3.9386206,3.7386713,3.4255435,3.8895764,3.8178966,4.1574326,4.564876,4.9119577,5.304311,5.1345425,6.0248823,6.043745,5.372218,6.2663302,6.579458,7.1566696,9.537196,12.691111,13.011784,12.630749,12.155397,9.563604,6.5266414,8.431817,9.175024,8.458225,7.752744,7.7640624,8.439363,8.503497,8.835487,9.258021,9.5183325,9.303293,9.288202,9.258021,9.695646,10.465261,10.853842,11.472552,11.495189,11.02361,10.47658,10.582213,9.937095,9.201432,8.737399,8.654402,8.809079,8.575176,8.197914,7.8432875,7.488661,6.94163,6.7341356,6.7680893,7.066127,7.3490734,7.0284004,6.8737226,7.5263867,7.967784,8.001738,8.2507305,8.197914,8.695901,9.186342,9.378746,9.26934,8.892077,9.242931,9.574923,9.831461,10.623712,10.521852,8.941121,10.197406,12.853333,9.725827,10.767072,14.0983,15.841252,15.011275,13.528633,12.155397,10.495442,10.005001,10.26154,8.956212,11.634775,10.069136,12.562841,20.560806,28.645542,27.92497,16.218515,10.657665,16.16947,25.46522,27.841972,22.232079,16.490145,13.86817,12.981603,9.7069645,7.756517,5.9682927,4.847823,6.5832305,6.7114997,6.7869525,6.8133607,6.700182,6.2625575,6.48137,6.8133607,7.1679873,7.1793056,6.224831,6.330465,6.752999,7.24344,7.4282985,6.8171334,6.749226,7.435844,8.0206,8.122461,7.8244243,7.8244243,7.5829763,7.3000293,6.990674,6.470052,5.9305663,5.8890676,6.1305156,6.405917,6.458734,6.900131,7.6697464,8.209232,8.507269,9.0957985,8.843033,8.941121,9.148616,9.4013815,9.820143,9.733373,9.914458,10.336992,10.638803,10.1294985,9.107117,7.937603,7.0849895,6.990674,8.050782,7.8395147,8.533678,9.6201935,10.238904,9.208978,8.428044,8.959985,9.854096,10.540714,10.819888,9.684328,8.986393,8.952439,9.522105,10.325675,10.623712,10.642575,10.435081,10.257768,10.597303,11.408418,11.563096,11.691365,12.042219,12.491161,12.393073,12.098808,11.959221,11.732863,10.612394,9.027891,8.416726,8.103599,7.914967,8.171506,8.68081,8.726082,8.231868,7.5603404,7.4999785,7.748972,7.816879,7.6207023,7.273621,7.0849895,7.643338,7.5527954,6.9491754,6.168242,5.7494807,5.0251365,5.3571277,6.0814714,6.436098,5.587258,5.413717,5.9909286,7.0359454,8.182823,9.009028,8.922258,8.820397,8.816625,8.89585,8.944894,9.42779,9.808825,9.88805,9.778644,9.903141,9.665465,9.431562,8.963757,8.586494,9.190115,10.310584,10.93684,11.046246,10.691619,10.005001,9.073163,8.484633,8.469543,8.929804,9.424017,14.641558,14.015302,14.1926155,14.196388,13.577678,12.434572,10.70671,10.065364,9.65792,9.261794,9.265567,9.635284,10.163452,10.453944,10.216269,9.273112,8.677037,8.744945,9.009028,9.291975,9.733373,10.050273,9.710737,9.190115,8.892077,9.159933,8.412953,8.14887,8.288457,8.790216,9.654147,10.514306,10.725573,11.016065,11.2801485,10.582213,10.393582,10.231359,10.212496,10.238904,9.982366,9.597558,9.457971,9.22784,8.933576,8.941121,9.035437,9.420244,10.035183,10.552032,10.370946,9.7069645,9.439108,9.646602,10.065364,10.133271,10.797253,10.574668,10.295494,10.223814,10.042727,9.559832,9.435335,9.748463,10.355856,10.887795,9.359882,10.578441,11.016065,11.710228,18.285913,23.465727,17.689838,8.76758,2.142851,0.87147635,0.59607476,0.3772625,0.23767537,0.13958712,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.0150905,0.0,0.0,0.018863125,0.02263575,0.11317875,0.211267,0.049044125,0.030181,0.10186087,0.16222288,0.16976812,0.150905,0.13204187,0.08299775,0.056589376,0.056589376,0.0452715,0.00754525,0.0150905,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24899325,0.4979865,0.6073926,0.5357128,0.935611,0.94315624,1.0789708,1.4071891,1.5505489,0.91674787,1.1091517,1.1808317,0.9922004,1.2034674,1.327964,1.4260522,1.5618668,1.6410918,1.4222796,1.5807298,1.3996439,1.569412,1.991946,1.7580433,2.2598023,2.6446102,2.938875,3.0181,2.6144292,3.2972744,4.0895257,4.274384,4.0404816,4.496969,4.666737,5.59103,6.2927384,6.2889657,5.572167,6.3342376,6.439871,6.537959,6.858632,7.201941,6.598321,6.9152217,7.4999785,7.9338303,8.028146,9.0957985,9.435335,9.416472,9.35611,9.533423,9.676784,9.733373,9.416472,9.148616,10.069136,10.159679,10.125726,10.076681,10.03141,9.9257765,10.567122,10.963248,11.208468,11.272603,10.997202,10.33322,10.099318,10.050273,10.012547,9.880505,9.442881,9.608876,9.782416,9.81637,10.005001,9.378746,9.390063,9.906913,10.650121,11.208468,12.30253,12.291212,12.50248,13.075918,12.970284,13.060828,12.725064,12.464753,12.566614,13.106099,13.58145,14.724555,16.33924,17.901106,18.561316,17.991648,17.463482,16.859861,16.222288,15.769572,17.312576,17.96524,18.4255,18.68204,17.991648,18.640541,20.010002,20.4514,20.017548,20.455173,21.153109,21.364376,21.541689,22.009495,22.963968,22.084948,19.296976,17.45971,17.591751,18.832945,20.104319,20.209951,19.07062,17.444618,16.920223,15.226315,14.456699,14.068119,13.936077,14.377474,14.539697,14.324657,13.494679,12.336484,11.649866,10.891568,9.167479,7.986647,7.911195,8.567632,9.544742,10.831206,11.555551,11.3971,10.56335,10.03141,9.771099,9.529651,9.491924,10.272858,11.32542,11.710228,11.691365,11.781908,12.762791,16.471281,15.509261,11.09529,6.462507,6.8661776,6.017337,5.3684454,4.8025517,4.146115,3.1576872,3.942393,4.7346444,4.3875628,3.3651814,3.7613072,2.3390274,2.867195,4.1498876,4.8742313,3.6292653,5.7494807,6.670001,7.4735703,8.52236,9.454198,11.442371,12.174261,12.3289385,12.294985,12.204442,12.366665,12.479843,12.928786,13.487134,13.324911,12.868423,11.480098,9.955957,8.646856,7.4735703,6.5002327,6.145606,6.3116016,6.749226,7.0812173,7.567886,7.779153,7.61693,7.2170315,6.952948,7.4773426,7.888559,7.748972,7.1302614,6.651138,7.0284004,7.3490734,7.4509344,7.3490734,7.232122,7.5263867,7.9791017,8.265821,8.182823,7.654656,8.231868,8.884532,9.175024,8.854351,7.865923,8.36391,9.122208,9.114662,8.122461,6.749226,6.730363,6.8058157,6.930312,7.0887623,7.3188925,7.9451485,8.495952,8.567632,8.160188,7.6622014,7.809334,7.8923316,8.299775,8.707218,8.080963,6.828451,6.1418333,5.8098426,5.824933,6.3644185,6.9227667,7.567886,8.420499,9.552286,10.989656,11.408418,12.215759,13.128735,13.8870325,14.252977,14.3095665,13.622949,12.702429,11.936585,11.634775,12.332711,12.47607,12.419481,12.408164,12.559069,13.140053,12.89106,12.857106,13.181552,13.113645,12.902377,12.826925,11.498961,9.288202,8.322411,8.243186,7.745199,7.322665,7.1000805,6.8435416,7.9036493,8.394091,9.073163,9.669238,8.888305,8.160188,8.29223,7.986647,7.0510364,6.4134626,7.960239,10.110635,11.559323,11.649866,10.382264,9.14107,9.058073,9.046755,8.801534,8.812852,8.91094,8.371455,8.367682,8.873214,8.650629,8.028146,7.273621,7.2660756,8.073418,8.967529,7.997965,7.594294,7.533932,7.9413757,9.239159,8.231868,7.496206,6.858632,6.2436943,5.6778007,6.168242,5.149633,4.191386,3.6556737,2.6898816,2.6974268,2.5993385,2.6068838,2.916239,3.6934,3.3689542,3.4670424,3.7235808,4.093298,4.749735,4.779916,6.2625575,6.8133607,6.198423,6.3455553,6.930312,7.141579,8.073418,9.952185,12.121444,15.245177,14.7170105,12.030901,8.816625,6.8397694,8.888305,8.9788475,8.409182,8.024373,8.194141,8.605357,8.933576,9.0543,9.001483,8.967529,9.405154,9.1976595,9.26934,9.839006,10.416218,10.868933,10.789707,10.393582,9.944639,9.733373,9.325929,9.21275,9.061845,8.926031,9.208978,9.065618,8.733627,8.495952,8.311093,7.828197,7.4169807,7.5075235,7.567886,7.4018903,7.149124,6.730363,7.020855,7.4811153,7.8810134,8.345046,8.099826,8.160188,8.088508,7.8734684,7.9262853,7.798016,8.175279,8.586494,8.89585,9.291975,9.786189,8.333729,8.386545,9.563604,7.6320205,8.492179,9.906913,11.114153,11.864905,12.393073,13.143826,12.47607,11.932813,11.732863,10.751981,13.219278,10.33322,13.687083,23.220507,27.223263,19.606333,10.484125,8.397863,13.264549,16.380737,13.045737,10.917976,10.804798,11.981857,12.200669,8.537451,8.190369,6.741681,4.659192,7.2962565,7.220804,6.888813,6.670001,6.63982,6.590776,6.881268,6.9567204,7.2094865,7.364164,6.462507,5.8588867,6.3153744,7.0812173,7.4509344,6.7643166,6.458734,6.7680893,7.3905725,7.9753294,8.118689,8.122461,7.9526935,7.6395655,7.2094865,6.696409,6.0776987,6.0022464,6.579458,7.3113475,7.073672,6.9491754,7.462252,8.065872,8.669493,9.64283,9.065618,9.016574,9.367428,9.87296,10.186088,10.170997,10.121953,10.393582,10.653893,9.884277,8.296002,7.3000293,6.8171334,6.8661776,7.575431,7.4169807,8.209232,9.2995205,10.038955,9.789962,9.0807085,9.193887,9.808825,10.446399,10.495442,9.578695,8.827943,8.590267,8.892077,9.439108,10.023865,10.250222,10.250222,10.257768,10.616167,11.299012,11.370691,11.378237,11.68382,12.479843,11.883769,11.3971,11.34051,11.299012,10.137043,8.744945,8.054554,7.6207023,7.383027,7.6886096,7.816879,7.858378,7.533932,7.0849895,7.281166,7.515069,7.5716586,7.4773426,7.326438,7.3000293,7.7112455,7.220804,6.398372,5.6815734,5.3910813,4.878004,5.6853456,6.375736,6.3945994,6.058836,6.1003346,6.4926877,7.277394,8.141325,8.409182,8.20546,8.258276,8.480861,8.76758,8.956212,9.190115,9.548513,9.771099,9.7220545,9.371201,8.907167,8.733627,8.52236,8.371455,8.809079,9.929549,10.382264,10.378491,10.023865,9.329701,8.688355,8.394091,8.52236,8.929804,9.216523,13.777626,13.094781,13.226823,12.97783,12.136535,11.491416,10.567122,10.095545,9.597558,8.975075,8.492179,9.092027,9.627739,9.81637,9.673011,9.495697,8.941121,8.756263,9.001483,9.556059,10.137043,10.344538,9.880505,9.167479,8.484633,7.956466,7.9036493,8.0206,8.382772,9.001483,9.797507,10.227587,10.461489,10.435081,10.197406,9.891823,10.336992,10.340765,10.159679,10.061591,10.310584,9.442881,8.786444,8.741172,9.076936,8.948667,9.261794,9.420244,9.559832,9.786189,10.163452,9.4013815,9.446653,10.182315,11.076427,11.185833,11.668729,10.702937,9.8239155,9.473062,9.005256,8.827943,9.574923,10.050273,10.178542,10.982111,10.419991,11.8045435,12.276122,12.664702,17.467255,20.29295,14.815099,7.375482,2.0636258,0.70170826,0.3961256,0.21503963,0.14713238,0.13958712,0.10186087,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.030181,0.003772625,0.011317875,0.05281675,0.056589376,0.03772625,0.02263575,0.02263575,0.018863125,0.08677038,0.15467763,0.1659955,0.1056335,0.09808825,0.06413463,0.033953626,0.0150905,0.0,0.003772625,0.030181,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.21503963,0.3470815,0.44894236,0.70170826,0.6073926,0.73566186,1.1053791,1.1808317,0.97710985,0.8337501,0.845068,1.0223814,1.2826926,1.6335466,1.3958713,1.267602,1.3807807,1.327964,1.629774,1.6335466,1.7693611,2.1768045,2.7125173,2.5276587,2.8445592,2.886058,2.6295197,2.7879698,3.5764484,3.663219,3.5387223,3.62172,4.2328854,4.0895257,4.38379,4.4177437,4.1762958,4.353609,5.6098933,5.666483,5.66271,6.145606,7.066127,6.903904,7.232122,7.5075235,7.6886096,8.243186,8.993938,9.593785,9.869187,9.880505,9.933322,10.291721,10.393582,10.272858,9.993684,9.627739,9.167479,9.061845,9.0807085,9.167479,9.42779,9.774872,10.050273,10.197406,10.197406,10.072908,10.453944,10.910432,10.559577,9.748463,10.050273,9.669238,9.627739,9.725827,9.835234,9.922004,8.971302,8.729855,9.273112,10.201178,10.665211,12.351574,12.898605,13.170234,13.43809,13.373956,13.057055,12.245941,11.695138,11.781908,12.528888,13.36641,14.637785,16.06761,17.384256,18.316093,17.761518,16.720274,15.788436,15.354584,15.588487,17.37671,18.45568,19.232841,19.342249,17.64834,16.950403,16.87118,16.874952,16.984358,17.753973,20.070366,20.692848,20.662666,21.043703,22.930016,21.964222,19.40261,17.591751,17.395575,18.221779,18.485863,18.13878,17.286167,16.135517,14.984866,14.901869,14.947141,14.535924,13.932304,14.245432,13.788944,14.015302,13.743673,12.615658,11.099063,10.499215,9.337247,8.601585,8.544995,8.6581745,9.133525,10.284176,11.23865,11.480098,10.846297,9.997457,9.593785,9.307066,9.167479,9.582467,11.068882,12.366665,12.966512,12.90615,12.774108,17.384256,16.818363,12.37421,7.032173,5.4288073,3.832987,3.0822346,3.5123138,4.4630156,4.315883,3.6556737,4.485651,3.9725742,2.4107075,3.2331395,2.9766011,4.8553686,6.673774,6.7869525,4.0706625,5.9418845,7.4773426,8.446907,9.125979,10.291721,12.076173,12.325166,12.196897,12.385528,13.102326,12.506252,13.132507,13.766309,13.800262,13.249459,12.872196,11.59705,10.378491,9.457971,8.3525915,7.0887623,6.7869525,7.0170827,7.432071,7.786698,8.099826,8.0206,7.8508325,7.7904706,7.960239,8.213005,8.307321,7.9338303,7.2962565,7.115171,7.643338,8.009283,8.224322,8.179051,7.6508837,7.888559,8.062099,8.269594,8.431817,8.288457,8.971302,9.906913,9.597558,8.52236,9.133525,9.137298,10.201178,10.759526,9.808825,6.911449,6.8925858,6.8699503,6.971811,7.254758,7.7150183,7.696155,7.8696957,8.013056,8.054554,8.043237,8.013056,8.333729,8.782671,8.963757,8.299775,7.0887623,6.3116016,5.832478,5.5457587,5.372218,5.934339,7.1679873,8.29223,9.175024,10.303039,10.95193,11.91395,12.630749,13.13628,14.04171,15.399856,15.060319,14.030393,13.192869,13.317367,13.45318,12.955194,12.491161,12.310076,12.2270775,13.456953,13.528633,13.230596,13.151371,13.6833105,14.196388,13.505998,11.925267,10.20495,9.525878,9.390063,8.914713,8.631766,8.409182,7.435844,8.043237,8.695901,9.540969,10.091772,9.220296,8.035691,8.299775,8.216777,7.4169807,6.9755836,8.420499,10.484125,12.347801,13.087236,11.7026825,9.654147,9.005256,8.89585,8.907167,9.0543,9.457971,9.246704,9.046755,8.89585,8.228095,7.911195,7.575431,7.4811153,8.00551,9.646602,8.578949,7.84706,7.250985,7.2094865,8.778898,8.5563135,7.7150183,6.862405,6.224831,5.6476197,5.9532022,4.8025517,3.4594972,2.5578396,2.1013522,2.1541688,1.6788181,1.7580433,2.4408884,2.7389257,2.5238862,3.0671442,3.4594972,3.5575855,3.9989824,4.779916,6.6549106,7.635793,7.2472124,6.541732,7.0887623,8.039464,7.7640624,6.6134114,6.911449,15.237633,15.049001,14.264296,13.555041,6.330465,6.8699503,8.167733,9.26934,9.623966,9.103344,8.914713,8.865668,8.835487,8.737399,8.529905,9.178797,9.1825695,8.8618965,8.714764,9.450426,10.005001,9.861642,9.737145,9.691874,9.137298,8.635539,9.310839,9.4013815,8.793989,9.024119,9.235386,9.110889,9.005256,8.892077,8.379,8.171506,8.507269,8.465771,7.937603,7.624475,7.043491,6.7114997,6.8774953,7.4811153,8.122461,8.047009,8.047009,7.3415284,6.3342376,6.598321,6.5455046,6.3342376,6.9227667,8.080963,8.409182,8.820397,7.7904706,6.0248823,4.90064,6.462507,9.001483,11.159425,12.294985,12.336484,11.785681,12.359119,13.355092,13.155144,12.102581,12.494934,12.97783,10.238904,11.574413,17.603067,22.269806,8.062099,6.2323766,12.0233555,17.70493,12.54775,7.0963078,11.272603,17.278622,19.810055,16.06761,9.899368,9.544742,8.246958,5.560849,7.352846,7.281166,7.1378064,6.9454026,6.8850408,7.2962565,7.8998766,7.6923823,7.586749,7.598067,6.8473144,5.9532022,6.2323766,6.6813188,6.7831798,6.5228686,6.7152724,6.8737226,7.281166,7.9451485,8.578949,8.933576,8.7600355,8.375228,7.809334,6.8133607,5.8664317,5.794752,6.5455046,7.496206,7.4773426,6.983129,7.17176,7.854605,8.790216,9.695646,8.963757,9.22784,9.948412,10.529396,10.344538,10.012547,9.842778,9.857869,9.922004,9.740918,8.318638,7.2962565,6.7039547,6.466279,6.3644185,6.2625575,7.115171,8.171506,9.024119,9.639057,10.178542,9.937095,9.740918,9.831461,9.842778,9.107117,8.499724,8.231868,8.3525915,8.733627,9.525878,10.016319,10.201178,10.329447,10.917976,11.219787,11.52537,11.351829,11.000975,11.551778,11.212241,10.77839,10.589758,10.401127,9.382519,8.382772,7.8206515,7.3490734,6.9755836,7.0510364,6.911449,7.1906233,7.5603404,7.77538,7.6886096,7.707473,7.488661,7.2887115,7.183078,7.069899,7.0548086,6.5002327,5.824933,5.3156285,5.13077,5.221313,6.9982195,8.028146,7.7829256,7.647111,7.277394,6.8133607,6.858632,7.3113475,7.375482,7.567886,7.997965,8.386545,8.692128,9.0957985,9.239159,9.159933,9.495697,10.035183,9.703192,8.843033,8.412953,8.329956,8.5563135,9.088254,9.839006,10.080454,10.0465,9.7069645,8.744945,8.612903,8.741172,8.8618965,8.827943,8.620448,11.261286,11.419736,11.77059,11.5857315,11.140562,11.6875925,11.359374,10.910432,10.11818,9.152389,8.590267,9.2995205,9.895596,10.061591,9.827688,9.582467,9.337247,9.386291,9.820143,10.453944,10.834979,10.699164,9.842778,8.967529,8.492179,8.529905,7.9791017,8.518587,8.899622,8.869441,9.186342,10.016319,9.940866,9.793735,9.831461,9.718282,9.756008,9.325929,9.333474,9.87296,10.238904,8.918486,8.443134,8.677037,9.205205,9.337247,9.533423,10.095545,10.291721,10.295494,11.200924,10.819888,11.348056,12.064855,12.393073,11.917723,11.955449,10.076681,8.477088,8.054554,8.409182,9.567377,10.552032,10.985884,11.140562,11.947904,11.23865,11.895086,12.287439,12.46098,14.143571,15.977067,11.216014,5.4665337,1.7769064,0.6413463,0.27540162,0.10940613,0.10940613,0.23767537,0.45648763,0.116951376,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.071679875,0.030181,0.0,0.0,0.0,0.011317875,0.05281675,0.120724,0.150905,0.030181,0.1056335,0.06790725,0.030181,0.02263575,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026408374,0.26031113,0.6073926,0.7167987,0.5696664,0.663982,0.76584285,0.76584285,0.65643674,0.76584285,0.91297525,1.0148361,1.1091517,1.3430545,1.4901869,1.5165952,1.5241405,1.50905,1.388326,1.388326,1.6448646,1.7354075,1.7354075,2.2107582,2.2107582,2.5616124,2.8785129,3.2029586,3.983892,4.1272516,3.7462165,3.6669915,4.0480266,4.3800178,3.6707642,3.8593953,3.8669407,3.5236318,3.5689032,4.7308717,5.20245,5.8437963,6.677546,6.8963585,6.273875,7.043491,7.6848373,7.7904706,8.073418,8.254503,9.0957985,10.152134,10.789707,10.178542,10.005001,10.103089,10.265312,10.34831,10.238904,9.703192,8.714764,7.884786,7.484888,7.462252,8.669493,9.767326,9.982366,9.476834,9.352338,10.038955,10.948157,10.710483,9.548513,9.291975,9.488152,9.665465,9.65792,9.703192,10.419991,9.529651,9.25425,9.733373,10.518079,10.544487,12.14408,12.981603,13.407909,13.445636,12.785426,12.276122,11.796998,11.578186,11.747954,12.359119,13.751218,15.271586,16.784409,17.95015,18.218006,17.693611,16.856089,16.644821,17.395575,18.859352,21.153109,22.00195,22.03213,21.700138,21.28515,19.60256,18.301004,18.184053,18.889534,18.889534,20.111864,20.783392,21.23988,21.624687,21.881226,21.58696,19.813826,18.23687,18.150099,20.432537,20.530624,19.47429,18.312323,17.497435,16.874952,17.05981,17.206944,16.784409,16.18456,16.724047,15.516807,15.082954,14.724555,13.7851715,11.672502,10.880251,10.005001,9.582467,9.684328,9.903141,11.0613365,11.608367,11.6875925,11.332966,10.469034,9.307066,8.605357,8.4544525,8.654402,8.729855,9.81637,11.7894535,12.857106,12.687338,12.419481,17.206944,17.421982,12.992921,7.2585306,7.001992,4.878004,3.9914372,3.1010978,2.4597516,3.8141239,4.768598,4.236658,2.9124665,1.8636768,2.546522,2.305074,3.4783602,5.3269467,6.3531003,4.304565,4.8138695,7.3151197,9.431562,10.374719,10.925522,11.106608,10.933067,11.306557,12.332711,13.321139,12.58925,13.577678,14.426518,14.407655,13.932304,13.075918,11.902632,10.944386,10.220041,9.231613,7.888559,7.635793,7.6584287,7.624475,7.673519,8.028146,7.8810134,7.8734684,8.265821,8.926031,8.963757,8.835487,8.646856,8.5563135,8.790216,9.57115,9.948412,10.065364,9.835234,8.956212,8.541223,8.375228,8.307321,8.458225,9.216523,9.703192,10.540714,9.7220545,8.009283,8.926031,8.45068,10.582213,12.687338,12.58925,8.560086,6.6549106,6.270103,6.217286,6.1531515,6.590776,6.590776,6.8925858,7.2585306,7.492433,7.432071,7.5905213,8.186596,8.699674,8.8618965,8.66572,7.726336,6.620957,5.915476,5.7004366,5.613666,5.7381625,6.692637,7.914967,8.948667,9.461743,10.412445,11.676274,12.706201,13.407909,14.11339,14.566105,14.577423,14.181297,13.819125,14.34352,15.271586,14.147344,12.83447,12.178034,11.993175,12.483616,12.347801,12.079946,11.891314,11.717773,13.158916,12.687338,11.234878,9.748463,9.186342,8.941121,9.446653,9.820143,9.4013815,7.7678347,7.5716586,7.5792036,7.8017883,8.182823,8.560086,8.695901,9.303293,9.26934,8.4544525,7.7225633,8.197914,10.174769,11.619685,11.691365,10.725573,9.031664,8.578949,8.375228,8.235641,8.7751255,9.812597,9.714509,9.239159,8.52236,7.0812173,7.9941926,8.763808,8.7751255,8.280911,8.379,8.314865,8.394091,8.209232,7.997965,8.620448,9.024119,8.82417,8.073418,6.8699503,5.3571277,4.67051,4.346064,4.1272516,3.712263,2.746471,2.3314822,1.6863633,1.6750455,2.2409391,2.4107075,2.4484336,2.886058,3.1048703,3.2444575,4.195159,5.2099953,6.0286546,6.6850915,7.3490734,8.360137,6.983129,7.7187905,8.590267,8.145098,5.4476705,11.721546,16.51278,16.452417,12.521342,10.054046,8.201687,9.556059,10.86516,10.982111,10.910432,10.005001,9.012801,8.7600355,8.809079,7.432071,8.431817,8.918486,9.012801,8.914713,8.926031,9.144843,9.567377,10.020092,10.197406,9.673011,9.076936,9.510788,9.574923,9.073163,9.046755,9.133525,9.144843,9.171251,9.088254,8.575176,8.710991,9.061845,8.880759,8.024373,6.9869013,7.111398,6.903904,6.7680893,6.964266,7.598067,7.5490227,7.3075747,6.258785,5.1345425,6.013564,6.571913,6.541732,7.5226145,9.0807085,8.729855,6.72659,5.292993,4.2291126,3.8141239,4.7912335,5.6589375,8.035691,9.854096,10.442626,10.529396,11.589504,13.815352,14.7170105,14.317112,15.120681,14.158662,11.857361,9.933322,8.073418,3.92353,4.142342,7.6923823,13.973803,17.384256,7.326438,9.899368,23.186554,33.512226,33.206646,20.583443,15.47908,11.570641,8.329956,6.33801,7.277394,7.6093845,7.7187905,7.5603404,7.3453007,7.5527954,8.175279,8.122461,8.054554,8.069645,7.6886096,7.115171,6.964266,6.858632,6.571913,5.9984736,7.069899,7.4396167,7.865923,8.480861,8.7751255,8.748717,8.854351,8.601585,7.937603,7.2170315,6.228604,6.273875,6.72659,7.145352,7.2924843,6.8774953,7.1302614,7.7301087,8.341274,8.620448,8.329956,9.325929,10.552032,11.189606,10.650121,10.442626,10.253995,9.601331,8.714764,8.544995,8.326183,7.4471617,6.620957,6.1078796,5.7079816,5.87775,7.0548086,8.171506,8.858124,9.446653,10.238904,10.11818,9.6051035,9.159933,9.171251,8.669493,8.552541,8.926031,9.465516,9.431562,10.016319,10.465261,10.695392,10.782163,10.940613,11.5857315,12.600568,12.510024,11.246195,10.148361,10.453944,9.997457,9.276885,8.650629,8.329956,7.6848373,7.3868,6.934085,6.3417826,6.1342883,6.221059,6.72659,7.7150183,8.518587,7.7376537,7.6395655,7.2660756,6.9982195,6.9227667,6.851087,6.326692,5.4174895,4.847823,4.8365054,5.081726,6.3153744,7.786698,8.216777,7.6848373,7.598067,7.0246277,6.8435416,6.9680386,7.254758,7.5226145,8.194141,8.793989,9.250477,9.533423,9.64283,9.64283,8.756263,8.60913,9.461743,10.193633,9.937095,8.726082,8.416726,9.295748,10.103089,9.808825,9.808825,9.6201935,8.903395,7.4773426,8.514814,8.601585,8.9788475,9.684328,9.537196,8.892077,8.8769865,9.307066,9.922004,10.457717,10.676529,10.246449,9.64283,9.024119,8.537451,8.296002,8.333729,8.431817,8.507269,8.582722,8.790216,9.288202,9.578695,10.080454,10.816116,11.419736,10.710483,10.023865,9.239159,8.507269,8.262049,8.443134,8.360137,8.416726,8.75249,9.246704,9.733373,9.601331,9.661693,9.982366,9.903141,9.58624,9.186342,9.110889,9.250477,8.993938,8.76758,9.231613,9.529651,9.469289,9.544742,9.684328,9.952185,10.020092,10.065364,10.774617,12.377983,12.777881,13.287186,13.6833105,12.223305,11.370691,10.295494,9.831461,10.0465,10.26154,10.427535,10.906659,10.963248,11.378237,14.449154,13.340002,13.494679,13.562587,14.211478,18.112373,18.489635,11.431054,4.538468,1.1921495,0.55457586,0.3734899,0.17731337,0.06790725,0.0754525,0.12826926,0.15845025,0.10940613,0.071679875,0.06413463,0.03772625,0.0754525,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.00754525,0.02263575,0.09808825,0.24522063,0.060362,0.116951376,0.150905,0.08677038,0.041498873,0.056589376,0.08677038,0.094315626,0.06790725,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041498873,0.13204187,0.32821837,0.7432071,0.6526641,0.76584285,0.95447415,1.0450171,0.8262049,1.0148361,1.4147344,1.3543724,0.935611,1.0487897,1.841041,2.233394,1.9768555,1.5505489,2.1692593,1.6222287,1.7731338,1.9504471,2.142851,2.969056,3.1727777,2.8181508,2.9011486,3.380272,3.1765501,3.6669915,3.893349,4.115934,4.3686996,4.4516973,4.9760923,5.330719,4.8855495,4.142342,4.768598,5.270357,5.5457587,6.006019,6.6134114,6.8737226,6.4738245,7.175533,7.8131065,8.009283,8.194141,8.2507305,8.729855,9.563604,10.352083,10.397354,10.295494,10.61994,10.929295,11.136789,11.495189,11.291467,10.499215,9.593785,8.99771,9.073163,9.450426,9.58624,9.348565,9.012801,9.280658,9.808825,9.918231,10.061591,9.971047,8.669493,8.737399,9.050528,9.623966,10.442626,11.495189,11.3669195,11.551778,11.498961,11.246195,11.385782,11.706455,12.50248,13.253232,13.468271,12.702429,13.04951,12.823153,12.528888,12.619431,13.483362,14.279386,14.675511,15.539442,16.984358,18.376457,18.840488,19.18757,19.723284,20.511763,21.349285,22.179262,21.884998,20.677757,19.300749,19.040438,18.976303,17.757746,17.180534,17.912424,19.512016,20.100546,20.357084,20.764528,21.462463,22.24717,22.141537,21.360603,20.085455,19.074392,19.685556,20.741892,20.575897,19.666695,18.795218,19.059301,19.059301,18.323639,17.89356,18.010511,18.127462,16.878725,16.418465,15.886524,14.947141,13.773854,13.155144,12.2270775,11.763044,11.812089,11.710228,12.743927,12.728837,12.027128,11.000975,10.0276375,9.065618,8.314865,7.7678347,7.5112963,7.752744,8.944894,10.748209,12.121444,12.709973,12.860879,17.342756,15.350811,11.532914,8.43559,6.541732,5.304311,4.3007927,3.0633714,2.305074,3.92353,4.104616,3.7462165,3.380272,3.4142256,4.146115,3.1237335,3.470815,4.0404816,4.3611546,4.644101,5.5193505,7.484888,9.623966,11.140562,11.378237,11.197151,11.812089,12.702429,13.600313,14.494425,13.875714,13.102326,13.015556,13.321139,12.551523,11.1782875,10.929295,10.676529,9.876732,8.597813,7.322665,6.9982195,7.0849895,7.33021,7.7602897,8.145098,8.280911,8.3525915,8.499724,8.827943,8.68081,8.884532,9.344792,9.767326,9.669238,10.401127,11.00852,11.1782875,10.808571,10.020092,9.058073,8.45068,8.137552,8.235641,9.06939,10.133271,10.974566,10.702937,9.26934,7.4509344,7.492433,8.816625,12.004493,15.924251,17.727566,8.216777,5.9230213,6.2135134,6.5832305,6.651138,6.692637,7.2585306,7.5226145,7.333983,7.2358947,7.326438,7.8395147,8.416726,8.865668,9.178797,8.590267,7.3490734,6.307829,5.8211603,5.7381625,5.9192486,6.696409,7.5905213,8.375228,9.0957985,9.80128,10.733118,11.77059,12.626976,12.845788,12.585477,12.887287,13.29473,13.649357,14.075664,15.128226,15.230087,14.313339,12.683565,11.016065,11.721546,12.291212,12.479843,12.166716,11.351829,11.502733,11.69891,10.997202,9.631512,9.001483,8.809079,9.163706,9.288202,8.884532,8.156415,7.462252,7.4697976,7.4773426,7.484888,8.20546,9.220296,10.223814,10.487898,9.854096,8.771353,8.231868,9.35611,10.201178,10.069136,9.507015,8.60913,7.677292,7.5188417,8.047009,8.262049,9.710737,9.714509,9.457971,9.280658,8.68081,8.597813,8.254503,7.967784,7.865923,7.877241,7.3453007,7.6282477,8.20546,8.703445,8.8769865,8.918486,8.420499,7.4509344,6.326692,5.624984,4.7648253,4.0291634,3.7537618,3.6292653,2.674791,2.9313297,2.2598023,1.9579924,2.4031622,3.0331905,3.1765501,3.308592,3.2972744,3.4330888,4.4177437,4.659192,5.379763,5.783434,6.1116524,7.654656,7.786698,7.466025,8.035691,8.993938,7.9753294,7.696155,9.378746,12.657157,15.961976,16.524097,12.50248,10.7557535,9.910686,9.703192,10.948157,10.940613,9.359882,8.907167,9.646602,8.967529,8.397863,8.771353,9.201432,9.242931,8.914713,8.782671,9.457971,10.106862,10.253995,9.797507,10.223814,10.163452,9.774872,9.4127,9.623966,9.484379,9.688101,9.767326,9.435335,8.601585,8.899622,8.737399,8.345046,7.6923823,6.488915,6.375736,6.571913,6.820906,7.1604424,7.8923316,7.5792036,7.066127,6.330465,5.8437963,6.587003,6.7680893,7.6131573,8.213005,8.243186,7.9451485,4.98741,3.1954134,2.546522,3.6141748,7.598067,4.930821,6.4549613,8.529905,9.861642,11.480098,12.113899,13.381501,13.732355,13.011784,12.46098,12.140307,8.179051,6.3455553,7.6584287,8.3525915,8.552541,8.790216,8.741172,7.707473,4.5912848,15.0376835,26.87618,31.018522,25.329405,14.641558,18.568861,12.762791,7.5263867,6.7379084,7.865923,7.598067,7.5226145,7.1264887,6.7077274,7.394345,7.8017883,7.7376537,7.91874,8.416726,8.654402,8.099826,7.111398,6.730363,7.020855,7.069899,7.394345,7.2962565,7.326438,7.6207023,7.8810134,7.33021,7.7414265,8.062099,8.0206,8.122461,7.6697464,7.745199,7.7301087,7.3415284,6.647365,6.5341864,6.8925858,7.564113,8.246958,8.499724,9.027891,10.250222,11.117926,11.11038,10.26154,10.080454,9.5183325,8.703445,7.8432875,7.201941,7.1793056,7.0057645,7.111398,7.3151197,6.85486,7.0548086,7.4773426,7.828197,8.126234,8.699674,9.661693,10.238904,10.18986,9.635284,9.073163,8.688355,8.654402,9.193887,9.97482,10.114408,10.435081,10.453944,10.231359,10.008774,10.208723,11.529142,12.7477,12.928786,11.966766,10.585986,10.27663,9.616421,8.975075,8.552541,8.394091,7.9489207,7.3868,6.696409,6.096562,6.0362,6.356873,7.0963078,7.6810646,7.8961043,7.907422,7.273621,6.903904,6.7680893,6.6813188,6.326692,5.6363015,4.9119577,4.82896,5.515578,6.571913,8.07719,8.284684,7.6508837,6.8058157,6.5228686,7.0246277,7.466025,7.748972,8.024373,8.68081,9.2844305,9.193887,9.107117,9.190115,9.046755,9.582467,10.250222,10.672756,10.61994,9.986138,9.563604,8.66572,8.228095,8.710991,10.103089,9.242931,8.990166,9.050528,8.8769865,7.6848373,8.047009,8.382772,8.869441,9.235386,8.756263,8.088508,8.733627,8.858124,9.125979,9.480607,9.167479,9.016574,8.541223,7.99042,7.5565677,7.383027,7.2698483,7.069899,7.2585306,7.84706,8.360137,9.016574,9.597558,10.299266,10.963248,11.080199,10.525623,9.590013,8.703445,8.175279,8.201687,8.216777,7.5565677,7.594294,8.514814,9.318384,9.676784,9.371201,9.1976595,9.22784,8.793989,9.265567,9.703192,9.827688,9.582467,9.129752,9.771099,10.574668,11.050018,11.212241,11.61214,11.646093,11.400873,11.208468,11.268831,11.664956,11.910177,11.838497,12.053536,12.117672,10.540714,10.054046,9.782416,9.955957,10.518079,11.148107,10.997202,11.027383,11.487643,12.37421,13.426772,14.022847,15.120681,15.082954,15.720529,22.299986,21.768045,13.132507,4.851596,0.8111144,0.31312788,0.18863125,0.07922512,0.02263575,0.0150905,0.018863125,0.08299775,0.09808825,0.09808825,0.124496624,0.26408374,0.27917424,0.17731337,0.08677038,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.181086,0.2263575,0.20372175,0.08299775,0.08299775,0.08677038,0.056589376,0.0452715,0.060362,0.094315626,0.10186087,0.06790725,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.06413463,0.14335975,0.090543,0.018863125,0.033953626,0.094315626,0.23767537,0.5998474,0.66020936,0.7884786,1.0072908,1.1883769,1.0525624,1.478869,1.9730829,1.8221779,1.1883769,1.0676528,1.6410918,2.335255,2.4522061,2.0862615,2.1353056,1.7957695,1.780679,2.142851,2.686109,2.9464202,3.6368105,2.8181508,2.7238352,3.6669915,4.0291634,4.0103,4.5007415,4.779916,4.851596,5.4401255,5.6476197,6.4738245,6.432326,5.692891,6.0739264,5.8966126,6.168242,6.1644692,6.0324273,6.828451,7.1038527,7.2924843,7.575431,7.8923316,7.9489207,8.318638,8.428044,8.918486,9.786189,10.38981,10.412445,10.876478,11.6008215,12.298758,12.562841,12.140307,10.687846,10.152134,10.718028,10.785934,10.691619,9.978593,9.208978,8.884532,9.416472,10.140816,9.967276,9.559832,9.14107,8.477088,9.805053,10.20495,10.544487,11.204697,12.076173,12.208215,12.642066,12.698656,12.464753,12.796744,12.811834,12.943876,13.468271,14.1058445,14.015302,13.619176,13.943622,14.11339,14.120935,14.807553,14.509516,14.283158,14.7170105,15.954432,17.72002,19.146072,20.179771,21.21347,22.035902,21.817091,19.481836,17.780382,16.33924,15.430037,15.988385,16.776863,16.720274,16.825907,17.565342,18.863125,19.568605,20.153362,20.545715,20.919205,21.688822,21.802,21.62846,21.145563,20.662666,20.802254,21.45869,21.130472,20.243906,19.410156,19.451654,19.33093,18.7839,18.327412,18.12369,18.010511,17.501207,17.316349,16.795727,16.06761,16.075155,14.981093,14.037937,13.36641,13.094781,13.35132,13.958713,13.777626,13.072145,12.034674,10.770844,9.839006,9.405154,8.918486,8.337502,8.122461,9.159933,10.627484,11.98563,13.241914,14.954685,18.689585,16.908905,13.494679,10.370946,7.4773426,4.9685473,4.5422406,4.402653,4.217795,5.0968165,4.4705606,4.7044635,4.5196047,4.3686996,6.4247804,4.4931965,3.8480775,4.164978,4.870459,5.149633,6.760544,8.262049,9.544742,10.487898,10.940613,10.759526,11.608367,12.442118,13.091009,14.264296,14.637785,13.268322,12.525115,12.709973,12.079946,10.853842,10.668983,10.303039,9.397609,8.465771,7.537705,7.1906233,7.2094865,7.3905725,7.533932,7.537705,7.8621507,8.311093,8.76758,9.190115,9.431562,9.635284,9.967276,10.386037,10.61994,11.619685,12.347801,12.513797,11.796998,9.87296,8.643084,8.431817,8.631766,8.83926,8.850578,10.423763,10.974566,10.827434,9.880505,7.5829763,6.5832305,6.5341864,8.801534,13.196642,17.987877,13.162688,8.099826,6.138061,7.0284004,6.9227667,7.2660756,7.7829256,7.7829256,7.2396674,6.7944975,6.7114997,6.722818,7.0812173,7.696155,8.137552,8.141325,7.7037,7.0170827,6.2436943,5.5306683,5.7117543,6.5341864,7.5263867,8.333729,8.729855,9.148616,9.861642,10.751981,11.4838705,11.54046,11.363147,11.5857315,12.091263,12.706201,13.174006,13.705947,14.490653,14.70192,13.788944,11.495189,11.16697,11.853588,12.536433,12.593022,11.800771,10.906659,11.129244,11.133017,10.408672,9.276885,8.631766,8.684583,8.888305,8.692128,7.541477,7.6886096,7.537705,7.5829763,8.118689,9.224068,9.748463,10.423763,10.597303,10.099318,9.235386,8.60913,9.590013,10.416218,10.193633,8.880759,8.726082,8.111144,8.152642,8.76758,8.68081,9.544742,9.665465,9.563604,9.631512,10.148361,9.118435,7.9300575,7.2660756,7.364164,8.016829,7.6622014,7.8319697,8.047009,8.141325,8.246958,8.175279,8.080963,7.1981683,5.73439,4.878004,5.1232247,4.847823,4.7308717,4.5837393,3.3236825,3.127506,2.655928,2.463524,2.7992878,3.572676,3.1350515,3.0897799,3.1199608,3.240685,3.821669,4.191386,5.4212623,6.047518,6.066381,6.9189944,7.254758,6.802043,6.7756343,7.5112963,8.458225,8.929804,7.865923,8.096053,10.631257,14.683057,12.789199,10.680302,8.68081,7.333983,7.413208,10.408672,11.053791,10.223814,9.14107,9.382519,8.975075,8.748717,8.918486,9.367428,9.669238,9.2844305,9.57115,9.797507,9.81637,10.065364,11.144334,10.967021,10.340765,9.899368,10.121953,9.714509,9.937095,10.235131,10.197406,9.574923,9.201432,8.692128,8.360137,7.9753294,6.7643166,5.885295,6.3531003,6.9982195,7.4169807,7.9941926,7.6584287,7.3075747,7.3905725,7.8810134,8.303548,8.820397,9.7296,9.797507,9.1825695,9.435335,5.168496,4.3724723,3.3538637,2.727608,7.413208,5.3684454,6.5002327,7.914967,8.83926,10.61994,11.189606,11.714001,12.570387,13.098554,11.5857315,10.970794,7.01331,6.368191,9.148616,8.892077,8.379,8.13378,8.379,7.956466,4.327201,20.375948,33.180237,34.549698,24.55979,11.54046,19.364883,12.3893,6.549277,6.9491754,7.8734684,7.2623034,7.4509344,7.009537,6.273875,7.3717093,7.009537,7.1566696,7.5792036,8.050782,8.382772,8.288457,7.277394,6.881268,7.326438,7.5490227,7.383027,7.1264887,7.175533,7.435844,7.3377557,6.677546,7.352846,8.016829,8.3525915,9.061845,8.054554,7.9828744,7.8131065,7.0887623,5.945657,6.466279,6.571913,6.8359966,7.4094353,8.0206,8.8769865,10.33322,11.117926,10.86516,10.106862,9.774872,8.748717,7.9338303,7.5905213,7.322665,7.1793056,7.2283497,7.3377557,7.281166,6.7114997,6.990674,7.284939,7.707473,8.2507305,8.778898,9.582467,10.299266,10.355856,9.763554,9.122208,9.193887,9.74469,10.231359,10.495442,10.751981,10.684074,10.736891,10.31813,9.563604,9.348565,10.499215,11.608367,12.37421,12.438345,11.3820095,10.106862,8.933576,8.265821,8.096053,7.9941926,7.413208,6.952948,6.428553,5.994701,6.1418333,6.9491754,7.3151197,7.149124,6.8246784,7.17176,6.752999,6.6662283,6.5568223,6.2097406,5.564622,4.949684,5.0741806,5.4740787,6.0776987,7.2170315,7.643338,7.484888,7.111398,6.7831798,6.6586833,7.281166,7.805561,8.00551,8.111144,8.816625,9.144843,9.129752,9.046755,9.005256,8.952439,9.665465,10.589758,11.117926,10.948157,10.080454,9.623966,9.386291,8.933576,8.529905,9.129752,8.526133,8.484633,8.737399,8.805306,8.0206,8.443134,8.548768,8.5563135,8.480861,8.130007,7.8998766,8.805306,8.718536,8.59404,8.646856,8.348819,8.397863,8.039464,7.6508837,7.3717093,7.1076255,6.9454026,6.6813188,6.8661776,7.5188417,8.130007,8.83926,9.408927,9.903141,10.26154,10.306811,10.020092,9.103344,8.401636,8.201687,8.231868,8.14887,7.77538,8.065872,9.031664,9.74469,9.9257765,9.42779,8.873214,8.480861,8.043237,9.2844305,10.023865,10.106862,9.767326,9.6051035,10.638803,11.476325,12.068627,12.396846,12.442118,12.170488,11.710228,11.351829,11.185833,11.083972,10.272858,10.054046,10.201178,10.27663,9.661693,9.276885,9.363655,9.827688,10.514306,11.227332,10.718028,10.8576145,12.166716,13.72481,13.177779,14.445381,16.25624,15.950659,15.950659,23.775084,23.084692,14.071891,5.3080835,0.8337501,0.150905,0.0452715,0.00754525,0.0,0.0,0.0,0.0150905,0.0754525,0.32821837,0.7469798,1.1393328,0.83752275,0.44139713,0.20372175,0.13958712,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.181086,0.29426476,0.28294688,0.271629,0.124496624,0.05281675,0.05281675,0.08677038,0.10186087,0.0754525,0.06790725,0.056589376,0.03772625,0.0,0.0,0.026408374,0.026408374,0.0,0.0,0.0,0.03772625,0.1358145,0.21881226,0.09808825,0.116951376,0.06413463,0.071679875,0.20372175,0.45648763,0.7582976,0.86770374,1.0186088,1.2336484,1.3392819,1.871222,2.3428001,2.2107582,1.5769572,1.2147852,1.6976813,2.5238862,2.7917426,2.3880715,1.9730829,1.9164935,2.1466236,2.5238862,2.867195,2.9766011,3.6896272,2.8936033,2.7653341,3.682082,4.217795,4.315883,4.7572803,5.028909,5.2250857,6.058836,5.5759397,6.2927384,6.579458,6.247467,6.549277,6.3945994,6.4210076,6.247467,6.115425,6.9152217,7.284939,7.3717093,7.466025,7.6018395,7.5716586,7.8961043,8.156415,8.567632,9.318384,10.578441,10.419991,10.834979,11.672502,12.479843,12.525115,12.291212,10.846297,10.536942,11.502733,11.668729,11.23865,10.374719,9.64283,9.378746,9.699419,10.250222,10.291721,9.906913,9.465516,9.623966,10.804798,11.170743,11.216014,11.355601,11.947904,12.415709,13.094781,13.671993,14.056801,14.388792,13.845533,13.521088,13.909668,14.894323,15.754482,14.781145,14.950912,15.211224,15.339493,15.916705,15.23386,14.452927,14.203933,14.766054,16.048746,18.319866,19.870417,20.99843,21.307787,19.70442,16.546734,14.856597,13.9888935,13.800262,14.652876,15.343266,16.376965,17.191853,17.686066,18.229324,18.617905,19.372429,20.289177,21.145563,21.688822,22.133991,22.232079,22.096264,22.160398,23.182781,23.797718,23.216734,22.126446,20.990885,20.06282,19.01403,18.71222,18.674494,18.621677,18.470772,18.074646,18.304777,18.119919,17.550251,17.697384,16.22606,15.354584,14.856597,14.705692,15.082954,15.24895,15.23386,14.86037,13.890805,12.027128,11.004747,10.744436,10.582213,10.246449,9.876732,10.446399,11.593277,13.004238,14.7736,17.384256,20.704166,19.436563,16.060064,12.287439,9.0807085,4.6742826,3.802806,4.134797,4.459243,4.6931453,4.7836885,5.372218,5.2628117,5.409944,8.888305,6.8171334,5.6325293,5.613666,6.198423,5.9796104,7.4396167,8.526133,9.325929,9.846551,10.023865,9.982366,11.034928,11.751727,11.989402,12.89106,13.917213,13.479589,13.045737,12.951422,12.385528,11.404645,10.748209,9.842778,8.733627,8.058327,7.432071,7.2170315,7.3000293,7.496206,7.564113,7.5527954,8.080963,8.816625,9.510788,9.993684,10.774617,10.801025,10.63503,10.578441,10.650121,11.434827,12.298758,12.679792,12.0233555,9.805053,8.6581745,8.929804,9.533423,9.725827,9.110889,10.235131,10.7557535,10.861387,10.193633,7.8810134,6.579458,6.156924,7.1340337,10.148361,15.965749,16.516552,11.310329,8.333729,8.7600355,6.930312,6.4964604,7.3000293,7.8810134,7.699928,7.141579,7.122716,6.6549106,6.6586833,7.1604424,7.2887115,7.564113,7.6093845,7.284939,6.5756855,5.5797124,5.715527,6.300284,7.1981683,8.07719,8.386545,8.458225,9.009028,9.597558,9.9257765,9.842778,10.197406,10.299266,10.846297,11.895086,12.864652,12.642066,13.272095,13.917213,13.902123,12.717519,11.495189,11.706455,12.261031,12.427027,11.812089,10.684074,10.944386,11.446144,11.223559,9.525878,8.424272,8.337502,8.756263,8.892077,7.7112455,8.07719,7.8395147,7.914967,8.597813,9.58624,9.933322,10.367173,10.336992,9.7296,8.869441,8.756263,9.789962,10.465261,10.050273,8.605357,8.639311,8.812852,9.084481,9.220296,8.805306,9.061845,9.533423,9.857869,10.03141,10.419991,9.465516,8.269594,7.5490227,7.537705,7.9791017,8.130007,8.345046,8.156415,7.6282477,7.3679366,7.141579,7.462252,7.17176,6.017337,4.644101,5.311856,5.481624,5.6325293,5.5382137,4.2819295,3.6066296,3.2482302,3.1199608,3.2444575,3.7613072,3.0143273,2.7087448,2.7691069,3.1237335,3.7235808,4.293247,5.4740787,6.2927384,6.462507,6.3945994,6.2663302,6.25124,6.1795597,6.2097406,6.8246784,9.092027,8.14887,6.790725,6.9755836,9.835234,10.238904,10.552032,9.5032425,7.254758,5.4174895,7.9300575,10.446399,10.61994,9.016574,9.088254,9.1976595,8.7751255,8.771353,9.386291,10.099318,9.612649,9.363655,9.310839,9.473062,9.940866,11.314102,11.68382,11.223559,10.502988,10.495442,10.0465,10.012547,10.223814,10.416218,10.197406,9.318384,8.601585,8.171506,7.7904706,6.8774953,5.8136153,6.187105,6.7831798,7.1038527,7.364164,7.322665,7.647111,8.2507305,8.986393,9.65792,10.831206,10.929295,10.423763,10.450171,12.800517,5.9418845,10.423763,9.337247,2.3163917,5.5457587,5.3458095,6.537959,7.7640624,8.782671,10.442626,11.3971,11.5857315,12.593022,13.649357,11.627231,10.295494,7.654656,7.4396167,9.348565,9.039209,8.620448,8.4544525,9.661693,10.355856,5.66271,26.857317,40.385952,37.692295,21.884998,7.7338815,14.913187,9.763554,5.8890676,7.073672,7.2924843,7.043491,7.624475,7.201941,6.258785,7.5792036,6.458734,6.779407,7.33021,7.6131573,7.828197,7.9828744,7.4169807,7.405663,7.77538,6.9152217,6.647365,6.5040054,6.760544,7.232122,7.284939,6.8133607,7.805561,8.4544525,8.477088,9.152389,7.8621507,7.696155,7.5829763,6.9189944,5.572167,6.579458,6.515323,6.4134626,6.8359966,7.884786,9.06939,10.159679,10.450171,9.993684,9.601331,9.737145,8.944894,8.280911,8.137552,8.258276,7.8696957,7.835742,7.586749,7.0510364,6.673774,7.066127,7.586749,8.099826,8.582722,9.14107,9.635284,10.374719,10.63503,10.242677,9.578695,9.952185,10.718028,10.785934,10.378491,10.997202,10.661438,10.367173,9.922004,9.386291,9.0957985,9.688101,10.336992,11.140562,11.868678,11.962994,10.665211,9.159933,7.986647,7.3490734,7.0849895,6.6322746,6.307829,6.0248823,5.8890676,6.19465,6.911449,6.8246784,6.428553,6.1644692,6.4021444,6.255012,6.2399216,6.066381,5.666483,5.1798143,5.0968165,5.7872066,6.5040054,6.952948,7.3075747,6.7567716,6.5341864,6.5530496,6.749226,7.0812173,7.24344,7.537705,7.6886096,7.756517,8.126234,8.477088,8.884532,9.042982,8.963757,8.993938,9.288202,9.876732,10.310584,10.378491,10.091772,9.612649,9.469289,9.125979,8.578949,8.397863,8.529905,8.526133,8.526133,8.412953,7.805561,8.058327,8.182823,8.031919,7.7716074,7.865923,7.4697976,8.043237,8.088508,8.031919,8.130007,8.443134,8.548768,8.326183,8.175279,8.084735,7.6207023,7.3113475,7.1604424,7.17176,7.364164,7.7376537,8.518587,8.941121,9.039209,9.012801,9.208978,8.944894,8.473316,8.36391,8.544995,8.307321,8.529905,9.001483,9.540969,9.97482,10.133271,10.065364,9.540969,8.786444,8.160188,8.141325,9.310839,9.57115,9.416472,9.303293,9.665465,10.567122,11.2650585,11.766817,11.857361,11.087745,10.589758,10.355856,9.997457,9.476834,9.110889,8.778898,8.869441,9.193887,9.635284,10.137043,9.608876,9.763554,10.216269,10.695392,11.042474,10.235131,11.0613365,12.845788,14.64533,15.237633,15.154634,16.98813,17.346529,17.25976,22.183035,21.183289,13.328684,5.560849,1.237421,0.150905,0.05281675,0.011317875,0.0,0.0,0.0,0.0,0.06790725,0.6526641,1.6637276,2.474842,1.6335466,0.754525,0.33576363,0.3055826,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.18485862,0.25276586,0.23013012,0.45648763,0.31312788,0.1358145,0.06790725,0.120724,0.15845025,0.071679875,0.018863125,0.0,0.0,0.0,0.033953626,0.120724,0.12826926,0.060362,0.06413463,0.0452715,0.1056335,0.17354076,0.17731337,0.011317875,0.22258487,0.11317875,0.05281675,0.18485862,0.392353,0.87902164,0.9808825,1.0450171,1.2487389,1.6373192,2.0787163,2.474842,2.4220252,1.9202662,1.3468271,2.0183544,2.7351532,2.8030603,2.2786655,1.9278114,2.0560806,2.6710186,2.8143783,2.5767028,3.0860074,3.4179983,3.0822346,3.006782,3.3236825,3.361409,4.2102494,4.564876,4.8063245,5.160951,5.7079816,4.9157305,5.1156793,5.3986263,5.564622,6.126743,6.5455046,6.296511,6.2323766,6.571913,6.8925858,6.9680386,7.405663,7.605612,7.4471617,7.254758,7.111398,7.8621507,8.503497,9.103344,10.77839,10.514306,10.774617,11.23865,11.6008215,11.578186,12.162943,11.581959,11.219787,11.510279,11.925267,11.2650585,10.672756,10.423763,10.412445,10.148361,10.197406,10.627484,10.982111,11.208468,11.642321,11.23865,11.449917,11.3971,11.083972,11.419736,12.261031,13.162688,14.245432,15.230087,15.426264,14.234114,13.902123,14.396337,15.531898,16.957949,16.35433,15.848798,15.731846,16.048746,16.569368,16.173243,14.958458,13.917213,13.592768,14.0983,16.731592,18.606586,19.54597,19.051756,16.301512,15.147089,14.93205,14.913187,14.886778,15.173498,15.222542,16.644821,17.712475,17.946377,18.135008,17.716248,18.16519,19.681786,21.507734,21.941587,22.745155,23.09601,22.990377,23.262005,25.578398,26.381968,26.023567,25.144547,23.892035,21.881226,19.50447,19.21398,19.855326,20.602304,20.975796,19.87796,20.104319,20.145817,19.534653,18.844261,17.30503,16.429781,16.25624,16.52787,16.697638,16.36942,16.55428,16.478827,15.584714,13.539951,12.340257,11.861133,11.91395,12.162943,12.136535,12.174261,12.966512,14.5132885,16.65614,19.089483,22.40562,21.402102,17.897333,13.532406,9.763554,5.142088,3.2482302,2.9954643,3.3161373,3.1350515,4.957229,5.6061206,5.956975,7.250985,11.102836,10.076681,8.952439,8.27714,7.8432875,6.7114997,7.2472124,8.080963,9.039209,9.64283,9.110889,9.295748,10.578441,11.283921,11.170743,11.389555,12.513797,13.494679,13.834216,13.498452,12.940104,12.2270775,11.083972,9.699419,8.382772,7.54525,6.900131,6.8171334,7.043491,7.3981175,7.748972,8.182823,8.899622,9.695646,10.38981,10.838752,11.944131,11.838497,11.25374,10.61994,10.038955,10.0276375,10.887795,11.608367,11.498961,10.212496,9.476834,9.869187,10.325675,10.253995,9.5032425,9.590013,10.340765,10.831206,10.208723,7.673519,7.250985,7.4471617,7.533932,8.695901,14.003984,16.018566,13.472044,11.457462,10.676529,7.424526,5.594803,6.3417826,7.6320205,8.27714,7.9338303,8.262049,7.6848373,7.424526,7.635793,7.4018903,7.4282985,7.24344,6.9265394,6.470052,5.783434,5.847569,5.904158,6.375736,7.17176,7.707473,7.564113,8.080963,8.416726,8.314865,8.122461,9.065618,9.231613,10.087999,11.781908,13.13628,12.381755,12.370438,12.577931,12.868423,13.502225,12.196897,11.778135,11.846043,11.891314,11.2801485,10.672756,11.050018,11.710228,11.736636,10.005001,8.303548,8.152642,8.771353,9.352338,9.088254,8.646856,8.329956,8.322411,8.6581745,9.21275,9.710737,10.140816,10.163452,9.578695,8.345046,8.827943,9.782416,10.050273,9.4127,8.601585,8.420499,9.065618,9.303293,8.831716,8.296002,8.5563135,9.42779,10.121953,10.140816,9.288202,9.156161,8.692128,8.416726,8.348819,7.9753294,8.390318,8.695901,8.420499,7.6395655,6.9944468,6.590776,6.85486,7.118943,6.752999,5.194905,5.4250345,5.692891,6.0211096,6.066381,5.1269975,4.4516973,4.0782075,3.8405323,3.6858547,3.6745367,3.1010978,2.6521554,2.6597006,3.240685,4.2781568,4.8025517,5.2628117,6.013564,6.670001,6.1078796,5.666483,6.0248823,6.398372,6.198423,5.036454,6.9869013,7.9753294,8.269594,7.8319697,6.3229194,6.7077274,10.7218,12.457208,10.193633,6.398372,5.553304,7.888559,9.593785,9.416472,8.66572,8.643084,8.590267,8.793989,9.276885,9.80128,9.333474,8.8769865,9.001483,9.574923,9.793735,10.95193,11.959221,11.91395,11.042474,10.718028,10.3634,9.918231,9.774872,9.948412,10.065364,9.186342,8.428044,7.752744,7.1793056,6.7869525,6.300284,6.2021956,6.3342376,6.48137,6.387054,6.7039547,7.7414265,8.492179,9.050528,10.623712,11.2650585,10.846297,10.457717,11.348056,14.9358225,5.832478,14.649103,14.0983,2.5502944,4.014073,4.6931453,5.926794,7.488661,9.167479,10.759526,12.657157,12.951422,13.43809,13.924759,12.2270775,10.736891,9.688101,8.797762,8.533678,10.140816,10.163452,9.491924,10.084227,11.125471,9.046755,29.143528,42.37035,36.300198,16.078928,4.4139714,8.341274,6.643593,5.8928404,7.254758,6.470052,7.1076255,7.8923316,7.413208,6.4134626,7.786698,6.3908267,6.6850915,7.1302614,7.2472124,7.594294,7.7301087,7.635793,8.058327,8.182823,5.66271,5.5268955,5.5382137,5.956975,6.7077274,7.394345,7.383027,8.571404,8.816625,8.039464,8.209232,7.3868,7.3377557,7.5075235,7.322665,6.187105,7.0472636,6.8359966,6.696409,7.2094865,8.409182,9.691874,9.854096,9.420244,8.907167,8.83926,9.714509,9.714509,9.34102,9.065618,9.310839,8.6581745,8.390318,7.779153,7.01331,7.1906233,7.7037,8.3525915,8.597813,8.60913,9.250477,9.540969,10.359629,11.000975,11.019837,10.223814,10.355856,10.608622,10.095545,9.424017,10.714255,10.427535,9.5032425,9.073163,9.273112,9.239159,9.397609,9.416472,9.57115,10.155907,11.476325,11.283921,10.1294985,8.465771,6.9152217,6.2851934,6.2323766,5.80607,5.511805,5.5985756,6.0626082,6.300284,6.017337,5.8928404,6.0211096,5.938112,5.938112,5.772116,5.4891696,5.292993,5.564622,6.126743,6.692637,7.3000293,7.6131573,6.911449,6.3417826,6.1908774,6.3116016,6.651138,7.284939,6.72659,6.6360474,6.8435416,7.1076255,7.1000805,7.6282477,8.239413,8.631766,8.809079,9.058073,8.631766,8.710991,8.967529,9.2995205,9.842778,9.439108,8.922258,8.612903,8.518587,8.296002,8.926031,8.733627,8.337502,7.9225125,7.2623034,7.0472636,7.496206,7.5829763,7.3490734,7.854605,6.043745,6.519096,7.0849895,7.4697976,7.8206515,8.710991,9.042982,9.333474,9.250477,8.718536,7.9489207,7.435844,7.4018903,7.326438,7.032173,6.651138,7.273621,8.088508,8.590267,8.45068,7.5226145,6.937857,6.971811,7.6207023,8.416726,8.4544525,9.088254,9.529651,9.812597,9.827688,9.337247,9.144843,9.058073,8.661947,8.167733,8.424272,8.152642,8.043237,8.073418,8.296002,8.835487,9.250477,9.6201935,9.661693,9.318384,8.744945,8.83926,9.058073,8.729855,8.171506,8.68081,9.231613,9.635284,10.133271,10.552032,10.284176,10.906659,11.5857315,11.676274,11.336739,11.521597,11.385782,13.008011,13.607859,13.95494,18.387774,16.06761,17.976559,22.50748,25.39354,19.73083,16.286423,11.32542,6.0286546,1.7995421,0.27540162,0.06790725,0.00754525,0.0,0.0,0.0,0.0,0.0452715,0.5998474,1.8033148,3.4632697,2.1956677,0.9808825,0.52062225,0.5885295,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.07922512,0.3961256,0.84884065,0.43007925,0.0452715,0.011317875,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.16976812,0.35085413,0.38858038,0.30935526,0.32067314,0.22258487,0.150905,0.13958712,0.1358145,0.0,0.120724,0.071679875,0.0754525,0.21881226,0.42630664,0.7205714,0.95824677,1.116697,1.3166461,1.8297231,2.1956677,2.4899325,2.5012503,2.1277604,1.358145,1.7957695,2.1466236,2.2560298,2.11267,1.8297231,2.3692086,2.4484336,2.2409391,2.0862615,2.4861598,2.8785129,3.1124156,3.0105548,2.7728794,3.006782,3.7877154,4.5120597,4.6252384,4.304565,4.485651,4.0970707,4.6026025,4.98741,5.0854983,5.5985756,6.1003346,6.417235,6.1418333,5.6589375,6.1342883,6.9152217,7.394345,7.7716074,7.877241,7.1566696,6.790725,7.4773426,8.367682,9.178797,10.193633,11.02361,11.283921,11.106608,10.834979,11.016065,12.528888,12.551523,12.185578,12.170488,12.879742,12.257258,11.219787,11.050018,11.514051,10.880251,10.891568,11.249968,11.857361,12.46098,12.679792,11.970539,11.978085,11.827179,11.3971,11.321648,11.970539,12.800517,13.728582,14.524607,14.815099,14.426518,14.181297,14.724555,15.882751,16.678776,17.176762,16.837225,16.603323,16.716501,16.693865,15.973294,15.015047,13.781399,12.879742,13.551269,15.441354,17.040947,17.87847,17.354074,14.739646,15.350811,16.463736,16.70141,15.943113,15.32063,15.173498,16.15438,17.191853,17.852062,18.342503,17.72002,17.663431,18.402864,19.598787,20.357084,21.296469,22.416937,23.262005,24.125937,26.076384,25.32186,25.834936,26.879953,27.166672,24.872917,22.465982,22.398075,23.103556,24.186298,26.397057,24.74842,23.631723,22.764019,21.896315,20.798481,19.149845,17.82188,17.150352,17.14658,17.501207,16.25624,16.13929,16.052519,15.675257,15.456445,14.04171,12.936331,12.562841,12.81938,13.075918,13.0646,13.215506,14.626467,17.123945,19.270569,22.382984,22.382984,19.191343,13.558814,7.066127,7.0170827,6.115425,5.4740787,5.100589,3.8895764,5.881522,6.8737226,8.375228,10.638803,12.664702,13.837989,13.057055,12.015811,10.484125,6.3342376,6.6624556,7.6508837,8.729855,9.303293,8.744945,9.390063,10.514306,11.125471,11.170743,11.536687,12.951422,13.45318,13.287186,12.879742,12.815607,12.815607,11.910177,10.661438,9.363655,8.058327,6.8473144,6.4549613,6.5643673,6.9189944,7.3075747,8.065872,8.805306,9.556059,10.291721,10.925522,11.864905,11.936585,11.506506,10.891568,10.329447,9.548513,9.831461,10.536942,11.016065,10.589758,10.49167,10.47658,10.250222,9.673011,8.7600355,8.903395,9.537196,10.038955,9.567377,7.066127,7.2962565,7.492433,7.009537,6.9491754,10.148361,12.162943,11.91395,10.469034,9.318384,10.38981,8.805306,7.1076255,6.7944975,7.594294,7.4471617,8.152642,8.073418,7.9526935,8.073418,8.254503,7.6697464,7.0284004,6.296511,5.624984,5.3571277,5.330719,5.0968165,5.1043615,5.462761,5.9494295,6.1078796,6.937857,7.462252,7.466025,7.4773426,8.612903,9.152389,10.604849,12.577931,12.770335,12.162943,12.027128,11.98563,11.966766,12.223305,11.5857315,11.2650585,11.661184,12.181807,11.231105,11.219787,11.261286,11.657412,12.102581,11.6875925,8.514814,7.8508325,8.5563135,9.733373,10.710483,9.623966,8.831716,8.722309,9.261794,9.993684,9.2995205,9.42779,10.246449,10.789707,9.261794,9.714509,10.303039,10.393582,9.835234,8.956212,8.98262,8.52236,7.964011,7.6282477,7.7376537,8.884532,9.6201935,9.6201935,8.82417,7.432071,7.322665,7.541477,8.175279,8.952439,9.231613,8.865668,8.616675,8.209232,7.8017883,7.9941926,7.726336,7.194396,6.6662283,6.1833324,5.523123,6.096562,6.304056,6.4511886,6.3719635,5.43258,5.1269975,4.8402777,4.561104,4.22534,3.7235808,3.2972744,3.4179983,3.4179983,3.4481792,4.485651,4.9119577,4.9119577,5.3910813,6.156924,5.873977,6.25124,5.9984736,6.3531003,7.2094865,7.111398,6.571913,6.670001,7.54525,8.409182,7.5075235,4.749735,10.676529,15.347038,14.211478,8.13378,7.8508325,7.745199,8.216777,8.937348,8.850578,7.4094353,7.726336,8.4544525,8.91094,9.0957985,8.605357,8.729855,9.367428,10.231359,10.880251,11.012292,11.34051,11.419736,11.155652,10.804798,10.20495,9.544742,9.291975,9.480607,9.673011,8.941121,8.409182,7.8131065,7.2887115,7.3868,7.435844,6.730363,6.488915,6.741681,6.3644185,6.5341864,7.3000293,8.458225,10.110635,12.649611,8.975075,10.729345,12.464753,11.921495,10.038955,3.1916409,2.0108092,2.1768045,2.6219745,5.5382137,4.696918,5.0439997,6.138061,7.515069,8.695901,12.2270775,12.943876,13.034419,13.377728,13.536179,13.8870325,12.989148,11.480098,10.446399,11.3971,9.748463,8.009283,7.888559,10.472807,16.233604,15.599804,28.588953,28.517273,13.713491,7.537705,8.869441,7.224577,6.779407,7.6886096,6.1041074,7.3490734,7.8508325,7.066127,6.043745,7.4471617,6.617184,6.647365,6.590776,6.6058664,7.9338303,8.326183,8.231868,8.280911,7.8961043,5.292993,5.111907,4.8930945,5.142088,5.9305663,6.881268,7.6508837,8.458225,8.028146,6.7680893,6.7454534,6.730363,7.115171,7.937603,8.7751255,8.726082,8.27714,7.4018903,7.6282477,8.888305,9.522105,9.718282,9.061845,8.748717,8.91094,8.605357,8.98262,9.261794,9.329701,9.348565,9.748463,8.82417,8.2507305,7.496206,6.907676,7.752744,8.360137,8.375228,8.096053,7.967784,8.590267,9.114662,9.933322,10.850069,11.299012,10.344538,9.393836,8.616675,7.8998766,7.8961043,9.993684,10.212496,9.408927,8.8769865,8.873214,8.590267,9.0543,8.650629,8.058327,7.914967,8.805306,9.880505,10.303039,9.522105,7.9338303,6.8963585,6.9227667,5.9192486,5.028909,4.90064,5.7079816,6.3153744,6.2323766,5.956975,5.7419353,5.583485,5.96452,5.8928404,5.5004873,5.4401255,6.881268,7.3075747,7.1868505,6.907676,6.5455046,5.873977,6.485142,6.8661776,7.111398,7.2358947,7.1868505,5.915476,5.3986263,5.6061206,6.19465,6.5002327,6.609639,6.462507,6.8963585,8.031919,9.276885,8.66572,8.194141,8.126234,8.548768,9.352338,9.439108,9.167479,8.465771,7.84706,8.409182,8.186596,8.141325,8.14887,8.0206,7.5075235,7.360391,7.84706,7.809334,7.3188925,7.6584287,6.72659,7.1906233,7.4773426,7.677292,7.8810134,8.186596,8.684583,8.75249,8.843033,8.91094,8.424272,8.597813,8.130007,7.5527954,7.2283497,7.3490734,7.2962565,7.4169807,7.326438,6.9944468,6.730363,6.7379084,6.8058157,7.201941,7.7678347,7.9413757,8.612903,8.948667,8.98262,8.865668,8.888305,8.533678,8.27714,7.8923316,7.3905725,7.032173,6.900131,6.8737226,7.360391,8.43559,9.812597,10.148361,9.918231,9.348565,8.903395,9.303293,9.129752,8.816625,8.560086,8.654402,9.49947,9.793735,10.661438,11.5857315,12.219532,12.370438,12.543978,12.626976,12.958967,13.20796,12.385528,11.940358,13.528633,14.607604,15.309312,18.470772,16.94286,20.50799,26.223516,27.849518,15.848798,10.49167,6.9189944,4.085753,1.7618159,0.52062225,0.1056335,0.0,0.0,0.0,0.0,0.030181,0.35462674,0.7469798,1.4977322,3.4029078,3.0822346,1.780679,0.79602385,0.43385187,0.026408374,0.06413463,0.13204187,0.10186087,0.018863125,0.08677038,0.018863125,0.0,0.06790725,0.19994913,0.32444575,0.5998474,0.36594462,0.1659955,0.16976812,0.16976812,0.033953626,0.0,0.0,0.0,0.0,0.033953626,0.071679875,0.362172,0.6752999,0.29426476,0.19994913,0.1659955,0.16222288,0.14713238,0.060362,0.20372175,0.09808825,0.0150905,0.13204187,0.52439487,0.70170826,0.83752275,1.0186088,1.2826926,1.599593,1.8787673,2.2371666,2.161714,1.7278622,1.6146835,1.8184053,1.9768555,1.750498,1.4826416,2.1956677,1.8863125,1.9051756,2.4559789,3.2444575,3.500996,3.6971724,3.2520027,3.0407357,3.108643,2.674791,3.5953116,3.953711,3.8895764,3.7801702,4.217795,4.3347464,4.6742826,4.776143,4.5799665,4.429062,4.7233267,4.7044635,4.5799665,4.6026025,5.05909,5.783434,7.0812173,8.179051,8.563859,8.009283,7.7829256,8.303548,8.952439,9.65792,10.925522,11.121698,11.291467,11.5857315,11.815862,11.442371,11.932813,11.77059,11.593277,11.653639,11.8045435,11.502733,11.332966,11.480098,11.68382,11.234878,10.827434,10.868933,12.068627,13.532406,12.766563,12.340257,12.404391,12.513797,12.445889,12.178034,12.958967,13.298503,13.230596,13.124963,13.679539,13.52486,13.743673,14.867915,16.293968,16.275105,16.833452,16.939087,16.927769,17.025856,17.354074,16.935314,16.388283,15.807299,15.418718,15.611122,16.52787,17.297485,18.153872,18.493408,16.890041,17.57666,18.572634,18.595268,17.508753,16.320375,16.622187,17.225805,17.987877,18.636768,18.742401,18.142553,17.4333,17.23335,17.77661,18.915941,19.542198,20.975796,22.711203,24.35984,25.63876,22.63575,21.609596,22.33394,23.654358,23.4695,23.45441,24.914415,26.31406,27.023314,27.287397,26.09902,24.307022,22.60557,21.115381,19.379974,18.614132,18.45568,18.018057,17.120173,16.293968,16.16947,17.04472,17.757746,17.916197,17.874697,16.546734,15.339493,14.762281,14.871688,15.275358,15.271586,15.199906,16.13929,18.063328,19.821371,21.002203,20.979568,19.881733,17.139036,11.4838705,7.911195,6.8171334,6.156924,5.4174895,5.624984,5.621211,5.764571,7.699928,11.170743,14.007756,14.984866,14.596286,14.226569,13.630494,10.948157,8.914713,9.646602,11.068882,11.732863,10.831206,10.091772,9.616421,9.548513,10.038955,11.25374,12.057309,12.276122,12.525115,12.974057,13.392818,13.185325,12.404391,11.495189,10.514306,9.118435,7.726336,7.2057137,6.9869013,6.8850408,7.1000805,7.3490734,8.065872,9.14107,10.253995,10.838752,11.193378,11.204697,10.948157,10.529396,10.084227,9.450426,9.367428,9.623966,9.982366,10.163452,10.963248,11.378237,11.487643,11.02361,9.35611,9.325929,9.5183325,9.205205,8.43559,8.054554,7.756517,6.9189944,6.3832817,6.820906,8.729855,12.66093,11.521597,9.122208,7.484888,6.851087,7.726336,9.039209,9.152389,7.6697464,5.43258,6.4436436,6.79827,7.0585814,7.5075235,8.167733,7.9828744,7.443389,6.6134114,5.7306175,5.2099953,5.1081343,4.889322,4.6818275,4.568649,4.606375,5.402399,6.270103,6.862405,7.254758,7.9413757,8.469543,8.677037,9.601331,10.929295,10.978339,11.159425,11.317875,11.136789,10.902886,11.491416,10.846297,10.220041,10.3634,11.038701,11.02361,11.185833,11.00852,10.812344,10.891568,11.529142,9.597558,8.054554,8.141325,9.2995205,9.175024,8.986393,8.4544525,8.394091,8.941121,9.556059,10.412445,9.49947,8.627994,8.499724,8.699674,9.065618,9.484379,10.386037,11.1631975,10.163452,8.578949,7.8696957,7.515069,7.4773426,8.213005,9.2995205,9.767326,9.654147,8.956212,7.6018395,7.960239,8.122461,8.062099,7.967784,8.231868,7.7187905,8.013056,8.171506,7.914967,7.643338,8.262049,7.914967,7.118943,6.4926877,6.730363,6.688864,7.3905725,7.8621507,7.635793,6.72659,6.5756855,5.8173876,5.0515447,4.5309224,4.13857,3.7613072,3.7537618,3.802806,3.8292143,3.9989824,4.696918,5.1534057,5.8966126,6.730363,6.7039547,6.888813,6.48137,5.9305663,5.704209,6.330465,7.069899,7.2585306,7.6848373,8.533678,9.386291,7.986647,7.5905213,9.650374,12.694883,12.306303,9.058073,9.103344,8.699674,7.8206515,10.155907,8.529905,8.235641,8.586494,9.024119,9.129752,8.858124,8.75249,9.337247,10.453944,11.246195,11.544232,11.283921,10.680302,10.050273,9.80128,9.710737,9.039209,8.507269,8.397863,8.526133,8.303548,8.314865,8.439363,8.560086,8.567632,8.307321,7.7225633,7.375482,7.2623034,6.8133607,7.062354,7.7037,8.68081,9.835234,10.891568,10.702937,10.759526,10.725573,10.355856,9.491924,3.8254418,2.3880715,3.85185,6.0286546,5.881522,3.99521,5.142088,6.851087,7.7829256,7.745199,10.510533,11.257513,11.638548,12.170488,12.242168,14.019074,13.9888935,12.951422,12.178034,13.422999,11.872451,11.148107,10.899114,11.370691,13.404137,13.109872,13.170234,11.050018,7.605612,7.073672,6.960493,6.470052,6.579458,7.073672,6.541732,7.496206,7.8432875,7.5829763,7.0849895,7.092535,6.779407,6.937857,6.9491754,7.043491,8.326183,8.382772,8.3525915,8.488406,8.145098,5.7570257,5.292993,4.7233267,4.9345937,6.1833324,8.103599,8.137552,7.756517,6.900131,6.089017,6.428553,6.270103,7.3000293,8.511042,9.378746,9.88805,9.593785,9.009028,8.963757,9.314611,8.922258,9.031664,8.420499,8.420499,9.039209,8.959985,8.567632,8.884532,9.027891,8.9788475,9.616421,9.224068,8.495952,7.9300575,7.809334,8.190369,8.360137,7.7338815,7.3490734,7.575431,8.088508,8.088508,8.231868,8.854351,9.680555,9.820143,8.869441,8.096053,7.4169807,7.273621,8.650629,9.261794,8.801534,8.239413,7.907422,7.5301595,7.9451485,7.9413757,7.9225125,8.016829,8.096053,8.213005,9.469289,10.220041,9.703192,8.0206,8.084735,7.4811153,6.19465,5.0025005,5.485397,5.5495315,5.3344917,5.5457587,5.926794,5.2779026,5.2288585,5.081726,5.081726,5.300538,5.6476197,5.8136153,5.983383,6.1041074,6.25124,6.6549106,6.8473144,7.0284004,6.700182,5.9192486,5.2967653,5.2250857,5.3609,5.617439,5.994701,6.571913,6.047518,5.7004366,6.439871,8.050782,9.178797,8.688355,8.439363,8.714764,9.386291,9.940866,9.310839,8.782671,8.280911,7.884786,7.8206515,7.5037513,7.586749,7.8244243,7.9036493,7.4697976,7.960239,8.228095,7.911195,7.5792036,8.771353,7.3000293,7.6622014,7.8961043,7.9753294,7.8923316,7.654656,7.6697464,7.4584794,7.3981175,7.605612,7.9300575,8.926031,8.8618965,8.239413,7.6131573,7.5792036,7.665974,7.4396167,7.066127,6.7114997,6.549277,6.7454534,6.7039547,6.8058157,7.01331,6.8699503,7.281166,7.496206,7.6131573,7.786698,8.186596,7.496206,7.2585306,7.3113475,7.462252,7.5075235,7.3792543,7.454707,8.099826,9.337247,10.853842,11.295239,11.133017,10.386037,9.623966,9.986138,9.329701,9.484379,9.933322,10.63503,12.030901,12.298758,13.030646,13.58145,13.781399,13.966258,14.200161,13.815352,13.449409,13.106099,12.155397,12.185578,13.856852,15.641303,17.28994,19.859098,19.817598,24.363613,27.747658,26.07261,17.312576,9.450426,5.040227,2.565385,1.1091517,0.36971724,0.10186087,0.026408374,0.02263575,0.124496624,0.5017591,1.2638294,1.9881734,2.2183034,2.2899833,3.3425457,4.055572,2.637065,1.5203679,1.2600567,0.543258,0.452715,0.32067314,0.150905,0.00754525,0.041498873,0.03772625,0.049044125,0.071679875,0.1056335,0.15845025,0.23013012,0.14713238,0.120724,0.1659955,0.124496624,0.026408374,0.0,0.0,0.0,0.0,0.15467763,0.25276586,0.63002837,0.9280658,0.116951376,0.0754525,0.13204187,0.17731337,0.14713238,0.030181,0.3470815,0.33953625,0.25276586,0.21881226,0.2565385,0.41121614,0.5696664,0.754525,0.9997456,1.3845534,1.750498,1.9957186,1.9655377,1.7316349,1.5580941,1.7882242,1.7731338,1.5769572,1.4826416,2.022127,1.4750963,1.9278114,2.6144292,3.1652324,3.5877664,3.4368613,3.3576362,3.4783602,3.5387223,2.9049213,3.006782,3.7763977,4.1536603,4.093298,4.534695,4.353609,4.2781568,4.2328854,4.0895257,3.6669915,4.496969,4.447925,4.406426,4.817642,5.6778007,5.617439,7.0057645,8.424272,9.216523,9.488152,9.167479,9.205205,9.26934,9.612649,11.091517,11.480098,12.351574,12.981603,13.041965,12.604341,13.04951,12.725064,12.536433,12.581704,12.140307,12.00072,12.076173,12.027128,11.706455,11.155652,11.121698,11.114153,11.966766,13.053283,12.310076,12.102581,12.019584,12.336484,12.811834,12.683565,13.502225,13.675766,13.456953,13.192869,13.324911,13.079691,13.2607765,14.151116,15.411173,16.056292,16.576914,16.705183,16.784409,16.957949,17.16167,17.237123,17.033401,16.686321,16.505234,16.980585,17.761518,18.493408,19.304522,19.908142,19.58747,20.57967,21.21347,21.14179,20.443855,19.647831,19.198889,19.455427,19.960958,20.22127,19.715738,18.99894,18.206688,17.120173,16.335466,17.255987,18.565088,20.26277,22.17549,23.790173,24.220253,21.503962,19.738375,19.613878,20.68153,21.330421,22.284895,23.073374,23.284641,23.163918,23.601542,23.737356,22.284895,20.964478,20.160908,18.92726,17.572887,17.53139,17.780382,17.799244,17.557796,17.20317,17.716248,18.995167,20.26277,20.081682,19.089483,18.082191,17.467255,17.467255,18.150099,17.901106,17.610613,18.233097,19.700647,20.919205,21.636003,21.636003,21.043703,19.67424,17.01831,11.853588,7.8961043,5.081726,3.7990334,4.9044123,4.798779,5.2326307,6.9567204,9.880505,13.087236,13.717264,13.86817,14.32843,14.66042,13.189097,10.601076,10.001229,11.193378,13.098554,13.777626,10.948157,9.654147,9.7069645,10.536942,11.212241,12.355347,12.958967,13.204187,13.317367,13.562587,13.460726,12.872196,11.951676,10.770844,9.35611,7.960239,7.24344,6.809588,6.6549106,7.1793056,7.643338,8.367682,9.378746,10.461489,11.129244,11.491416,11.427281,11.249968,10.993429,10.408672,9.952185,9.582467,9.390063,9.476834,9.97482,10.450171,10.552032,10.593531,10.518079,9.899368,9.469289,9.250477,9.092027,9.042982,9.371201,6.900131,5.8588867,5.8400235,6.255012,6.3644185,9.450426,10.699164,9.793735,7.643338,6.360646,6.809588,8.103599,8.601585,7.707473,5.8702044,5.704209,5.8136153,6.2097406,6.8058157,7.3981175,7.488661,7.3000293,6.858632,6.247467,5.6476197,5.4250345,5.3948536,5.3080835,5.05909,4.6856003,5.270357,5.907931,6.2625575,6.519096,7.3868,7.8923316,7.911195,8.458225,9.378746,9.374973,10.506761,10.631257,10.521852,10.725573,11.570641,11.23865,10.940613,10.933067,11.223559,11.574413,11.91395,11.695138,11.148107,10.536942,10.133271,8.922258,7.635793,7.707473,8.880759,9.220296,8.722309,7.9715567,8.09228,9.012801,9.473062,9.808825,8.865668,8.269594,8.461998,8.714764,8.507269,8.586494,9.273112,10.072908,9.661693,8.492179,8.028146,7.997965,8.345046,9.239159,9.710737,10.220041,10.49167,10.178542,8.873214,8.718536,8.888305,8.5563135,7.8696957,7.9338303,7.5829763,7.84706,8.084735,8.065872,7.9753294,8.371455,7.665974,7.009537,6.934085,7.352846,7.2623034,7.4094353,7.484888,7.2358947,6.462507,6.7341356,6.375736,5.4174895,4.4101987,4.3875628,4.123479,3.9197574,3.8367596,3.8593953,3.9122121,4.719554,5.3344917,5.9909286,6.48137,6.1531515,6.515323,6.771862,6.617184,6.2097406,6.1795597,6.9869013,7.707473,8.394091,8.907167,8.941121,9.623966,9.318384,9.009028,10.042727,14.120935,12.67602,11.249968,8.805306,6.971811,10.023865,8.4544525,8.009283,8.405409,9.107117,9.295748,9.178797,8.993938,9.473062,10.525623,11.25374,11.774363,11.449917,10.714255,9.982366,9.699419,9.318384,8.710991,8.14887,7.865923,8.047009,8.431817,8.5563135,8.918486,9.442881,9.450426,8.8618965,8.439363,8.001738,7.605612,7.515069,8.243186,9.220296,10.155907,11.106608,12.457208,12.487389,11.649866,10.93684,11.476325,14.498198,6.3229194,3.0520537,5.2326307,8.986393,6.013564,4.881777,5.715527,7.326438,9.242931,11.729091,10.70671,10.144588,9.540969,9.337247,10.899114,13.272095,14.4152,14.347293,13.890805,14.671739,13.257004,13.389046,12.872196,11.32542,10.167224,9.265567,8.477088,8.269594,8.382772,7.828197,6.903904,6.5756855,6.168242,5.802297,6.368191,7.6282477,7.673519,7.3000293,6.8058157,5.987156,6.609639,7.322665,7.533932,7.4697976,8.175279,7.118943,7.4811153,8.379,8.639311,6.79827,6.1305156,5.0779533,5.251494,6.8925858,8.892077,8.096053,7.122716,6.089017,5.4250345,5.881522,5.753253,7.6018395,9.152389,9.574923,9.491924,9.997457,9.703192,9.390063,9.148616,8.360137,8.835487,8.360137,8.484633,9.2995205,9.405154,8.394091,8.552541,8.643084,8.537451,9.224068,8.903395,8.650629,8.43559,8.246958,8.088508,7.5075235,7.462252,7.786698,8.028146,7.462252,7.1076255,7.0849895,7.3981175,7.9526935,8.544995,7.835742,7.443389,7.3490734,7.5565677,8.122461,8.590267,8.201687,7.5603404,7.149124,7.3188925,7.201941,7.1604424,7.492433,7.9753294,7.8734684,7.8621507,8.884532,10.182315,10.884023,9.993684,10.412445,9.507015,7.3151197,5.040227,5.0553174,4.881777,5.070408,5.692891,6.2436943,5.643847,5.6513925,5.27413,5.1458607,5.2288585,4.817642,4.6290107,5.247721,6.013564,6.6247296,7.145352,6.247467,5.9305663,5.6551647,5.2175403,4.749735,5.3156285,5.6098933,5.723072,5.8626595,6.326692,6.1644692,6.40969,7.115171,8.111144,9.027891,8.6732645,8.477088,8.616675,9.042982,9.5183325,9.216523,8.737399,8.2507305,7.911195,7.858378,7.6697464,7.91874,8.069645,7.9225125,7.61693,8.703445,8.503497,7.798016,7.4094353,8.20546,7.99042,7.997965,8.07719,7.9526935,7.5075235,6.7567716,6.436098,6.0626082,5.9909286,6.3417826,6.971811,8.035691,8.533678,8.239413,7.4999785,7.24344,7.3113475,7.0812173,6.700182,6.3531003,6.2361493,6.3832817,6.462507,6.5228686,6.458734,5.9984736,6.560595,6.749226,6.8925858,7.149124,7.4999785,6.9793563,6.8661776,7.115171,7.5829763,8.013056,7.515069,8.171506,9.22784,10.340765,11.59705,11.717773,11.940358,11.732863,11.302785,11.608367,11.408418,11.653639,12.140307,13.023102,14.856597,15.109364,14.950912,14.57365,14.252977,14.34352,14.347293,13.777626,13.023102,12.294985,11.653639,12.00072,13.630494,16.478827,19.327158,19.83269,21.74541,25.491627,26.208426,23.073374,19.300749,11.400873,5.3156285,1.8033148,0.5772116,0.32821837,0.27540162,0.47912338,0.41498876,0.24899325,0.8337501,1.7542707,2.6295197,2.7615614,2.3654358,2.5540671,4.3649273,3.6707642,2.8785129,2.6710186,2.0070364,0.95447415,0.38480774,0.1056335,0.0,0.0,0.030181,0.060362,0.049044125,0.0150905,0.03772625,0.0150905,0.011317875,0.0452715,0.09808825,0.120724,0.02263575,0.0,0.0,0.0,0.0,0.15467763,0.25276586,0.48666862,0.62248313,0.0,0.23013012,0.181086,0.120724,0.12826926,0.07922512,0.36971724,0.47912338,0.6073926,0.6375736,0.120724,0.17731337,0.32821837,0.5470306,0.875249,1.4524606,1.9391292,2.1654868,2.0183544,1.6410918,1.4600059,1.5920477,1.6373192,1.5430037,1.4147344,1.5241405,1.5656394,2.071171,2.4333432,2.625747,3.1916409,3.218049,3.199186,3.410453,3.7084904,3.519859,2.8294687,3.6707642,4.2064767,4.115934,4.6026025,4.063117,4.1272516,4.3007927,4.191386,3.4972234,4.5309224,4.776143,4.919503,5.515578,6.9491754,6.4964604,7.375482,8.718536,9.842778,10.220041,9.918231,9.786189,9.684328,9.978593,11.510279,12.14408,13.389046,14.147344,14.249205,14.441608,14.460471,13.717264,13.36641,13.539951,13.343775,13.030646,13.113645,12.706201,11.830952,11.408418,11.664956,11.796998,12.170488,12.54775,12.102581,12.162943,12.2270775,12.434572,12.728837,12.83447,13.970031,14.1926155,14.237886,14.260523,13.830443,13.50977,13.2607765,13.562587,14.6151495,16.343012,17.13149,17.003222,16.90136,17.199398,17.708702,17.701157,17.425755,17.105082,17.022083,17.523844,18.289686,19.444109,20.357084,20.775846,20.82489,21.824636,22.454664,22.775337,22.782883,22.443346,21.900087,21.639776,21.598278,21.568098,21.228561,21.209698,20.594759,18.92726,16.912678,16.45619,17.440845,19.240387,21.541689,23.477045,23.601542,21.907633,19.87419,18.704676,18.795218,19.727057,21.175745,20.806026,19.885506,19.451654,20.311813,21.334194,20.496672,19.825144,19.791191,19.300749,17.120173,16.51278,16.90136,17.803017,18.836716,18.523588,18.776354,20.470263,22.741383,22.97906,21.696367,20.82489,20.319359,20.168453,20.406128,19.65915,19.11589,19.534653,20.794708,21.888771,23.624178,24.405111,23.68454,22.481071,23.371412,16.444872,9.748463,4.6516466,2.335255,3.7763977,3.9989824,5.2175403,7.1000805,9.34102,11.691365,12.034674,12.66093,13.705947,14.777372,14.954685,12.287439,11.09529,11.634775,13.377728,14.973549,12.034674,10.646348,10.469034,10.970794,11.449917,12.770335,13.664448,13.951167,13.841762,13.958713,13.841762,13.234368,12.2270775,10.925522,9.465516,8.099826,7.0246277,6.470052,6.4964604,6.971811,7.726336,8.45068,9.224068,10.050273,10.853842,11.246195,11.234878,11.148107,11.02361,10.582213,10.423763,9.948412,9.476834,9.303293,9.691874,9.650374,9.4013815,9.310839,9.491924,9.831461,9.49947,9.020347,8.880759,8.884532,8.175279,6.1229706,5.8098426,6.175787,6.300284,5.372218,6.5341864,8.858124,9.948412,8.91094,6.379509,6.017337,6.587003,6.888813,6.670001,6.609639,5.873977,5.119452,5.1571784,5.904158,6.3719635,6.828451,7.066127,7.0057645,6.700182,6.3455553,5.987156,5.934339,5.994701,5.9607477,5.6363015,5.572167,5.9984736,6.270103,6.417235,7.115171,7.8810134,8.062099,8.431817,8.937348,8.714764,9.876732,9.937095,10.057818,10.63503,11.261286,10.95193,11.080199,11.125471,11.019837,11.170743,11.815862,11.7894535,11.299012,10.453944,9.288202,8.484633,7.726336,7.537705,8.099826,9.242931,8.446907,7.8432875,8.141325,9.06939,9.393836,9.016574,8.424272,8.114917,8.22055,8.477088,8.024373,8.111144,8.582722,8.959985,8.446907,8.771353,8.624221,8.797762,9.461743,10.148361,9.64283,9.80128,10.106862,10.167224,9.688101,9.061845,9.246704,8.929804,8.016829,7.6282477,7.6131573,7.7150183,7.888559,8.16396,8.639311,8.801534,8.096053,7.4999785,7.364164,7.4018903,7.6320205,7.4207535,7.164215,6.8397694,5.9682927,6.039973,6.3153744,5.855114,4.7912335,4.315883,4.168751,4.025391,3.9197574,3.8971217,3.983892,5.0779533,5.59103,6.0550632,6.5266414,6.590776,6.971811,7.356619,7.360391,6.9869013,6.5945487,7.394345,8.311093,9.039209,9.205205,8.386545,9.669238,10.638803,9.778644,8.616675,11.747954,13.072145,10.397354,7.3792543,6.349328,8.341274,7.2396674,7.3113475,7.956466,8.563859,8.533678,9.031664,9.484379,10.167224,10.989656,11.487643,12.0233555,11.876224,11.219787,10.34831,9.691874,9.073163,8.688355,8.416726,8.326183,8.688355,8.975075,8.850578,9.0957985,9.684328,9.756008,9.454198,9.265567,8.805306,8.326183,8.710991,9.390063,10.061591,10.427535,11.619685,16.192106,12.249713,11.02361,10.902886,11.747954,14.871688,6.598321,3.6141748,5.9494295,9.986138,8.4544525,8.216777,6.9944468,7.3792543,9.623966,11.631002,8.812852,7.8923316,8.480861,9.81637,10.770844,13.132507,14.913187,15.720529,15.629986,15.173498,14.1926155,14.154889,13.155144,10.759526,7.99042,7.7112455,8.307321,8.971302,9.318384,9.367428,7.9451485,6.820906,5.8664317,5.4401255,6.379509,7.224577,7.164215,6.903904,6.5455046,5.572167,6.439871,7.201941,7.533932,7.6923823,8.503497,6.4511886,6.417235,7.352846,8.062099,7.1793056,6.820906,5.775889,5.885295,7.303802,8.484633,7.3717093,6.6020937,5.73439,5.040227,5.4665337,5.5004873,7.5792036,9.420244,10.020092,9.661693,9.767326,9.435335,8.933576,8.428044,7.960239,8.307321,8.114917,8.560086,9.514561,9.552286,8.228095,8.280911,8.552541,8.714764,9.291975,8.756263,8.741172,8.669493,8.239413,7.424526,6.5643673,7.1000805,8.00551,8.367682,7.4018903,6.7039547,6.507778,6.530414,6.7341356,7.322665,7.115171,7.1038527,7.3075747,7.654656,7.9828744,8.0206,7.624475,7.0359454,6.677546,7.122716,6.670001,6.5568223,6.888813,7.364164,7.2698483,7.2358947,7.7678347,8.929804,10.201178,10.457717,11.623458,10.782163,8.152642,5.2326307,4.7836885,4.478106,5.2250857,5.9003854,5.9720654,5.485397,5.9984736,5.523123,5.1760416,5.089271,4.432834,4.647874,5.379763,5.9305663,6.175787,6.5455046,5.2779026,4.817642,4.749735,4.798779,4.821415,5.4740787,5.5382137,5.485397,5.6400743,6.1606965,6.217286,6.6058664,7.122716,7.6131573,8.001738,8.228095,8.548768,8.68081,8.692128,9.005256,9.156161,8.880759,8.424272,8.084735,8.231868,7.9262853,7.9753294,8.107371,8.141325,7.9828744,8.29223,8.14887,7.8432875,7.635793,7.752744,8.231868,7.967784,7.77538,7.4471617,6.8133607,5.7796617,5.3948536,5.089271,5.243949,5.783434,6.156924,6.6058664,7.281166,7.375482,6.8473144,6.4134626,6.126743,6.0814714,5.885295,5.541986,5.4401255,5.4174895,5.775889,6.006019,5.9003854,5.5495315,6.439871,6.617184,6.6360474,6.719045,6.7643166,7.020855,7.0510364,7.0887623,7.2962565,7.8017883,6.9982195,8.337502,9.884277,10.823661,11.487643,11.246195,11.785681,12.381755,12.785426,13.245687,14.083209,13.996439,13.958713,14.611377,16.260014,16.35433,15.241405,14.132254,13.607859,13.622949,13.117417,12.781653,12.196897,11.438599,11.076427,11.559323,12.989148,16.58446,20.142044,18.025602,22.17549,24.352295,23.601542,21.07011,20.028866,13.29473,6.043745,1.5807298,0.46026024,0.49421388,0.5055317,1.086516,1.0223814,0.452715,0.87902164,1.2110126,1.7769064,1.9089483,1.6071383,1.5241405,3.5877664,3.9008942,3.5839937,3.2520027,3.0256453,1.1280149,0.27917424,0.02263575,0.00754525,0.003772625,0.0,0.02263575,0.0754525,0.1358145,0.1358145,0.10186087,0.11317875,0.16222288,0.21503963,0.20372175,0.1358145,0.11317875,0.1056335,0.12826926,0.23013012,0.09808825,0.06413463,0.03772625,0.0,0.0,0.5281675,0.31312788,0.0754525,0.09808825,0.23013012,0.241448,0.4376245,0.80734175,0.97333723,0.19994913,0.17354076,0.22258487,0.46026024,0.91674787,1.5354583,2.173032,2.5087957,2.123988,1.3770081,1.3958713,1.388326,1.5845025,1.4901869,1.146878,1.1581959,1.9240388,2.0787163,2.082489,2.2371666,2.6483827,3.4632697,3.1539145,3.1425967,3.7537618,4.217795,3.2557755,3.5877664,3.8141239,3.7613072,4.478106,4.0480266,4.4818783,4.8365054,4.606375,3.7386713,4.3649273,5.0741806,5.704209,6.5228686,8.239413,8.043237,8.160188,9.009028,10.0465,9.759781,9.910686,9.895596,9.948412,10.416218,11.778135,12.623203,13.841762,14.683057,15.124454,15.863888,15.230087,13.932304,13.226823,13.419228,13.856852,13.407909,13.634267,13.170234,12.121444,12.064855,12.166716,12.362892,12.50248,12.46098,12.128989,12.498707,13.053283,12.947649,12.415709,12.774108,14.177525,14.566105,14.890551,15.218769,14.769827,14.747191,14.181297,14.1926155,15.377219,17.787928,18.949896,18.463226,17.716248,17.667202,18.859352,18.470772,17.969013,17.621931,17.565342,17.7917,18.26705,19.708193,20.806026,21.009748,20.534397,20.96825,21.771818,22.684793,23.38273,23.461954,23.631723,22.643295,21.817091,21.719002,22.167944,23.235598,23.099783,21.669958,19.462973,17.572887,16.965494,18.12369,20.519308,22.933788,23.461954,22.42071,20.68153,19.002712,18.187824,19.081938,20.689075,19.757236,18.629223,18.5085,19.440336,20.440083,20.243906,20.183544,20.50799,20.37972,17.82188,16.414692,16.105335,16.837225,18.519815,18.953669,19.61765,21.481327,23.975033,25.008732,23.243143,22.548979,22.137764,21.632233,21.09652,20.153362,19.48561,19.523335,20.477808,22.352802,25.419947,25.880207,24.393793,23.639269,28.294687,20.040184,12.019584,5.481624,2.04099,3.663219,3.7235808,5.353355,7.752744,9.948412,10.816116,11.117926,11.751727,12.664702,13.93985,15.788436,13.754991,13.36641,13.238141,13.20796,14.366156,13.4644985,12.310076,11.385782,11.200924,12.272349,13.230596,13.853079,14.1926155,14.388792,14.675511,14.230342,13.313594,12.170488,10.899114,9.450426,8.107371,6.85486,6.4021444,6.673774,6.79827,7.443389,8.0206,8.533678,9.065618,9.767326,10.121953,10.382264,10.574668,10.631257,10.374719,10.4049,9.944639,9.424017,9.133525,9.224068,8.937348,8.718536,8.639311,8.771353,9.186342,9.314611,8.89585,8.544995,7.9828744,6.043745,5.975838,6.4021444,6.6850915,6.5228686,5.9494295,5.9532022,7.3151197,9.446653,10.740664,8.560086,6.4436436,6.0362,5.772116,5.511805,6.530414,6.5756855,4.927048,4.172523,4.881777,5.613666,6.466279,6.9793563,7.1378064,7.0774446,7.069899,6.696409,6.4436436,6.466279,6.692637,6.820906,6.175787,6.40969,6.771862,7.039718,7.5188417,8.473316,8.975075,9.239159,9.239159,8.714764,9.122208,9.291975,9.725827,10.340765,10.499215,9.827688,10.042727,10.170997,9.937095,9.786189,10.627484,10.997202,10.989656,10.597303,9.688101,8.843033,8.348819,7.7414265,7.4471617,8.778898,8.171506,8.062099,8.367682,8.801534,8.907167,8.439363,8.224322,7.7602897,7.3000293,7.865923,7.5075235,7.8961043,8.552541,8.809079,7.798016,8.956212,8.9788475,9.208978,9.918231,10.295494,9.061845,8.601585,8.567632,8.869441,9.684328,9.061845,9.114662,8.827943,7.967784,7.0548086,7.4282985,7.6320205,7.8998766,8.360137,9.050528,9.250477,9.216523,8.782671,8.035691,7.3113475,7.748972,7.6320205,7.4094353,7.0849895,6.217286,5.4212623,5.8626595,6.1116524,5.5268955,4.2404304,4.036709,4.0895257,4.164978,4.1536603,4.063117,5.311856,5.7909794,6.330465,7.2396674,8.322411,8.507269,8.216777,7.7301087,7.322665,7.250985,8.27714,8.771353,9.092027,9.265567,8.948667,9.103344,9.940866,10.0276375,8.975075,7.4396167,9.971047,7.432071,5.613666,6.1795597,6.670001,5.8928404,6.3832817,7.1868505,7.699928,7.643338,8.75249,9.884277,10.846297,11.544232,12.0082655,12.291212,12.238396,11.695138,10.729345,9.650374,9.224068,9.122208,9.250477,9.556059,10.0465,9.699419,9.2844305,9.280658,9.597558,9.544742,9.940866,10.080454,9.756008,9.367428,9.918231,10.084227,10.106862,9.891823,11.200924,17.659658,10.061591,9.190115,10.472807,11.532914,12.208215,7.2472124,5.1043615,5.8098426,8.548768,11.668729,11.3971,8.024373,6.9869013,8.439363,7.277394,6.217286,6.277648,8.993938,12.453435,11.257513,13.302276,14.898096,16.143063,16.475054,14.66042,14.298248,13.151371,11.559323,9.608876,7.1340337,8.937348,9.012801,8.262049,8.073418,10.340765,8.771353,6.7756343,5.9003854,6.3116016,6.820906,6.590776,6.6549106,6.741681,6.6134114,6.096562,6.4511886,6.6549106,6.9680386,7.643338,8.933576,6.598321,5.6023483,5.726845,6.3719635,6.5643673,6.7944975,6.3153744,6.5568223,7.443389,7.3981175,6.519096,6.3531003,5.80607,5.010046,5.3344917,5.6551647,7.435844,9.397609,10.589758,10.370946,8.956212,8.409182,8.013056,7.647111,7.816879,7.6584287,7.805561,8.59404,9.5032425,9.133525,8.107371,8.394091,8.98262,9.439108,9.918231,9.239159,9.031664,8.763808,8.073418,6.790725,6.1795597,6.862405,7.8395147,8.397863,8.137552,7.183078,6.462507,6.0022464,5.9607477,6.63982,6.990674,7.1981683,7.3075747,7.4697976,7.9338303,7.594294,7.1793056,6.677546,6.2814207,6.3719635,6.168242,6.221059,6.3116016,6.296511,6.126743,6.0211096,6.2135134,6.903904,7.956466,8.903395,10.604849,10.27663,8.069645,5.323174,4.5799665,4.2706113,5.4401255,5.904158,5.2590394,4.889322,6.013564,5.674028,5.2326307,5.0251365,4.353609,5.304311,5.9418845,5.794752,5.2062225,5.3609,4.5988297,4.221567,4.195159,4.504514,5.172269,5.3609,5.0515447,4.9421387,5.3458095,6.1720147,6.0739264,6.0248823,6.3153744,6.749226,6.651138,7.726336,8.631766,8.809079,8.469543,8.601585,8.971302,8.918486,8.541223,8.228095,8.684583,8.156415,7.7338815,7.84706,8.258276,8.035691,7.0963078,7.3717093,7.9036493,8.141325,7.937603,6.6850915,7.01331,6.7643166,6.5266414,6.330465,5.6476197,4.938366,4.961002,5.304311,5.7306175,6.19465,6.379509,6.4247804,6.436098,6.228604,5.3269467,4.983638,5.0175915,5.040227,4.8025517,4.1800685,3.92353,4.217795,4.4743333,4.644101,5.2175403,5.4401255,5.3269467,5.292993,5.4476705,5.6287565,6.752999,6.8774953,6.590776,6.4926877,7.201941,7.2887115,8.20546,9.416472,10.216269,9.767326,10.510533,10.887795,11.370691,11.962994,12.208215,12.830698,13.2607765,13.664448,14.037937,14.222796,13.902123,13.347548,12.928786,12.770335,12.755245,12.3289385,12.751472,12.147853,10.56335,9.963503,11.3669195,12.577931,15.131999,17.757746,16.403374,22.945105,25.917934,24.76351,21.503962,20.73812,10.789707,4.1989317,1.1242423,0.60362,0.58098423,0.33576363,0.8978847,1.1883769,1.026154,1.0978339,0.9997456,0.7469798,0.9808825,1.6335466,1.9391292,1.6071383,1.2223305,0.8563859,0.56212115,0.36594462,0.29426476,0.12826926,0.03772625,0.041498873,0.0150905,0.003772625,0.0,0.27540162,0.6828451,0.67152727,0.5017591,0.52062225,0.77338815,0.9242931,0.29049212,0.5357128,0.5583485,0.5281675,0.6451189,1.1431054,0.4979865,0.32821837,0.19240387,0.0,0.0,0.35462674,0.41498876,0.24899325,0.094315626,0.35085413,0.071679875,0.38480774,0.49421388,0.24899325,0.1358145,0.4074435,0.30935526,0.39989826,0.72811663,0.83752275,1.7919968,2.1390784,1.8297231,1.2525115,1.2525115,1.5920477,1.5430037,1.2789198,1.1431054,1.6335466,1.6675003,1.8787673,2.203213,2.4295704,2.1956677,3.8707132,4.187614,4.1800685,4.327201,4.5460134,3.8895764,3.731126,3.712263,3.9688015,5.1269975,5.553304,5.1571784,4.6026025,4.191386,3.8593953,3.9574835,4.991183,6.6020937,8.27714,9.337247,9.435335,9.103344,8.98262,9.039209,8.575176,9.918231,9.669238,9.186342,9.288202,10.253995,11.876224,13.664448,14.924504,15.290449,14.739646,14.886778,13.411682,12.038446,11.415963,11.125471,11.465008,12.366665,12.725064,12.464753,12.528888,12.162943,11.9064045,11.996947,12.155397,11.581959,12.14408,13.143826,12.985375,12.064855,12.785426,13.347548,13.981348,14.226569,14.317112,15.196134,16.260014,16.388283,17.286167,19.289433,21.375692,22.194353,21.447372,19.372429,17.516298,18.738628,18.995167,19.01403,18.693357,18.414183,19.01403,18.85558,19.60256,20.643805,21.254969,20.583443,19.862871,20.051502,20.813572,21.888771,23.069601,23.182781,21.38701,19.964731,19.787418,20.323132,21.07011,22.096264,22.556524,22.24717,21.636003,19.670467,18.376457,18.632996,20.130728,21.360603,20.202406,19.84778,19.349794,18.72731,18.99894,19.70442,19.28566,18.689585,18.719765,20.051502,20.46649,21.183289,22.03213,22.56407,22.062311,19.73083,17.784155,16.399601,15.712983,15.82239,16.957949,18.414183,19.893051,21.175745,22.141537,21.45869,21.568098,20.900343,19.606333,19.606333,19.87796,19.606333,18.519815,18.229324,22.232079,24.623924,19.217752,15.354584,17.969013,27.589207,21.752956,13.619176,6.405917,2.8822856,5.3873086,4.4101987,4.991183,7.213259,9.910686,10.680302,11.314102,10.899114,10.435081,10.834979,12.909923,14.007756,15.335721,15.120681,13.8870325,14.449154,15.426264,14.049255,12.67602,12.638294,14.237886,14.68683,14.260523,14.173752,14.724555,15.275358,14.222796,12.864652,11.295239,9.756008,8.620448,7.364164,6.903904,7.020855,7.4471617,7.8734684,7.726336,7.752744,8.07719,8.461998,8.314865,8.963757,9.756008,10.646348,11.09529,10.069136,9.582467,9.058073,8.654402,8.503497,8.710991,8.345046,8.695901,8.858124,8.646856,8.575176,8.537451,8.722309,8.843033,8.865668,8.986393,6.156924,5.4288073,5.13077,4.98741,6.1342883,7.805561,9.276885,10.56335,12.90615,18.75372,10.31813,7.284939,7.039718,7.1906233,5.553304,7.141579,5.66271,4.055572,3.9688015,5.7381625,6.6662283,7.043491,7.4282985,7.828197,7.707473,7.643338,7.454707,7.175533,7.039718,7.492433,6.9567204,6.749226,6.9189944,7.4207535,8.118689,8.729855,9.144843,9.046755,8.52236,8.058327,8.288457,8.869441,9.533423,10.084227,10.374719,9.374973,8.986393,8.786444,8.710991,9.0807085,9.420244,10.231359,11.0613365,11.457462,10.970794,9.125979,8.428044,8.2507305,8.280911,8.499724,8.29223,8.167733,8.118689,8.00551,7.5527954,7.356619,7.4811153,7.4282985,7.2283497,7.462252,6.752999,7.0887623,8.13378,9.201432,9.261794,8.07719,8.122461,8.443134,8.68081,9.046755,8.3525915,8.013056,8.039464,8.52236,9.65792,9.378746,8.922258,8.280911,7.4471617,6.40969,7.1038527,8.047009,8.816625,9.039209,8.394091,8.367682,9.405154,10.065364,9.593785,7.9338303,7.677292,7.432071,7.394345,7.5829763,7.828197,6.300284,5.66271,5.492942,5.3910813,4.9760923,4.2404304,4.06689,4.3800178,4.6856003,4.074435,4.3686996,5.5382137,6.937857,8.262049,9.567377,9.763554,8.812852,7.8961043,7.5301595,7.567886,8.507269,8.194141,8.152642,9.0807085,10.86516,9.876732,9.1976595,9.540969,9.891823,7.537705,8.477088,7.8961043,7.0812173,6.9869013,8.269594,6.3908267,5.406172,5.96452,7.707473,9.291975,9.559832,9.510788,9.95973,11.080199,12.37421,12.215759,11.857361,11.434827,10.917976,10.103089,10.212496,10.201178,10.34831,10.657665,10.86516,10.499215,10.295494,10.242677,10.054046,9.201432,9.676784,10.253995,10.370946,10.054046,9.918231,10.163452,10.891568,11.793225,11.812089,9.125979,8.160188,9.137298,11.536687,15.116908,19.911915,17.554024,9.97482,4.7836885,5.2137675,10.069136,8.360137,6.688864,6.2814207,6.9982195,7.3377557,9.7069645,10.555805,10.427535,9.963503,9.903141,11.68382,12.570387,13.717264,14.5132885,12.574159,12.525115,10.378491,8.379,7.3415284,6.6850915,10.272858,9.522105,7.564113,6.7152724,8.499724,7.5226145,6.307829,6.417235,7.515069,7.3717093,6.858632,7.01331,6.79827,6.2814207,6.620957,6.6850915,6.432326,6.677546,7.383027,7.673519,6.0626082,5.138315,4.7308717,4.817642,5.5382137,5.723072,5.8966126,6.903904,8.118689,7.4471617,6.7643166,6.647365,6.0776987,5.2250857,5.43258,6.1644692,7.986647,9.695646,10.382264,9.431562,7.3905725,7.092535,7.4169807,7.752744,8.009283,8.145098,8.416726,8.880759,9.073163,8.009283,8.341274,9.5032425,10.005001,9.857869,10.589758,10.370946,10.020092,9.307066,8.303548,7.4018903,6.888813,7.647111,8.345046,8.688355,9.446653,8.616675,6.8435416,5.27413,4.919503,6.651138,7.1906233,7.515069,7.7414265,7.8734684,7.8131065,7.567886,7.066127,6.330465,5.481624,4.7610526,5.492942,6.096562,6.0286546,5.406172,5.0062733,5.149633,5.1873593,5.4703064,6.047518,6.670001,7.413208,7.1302614,6.0022464,4.606375,3.9197574,3.9348478,5.191132,5.6476197,5.1081343,5.2175403,6.4511886,6.3644185,5.96452,5.455216,4.255521,4.610148,5.6778007,6.1795597,5.836251,5.3873086,4.9345937,3.9688015,3.6330378,4.353609,5.8437963,5.0251365,4.5761943,4.6252384,5.1835866,6.1342883,6.19465,6.119198,6.1908774,6.4926877,6.8963585,8.299775,8.439363,7.9413757,7.4811153,7.798016,8.371455,8.412953,8.00551,7.7942433,9.001483,8.903395,8.296002,7.865923,7.5829763,6.670001,7.1566696,7.1038527,7.322665,7.865923,8.009283,6.0626082,6.273875,6.247467,6.119198,5.9192486,5.5495315,5.0741806,4.90064,4.9949555,5.3269467,5.8890676,6.198423,6.085244,5.674028,5.1232247,4.6290107,4.5007415,4.5988297,4.538468,4.29702,4.1800685,4.1310244,4.195159,4.3007927,4.515832,5.05909,5.3759904,5.534441,5.7079816,6.149379,7.1793056,7.5603404,6.9680386,6.620957,6.9982195,7.8131065,8.201687,8.601585,9.186342,9.842778,10.182315,9.616421,9.695646,10.26154,11.09529,11.91395,12.966512,12.894833,12.664702,12.853333,13.671993,13.109872,13.147598,13.091009,12.823153,12.792972,12.785426,12.90615,12.113899,10.846297,10.989656,12.608112,13.63804,14.569878,15.501716,16.146835,22.552752,26.310287,27.543936,26.921452,25.642532,13.098554,5.5306683,3.5424948,4.636556,3.2029586,1.8070874,0.80734175,0.33953625,0.30935526,0.392353,1.3091009,1.3241913,1.1242423,1.0072908,0.8639311,0.6413463,0.6149379,1.237421,1.8900851,0.8526133,1.8863125,1.4977322,0.72811663,0.17731337,0.0150905,0.011317875,0.011317875,0.06790725,0.15467763,0.16976812,0.15467763,0.2678564,0.32444575,0.3055826,0.362172,0.6187105,0.41121614,0.32067314,0.5470306,0.91297525,0.5394854,0.39989826,0.35462674,0.38480774,0.6111652,0.19240387,0.08299775,0.049044125,0.018863125,0.071679875,0.16976812,0.43385187,0.7809334,1.0638802,1.0525624,0.8224323,0.73188925,0.694163,0.70170826,0.83752275,1.1280149,1.3317367,1.3505998,1.2562841,1.2751472,1.599593,1.871222,2.0485353,2.11267,2.071171,2.3126192,2.11267,2.1994405,2.746471,3.3915899,4.7346444,5.66271,6.0814714,6.1418333,6.2436943,5.643847,5.040227,5.6325293,6.6624556,5.4212623,6.4436436,5.945657,5.6098933,5.745708,5.2892203,5.2779026,6.0286546,7.326438,8.5563135,8.68081,8.98262,9.042982,9.26934,9.6051035,9.540969,10.510533,11.25374,11.287694,10.733118,10.303039,10.608622,11.751727,12.932558,13.732355,14.128481,13.611631,12.325166,11.672502,11.883769,11.989402,11.981857,11.92904,12.344029,12.785426,11.879996,11.944131,12.00072,12.2270775,12.566614,12.717519,12.468526,12.717519,12.864652,13.0646,14.215251,14.592513,14.667966,15.07541,16.078928,17.554024,18.1086,17.689838,18.168962,19.455427,19.523335,19.647831,19.180025,18.157644,17.184307,17.41821,17.95015,18.814081,19.395065,19.57615,19.74592,19.840235,19.889278,19.836462,19.65915,19.38752,19.372429,19.798737,19.557287,18.89708,19.447882,20.013775,19.889278,20.111864,20.689075,20.594759,21.122927,21.994404,22.594252,22.458437,21.27006,19.108345,18.350048,18.708447,19.83269,21.300241,20.541943,19.519562,18.621677,18.21046,18.606586,18.991394,19.195116,19.31584,19.512016,20.013775,19.979822,20.217497,20.504217,20.832436,21.405874,20.723028,19.979822,18.806536,17.557796,17.335213,17.399347,18.270823,19.093256,19.542198,19.821371,20.349539,20.919205,20.232588,18.75372,18.715992,19.296976,19.112118,18.92726,19.644058,22.281124,23.277096,17.969013,14.460471,16.437326,23.156372,17.176762,12.498707,8.627994,6.1041074,6.4964604,6.1342883,5.3759904,6.5341864,9.205205,10.265312,11.321648,11.125471,10.419991,10.303039,12.2119875,13.52486,14.211478,13.694629,12.649611,12.985375,13.219278,13.328684,13.230596,13.306048,14.407655,14.603831,14.400109,14.68683,15.430037,15.675257,15.086727,13.751218,12.140307,10.54826,9.122208,8.126234,7.7678347,7.5829763,7.4207535,7.4471617,7.3490734,7.1981683,7.394345,7.9338303,8.412953,8.846806,9.850324,10.676529,10.804798,9.9257765,9.718282,9.344792,8.922258,8.428044,7.699928,8.114917,8.394091,8.495952,8.416726,8.197914,7.9262853,7.7150183,8.016829,8.495952,8.024373,7.3490734,6.1720147,4.6629643,3.4670424,3.7160356,5.0854983,7.0170827,10.27663,14.25675,16.957949,13.826671,10.412445,8.59404,8.22055,7.092535,7.858378,7.322665,5.9230213,4.776143,5.6778007,7.0246277,7.4773426,7.7602897,7.9828744,7.643338,7.3490734,7.33021,7.364164,7.3000293,7.039718,6.8171334,6.907676,6.9680386,6.964266,7.141579,8.307321,8.710991,8.382772,7.6622014,7.1793056,7.3792543,7.9225125,8.379,8.590267,8.68081,8.45068,8.299775,8.009283,7.752744,8.088508,9.359882,10.310584,10.812344,10.653893,9.578695,8.869441,8.379,8.145098,8.262049,8.903395,8.031919,7.7037,7.8621507,8.047009,7.383027,6.971811,6.983129,7.062354,7.254758,8.024373,7.665974,7.356619,7.748972,8.684583,9.21275,8.262049,7.54525,7.7904706,8.688355,8.8769865,8.68081,8.582722,8.620448,8.744945,8.816625,8.563859,8.29223,7.7716074,7.115171,6.79827,7.2396674,7.484888,8.050782,8.718536,8.488406,8.337502,8.567632,9.046755,9.178797,7.911195,7.7716074,7.7150183,7.673519,7.6923823,7.9262853,7.141579,6.168242,5.6363015,5.458988,4.8402777,4.7044635,4.3649273,4.3724723,4.851596,5.4891696,5.5797124,6.4210076,7.594294,8.616675,8.944894,8.76758,8.333729,8.386545,8.888305,9.031664,9.046755,9.295748,9.480607,9.903141,11.498961,10.529396,10.529396,11.193378,11.461235,9.514561,8.82417,9.125979,9.378746,9.65792,11.1631975,10.016319,9.574923,8.428044,7.4999785,10.072908,9.725827,9.42779,9.718282,10.668983,11.887542,11.434827,11.0613365,10.555805,9.944639,9.480607,9.688101,10.061591,10.612394,11.302785,12.049765,11.819634,11.608367,11.3971,11.18206,10.970794,11.065109,11.299012,11.053791,10.287949,9.525878,9.6051035,10.423763,11.457462,11.921495,10.808571,8.182823,7.786698,10.091772,15.0376835,22.013268,25.963205,17.350302,7.997965,5.191132,11.668729,9.480607,6.8699503,5.7494807,6.387054,7.413208,9.567377,10.895341,11.246195,10.921749,10.684074,10.767072,10.408672,10.79348,11.661184,11.302785,10.220041,9.491924,8.130007,6.7454534,7.5490227,9.175024,8.088508,6.6813188,6.145606,6.4738245,6.571913,6.752999,6.730363,6.439871,6.039973,6.3945994,6.477597,6.3832817,6.4474163,7.220804,7.0472636,6.9227667,6.94163,6.8963585,6.270103,5.4401255,5.2892203,5.2175403,5.2099953,5.832478,6.258785,6.19465,6.511551,7.0963078,6.8359966,6.79827,6.9227667,6.5341864,5.802297,5.726845,6.2021956,7.537705,8.661947,8.922258,8.088508,7.201941,7.145352,7.092535,6.937857,7.2924843,8.273367,8.809079,9.137298,9.0957985,8.122461,8.733627,9.533423,9.937095,9.81637,9.5032425,9.616421,9.454198,9.020347,8.424272,7.8508325,7.9338303,7.986647,8.239413,8.835487,9.846551,8.948667,7.333983,6.0626082,5.696664,6.2851934,6.832224,7.3075747,7.3868,7.1868505,7.2623034,7.0887623,6.63982,5.9607477,5.353355,5.383536,6.2323766,6.4926877,6.006019,5.089271,4.52715,4.5497856,4.7648253,5.0251365,5.3156285,5.753253,6.8473144,6.273875,5.194905,4.2102494,3.3727267,3.802806,4.6742826,5.485397,5.983383,6.1833324,6.3116016,6.0739264,5.8173876,5.481624,4.5988297,4.142342,4.678055,5.3986263,5.7306175,5.3382645,5.13077,4.8063245,4.7610526,4.949684,4.8553686,3.9122121,3.9386206,4.38379,4.82896,4.9987283,5.6061206,5.511805,5.934339,6.971811,7.6282477,8.605357,8.8769865,8.782671,8.616675,8.639311,8.382772,7.9413757,7.809334,7.9753294,7.9036493,7.3000293,7.2358947,7.3981175,7.5188417,7.364164,7.069899,6.990674,7.3377557,7.956466,8.314865,5.9230213,5.6363015,5.6815734,5.6513925,5.4250345,5.149633,4.8440504,4.6931453,4.8063245,5.1647234,5.613666,5.6476197,5.4703064,5.353355,5.2628117,4.8855495,4.6516466,4.5950575,4.478106,4.349837,4.538468,4.538468,4.678055,4.7912335,4.9044123,5.2590394,5.783434,5.8966126,6.1644692,6.802043,7.6886096,7.84706,7.3868,7.2924843,7.907422,8.918486,8.918486,9.1976595,9.480607,9.65792,9.763554,9.133525,9.06939,9.1976595,9.540969,10.502988,12.178034,12.377983,12.08749,11.981857,12.453435,12.219532,12.540206,12.498707,12.132762,12.427027,12.200669,11.834724,11.427281,11.291467,11.959221,13.909668,16.290195,16.35433,15.286676,18.206688,22.315077,25.457674,27.80802,28.781357,27.027086,12.630749,5.455216,3.399135,3.561358,2.2409391,2.5389767,1.7089992,0.98465514,0.7469798,0.51684964,0.9997456,0.84884065,0.56212115,0.38103512,0.30181,0.36971724,0.7167987,1.3392819,1.720317,0.8224323,2.7804246,1.841041,0.58098423,0.10186087,0.0150905,0.0150905,0.011317875,0.00754525,0.011317875,0.026408374,0.06790725,0.120724,0.12826926,0.120724,0.23390275,0.44139713,0.29426476,0.35085413,0.73566186,1.146878,0.5055317,0.28294688,0.2867195,0.35839936,0.4074435,0.116951376,0.0452715,0.19994913,0.362172,0.08299775,0.1659955,0.35085413,0.79602385,1.2713746,1.1355602,1.2487389,1.4600059,1.629774,1.6335466,1.3619176,1.3204187,1.2751472,1.2034674,1.1544232,1.2449663,1.6939086,2.2296214,2.2107582,1.8599042,2.2371666,2.4069347,2.9954643,3.3350005,3.500996,4.323428,6.85486,7.24344,7.039718,6.9869013,6.9793563,6.722818,6.273875,6.881268,7.8244243,6.398372,7.432071,6.9869013,6.628502,6.673774,6.187105,6.25124,6.7680893,7.333983,7.9941926,9.239159,10.087999,10.272858,10.917976,11.895086,11.785681,12.095036,12.751472,12.721292,11.940358,11.348056,11.566868,11.740409,12.691111,14.030393,14.151116,13.773854,12.89106,12.272349,12.291212,12.902377,12.1252165,11.895086,12.245941,12.642066,11.993175,11.857361,11.676274,12.08749,13.045737,13.841762,13.894578,13.6833105,13.630494,13.924759,14.509516,14.434063,15.086727,16.097792,17.33144,18.912169,19.293203,18.244415,17.380484,17.184307,16.980585,17.320122,17.953922,18.274595,18.150099,17.931286,18.72731,19.927006,20.768301,20.900343,20.413673,19.787418,19.232841,18.53868,18.184053,19.31584,19.651604,20.232588,19.610106,18.070873,17.63325,18.03692,18.297232,19.312067,20.677757,20.670212,20.477808,21.149336,21.934042,22.081175,20.858843,18.599041,17.625704,17.686066,18.61036,20.30804,20.613623,20.130728,19.398838,18.742401,18.289686,18.52736,18.964987,19.093256,18.980076,19.281887,19.48561,19.678013,20.093,20.802254,21.688822,21.647322,20.938068,19.783646,18.68204,18.391546,18.040693,19.097027,20.145817,20.719257,21.319103,21.620914,21.560553,20.560806,19.462973,20.496672,20.68153,20.198635,20.217497,20.938068,21.605824,22.677248,20.100546,18.214233,19.130981,22.733839,16.452417,13.434318,10.910432,8.386545,7.598067,6.2323766,5.4250345,6.40969,8.537451,9.2844305,10.287949,10.978339,11.664956,12.525115,13.585222,14.6151495,15.128226,14.332202,12.577931,11.363147,11.261286,11.721546,12.279895,12.913695,14.064346,14.418973,14.43029,14.713238,15.256495,15.411173,15.731846,15.045229,13.604086,11.7894535,10.087999,8.771353,8.29223,8.058327,7.8244243,7.7150183,7.586749,7.594294,7.8621507,8.254503,8.394091,8.89585,9.367428,9.64283,9.740918,9.850324,9.782416,9.665465,9.616421,10.076681,11.812089,8.246958,7.1264887,7.069899,7.3000293,7.635793,8.065872,7.9451485,7.752744,7.91874,8.835487,8.160188,6.771862,5.3344917,4.406426,4.459243,4.6554193,5.7192993,7.6584287,10.47658,14.203933,11.027383,8.98262,7.8621507,7.352846,7.009537,6.903904,6.7341356,5.802297,4.7572803,5.613666,7.032173,7.7414265,7.9828744,7.964011,7.865923,7.33021,7.118943,6.990674,6.8699503,6.862405,6.651138,7.183078,7.598067,7.533932,7.145352,7.8508325,7.9300575,7.6282477,7.2170315,6.9869013,6.858632,7.0963078,7.4207535,7.575431,7.3377557,7.1340337,7.3075747,7.284939,7.118943,7.4773426,9.21275,10.265312,10.612394,10.238904,9.148616,8.699674,8.439363,8.265821,8.318638,8.98262,8.307321,7.533932,7.4169807,7.7942433,7.5792036,6.9152217,6.7454534,6.8171334,7.066127,7.6320205,7.4282985,7.2887115,7.677292,8.59404,9.574923,9.774872,8.737399,8.179051,8.6581745,9.593785,9.163706,8.224322,8.009283,8.511042,8.469543,8.107371,7.752744,7.062354,6.3116016,6.4134626,7.062354,6.779407,6.8737226,7.6697464,8.514814,9.144843,9.171251,9.125979,8.993938,8.224322,7.756517,7.8395147,7.8131065,7.5905213,7.647111,7.5263867,6.749226,5.9682927,5.281675,4.2291126,4.402653,4.719554,4.7120085,4.5761943,5.1760416,6.1116524,6.862405,7.4584794,7.9828744,8.560086,8.239413,7.9715567,8.348819,9.031664,8.741172,8.6732645,9.276885,9.639057,9.914458,11.317875,10.940613,11.257513,12.0082655,12.381755,10.997202,10.303039,10.272858,9.861642,9.405154,10.623712,14.535924,12.615658,8.990166,6.617184,7.284939,7.647111,8.231868,9.016574,9.914458,10.767072,11.038701,10.993429,10.525623,9.865415,9.559832,9.507015,9.616421,10.20495,11.129244,11.766817,11.925267,11.634775,11.661184,12.049765,12.117672,11.438599,11.664956,11.876224,11.642321,11.050018,10.412445,10.834979,11.529142,12.0082655,12.064855,10.3634,10.442626,11.344283,13.20796,17.255987,26.32915,19.263023,9.246704,4.4743333,8.114917,9.390063,8.345046,7.24344,7.111398,7.7150183,8.533678,8.495952,7.91874,7.598067,8.809079,8.601585,8.375228,9.371201,11.121698,11.434827,9.914458,8.345046,6.8850408,6.2361493,7.6584287,7.5188417,6.0324273,4.957229,4.8666863,5.149633,5.511805,6.670001,7.01331,6.307829,5.73439,5.8966126,5.934339,6.1795597,6.8359966,7.956466,7.4169807,7.152897,6.8133607,6.1644692,5.070408,4.82896,4.9157305,5.2364035,5.7381625,6.417235,6.790725,6.6247296,6.4964604,6.6322746,6.911449,6.952948,6.9227667,6.8850408,6.643593,5.73439,5.621211,6.428553,7.213259,7.5226145,7.3679366,7.24344,7.3717093,7.1604424,6.779407,7.118943,7.907422,8.371455,8.695901,8.83926,8.533678,9.0543,9.582467,10.208723,10.536942,9.661693,9.235386,8.797762,8.367682,8.126234,8.412953,8.397863,8.13378,8.0206,8.265821,8.8769865,8.329956,7.201941,6.349328,6.1003346,6.258785,6.677546,7.2396674,7.2283497,6.7341356,6.63982,6.541732,6.1116524,5.6061206,5.300538,5.485397,6.356873,6.647365,6.1531515,5.191132,4.6290107,4.425289,4.564876,4.67051,4.708236,4.983638,6.3153744,5.934339,5.1269975,4.4743333,3.8669407,4.5422406,5.1647234,5.7872066,6.2889657,6.379509,6.2097406,5.8098426,5.3571277,4.908185,4.38379,4.323428,4.508287,4.908185,5.270357,5.1345425,5.515578,5.3986263,4.9647746,4.3422914,3.6292653,3.640583,4.104616,4.5837393,4.8440504,4.8327327,5.409944,5.7419353,6.3116016,7.164215,7.9225125,8.480861,8.6581745,8.684583,8.646856,8.465771,8.337502,7.9338303,7.7338815,7.756517,7.5565677,6.7944975,6.6020937,6.9152217,7.383027,7.383027,7.5301595,7.9338303,8.0206,7.854605,8.145098,5.4703064,4.98741,4.908185,4.8025517,4.617693,4.696918,4.5724216,4.496969,4.715781,5.1534057,5.3986263,5.3986263,5.3910813,5.4778514,5.5004873,5.0251365,4.8930945,4.8440504,4.7950063,4.772371,4.9157305,4.9459114,5.089271,5.198677,5.281675,5.5080323,5.994701,5.945657,6.1908774,6.900131,7.594294,7.533932,7.5490227,8.031919,9.020347,10.212496,10.095545,10.216269,10.152134,9.752235,9.110889,8.60913,8.552541,8.601585,8.771353,9.435335,11.09529,11.627231,11.461235,11.148107,11.32542,11.548005,11.778135,11.487643,10.861387,10.808571,10.461489,10.303039,10.499215,11.121698,12.117672,14.943368,18.776354,18.8254,16.90136,21.398329,23.450638,24.024076,24.48811,24.367384,21.334194,9.114662,3.6254926,1.7919968,1.3166461,0.70170826,1.7052265,1.4222796,0.94315624,0.694163,0.4376245,0.452715,0.26408374,0.09808825,0.041498873,0.06413463,0.23013012,0.7205714,1.3468271,1.6825907,1.0601076,2.3692086,1.6071383,0.56212115,0.071679875,0.0150905,0.0150905,0.00754525,0.0,0.0,0.00754525,0.03772625,0.041498873,0.0452715,0.06790725,0.08677038,0.24899325,0.2263575,0.34330887,0.663982,0.9997456,0.543258,0.3055826,0.30935526,0.4376245,0.41121614,0.36971724,0.24899325,0.48666862,0.86770374,0.51684964,0.44894236,0.35839936,0.5319401,0.875249,0.9205205,1.599593,1.8561316,1.9391292,1.9127209,1.6712729,1.4373702,1.1204696,0.8865669,0.94315624,1.5618668,2.1088974,2.4899325,2.1805773,1.6524098,2.3465726,2.6672459,3.7650797,4.406426,4.644101,5.832478,7.914967,8.043237,7.8432875,7.911195,7.8206515,7.911195,7.3792543,7.5037513,7.9941926,7.001992,7.8017883,8.167733,8.114917,7.7602897,7.3377557,7.5565677,7.6508837,7.5905213,7.805561,9.159933,10.3634,10.985884,12.132762,13.468271,13.226823,13.739901,13.894578,13.573905,12.898605,12.253486,12.626976,12.615658,13.373956,14.690601,15.022593,15.067864,14.852824,14.434063,14.037937,14.030393,12.3893,11.932813,12.091263,12.355347,12.279895,12.079946,11.710228,11.9064045,12.808062,13.947394,14.154889,13.9888935,14.211478,14.728328,14.603831,14.5283785,15.460217,16.576914,17.67852,19.206434,19.772327,18.851807,17.112627,15.403628,14.747191,15.792209,17.37671,18.678267,19.25925,19.055529,19.549744,20.85507,21.964222,22.288668,21.681276,20.48158,19.225298,18.052011,17.723793,19.591242,19.964731,20.37972,19.595015,17.844517,16.84477,17.025856,17.584206,18.72731,20.043957,20.504217,19.817598,19.821371,20.48158,21.119154,20.421219,18.399092,16.837225,16.260014,16.833452,18.376457,19.54597,20.055275,19.953413,19.353567,18.421728,18.448135,18.470772,18.576405,18.885761,19.557287,20.258997,20.907888,21.964222,23.288414,24.137255,23.495909,22.303759,20.839981,19.58747,19.25925,18.568861,19.338476,20.700394,22.107582,23.32614,23.32614,22.42071,20.934296,20.051502,21.798227,21.326649,20.647577,20.564579,20.82489,20.100546,21.692595,21.900087,21.817091,22.277351,23.835445,16.874952,14.517061,12.909923,10.370946,7.3905725,6.0324273,4.727099,5.6363015,8.103599,8.661947,9.548513,10.47658,11.812089,13.185325,13.4644985,14.441608,15.490398,15.554533,14.305794,12.128989,10.782163,10.7557535,11.514051,12.604341,13.645585,14.3095665,14.302021,14.260523,14.452927,14.777372,15.792209,15.596032,14.252977,12.340257,10.948157,9.310839,8.597813,8.348819,8.171506,7.7338815,7.462252,7.515069,7.6810646,7.835742,7.9451485,8.7751255,9.073163,9.076936,9.137298,9.710737,9.529651,9.688101,10.038955,10.657665,11.819634,8.175279,6.5568223,6.1342883,6.349328,6.8963585,7.9828744,8.145098,7.786698,7.654656,8.827943,8.054554,6.9491754,5.934339,5.409944,5.745708,5.6589375,5.96452,6.3531003,7.3151197,10.152134,8.669493,8.028146,7.356619,6.692637,6.990674,6.0324273,5.6891184,5.0854983,4.6856003,6.2927384,6.8699503,8.099826,8.5563135,8.107371,7.9225125,7.2283497,6.8963585,6.537959,6.2135134,6.4134626,6.25124,6.488915,6.790725,6.937857,6.8133607,7.352846,7.2887115,7.1378064,7.0887623,7.001992,6.2851934,6.092789,6.458734,6.9793563,6.809588,6.2323766,6.477597,6.6247296,6.5228686,6.8058157,8.29223,9.295748,9.676784,9.420244,8.654402,8.465771,8.405409,8.424272,8.563859,8.922258,8.401636,7.7376537,7.515069,7.7338815,7.8017883,7.1264887,6.6586833,6.6247296,6.9227667,7.118943,6.911449,6.983129,7.5112963,8.488406,9.710737,10.585986,9.556059,8.333729,8.069645,9.352338,9.065618,8.235641,7.8734684,8.107371,8.156415,7.2698483,7.0057645,6.4247804,5.583485,5.5193505,6.349328,6.439871,6.7944975,7.673519,8.586494,8.963757,9.193887,9.084481,8.677037,8.280911,7.7942433,7.7904706,7.858378,7.828197,7.752744,7.7187905,6.8359966,5.828706,4.991183,4.22534,4.217795,4.983638,5.1269975,4.6856003,5.1269975,6.5756855,7.432071,7.586749,7.405663,7.7225633,7.858378,7.533932,7.756517,8.439363,8.405409,8.314865,8.677037,8.9788475,9.2844305,10.220041,10.785934,11.710228,12.325166,12.400619,12.162943,11.69891,11.3971,10.423763,9.0543,8.68081,13.3626375,12.155397,9.378746,7.2623034,5.9494295,6.8133607,7.786698,8.480861,8.869441,9.276885,10.435081,10.8576145,10.604849,10.008774,9.688101,9.49947,9.420244,9.986138,10.929295,11.204697,11.725319,11.657412,11.879996,12.453435,12.638294,11.834724,12.00072,12.408164,12.626976,12.498707,11.283921,11.495189,12.238396,12.842015,12.864652,12.683565,13.664448,13.743673,13.045737,13.909668,19.889278,14.1926155,7.6810646,5.0213637,4.696918,8.677037,9.408927,9.310839,8.82417,6.4210076,7.567886,6.8661776,5.696664,5.4665337,7.6093845,7.2358947,7.0284004,8.22055,10.103089,10.020092,8.529905,6.7869525,5.5570765,5.553304,7.443389,7.039718,5.5683947,4.504514,4.466788,5.2250857,5.5495315,6.749226,7.273621,6.8246784,6.3455553,6.0814714,6.1418333,6.5266414,7.17176,7.9262853,7.5226145,7.0887623,6.439871,5.583485,4.749735,4.5233774,4.5724216,5.0553174,5.783434,6.228604,6.7756343,6.7454534,6.5040054,6.466279,7.1076255,7.183078,6.9265394,6.9491754,6.9491754,5.7079816,5.3344917,5.9117036,6.368191,6.4436436,6.688864,6.9189944,7.0963078,7.020855,6.8435416,7.0585814,7.533932,7.986647,7.986647,7.7904706,8.329956,9.06939,9.756008,10.446399,10.733118,9.752235,9.5183325,8.714764,8.039464,7.9225125,8.529905,8.4544525,8.386545,8.065872,7.6207023,7.5829763,7.488661,6.851087,6.5228686,6.8359966,7.5716586,7.333983,7.7225633,7.8244243,7.383027,6.7756343,6.4021444,5.8664317,5.617439,5.696664,5.73439,5.987156,6.1606965,5.934339,5.3382645,4.7648253,4.346064,4.38379,4.478106,4.4630156,4.4101987,5.4212623,5.3194013,4.9459114,4.738417,4.719554,5.43258,5.6476197,5.7872066,6.096562,6.6850915,6.379509,5.934339,5.1571784,4.29702,4.0480266,4.7006907,4.8365054,4.8063245,4.8100967,4.908185,5.50426,5.1156793,4.3121104,3.5236318,3.0407357,3.7537618,4.2630663,4.719554,5.05909,4.9987283,5.0138187,5.4891696,6.066381,6.730363,7.805561,8.375228,8.371455,8.473316,8.646856,8.122461,8.080963,7.937603,7.7150183,7.515069,7.5263867,7.115171,6.8397694,6.851087,7.0774446,7.1981683,7.5226145,8.356364,8.514814,8.050782,8.243186,4.644101,4.3385186,4.0970707,3.874486,3.821669,4.285702,4.38379,4.353609,4.5724216,4.9723196,5.0666356,5.3646727,5.613666,5.7004366,5.515578,4.957229,5.142088,5.240176,5.292993,5.270357,5.093044,5.1345425,5.1798143,5.3080835,5.5004873,5.6325293,5.7306175,5.670255,5.975838,6.719045,7.5075235,7.273621,7.6207023,8.526133,9.80128,11.102836,11.283921,11.11038,10.597303,9.733373,8.480861,7.986647,8.09228,8.511042,9.009028,9.405154,10.303039,10.774617,10.676529,10.306811,10.401127,10.978339,10.899114,10.38981,9.58624,8.529905,8.60913,9.261794,9.895596,10.695392,12.657157,15.950659,19.693102,20.108091,18.863125,23.065828,23.473272,20.647577,17.538933,14.769827,10.63503,4.146115,1.1091517,0.10940613,0.02263575,0.011317875,0.071679875,0.049044125,0.0150905,0.003772625,0.011317875,0.018863125,0.00754525,0.0,0.0,0.0,0.03772625,0.38103512,1.1355602,1.8938577,1.7165444,1.4713237,1.4109617,0.94315624,0.20372175,0.03772625,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.12826926,0.17354076,0.21881226,0.30935526,0.4678055,0.73188925,0.6375736,0.7054809,0.94692886,0.875249,0.9016574,0.5696664,0.7469798,1.2751472,1.0148361,0.7922512,0.5394854,0.35839936,0.40367088,0.8639311,1.6071383,1.6524098,1.4335974,1.2940104,1.5052774,1.1883769,0.8224323,0.66775465,1.0299267,2.2484846,2.4220252,2.3277097,2.022127,1.8221779,2.323937,2.9086938,3.9499383,5.028909,6.115425,7.564113,7.858378,8.122461,8.624221,9.14107,8.990166,9.027891,8.243186,7.8131065,7.748972,6.8699503,7.164215,8.52236,9.137298,8.695901,8.375228,8.484633,8.326183,8.329956,8.597813,8.892077,9.64283,10.627484,12.272349,13.849306,13.494679,14.70192,14.268067,13.72481,13.494679,12.898605,13.324911,13.702174,14.196388,14.947141,16.06761,16.188334,16.603323,16.791954,16.358103,15.0376835,13.166461,12.30253,12.128989,12.249713,12.178034,12.204442,12.004493,11.838497,12.102581,13.313594,13.158916,13.336229,14.219024,15.181043,14.618922,14.883006,15.437581,16.25624,17.40312,19.01403,19.783646,19.48561,17.908651,15.62244,13.996439,15.252723,16.991903,18.576405,19.598787,19.893051,20.115637,21.477554,22.696112,23.26955,23.4695,22.266033,20.700394,19.628967,19.591242,20.802254,20.29295,20.104319,19.300749,17.855835,16.65614,16.724047,17.618158,18.421728,18.949896,19.757236,19.406384,18.666948,18.700903,19.417702,19.4592,18.13878,16.516552,15.430037,15.384765,16.520325,17.87847,19.01403,19.527107,19.372429,18.832945,18.7839,18.202915,18.48209,19.7761,20.987112,22.10381,23.43932,25.054003,26.551735,27.07613,25.570852,23.982576,22.152855,20.557034,20.285404,19.349794,19.093256,20.22127,22.326395,23.869398,24.008986,22.948877,21.19838,19.91946,20.930523,20.160908,19.791191,19.74592,19.625195,18.69713,20.492899,21.915178,22.948877,23.94485,25.589716,17.316349,14.762281,13.483362,10.906659,6.330465,5.9494295,3.874486,4.5196047,7.6697464,8.499724,9.446653,9.680555,10.336992,11.351829,11.45369,12.577931,14.464244,16.26756,16.995676,15.513034,12.46098,11.351829,11.744182,12.755245,13.068373,13.985121,13.95494,13.59654,13.43809,13.902123,15.011275,14.928277,13.690856,12.034674,11.363147,9.763554,8.89585,8.590267,8.36391,7.4509344,6.983129,6.8435416,6.7341356,6.760544,7.443389,8.499724,8.98262,9.046755,8.959985,9.114662,9.416472,9.918231,10.208723,9.673011,7.492433,7.250985,6.255012,5.7494807,5.938112,5.9909286,7.2472124,7.7037,7.888559,7.937603,7.586749,7.1038527,6.5266414,5.87775,5.511805,6.1041074,6.515323,6.673774,6.7039547,6.670001,6.571913,8.616675,8.858124,8.118689,7.2358947,7.0774446,6.5040054,5.794752,5.160951,5.353355,7.6886096,7.111398,8.428044,8.937348,8.096053,7.5112963,6.7114997,6.515323,6.25124,5.855114,5.855114,5.9305663,5.462761,5.1269975,5.240176,5.745708,6.488915,6.6360474,6.688864,6.752999,6.537959,5.5495315,5.100589,5.4778514,6.2814207,6.428553,5.696664,5.7796617,5.847569,5.726845,5.8928404,6.771862,7.643338,8.114917,8.107371,7.8508325,8.152642,8.224322,8.488406,8.8769865,8.805306,8.197914,8.175279,8.197914,8.07719,8.00551,7.541477,6.741681,6.519096,6.8737226,6.858632,6.6662283,6.651138,7.1038527,8.058327,9.273112,9.635284,8.918486,7.997965,7.6207023,8.409182,8.4544525,8.567632,8.231868,7.654656,7.752744,6.2135134,6.1606965,6.0626082,5.455216,4.927048,5.594803,6.33801,7.394345,8.488406,8.820397,7.9300575,8.22055,8.367682,8.058327,7.9791017,7.91874,7.654656,7.8734684,8.428044,8.348819,8.073418,6.7567716,5.4891696,4.8553686,4.930821,4.4215164,5.1571784,5.5193505,5.2892203,5.66271,6.9567204,7.8961043,7.8696957,7.0963078,6.590776,7.2358947,6.9680386,6.934085,7.492433,8.197914,7.9828744,7.9451485,8.228095,8.771353,9.318384,10.506761,11.996947,12.283667,11.714001,12.491161,12.185578,12.2119875,11.680047,10.212496,7.9791017,8.303548,9.612649,10.174769,9.424017,7.9451485,8.296002,8.571404,8.480861,8.179051,8.27714,9.563604,10.457717,10.612394,10.148361,9.654147,9.597558,9.556059,10.1294985,11.042474,11.121698,11.608367,11.951676,12.189351,12.377983,12.596795,12.404391,12.283667,12.242168,12.279895,12.377983,11.355601,11.495189,12.577931,13.607859,12.811834,13.95494,15.313085,15.901614,15.539442,14.84528,13.200415,8.75249,7.5829763,8.590267,3.5047686,7.2660756,9.688101,11.653639,11.54046,5.198677,7.1868505,7.175533,6.439871,6.3116016,8.175279,7.3792543,6.7869525,7.6207023,9.088254,8.360137,6.8925858,5.9230213,5.0854983,4.9760923,7.1264887,7.515069,6.3945994,5.281675,5.1269975,6.3153744,6.719045,7.2698483,7.6018395,7.5716586,7.273621,6.628502,6.7341356,7.0246277,7.2472124,7.4584794,7.515069,6.858632,5.9909286,5.353355,5.323174,4.6742826,4.606375,4.9232755,5.3080835,5.3156285,6.2361493,6.477597,6.319147,6.2361493,6.8699503,7.1378064,6.7869525,6.722818,6.8661776,6.156924,5.8664317,6.2323766,6.156924,5.6551647,5.885295,6.4926877,6.617184,6.5832305,6.609639,6.820906,7.2887115,7.7716074,7.3075747,6.549277,7.786698,8.89585,9.831461,10.359629,10.310584,9.574923,10.023865,9.103344,8.262049,8.103599,8.375228,8.409182,8.616675,8.084735,6.983129,6.5568223,6.9454026,6.8133607,7.001992,7.884786,9.371201,8.367682,8.254503,8.548768,8.586494,7.515069,6.7039547,6.085244,5.9984736,6.25124,6.1078796,5.481624,5.379763,5.4476705,5.353355,4.7610526,4.2328854,4.266839,4.5007415,4.5950575,4.255521,4.768598,4.991183,5.0854983,5.191132,5.413717,5.764571,5.511805,5.300538,5.6400743,6.907676,6.6020937,6.296511,5.2967653,4.006528,3.9122121,5.0251365,5.2967653,4.9685473,4.5120597,4.6214657,5.028909,4.376245,3.651901,3.3425457,3.4142256,3.9763467,4.247976,4.738417,5.3344917,5.27413,4.5837393,4.7308717,5.160951,5.836251,7.2472124,8.20546,8.054554,8.22055,8.643084,7.798016,7.492433,7.5527954,7.515069,7.3377557,7.4018903,7.6848373,7.6886096,7.322665,6.907676,7.1793056,7.1679873,8.088508,8.684583,8.695901,8.873214,4.1197066,3.863168,3.7462165,3.7990334,3.9197574,3.8443048,4.1989317,4.195159,4.104616,4.0895257,4.2102494,4.689373,4.870459,5.2967653,5.8098426,5.553304,5.7494807,5.73439,5.6476197,5.458988,4.961002,4.8742313,5.0251365,5.4288073,5.80607,5.583485,5.0968165,5.534441,6.379509,7.3113475,8.179051,8.424272,8.503497,8.729855,9.382519,10.710483,10.944386,10.56335,9.752235,8.737399,7.798016,7.6131573,8.024373,8.586494,9.246704,10.344538,10.33322,10.182315,9.963503,9.654147,9.156161,9.948412,9.718282,9.540969,9.288202,7.6131573,8.835487,9.861642,10.310584,11.544232,16.708956,17.757746,18.002966,18.101055,18.4255,19.074392,16.180788,11.944131,7.9489207,4.9119577,2.6408374,1.1996948,0.392353,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.02263575,0.00754525,0.0,0.0,0.0,0.00754525,0.271629,0.9808825,2.2899833,2.3390274,2.0183544,1.3053282,0.47535074,0.120724,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.03772625,0.090543,0.18485862,0.38103512,1.0789708,1.3241913,1.7014539,2.0108092,1.267602,1.388326,0.84129536,0.8601585,1.3166461,0.73188925,0.36594462,0.8526133,1.0450171,0.875249,1.327964,0.8526133,0.94315624,0.98465514,0.88279426,1.0525624,0.94315624,1.116697,1.569412,2.2258487,2.9464202,1.5656394,1.2298758,1.448688,1.7769064,1.7995421,2.033445,3.3350005,5.6287565,7.858378,7.9791017,8.907167,8.4544525,8.850578,10.076681,9.857869,8.918486,8.66572,8.409182,7.699928,6.3342376,5.455216,6.205968,7.383027,8.09228,7.752744,6.9454026,7.677292,9.039209,10.355856,11.200924,10.016319,9.865415,11.857361,14.543469,13.947394,14.4114275,13.298503,12.830698,13.521088,14.2077055,14.864142,14.671739,14.460471,14.735873,15.701665,14.8339615,15.196134,16.018566,16.358103,15.07541,14.747191,13.849306,13.20796,12.679792,11.155652,11.227332,11.604594,11.857361,12.2119875,13.521088,12.992921,13.185325,13.947394,14.581196,13.822898,13.8870325,14.102073,15.316857,17.463482,19.57615,19.844007,19.270569,18.65563,17.912424,16.0827,15.482853,16.26756,17.399347,18.500954,19.866644,21.624687,23.069601,23.254461,23.005466,24.94837,24.05803,23.733583,24.484337,25.548216,24.903097,21.337967,20.100546,19.68933,18.938578,16.999449,16.852316,17.172989,17.380484,17.425755,17.7917,19.123436,18.742401,17.599297,16.675003,16.969267,16.822134,17.086218,16.524097,15.656394,16.754227,17.584206,18.104828,18.312323,18.406637,18.7839,19.466745,19.24416,19.670467,20.99843,22.171717,23.356321,24.97855,26.07261,26.295197,25.940569,25.499172,24.118391,22.598024,21.651094,21.896315,21.420965,20.11941,19.979822,21.221016,22.307531,22.699884,23.126192,22.01704,19.553514,17.686066,17.73511,18.542452,19.123436,19.236614,19.395065,20.55326,20.979568,21.768045,24.00144,28.762493,18.251959,14.079436,10.691619,7.0510364,6.620957,5.5004873,4.485651,4.878004,6.571913,8.073418,9.34102,8.688355,8.537451,9.488152,10.329447,11.012292,12.989148,15.728074,18.319866,19.455427,16.403374,13.837989,12.89106,12.970284,11.747954,12.67602,13.283413,13.230596,12.770335,12.755245,13.268322,13.234368,12.577931,11.657412,11.231105,10.155907,9.5032425,9.137298,8.718536,7.707473,7.1302614,6.7680893,6.587003,6.809588,7.91874,8.420499,8.360137,8.167733,7.9300575,7.432071,10.593531,11.729091,10.86516,8.89585,7.6131573,4.745962,3.7084904,4.4705606,5.73439,4.927048,5.9909286,6.7152724,7.8810134,8.710991,6.8661776,5.96452,5.4363527,5.198677,5.149633,5.1873593,4.8968673,5.1043615,5.745708,6.609639,7.352846,7.854605,9.050528,9.718282,8.846806,5.66271,9.092027,8.484633,7.3792543,7.5527954,9.016574,8.726082,8.22055,7.598067,6.971811,6.485142,5.4703064,5.6400743,6.126743,6.368191,6.089017,6.5040054,6.488915,5.7909794,4.7836885,4.4403796,4.587512,5.1647234,5.4740787,5.2552667,4.67051,4.8629136,4.8138695,4.647874,4.485651,4.425289,4.6327834,4.6856003,4.587512,4.5120597,4.8063245,5.6853456,6.5568223,6.9152217,6.900131,7.277394,7.8998766,8.001738,8.379,8.926031,8.620448,8.167733,8.495952,8.793989,8.726082,8.409182,8.103599,7.1566696,6.6360474,6.7379084,6.7756343,6.934085,6.617184,6.56814,7.122716,8.209232,6.85486,6.828451,7.914967,9.216523,9.156161,8.201687,7.809334,7.432071,7.1076255,7.462252,6.009792,5.7381625,6.1041074,6.4436436,5.96452,5.9796104,5.7079816,6.3116016,7.854605,9.307066,8.122461,7.435844,7.1038527,7.149124,7.7376537,8.016829,7.6093845,7.9413757,8.91094,8.91094,9.046755,7.7150183,6.1644692,5.2628117,5.492942,4.7006907,5.4174895,5.9532022,5.7607985,5.43258,6.628502,7.2094865,7.039718,6.432326,6.1644692,5.9192486,6.3455553,6.5530496,6.4511886,6.7454534,6.7944975,7.4471617,8.495952,9.733373,10.940613,11.332966,12.004493,11.846043,10.978339,10.7557535,11.332966,12.068627,12.936331,13.264549,11.763044,9.578695,10.223814,10.838752,10.861387,12.0082655,10.751981,9.688101,9.125979,9.06939,9.216523,8.91094,10.18986,10.940613,10.506761,9.688101,9.846551,9.6051035,10.140816,11.351829,11.84227,11.438599,11.759273,12.019584,12.0233555,12.147853,12.400619,11.84227,10.982111,10.193633,9.703192,10.20495,9.635284,10.340765,11.9064045,11.140562,13.837989,14.520834,16.58446,19.240387,17.53139,18.142553,17.663431,18.376457,16.746683,3.4179983,4.406426,10.11818,15.147089,15.62244,9.201432,7.4811153,8.284684,8.631766,8.213005,9.382519,8.382772,7.914967,9.352338,11.793225,12.0233555,9.763554,8.111144,6.4210076,5.3194013,6.700182,6.749226,5.6778007,5.0854983,5.621211,6.9869013,7.8810134,8.122461,8.137552,8.00551,7.432071,6.1720147,6.224831,6.5228686,6.907676,8.118689,7.960239,6.730363,5.6853456,5.4703064,6.1041074,5.2967653,5.1798143,5.081726,4.851596,4.851596,5.7419353,6.085244,5.8664317,5.4665337,5.66271,6.1720147,5.934339,6.368191,7.4735703,7.828197,7.352846,6.620957,5.624984,4.8327327,5.1873593,7.1038527,7.1981683,6.2663302,5.455216,6.270103,6.94163,7.092535,6.8359966,6.8473144,8.360137,9.009028,9.242931,9.74469,10.340765,10.023865,9.597558,9.114662,8.797762,8.729855,8.850578,8.692128,8.2507305,7.1264887,5.8626595,5.934339,6.9982195,7.7678347,8.216777,8.503497,8.956212,8.284684,7.4018903,7.586749,8.409182,7.7376537,7.039718,6.730363,6.405917,6.0211096,5.873977,5.4363527,5.406172,5.4212623,5.247721,4.821415,4.38379,4.5196047,4.776143,4.9157305,4.927048,5.9305663,6.8661776,7.2698483,6.8661776,5.583485,4.8402777,4.534695,4.7535076,5.3194013,5.783434,6.2097406,6.198423,5.3609,4.217795,4.1800685,5.2552667,5.4967146,5.0515447,4.3385186,4.0593443,4.534695,4.6554193,4.606375,4.52715,4.5007415,4.2328854,4.5233774,5.05909,5.5797124,5.8588867,5.0553174,4.7610526,4.779916,5.149633,6.149379,7.3717093,7.1906233,7.232122,7.6282477,7.001992,6.5040054,6.4436436,6.7152724,7.01331,6.8058157,7.624475,8.194141,8.096053,7.5792036,7.567886,7.7150183,8.382772,9.110889,9.616421,9.812597,3.350091,3.3689542,3.572676,3.5651307,3.440634,3.7952607,3.9763467,4.0216184,3.9914372,3.9763467,4.13857,4.508287,4.772371,5.1081343,5.43258,5.4212623,5.2062225,5.1156793,5.349582,5.794752,6.043745,6.1644692,5.994701,5.828706,5.824933,6.0362,6.1720147,6.771862,7.364164,7.7716074,8.141325,8.084735,8.122461,8.367682,8.884532,9.688101,10.152134,9.989911,9.34102,8.465771,7.7602897,7.7037,8.296002,8.899622,9.35611,9.967276,10.054046,10.016319,9.635284,9.009028,8.5563135,9.261794,8.82417,8.213005,7.77538,7.2358947,8.028146,8.771353,9.8239155,11.917723,16.18456,16.090246,16.810818,17.708702,18.49718,19.232841,19.229069,15.143317,9.612649,4.847823,2.6144292,1.2826926,0.5357128,0.19240387,0.07922512,0.03772625,0.026408374,0.011317875,0.003772625,0.011317875,0.0,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.05281675,0.3055826,1.0072908,1.5731846,1.50905,1.1506506,0.7394345,0.41498876,0.19994913,0.094315626,0.0452715,0.02263575,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.14713238,0.08677038,0.033953626,0.060362,0.10186087,0.24899325,0.30181,0.38103512,0.452715,0.30181,0.35462674,0.38480774,0.66775465,1.0336993,0.86770374,0.5394854,0.8526133,1.2864652,1.3656902,0.65643674,0.43385187,0.77338815,0.845068,0.58098423,0.6752999,1.0412445,1.4826416,1.8599042,2.1013522,2.1881225,1.3958713,1.7995421,1.7391801,1.2034674,1.81086,2.9049213,3.5500402,5.1458607,7.484888,8.748717,9.393836,9.616421,9.4013815,9.092027,9.367428,8.967529,7.9828744,7.232122,6.8246784,6.1606965,7.118943,7.303802,7.567886,8.035691,8.09228,8.567632,9.574923,10.408672,10.95193,11.6875925,11.234878,11.54046,12.917468,14.452927,14.030393,14.136025,13.732355,13.856852,14.517061,14.694374,14.622695,15.746937,16.143063,15.565851,15.456445,14.377474,14.769827,15.592259,15.690348,13.792717,13.336229,12.857106,13.060828,13.611631,13.12119,13.27964,12.438345,11.872451,12.189351,13.347548,13.430545,14.1926155,14.747191,14.837734,14.86037,14.249205,14.339747,14.984866,16.22606,18.319866,18.881989,19.478064,19.942095,19.719511,17.87847,16.946632,17.040947,17.482344,18.244415,19.964731,21.70391,22.439573,22.526344,22.465982,22.933788,22.786655,25.080412,27.823109,28.660633,24.891779,19.636513,19.478064,20.69662,21.066338,19.817598,19.1423,18.85558,18.840488,18.949896,19.025349,19.263023,19.168707,18.21046,16.935314,16.991903,17.052265,16.97304,16.678776,16.309057,16.218515,17.184307,18.285913,19.338476,20.142044,20.48158,21.164427,21.058792,21.337967,22.122673,22.4773,21.941587,22.19058,22.46221,22.552752,22.816835,22.258488,21.688822,21.405874,21.187061,20.30804,20.157135,19.281887,18.915941,19.481836,20.587215,20.821117,20.29295,18.738628,16.897587,16.524097,16.165699,16.803272,18.331184,19.885506,19.859098,21.281378,21.900087,23.246916,25.19359,25.92925,14.747191,11.759273,9.937095,7.284939,6.8171334,6.1041074,5.553304,5.251494,5.451443,6.5832305,8.224322,8.254503,8.216777,8.869441,10.208723,11.155652,12.419481,13.93985,15.328176,15.878979,15.256495,15.388537,15.935568,16.052519,14.362384,14.18507,14.166207,14.1058445,13.943622,13.758763,13.419228,12.879742,12.245941,11.680047,11.389555,10.970794,10.518079,10.023865,9.35611,8.254503,7.2623034,6.771862,6.549277,6.6134114,7.2358947,7.8923316,8.231868,8.390318,8.284684,7.624475,12.925014,14.400109,14.034165,12.551523,9.446653,6.6850915,4.3196554,2.8596497,2.957738,5.3910813,4.708236,5.300538,6.119198,6.462507,5.975838,5.6476197,5.0439997,4.9044123,5.1458607,4.870459,4.5196047,4.406426,4.52715,5.2854476,7.515069,9.80128,11.34051,12.283667,11.408418,6.1116524,9.846551,10.989656,9.910686,7.84706,6.930312,9.129752,9.684328,9.050528,8.265821,8.99771,10.182315,8.66572,7.4509344,7.3000293,6.749226,6.4511886,6.541732,6.1720147,5.2665844,4.5120597,4.221567,4.4818783,4.851596,4.9232755,4.327201,4.436607,4.6742826,4.7912335,4.557331,3.802806,3.610402,3.6141748,3.7235808,3.9801195,4.538468,5.3684454,5.6098933,5.696664,5.832478,5.983383,6.881268,7.6282477,8.13378,8.4544525,8.790216,9.258021,9.352338,9.163706,8.858124,8.677037,8.156415,7.756517,7.3490734,6.930312,6.6058664,6.507778,6.0550632,5.772116,6.0324273,7.0510364,6.2021956,6.089017,6.6247296,7.4811153,8.09228,7.854605,7.0887623,6.802043,6.8963585,6.156924,6.089017,6.039973,6.2097406,6.4134626,6.0626082,6.5341864,7.1906233,7.213259,6.8397694,7.356619,6.677546,6.224831,6.417235,7.0284004,7.175533,6.760544,6.6020937,6.934085,7.6622014,8.326183,8.75249,7.8244243,6.6360474,5.8136153,5.5193505,5.87775,5.8626595,6.009792,6.228604,5.8211603,6.4436436,7.5905213,7.6207023,6.519096,5.907931,6.228604,7.0887623,7.8923316,8.36391,8.537451,8.137552,8.6581745,9.476834,10.299266,11.136789,11.400873,11.498961,11.3820095,11.151879,11.099063,11.272603,11.751727,12.253486,12.551523,12.434572,11.072655,10.484125,9.933322,9.616421,10.665211,11.057564,9.359882,8.809079,9.684328,9.314611,9.593785,10.733118,11.332966,11.23865,11.544232,11.604594,11.623458,12.061082,12.762791,12.940104,12.30253,11.559323,11.227332,11.261286,11.072655,10.887795,10.578441,9.993684,10.838752,16.697638,13.547497,10.63503,9.718282,11.174516,14.019074,12.351574,13.283413,15.128226,15.939341,13.517315,18.187824,20.089228,20.394812,17.395575,6.458734,5.5306683,7.8508325,14.947141,21.337967,14.535924,7.9715567,8.326183,9.231613,8.503497,8.152642,7.424526,7.1604424,9.042982,11.819634,11.329193,11.02361,7.798016,6.0022464,6.790725,8.137552,7.250985,6.5832305,6.2135134,6.1908774,6.560595,7.805561,8.360137,8.111144,7.5112963,7.6018395,6.7944975,6.5568223,6.6247296,7.0472636,8.179051,8.254503,7.0887623,6.2021956,5.987156,5.7117543,5.0251365,4.878004,4.817642,4.776143,5.05909,5.6476197,5.7607985,5.617439,5.5080323,5.772116,5.836251,5.511805,6.089017,7.352846,7.6093845,6.9869013,6.48137,5.704209,4.938366,5.1156793,6.326692,6.628502,6.300284,6.0512905,7.0170827,6.8963585,6.730363,6.398372,6.217286,6.971811,8.299775,9.035437,9.484379,9.608876,9.046755,8.89585,8.729855,8.748717,8.741172,8.09228,8.197914,8.028146,7.484888,6.9152217,7.1076255,8.258276,8.937348,8.827943,8.401636,8.918486,7.5263867,6.5455046,6.6624556,7.435844,7.273621,6.5568223,6.1305156,5.9230213,5.7607985,5.3609,5.379763,5.3646727,5.4778514,5.564622,5.1760416,4.9987283,5.028909,5.05909,5.221313,5.96452,6.7039547,7.6848373,7.877241,6.9227667,5.1345425,4.7308717,4.957229,5.2552667,5.4363527,5.6853456,6.5040054,6.187105,5.2552667,4.346064,4.1800685,4.45547,4.5837393,4.4743333,4.2291126,4.1310244,4.1310244,4.247976,4.496969,4.6856003,4.429062,4.696918,4.90064,5.036454,4.979865,4.4818783,3.9876647,3.9914372,4.293247,4.8440504,5.745708,6.673774,7.352846,7.7942433,7.798016,6.930312,6.7831798,6.700182,7.032173,7.5829763,7.6093845,7.8923316,8.465771,8.424272,7.9753294,8.473316,8.616675,9.016574,9.386291,9.7069645,10.227587,2.7841973,3.029418,3.2142766,3.2255943,3.1652324,3.3350005,3.4783602,3.6330378,3.7198083,3.7650797,3.9008942,4.1989317,4.3875628,4.5309224,4.659192,4.7346444,4.8138695,4.8742313,5.13077,5.5495315,5.8136153,5.802297,5.7872066,5.6400743,5.5268955,5.9003854,6.19465,6.809588,7.164215,7.254758,7.6395655,7.4811153,7.5301595,8.062099,8.89585,9.393836,9.88805,9.891823,9.654147,9.310839,8.869441,8.571404,8.756263,8.888305,8.971302,9.533423,9.65792,9.559832,9.129752,8.461998,7.8395147,8.171506,7.654656,7.1981683,7.164215,7.3717093,8.001738,9.175024,10.974566,13.166461,15.199906,15.23386,17.195625,18.572634,18.51227,17.833199,18.795218,15.894069,10.8576145,5.7306175,2.867195,1.478869,0.76207024,0.45648763,0.33953625,0.19994913,0.15845025,0.120724,0.06790725,0.011317875,0.0,0.011317875,0.011317875,0.018863125,0.03772625,0.03772625,0.03772625,0.018863125,0.00754525,0.1659955,0.79602385,1.6184561,1.5052774,1.3317367,1.2600567,0.754525,0.55457586,0.35839936,0.18863125,0.071679875,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.071679875,0.041498873,0.00754525,0.0150905,0.02263575,0.018863125,0.018863125,0.049044125,0.08299775,0.02263575,0.0452715,0.34330887,0.5696664,0.663982,0.83752275,0.5394854,0.8111144,0.97710985,0.845068,0.67152727,0.4979865,0.5093044,0.49044126,0.38480774,0.29426476,0.724344,1.4034165,1.7731338,1.6561824,1.267602,1.4034165,1.5882751,1.4335974,1.2864652,2.2560298,3.1425967,3.4896781,4.6516466,6.730363,8.567632,9.163706,9.812597,9.420244,8.2507305,7.937603,7.677292,7.326438,7.232122,7.3868,7.4094353,7.6848373,8.09228,8.420499,8.643084,8.948667,8.956212,9.235386,9.797507,10.506761,11.0613365,11.363147,12.276122,13.472044,14.460471,14.558559,15.060319,14.226569,13.815352,14.369928,15.211224,15.267814,15.875206,15.950659,15.460217,15.403628,14.950912,15.596032,16.437326,16.637276,15.414946,14.728328,14.219024,14.079436,14.245432,14.369928,14.539697,14.011529,13.894578,14.490653,15.290449,14.584969,14.807553,15.147089,15.135772,14.64533,14.479335,14.505743,14.988639,16.078928,17.814335,18.821627,19.791191,20.534397,20.77962,20.175999,18.919714,18.055782,18.014284,19.078165,21.398329,22.582933,22.684793,22.39053,22.100037,21.918951,22.066084,24.808783,28.173964,28.57009,20.787165,16.36942,18.391546,21.4436,22.790428,22.382984,21.737865,20.783392,20.017548,19.73083,20.010002,19.945868,19.293203,18.206688,17.165443,16.98813,17.595524,17.99542,18.18028,18.070873,17.512526,17.953922,19.564833,21.466236,22.869654,23.084692,22.828154,22.616886,22.647068,22.760246,22.450891,20.074137,18.923487,19.251705,20.50799,21.35683,20.938068,20.756983,20.919205,20.994658,19.994913,19.31584,18.580177,18.12369,18.248188,19.240387,19.108345,18.044466,16.837225,16.29774,17.28994,16.678776,17.452164,19.338476,21.292696,21.511507,22.714975,21.986858,21.4851,22.096264,23.409138,14.781145,11.61214,9.756008,7.6207023,6.1606965,5.3684454,5.7306175,6.0739264,5.96452,5.73439,7.3075747,8.058327,8.443134,9.0957985,10.846297,12.291212,13.358865,14.019074,14.351066,14.57365,15.23386,16.044973,16.52787,16.233604,14.750964,13.815352,13.336229,13.313594,13.573905,13.751218,13.555041,13.215506,12.792972,12.3289385,11.830952,10.974566,10.487898,10.099318,9.461743,8.152642,7.2396674,6.8737226,6.5945487,6.4511886,7.020855,7.91874,8.465771,8.8618965,8.9788475,8.333729,10.880251,13.106099,13.468271,11.84227,9.537196,7.4396167,8.7751255,7.835742,4.8855495,6.1418333,5.572167,6.138061,6.647365,6.907676,7.7112455,6.911449,6.488915,5.9230213,5.1345425,4.4894238,4.5460134,5.587258,6.2135134,6.307829,7.0510364,9.058073,11.480098,13.732355,13.573905,7.122716,10.86516,14.777372,14.245432,10.005001,8.14887,9.439108,7.9300575,6.888813,7.575431,9.242931,8.993938,8.122461,7.2962565,6.6058664,5.594803,5.028909,5.515578,5.80607,5.4288073,4.7044635,4.0404816,3.5424948,3.2482302,3.0897799,2.8785129,3.0671442,3.4481792,3.5651307,3.3425457,3.1350515,2.9351022,3.006782,3.097325,3.240685,3.7462165,4.689373,5.1798143,5.198677,4.9157305,4.689373,5.5382137,6.8774953,7.835742,8.235641,8.605357,9.001483,9.208978,9.190115,9.092027,9.246704,8.805306,8.284684,7.7150183,7.1868505,6.85486,6.2927384,5.7570257,5.50426,5.6891184,6.3644185,5.915476,5.8437963,5.824933,5.983383,6.911449,7.1604424,6.719045,6.643593,6.72659,5.5080323,6.0022464,6.0324273,6.0701537,6.319147,6.719045,6.560595,7.7112455,8.001738,7.303802,7.5263867,6.8359966,6.096562,6.1720147,6.903904,7.069899,6.3153744,6.4964604,7.3490734,8.265821,8.296002,8.477088,7.5301595,6.7756343,6.398372,5.458988,5.666483,5.4665337,5.715527,6.168242,5.4703064,6.432326,7.7150183,8.152642,7.454707,6.247467,6.72659,7.7112455,8.8618965,9.695646,9.601331,8.816625,9.344792,10.087999,10.61994,11.174516,11.042474,11.555551,12.208215,12.555296,12.219532,11.868678,12.064855,12.313848,12.396846,12.366665,11.732863,11.053791,10.386037,9.81637,9.450426,10.423763,8.7751255,7.877241,8.318638,7.8810134,8.793989,9.854096,10.63503,11.359374,12.894833,12.800517,13.102326,13.532406,13.781399,13.498452,13.079691,12.034674,11.449917,11.227332,10.087999,9.635284,9.786189,9.461743,10.378491,17.048492,17.097536,15.354584,12.3893,9.827688,10.336992,12.7477,13.8870325,15.422491,15.958203,11.038701,14.449154,20.26277,24.99364,22.884743,5.881522,6.6020937,7.0585814,14.969776,24.854053,18.029375,9.167479,8.084735,9.544742,10.510533,10.121953,8.175279,7.7225633,8.397863,8.903395,7.0246277,6.930312,5.9418845,5.881522,7.1076255,8.507269,7.779153,7.2170315,6.5341864,5.9003854,5.9494295,6.9944468,7.6584287,7.605612,7.175533,7.3868,6.8699503,6.752999,6.930312,7.303802,7.7904706,7.8017883,7.073672,6.5568223,6.3417826,5.643847,4.82896,4.436607,4.3649273,4.5912848,5.194905,5.2364035,5.2590394,5.247721,5.3344917,5.798525,5.696664,5.43258,5.847569,6.7077274,6.673774,6.1116524,6.1078796,6.009792,5.7004366,5.6098933,5.745708,6.19465,6.6058664,6.8737226,7.1566696,7.1264887,7.066127,6.8058157,6.5228686,6.7680893,8.058327,9.273112,9.552286,8.952439,8.439363,8.99771,8.854351,8.548768,8.186596,7.4207535,8.050782,8.299775,8.3525915,8.296002,8.114917,8.801534,9.175024,8.918486,8.36391,8.499724,7.2094865,6.5266414,6.5756855,7.0170827,7.0359454,6.2663302,5.8211603,5.696664,5.704209,5.4438977,5.7381625,5.6853456,5.704209,5.7796617,5.4665337,5.515578,5.481624,5.455216,5.6061206,6.1606965,6.598321,7.462252,7.54525,6.4964604,4.798779,4.9459114,5.4363527,5.764571,5.7494807,5.5495315,6.1078796,5.6778007,4.7044635,3.7801702,3.6481283,3.6481283,3.8707132,4.08198,4.2328854,4.425289,4.4931965,4.640329,4.7535076,4.719554,4.398881,4.5120597,4.5837393,4.6516466,4.6026025,4.1612053,3.6368105,3.5689032,3.863168,4.504514,5.534441,6.2663302,7.039718,7.4282985,7.2962565,6.7831798,7.039718,7.062354,7.405663,7.9828744,8.069645,7.8621507,8.088508,8.224322,8.299775,8.899622,8.929804,9.224068,9.6201935,9.940866,9.989911,2.293756,2.5427492,2.6710186,2.7841973,2.9200118,3.0671442,3.0671442,3.1954134,3.4142256,3.6330378,3.7047176,3.7914882,3.8971217,4.032936,4.164978,4.1800685,4.4101987,4.61392,4.847823,5.119452,5.3759904,5.2590394,5.191132,5.0175915,4.908185,5.353355,5.6023483,6.1305156,6.4210076,6.5002327,6.937857,7.1264887,7.183078,7.8319697,8.91094,9.382519,9.971047,10.0465,9.937095,9.789962,9.559832,8.809079,8.616675,8.495952,8.439363,8.937348,9.0807085,8.639311,8.186596,7.77538,6.9491754,7.1340337,7.0963078,7.122716,7.3981175,8.00551,9.092027,10.827434,13.249459,15.339493,15.022593,14.607604,16.463736,17.557796,17.391802,18.040693,17.41821,13.13628,8.224322,4.4441524,2.305074,1.418507,0.9620194,0.68661773,0.46026024,0.24522063,0.1961765,0.13958712,0.06790725,0.00754525,0.0,0.011317875,0.018863125,0.033953626,0.049044125,0.041498873,0.041498873,0.030181,0.0150905,0.11317875,0.52062225,1.1959221,1.1619685,1.1280149,1.2034674,0.875249,0.69039035,0.513077,0.3470815,0.20372175,0.08677038,0.041498873,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.071679875,0.15467763,0.071679875,0.030181,0.29426476,0.5055317,0.6187105,0.90920264,0.68661773,0.8186596,0.79602385,0.56589377,0.55457586,0.4376245,0.3961256,0.40367088,0.40367088,0.32067314,0.7884786,1.2864652,1.50905,1.4147344,1.2487389,1.7127718,1.6033657,1.5543215,1.9051756,2.6823363,3.0030096,3.5538127,4.3385186,5.330719,6.4436436,7.8131065,8.590267,8.461998,7.696155,7.149124,7.3188925,7.3453007,7.745199,8.439363,8.75249,8.858124,9.49947,9.6201935,9.322156,9.88805,9.552286,9.420244,9.861642,10.657665,10.993429,11.714001,12.653384,13.415455,13.9888935,14.7170105,15.192361,14.483108,13.743673,13.890805,15.562078,15.611122,15.531898,15.501716,15.433809,14.977322,15.0905,15.7657995,16.520325,16.886269,16.4411,15.584714,15.335721,15.165953,15.015047,15.290449,15.313085,14.977322,15.279131,16.192106,16.667458,15.207452,14.762281,14.928277,15.256495,15.279131,15.32063,15.331948,15.818617,16.833452,17.991648,19.04421,19.84778,20.7268,21.4436,21.224789,20.52308,19.398838,19.153618,20.300495,22.575388,23.518545,23.514772,22.854563,21.949133,21.360603,21.424738,22.805517,24.99364,25.03514,17.520071,14.215251,17.086218,20.515535,22.14531,22.862108,23.548725,22.541435,21.179516,20.300495,20.247679,20.089228,19.296976,18.297232,17.48989,17.252214,17.67852,18.395319,19.059301,19.312067,18.79899,18.738628,20.23636,22.352802,24.167437,24.812555,24.182526,23.673222,22.828154,21.617142,20.4514,18.470772,17.799244,18.980076,21.236107,22.447119,21.722775,20.994658,20.670212,20.560806,19.855326,18.606586,17.73511,17.071129,16.7995,17.4333,17.486116,16.946632,16.55428,16.984358,18.836716,18.795218,19.534653,21.092747,22.790428,23.246916,23.854307,21.952906,19.681786,18.746174,20.421219,16.459963,12.638294,10.140816,8.280911,4.4894238,4.0178456,5.036454,6.115425,6.2097406,4.666737,5.6815734,7.194396,8.273367,9.035437,10.676529,12.691111,13.894578,14.241659,14.037937,13.951167,14.905642,15.629986,15.860115,15.362129,13.932304,12.909923,12.543978,12.5326605,12.694883,12.943876,13.166461,13.347548,13.200415,12.728837,12.245941,11.321648,10.63503,10.099318,9.461743,8.27714,7.696155,7.435844,7.073672,6.790725,7.360391,8.544995,9.201432,9.220296,8.76758,8.296002,8.495952,10.782163,11.710228,10.623712,9.646602,6.092789,8.941121,9.4127,6.2399216,5.6589375,5.643847,6.224831,7.4396167,9.024119,10.397354,7.5037513,6.9793563,6.5455046,5.4288073,4.3686996,4.7572803,6.187105,7.3490734,7.726336,7.605612,7.496206,9.2995205,11.747954,12.291212,7.092535,10.423763,15.882751,16.497688,11.872451,8.201687,8.756263,6.4247804,5.523123,6.990674,8.382772,7.273621,6.56814,5.828706,5.062863,4.689373,4.2064767,4.881777,5.409944,5.243949,4.640329,3.904667,2.9954643,2.1881225,1.7052265,1.7240896,1.9127209,2.214531,2.2371666,2.0598533,2.2371666,2.1843498,2.335255,2.425798,2.4710693,2.7653341,3.500996,4.3649273,4.4441524,3.802806,3.4934506,4.1498876,5.6551647,7.0359454,7.8621507,8.239413,8.099826,8.461998,8.873214,9.148616,9.374973,9.265567,8.469543,7.647111,7.1302614,6.903904,6.2399216,5.772116,5.583485,5.6891184,6.017337,5.5985756,5.5797124,5.4438977,5.3609,6.1908774,6.432326,6.2814207,6.360646,6.488915,5.666483,6.48137,6.458734,6.217286,6.330465,7.3113475,6.9567204,8.126234,8.492179,7.816879,7.99042,7.424526,6.598321,6.507778,7.073672,7.145352,6.722818,6.9189944,7.5905213,8.243186,8.065872,8.152642,7.2094865,6.719045,6.6662283,5.5570765,5.2665844,5.119452,5.587258,6.2021956,5.5759397,6.398372,7.2358947,7.8961043,7.964011,6.790725,7.039718,7.960239,9.084481,9.95973,10.163452,9.129752,9.544742,10.020092,10.212496,10.816116,10.465261,11.59705,13.079691,13.898351,13.158916,12.494934,12.683565,12.970284,12.909923,12.336484,12.004493,12.106354,11.706455,10.427535,8.473316,8.677037,7.7602897,7.2887115,7.435844,6.971811,7.964011,9.34102,10.657665,11.955449,13.773854,13.472044,13.702174,14.132254,14.34352,13.853079,13.936077,12.709973,11.6875925,11.000975,9.416472,9.148616,9.597558,9.578695,9.929549,13.521088,17.670975,16.886269,13.630494,9.639057,5.9117036,12.261031,13.011784,14.241659,15.362129,9.122208,10.559577,18.912169,27.642023,27.113855,4.5912848,10.001229,7.673519,12.585477,22.839472,19.647831,10.438853,7.5263867,8.537451,10.79348,11.317875,8.345046,7.643338,7.322665,6.228604,3.9386206,4.014073,5.0025005,6.0248823,6.8699503,8.001738,7.9338303,7.4735703,6.719045,5.983383,5.8173876,6.379509,6.9755836,7.1302614,6.881268,6.7643166,6.488915,6.477597,6.752999,7.1038527,7.0585814,6.9265394,6.485142,6.2323766,6.0814714,5.3759904,4.496969,3.8782585,3.893349,4.5233774,5.342037,4.949684,4.9157305,4.90064,4.991183,5.7117543,5.6891184,5.409944,5.6589375,6.255012,6.058836,5.73439,5.945657,6.0776987,5.994701,6.0248823,5.6589375,6.1908774,6.9227667,7.375482,7.273621,7.224577,7.122716,6.9944468,6.907676,6.9567204,7.9489207,9.393836,9.491924,8.405409,8.254503,8.963757,8.907167,8.43559,7.8206515,7.2358947,8.213005,8.737399,9.06939,9.1825695,8.748717,8.778898,8.990166,9.001483,8.748717,8.518587,7.3151197,6.643593,6.477597,6.598321,6.609639,6.228604,5.881522,5.7494807,5.7494807,5.5306683,5.59103,5.6778007,5.855114,6.006019,5.855114,5.881522,5.7306175,5.7494807,5.9796104,6.138061,6.2851934,7.062354,7.360391,6.790725,5.6778007,5.7306175,5.8664317,6.0814714,6.1418333,5.6061206,5.4401255,4.9534564,4.217795,3.5123138,3.308592,3.270866,3.640583,4.074435,4.4931965,5.0779533,5.2137675,5.2665844,5.0741806,4.719554,4.5120597,4.5120597,4.738417,4.7648253,4.478106,4.0480266,3.399135,3.410453,3.7348988,4.285702,5.2326307,5.983383,6.530414,6.72659,6.590776,6.300284,6.72659,7.1000805,7.5263867,7.911195,7.9526935,8.0206,8.054554,8.213005,8.507269,8.793989,8.6581745,9.148616,9.714509,9.978593,9.7296,1.9391292,2.052308,2.191895,2.354118,2.5767028,2.9501927,2.8596497,2.897376,3.169005,3.5424948,3.663219,3.4934506,3.531177,3.772625,4.032936,3.9348478,4.063117,4.349837,4.659192,4.9345937,5.194905,5.2099953,4.8666863,4.534695,4.515832,5.040227,5.2779026,5.6891184,6.0324273,6.2361493,6.428553,7.1566696,7.3075747,7.779153,8.631766,9.0807085,9.827688,9.948412,9.691874,9.2995205,9.020347,7.8998766,7.8131065,7.9526935,8.001738,8.182823,8.288457,7.515069,7.1000805,7.092535,6.360646,6.8435416,7.492433,7.854605,8.114917,9.073163,10.902886,12.800517,15.509261,17.712475,16.01102,14.441608,14.852824,15.211224,15.648849,18.448135,15.505488,8.405409,3.0935526,1.4034165,1.0412445,0.9808825,0.9205205,0.6828451,0.32444575,0.12826926,0.46026024,0.2678564,0.05281675,0.00754525,0.003772625,0.011317875,0.02263575,0.026408374,0.026408374,0.02263575,0.0150905,0.018863125,0.0150905,0.0,0.0,0.2678564,0.44516975,0.55080324,0.6149379,0.694163,0.5055317,0.4376245,0.39989826,0.32444575,0.15467763,0.08299775,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.08299775,0.1961765,0.15467763,0.060362,0.124496624,0.43385187,0.8262049,0.91297525,0.7696155,0.7054809,0.7432071,0.69793564,0.16976812,0.32821837,0.49044126,0.5885295,0.6073926,0.5998474,1.1883769,1.3468271,1.3732355,1.5241405,1.9994912,1.9730829,1.8825399,2.1541688,2.6898816,2.8558772,2.7351532,3.6783094,4.1536603,3.92353,4.0404816,5.9117036,6.5530496,6.8963585,7.2094865,7.092535,8.171506,7.997965,8.307321,9.25425,9.4127,10.087999,10.782163,10.650121,10.084227,10.70671,10.838752,11.080199,11.393328,11.747954,12.113899,12.958967,13.147598,13.057055,13.219278,14.335975,14.260523,14.475562,14.158662,13.924759,15.82239,15.573396,15.165953,15.214996,15.358356,14.234114,14.479335,14.766054,15.143317,15.430037,15.245177,14.7736,15.207452,15.675257,15.863888,16.033657,16.060064,15.573396,15.70921,16.52787,17.01831,15.961976,15.294222,15.192361,15.724301,16.848543,16.614641,16.750456,17.350302,18.168962,18.614132,19.496925,19.90437,20.673985,21.481327,20.817345,21.23988,20.760756,20.65135,21.45869,22.997923,23.97126,24.242887,23.48459,22.092491,21.19838,20.794708,20.247679,20.406128,20.274086,17.040947,14.490653,16.03743,17.999193,19.180025,20.858843,23.32614,23.250689,22.14531,20.934296,19.94964,19.58747,19.191343,18.557543,17.844517,17.57666,17.127718,17.674747,18.632996,19.364883,19.1423,18.65563,19.308294,20.900343,22.918697,24.556017,24.548471,24.005213,22.326395,19.851553,17.844517,17.761518,18.693357,20.790936,23.235598,24.261751,23.092237,21.420965,20.232588,19.708193,19.240387,17.931286,16.731592,15.675257,15.086727,15.565851,16.490145,17.067356,17.399347,18.052011,20.059048,20.719257,20.987112,21.575642,22.53389,23.254461,23.68454,21.692595,19.032892,17.395575,18.421728,18.048239,13.743673,10.616167,8.756263,3.259548,2.9803739,3.6481283,4.8063245,5.3382645,3.4594972,3.6066296,5.5382137,7.2094865,8.152642,9.480607,11.898859,13.36641,13.898351,13.6833105,13.102326,13.615403,14.400109,14.962231,14.800008,13.373956,12.800517,12.932558,12.808062,12.253486,11.910177,12.581704,13.196642,13.215506,12.770335,12.687338,12.079946,11.136789,10.253995,9.522105,8.748717,8.45068,8.096053,7.6622014,7.3490734,7.5905213,9.178797,10.087999,9.684328,8.412953,7.798016,7.4282985,9.1976595,10.419991,10.321902,10.012547,4.142342,5.8136153,8.201687,8.428044,7.567886,6.379509,5.7306175,7.594294,11.080199,12.438345,7.7112455,6.4021444,6.2625575,5.836251,4.4177437,4.7535076,5.4665337,6.900131,8.771353,10.133271,7.462252,6.9680386,7.7225633,8.126234,5.9192486,8.726082,13.389046,14.890551,11.823407,6.398372,7.2170315,6.205968,6.0286546,7.001992,7.1000805,6.7944975,5.5382137,4.798779,5.010046,5.5570765,5.4891696,5.8098426,5.594803,4.7610526,4.0517993,3.6141748,2.9351022,2.1466236,1.5052774,1.4147344,1.4373702,1.4864142,1.4411428,1.3355093,1.3694628,1.3694628,1.5316857,1.690136,1.7957695,1.9051756,2.1692593,3.0369632,3.1916409,2.5880208,2.4333432,2.938875,4.1536603,5.692891,7.043491,7.6093845,7.1302614,7.496206,8.29223,8.99771,8.990166,9.21275,8.394091,7.413208,6.7643166,6.5568223,6.217286,5.994701,5.8098426,5.7494807,6.0776987,5.353355,5.20245,5.27413,5.43258,5.73439,5.7909794,5.704209,5.8664317,6.228604,6.3153744,7.1000805,7.0548086,6.620957,6.477597,7.5301595,7.9338303,8.7600355,8.710991,7.937603,8.039464,7.707473,7.122716,7.145352,7.5905213,7.2283497,7.3868,7.435844,7.466025,7.5075235,7.533932,7.8131065,7.141579,6.598321,6.3455553,5.6098933,5.0779533,5.1043615,5.6778007,6.405917,6.530414,6.802043,7.0548086,7.454707,7.7187905,7.1000805,7.1604424,7.8734684,8.586494,9.190115,10.121953,9.318384,9.733373,9.952185,9.842778,10.574668,10.642575,11.970539,13.645585,14.611377,13.664448,12.928786,13.113645,13.498452,13.521088,12.751472,12.223305,13.109872,13.328684,11.978085,9.337247,7.352846,6.964266,7.5527954,8.186596,7.6207023,8.258276,9.933322,11.653639,13.038192,14.32843,13.615403,13.385274,13.875714,14.705692,14.875461,15.113135,13.728582,12.264804,11.117926,9.529651,9.612649,10.106862,10.555805,10.435081,9.129752,14.818871,14.916959,13.419228,10.955703,4.8063245,11.204697,11.551778,12.528888,14.011529,9.0807085,8.318638,15.173498,23.593996,24.310795,4.8100967,13.830443,8.75249,8.922258,17.097536,19.444109,11.747954,7.3868,7.0472636,9.457971,11.363147,7.6282477,6.5228686,6.115425,5.4174895,4.38379,4.3309736,5.330719,6.217286,6.6662283,7.213259,7.7187905,7.4773426,7.1076255,6.7756343,6.205968,6.1795597,6.677546,6.937857,6.63982,5.907931,5.643847,5.7117543,6.126743,6.530414,6.168242,5.907931,5.5004873,5.27413,5.1647234,4.7421894,4.025391,3.3689542,3.62172,4.6818275,5.492942,4.8553686,4.749735,4.6629643,4.696918,5.5797124,5.5495315,5.243949,5.50426,6.156924,6.0211096,5.9003854,6.017337,5.824933,5.5004873,5.945657,5.8702044,6.40969,6.934085,7.201941,7.33021,7.0510364,6.6850915,6.6020937,6.802043,6.937857,7.8696957,9.178797,9.250477,8.371455,8.722309,8.820397,8.959985,8.827943,8.36391,7.7225633,8.488406,8.956212,9.288202,9.378746,8.846806,8.503497,8.846806,9.273112,9.390063,9.016574,7.515069,6.609639,6.258785,6.224831,6.0701537,6.221059,6.0211096,5.9003854,5.8664317,5.515578,4.9534564,5.160951,5.6325293,6.0362,6.2361493,6.092789,5.96452,6.0550632,6.255012,6.1342883,5.9984736,6.643593,7.352846,7.6886096,7.4811153,6.7944975,6.1833324,6.119198,6.2927384,5.613666,4.768598,4.3121104,3.9763467,3.6254926,3.2746384,3.3840446,3.8895764,4.353609,4.7610526,5.534441,5.715527,5.6400743,5.2552667,4.8138695,4.878004,4.9534564,5.300538,5.191132,4.5422406,3.9159849,3.1954134,3.3689542,3.742444,4.115934,4.8025517,5.5759397,5.9909286,6.175787,6.1342883,5.726845,6.0512905,6.851087,7.33021,7.3490734,7.4207535,8.348819,8.495952,8.514814,8.620448,8.560086,8.409182,9.0543,9.688101,9.95973,9.97482,1.9542197,2.161714,2.2748928,2.1843498,2.0485353,2.305074,2.7200627,2.9615107,3.0709167,3.2331395,3.783943,3.6745367,3.572676,3.610402,3.7273536,3.6783094,4.08198,4.5007415,5.0439997,5.451443,5.0968165,5.523123,5.311856,5.1647234,5.4288073,6.089017,6.5530496,6.8963585,7.1604424,7.1868505,6.6360474,7.3453007,7.8810134,8.088508,7.9941926,7.8131065,8.52236,8.809079,8.661947,8.107371,7.201941,6.224831,7.0057645,7.786698,7.828197,7.4018903,7.303802,6.903904,6.749226,6.934085,7.0812173,8.228095,8.661947,8.526133,8.631766,10.453944,12.332711,13.472044,15.992157,18.806536,17.60684,15.777118,15.520579,15.777118,15.384765,13.075918,11.355601,5.836251,1.7165444,0.5772116,0.38103512,0.28294688,0.31312788,0.22258487,0.030181,0.030181,1.7882242,1.1016065,0.23013012,0.041498873,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.011317875,0.1358145,0.3169005,0.4376245,0.3055826,0.18485862,0.150905,0.18863125,0.21503963,0.1056335,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.056589376,0.033953626,0.34330887,0.7167987,0.23013012,0.056589376,0.0150905,0.15467763,0.3055826,0.060362,0.9393836,0.6828451,0.58475685,0.8186596,0.42630664,1.0374719,1.6033657,1.7655885,1.7165444,2.1805773,1.3656902,1.50905,2.2899833,3.0407357,2.746471,2.5880208,3.3350005,3.7801702,4.063117,5.6778007,4.979865,5.3269467,5.8966126,6.25124,6.349328,8.518587,8.52236,8.631766,9.303293,9.156161,8.533678,9.529651,10.804798,11.536687,11.41219,12.366665,13.3626375,13.321139,12.800517,14.007756,15.105591,14.124708,13.132507,13.087236,13.8719425,13.698401,14.452927,15.0376835,15.358356,16.31283,16.188334,15.188588,14.317112,13.951167,13.856852,13.951167,13.472044,12.955194,12.559069,12.068627,13.377728,14.4152,15.403628,16.24115,16.509007,17.37671,17.621931,17.225805,16.905132,18.127462,19.444109,19.11589,18.365139,17.799244,17.410664,17.312576,17.89356,18.844261,19.58747,19.270569,20.711712,20.798481,20.383493,20.085455,20.277859,20.92675,21.424738,21.839725,22.352802,23.254461,23.620405,23.75622,23.409138,22.639523,21.820864,20.489126,19.61765,19.202662,18.957441,18.312323,17.139036,15.965749,15.471535,15.965749,17.380484,19.651604,21.553007,22.281124,21.632233,20.036411,19.300749,18.79899,18.414183,17.976559,17.255987,16.392056,16.603323,17.527617,18.485863,18.5085,17.093763,16.4826,17.252214,19.308294,21.896315,22.873425,23.420456,22.797974,21.05502,19.029121,18.478317,18.742401,20.402355,22.443346,22.24717,21.820864,20.432537,19.240387,18.58395,17.961468,17.372938,15.826162,14.283158,13.743673,15.260268,17.248442,17.984104,18.131235,18.459454,19.851553,19.338476,18.632996,17.784155,17.482344,19.04421,21.190834,20.281631,18.742401,18.534906,21.134245,17.984104,13.762536,10.227587,7.8017883,5.553304,3.380272,1.9127209,2.2371666,3.5462675,3.1425967,2.4974778,3.7273536,5.20245,6.5040054,8.409182,10.725573,12.370438,13.290957,13.249459,11.796998,11.491416,13.072145,14.7170105,15.422491,14.984866,14.800008,15.0376835,14.532151,13.106099,11.581959,12.925014,13.487134,13.385274,13.113645,13.5663595,12.234623,11.140562,10.26154,9.556059,8.956212,8.492179,7.745199,7.33021,7.1264887,6.270103,8.601585,10.284176,11.09529,10.702937,8.650629,6.9567204,8.948667,10.355856,9.914458,9.352338,5.485397,9.533423,15.441354,19.553514,20.628714,13.671993,8.00551,7.303802,10.608622,12.3289385,10.374719,7.2962565,5.7570257,5.66271,4.1498876,3.9688015,4.3875628,6.273875,9.88805,14.890551,11.793225,9.001483,6.7454534,5.2967653,4.991183,7.8961043,9.42779,9.782416,8.763808,5.798525,5.994701,5.8588867,6.145606,6.5266414,5.5985756,5.723072,5.5683947,7.5226145,10.340765,9.171251,9.952185,9.159933,6.8699503,4.1008434,2.806833,2.9049213,2.8747404,2.5389767,1.9994912,1.6335466,1.4147344,1.2110126,1.1431054,1.1996948,1.237421,0.94315624,0.98842776,1.146878,1.3053282,1.4637785,1.5731846,1.8221779,1.9429018,1.8221779,1.478869,2.052308,2.8936033,4.1989317,5.643847,6.3644185,6.5568223,6.700182,7.6282477,8.880759,8.695901,8.782671,8.503497,7.6282477,6.507778,6.043745,6.006019,6.187105,5.945657,5.6778007,6.8359966,5.7872066,5.0213637,4.9534564,5.198677,4.561104,5.1345425,5.251494,5.5457587,6.145606,6.6850915,6.255012,6.5530496,6.6813188,6.651138,7.3717093,9.005256,9.378746,8.907167,8.209232,8.088508,7.4018903,6.8850408,7.3905725,8.254503,7.277394,7.0849895,7.5565677,8.197914,8.36391,7.277394,7.594294,7.4811153,6.530414,5.2326307,4.9760923,4.7044635,5.0779533,5.5985756,6.3342376,7.9338303,8.75249,9.333474,8.75249,7.3453007,6.700182,7.432071,7.7716074,7.7942433,7.9489207,9.046755,9.559832,10.834979,11.559323,11.551778,11.732863,13.29473,13.932304,14.452927,14.822643,14.173752,13.332457,12.691111,12.577931,12.996693,13.656902,12.619431,12.800517,14.622695,16.565596,15.135772,9.703192,7.8508325,8.718536,10.378491,9.842778,10.536942,11.299012,12.306303,13.547497,14.815099,13.204187,12.434572,13.223051,15.414946,17.991648,16.927769,15.803526,14.807553,13.570132,11.155652,10.884023,11.385782,12.66093,12.6345215,7.141579,10.816116,15.743164,16.45619,12.679792,9.322156,12.985375,14.603831,15.388537,15.588487,14.524607,7.6886096,6.587003,7.8998766,9.020347,8.054554,11.902632,8.488406,8.8769865,14.584969,17.56157,13.6682205,9.133525,7.7904706,10.167224,13.472044,7.699928,5.534441,5.4967146,6.56814,8.179051,5.481624,5.1458607,6.0550632,7.092535,7.141579,7.5565677,7.5603404,7.7112455,7.7414265,6.5455046,5.934339,6.541732,7.0057645,6.590776,5.1873593,4.2102494,4.772371,5.80607,6.3153744,5.3873086,4.9723196,4.6554193,4.2894745,3.9499383,3.9386206,3.6179473,3.2482302,3.8103511,5.0666356,5.553304,4.6629643,4.447925,4.5460134,4.859141,5.553304,4.821415,4.8025517,5.3458095,6.009792,6.058836,5.704209,5.934339,5.534441,4.7233267,5.1873593,5.7004366,6.149379,6.2399216,6.1833324,6.6850915,6.7077274,6.330465,5.975838,5.926794,6.3153744,7.9413757,8.741172,9.178797,9.601331,10.223814,9.552286,9.7220545,10.344538,10.518079,8.835487,8.503497,8.52236,8.986393,9.322156,8.284684,8.469543,9.163706,9.635284,9.601331,9.246704,7.1604424,6.5568223,6.56814,6.5341864,5.9984736,5.726845,5.5797124,5.772116,6.0776987,5.783434,4.7836885,4.447925,4.67051,5.3080835,6.2097406,6.187105,6.700182,6.8171334,6.379509,6.013564,5.534441,5.6551647,6.5228686,7.7716074,8.529905,7.3075747,6.3644185,5.9192486,5.6891184,4.881777,4.2102494,4.1083884,3.8405323,3.3123648,3.0671442,3.712263,4.323428,4.5120597,4.3875628,4.5460134,5.243949,5.379763,5.2137675,5.1345425,5.66271,5.4891696,4.961002,4.689373,4.647874,4.195159,3.4745877,3.2331395,3.3123648,3.6934,4.485651,4.6931453,5.4778514,6.1606965,6.3229194,5.798525,5.9682927,6.809588,6.9793563,6.5568223,7.020855,8.337502,8.677037,8.6581745,8.707218,9.046755,9.367428,9.307066,9.673011,10.521852,11.170743,1.8938577,1.9730829,2.093807,2.1277604,2.0975795,2.1579416,2.493705,2.7615614,2.8747404,2.9652832,3.3689542,3.259548,3.5462675,3.9650288,4.3007927,4.398881,4.4894238,4.647874,4.919503,5.243949,5.4740787,5.4250345,5.6551647,5.836251,5.9720654,6.405917,6.8397694,7.1868505,7.2698483,7.17176,7.1981683,7.6320205,7.748972,7.696155,7.677292,7.9225125,7.937603,7.9262853,7.6131573,7.020855,6.458734,6.330465,6.5643673,6.907676,7.2924843,7.7904706,7.4773426,7.2887115,7.24344,7.3151197,7.435844,8.160188,8.284684,8.439363,9.167479,10.929295,12.14408,14.1058445,16.67123,18.327412,16.192106,14.558559,13.970031,14.426518,13.88326,8.254503,5.975838,3.218049,1.4750963,0.94315624,0.5017591,0.44516975,0.5885295,0.9997456,1.2110126,0.21503963,0.4376245,0.27540162,0.09808825,0.041498873,0.0150905,0.026408374,0.026408374,0.018863125,0.003772625,0.00754525,0.0,0.00754525,0.00754525,0.0,0.0,0.003772625,0.1056335,0.15467763,0.120724,0.120724,0.17731337,0.3734899,0.4979865,0.42630664,0.13204187,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.0452715,0.06790725,0.060362,0.12826926,0.20372175,0.0452715,0.24522063,0.19994913,0.30181,0.48666862,0.24522063,0.6451189,0.7432071,0.8526133,1.0751982,1.3317367,1.4901869,1.7919968,1.9504471,1.8749946,1.6561824,1.8259505,1.9655377,2.1088974,2.3013012,2.625747,2.9728284,2.9615107,3.5538127,4.568649,4.689373,4.557331,4.8629136,5.4891696,6.466279,7.960239,9.25425,9.703192,9.627739,9.378746,9.337247,9.691874,10.035183,10.340765,10.827434,11.925267,12.525115,13.083464,13.558814,13.81158,13.604086,15.007503,14.34352,13.475817,13.128735,12.90615,14.913187,15.580941,15.46399,14.769827,13.358865,13.430545,14.128481,14.562332,14.569878,14.698147,13.690856,13.170234,12.842015,12.47607,11.898859,12.336484,13.415455,14.871688,16.26756,16.984358,17.316349,18.734856,19.270569,18.602814,18.055782,18.289686,18.025602,18.421728,19.54597,20.375948,20.52308,20.930523,21.115381,20.99843,20.89657,21.613369,21.436056,20.821117,20.243906,20.194862,20.341993,20.526854,21.583187,23.322369,24.548471,24.1448,23.646814,23.26955,22.790428,21.553007,19.478064,19.496925,19.87796,19.957186,20.130728,20.440083,18.666948,17.056038,16.592005,17.014538,17.840744,18.708447,18.912169,18.391546,17.738882,17.271078,16.776863,16.493916,16.59955,17.195625,16.641048,16.663685,17.40312,18.417955,18.65563,17.025856,15.863888,15.773345,16.87118,18.7839,20.093,21.205925,21.187061,20.14959,19.247932,18.765038,18.402864,18.549997,19.119663,19.549744,19.319613,18.900852,18.749947,18.58395,17.372938,17.335213,16.531643,15.543215,15.052773,15.845025,17.063583,17.904879,18.614132,19.255478,19.73083,18.172735,16.350557,15.784663,16.712729,18.078419,20.315586,20.387266,19.255478,18.304777,19.349794,19.180025,16.803272,11.84227,6.205968,4.0782075,2.6182017,1.8561316,2.052308,2.6031113,2.0447628,2.3956168,3.1312788,4.323428,5.7079816,6.722818,8.858124,10.95193,12.408164,12.955194,12.623203,12.808062,13.264549,13.671993,13.773854,13.373956,13.422999,13.875714,13.928532,13.411682,12.766563,13.023102,12.694883,12.068627,11.608367,11.955449,11.69891,11.083972,10.495442,9.914458,8.956212,9.099571,8.273367,7.4697976,7.183078,7.432071,8.627994,9.661693,9.6051035,8.586494,7.786698,8.431817,9.955957,10.521852,9.684328,8.390318,5.0553174,4.889322,7.1038527,9.808825,10.035183,10.506761,7.605612,7.254758,9.756008,9.778644,10.11818,6.609639,4.187614,4.06689,3.7235808,4.7120085,4.436607,5.081726,7.5603404,11.510279,12.50248,10.729345,8.122461,6.25124,6.307829,8.254503,11.050018,11.570641,9.559832,7.61693,8.262049,8.409182,8.537451,8.635539,8.175279,8.82417,8.152642,6.960493,5.9682927,5.802297,7.756517,10.469034,10.495442,7.4735703,4.13857,3.7763977,3.361409,2.5427492,1.5316857,1.0940613,0.91674787,0.90543,0.8299775,0.663982,0.5998474,0.6413463,0.8111144,0.98465514,1.1091517,1.20724,1.1242423,1.4600059,1.6561824,1.5958204,1.6260014,1.9278114,2.6521554,3.7877154,5.0477724,5.873977,6.138061,6.2097406,6.9567204,8.197914,8.695901,7.9338303,7.3075747,6.571913,5.7872066,5.3344917,5.160951,5.8437963,5.824933,5.247721,5.9682927,5.6815734,5.062863,4.7836885,4.7535076,4.112161,4.568649,4.7912335,5.3873086,6.405917,7.3415284,7.443389,7.8998766,8.141325,7.854605,7.001992,7.7301087,7.884786,7.677292,7.5037513,7.9300575,7.4396167,6.590776,6.7114997,7.877241,8.903395,7.9941926,6.85486,6.6624556,7.1378064,6.5228686,6.722818,7.6923823,7.643338,6.428553,5.534441,5.0515447,5.2552667,5.2892203,5.198677,5.907931,7.8998766,8.412953,7.865923,6.990674,6.832224,6.462507,6.8246784,7.5490227,8.356364,9.073163,8.431817,9.088254,9.771099,10.231359,11.246195,12.543978,12.925014,13.6682205,14.64533,14.320885,14.3095665,14.147344,13.9888935,13.819125,13.472044,13.20796,13.479589,13.732355,13.302276,11.41219,10.540714,9.024119,8.835487,10.080454,10.989656,11.966766,11.91395,12.66093,14.558559,16.452417,16.452417,15.486626,15.218769,16.248695,18.112373,17.497435,17.746428,17.708702,16.633503,14.158662,12.034674,11.415963,12.445889,12.996693,8.703445,11.917723,12.96274,12.434572,10.974566,9.239159,9.774872,14.385019,16.505234,14.490653,11.634775,10.393582,8.812852,8.360137,8.7751255,8.043237,9.352338,8.631766,8.8618965,11.510279,16.550507,12.019584,8.661947,7.9828744,10.336992,14.924504,10.929295,9.178797,7.435844,6.0701537,8.043237,6.255012,6.270103,6.1305156,5.798525,7.164215,6.5455046,6.6322746,7.149124,7.5263867,6.937857,5.8966126,6.2927384,6.790725,6.537959,5.1647234,4.508287,4.859141,5.624984,6.168242,5.7909794,4.515832,3.6254926,3.259548,3.3764994,3.7537618,3.640583,3.7462165,4.142342,4.640329,4.798779,4.6290107,4.8100967,4.930821,4.8440504,4.6516466,4.485651,5.304311,6.1116524,6.428553,6.300284,5.987156,5.451443,5.2137675,5.455216,6.006019,6.6850915,6.4511886,5.9192486,5.6061206,5.9003854,5.534441,5.572167,5.8928404,6.1908774,5.975838,7.394345,8.382772,9.092027,9.6051035,9.940866,8.578949,8.379,8.790216,9.288202,9.359882,8.669493,8.575176,8.75249,8.831716,8.420499,8.944894,9.529651,10.072908,10.159679,9.065618,6.8774953,6.696409,7.0170827,6.971811,6.326692,5.9494295,5.847569,5.715527,5.413717,4.9534564,4.5460134,4.504514,4.7610526,5.3156285,6.198423,5.764571,6.0022464,6.066381,5.80607,5.7306175,5.8136153,6.436098,7.069899,7.488661,7.786698,7.01331,6.428553,6.0701537,5.666483,4.6252384,4.715781,4.644101,4.2027044,3.6028569,3.4444065,4.014073,4.779916,5.2590394,5.3759904,5.485397,5.624984,5.594803,5.2590394,4.957229,5.4891696,5.66271,5.3269467,5.089271,5.0741806,4.9647746,4.304565,3.5839937,3.3764994,3.783943,4.447925,4.745962,5.281675,5.7306175,5.9192486,5.8211603,5.613666,5.7796617,6.013564,6.3417826,7.1302614,8.182823,8.601585,8.91094,9.291975,9.58624,9.608876,9.608876,9.688101,9.952185,10.510533,1.7127718,1.7391801,1.8448136,1.9202662,1.9844007,2.1956677,2.4899325,2.7540162,2.8332415,2.7917426,2.9464202,2.8558772,3.1765501,3.6179473,4.0706625,4.5761943,4.478106,4.617693,4.8025517,5.0251365,5.4778514,5.481624,5.666483,5.8588867,6.1116524,6.696409,7.277394,7.567886,7.5829763,7.4169807,7.2283497,7.194396,7.0510364,6.862405,6.79827,7.152897,6.9227667,6.9491754,6.779407,6.398372,6.25124,6.771862,7.001992,7.3453007,7.9036493,8.484633,8.050782,8.239413,8.326183,8.050782,7.594294,7.967784,8.156415,8.684583,9.6051035,10.480352,12.51757,15.271586,16.750456,16.418465,15.214996,14.268067,15.0905,15.63753,14.690601,11.872451,7.062354,5.6589375,5.9003854,5.5759397,2.0070364,1.1317875,1.1431054,1.7127718,1.9655377,0.5055317,0.24522063,0.11317875,0.049044125,0.0150905,0.00754525,0.011317875,0.018863125,0.0150905,0.00754525,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.041498873,0.08677038,0.10186087,0.056589376,0.18485862,0.38103512,0.52062225,0.49421388,0.17354076,0.06413463,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.026408374,0.060362,0.041498873,0.11317875,0.24522063,0.23767537,0.331991,0.211267,0.26031113,0.452715,0.3169005,0.91297525,1.1355602,1.1808317,1.1317875,0.9620194,1.4147344,1.6788181,1.6825907,1.539231,1.5731846,2.0447628,2.5087957,2.8030603,3.0633714,3.7009451,3.1614597,3.4066803,4.1989317,4.991183,4.927048,4.961002,5.119452,5.6363015,6.722818,8.571404,10.152134,10.767072,10.352083,9.684328,10.38981,10.9594755,11.536687,12.019584,12.687338,14.188843,14.252977,13.588995,13.347548,13.539951,13.038192,14.109617,14.022847,13.35132,12.47607,11.566868,12.785426,13.739901,14.154889,14.094527,13.973803,12.996693,12.921241,13.328684,13.864397,14.237886,12.913695,12.272349,12.58925,13.309821,13.0646,12.940104,13.573905,15.264041,17.271078,17.84829,16.957949,17.961468,18.915941,19.047983,18.76881,18.591496,18.632996,19.093256,19.855326,20.477808,20.764528,21.598278,22.137764,22.058538,21.537916,21.688822,21.334194,20.922977,20.658894,20.48158,19.94964,20.243906,21.251196,22.884743,25.054003,25.634987,25.39354,24.065575,22.062311,20.440083,18.848034,19.251705,20.051502,20.8513,22.450891,23.925987,22.284895,19.930779,18.297232,17.882242,18.119919,18.244415,18.02183,17.527617,17.157898,16.731592,16.376965,16.248695,16.478827,17.16167,16.935314,16.77309,16.984358,17.64834,18.599041,17.595524,16.984358,16.795727,16.980585,17.399347,18.221779,19.255478,19.934551,20.198635,20.48158,19.983595,19.28566,18.270823,17.384256,17.610613,18.146326,18.206688,18.41041,18.440592,17.025856,16.946632,16.58446,16.214743,16.052519,16.237377,16.158154,16.969267,18.278368,19.357338,19.176252,17.014538,15.875206,16.335466,17.667202,17.829426,20.07791,20.719257,19.685556,18.097282,18.23687,19.036665,17.580433,12.781653,6.530414,3.651901,3.4481792,2.6144292,2.203213,2.2069857,1.5580941,1.8334957,2.3805263,3.3878171,4.6214657,5.413717,7.039718,9.273112,11.321648,12.743927,13.4644985,13.777626,13.6682205,13.377728,12.996693,12.50248,12.97783,13.4644985,13.570132,13.275867,12.90615,13.332457,13.143826,12.483616,11.759273,11.615912,11.706455,11.408418,10.989656,10.446399,9.476834,9.016574,8.050782,7.1038527,6.741681,7.575431,8.7751255,9.6051035,9.857869,10.061591,11.487643,14.566105,15.071637,13.132507,9.948412,7.7829256,5.6098933,4.2328854,4.1574326,5.0439997,5.7004366,6.48137,5.583485,5.6023483,6.4436436,5.3609,8.763808,6.741681,4.323428,3.7499893,4.485651,5.1835866,6.0626082,7.5112963,9.627739,12.257258,13.422999,12.079946,9.152389,6.4436436,6.6549106,6.6813188,9.0543,9.9257765,8.477088,6.9567204,10.084227,11.970539,13.758763,14.739646,12.362892,10.808571,8.601585,6.013564,3.9989824,4.217795,6.0739264,9.107117,10.623712,10.352083,10.438853,8.631766,5.938112,3.874486,2.686109,1.3656902,0.6149379,0.45648763,0.422534,0.33576363,0.29426476,0.38103512,0.56589377,0.7507524,0.8941121,1.0072908,0.95447415,1.1129243,1.2449663,1.2487389,1.1883769,1.4411428,1.9693103,2.916239,4.093298,4.983638,5.5570765,5.7494807,6.221059,7.0472636,7.7187905,7.152897,6.3116016,5.6098933,5.240176,5.1760416,4.7044635,5.451443,5.692891,5.1269975,4.8742313,5.062863,4.708236,4.6327834,4.6856003,3.7688525,4.0216184,4.346064,5.010046,5.9984736,7.020855,7.496206,7.816879,7.9715567,7.937603,7.6810646,8.167733,7.865923,7.4509344,7.3113475,7.5603404,7.4207535,6.617184,6.3342376,6.9265394,7.9262853,8.575176,7.8923316,6.9491754,6.300284,5.983383,6.205968,6.862405,6.851087,6.156924,5.8702044,5.323174,5.0025005,4.919503,5.160951,5.87775,7.281166,7.7301087,7.4207535,6.8473144,6.802043,6.6247296,6.934085,8.228095,9.831461,9.922004,9.367428,9.574923,10.038955,10.570895,11.314102,12.2119875,13.04951,14.162435,15.022593,14.230342,13.45318,13.373956,13.70972,14.045483,13.849306,14.022847,14.290704,14.007756,12.200669,7.564113,10.174769,10.008774,9.850324,10.604849,11.302785,12.785426,13.517315,14.943368,17.063583,18.45568,19.221525,18.644312,18.62545,19.534653,20.202406,19.723284,20.179771,19.83269,18.568861,17.908651,14.852824,13.547497,13.215506,12.842015,11.1631975,13.898351,12.815607,12.789199,13.521088,9.556059,9.567377,12.483616,16.463736,18.621677,15.056546,12.800517,10.329447,9.997457,11.310329,10.914205,10.223814,9.808825,9.929549,10.93684,13.275867,10.725573,8.29223,8.782671,12.359119,16.524097,11.98563,11.004747,11.419736,11.170743,8.311093,7.5037513,7.9941926,8.137552,7.745199,8.096053,6.9755836,6.33801,6.3342376,6.6662283,6.5756855,6.673774,6.760544,6.643593,6.1720147,5.2288585,4.9119577,4.938366,5.13077,5.2854476,5.1571784,4.014073,3.078462,2.776652,3.138824,3.7990334,3.893349,4.1083884,4.3347464,4.4705606,4.425289,4.5120597,4.817642,4.889322,4.6516466,4.406426,4.7346444,5.1081343,5.7117543,6.368191,6.5643673,6.398372,6.1644692,6.217286,6.4738245,6.4134626,6.722818,6.4210076,6.33801,6.6134114,6.696409,6.1003346,5.855114,6.119198,6.5228686,6.156924,6.964266,7.7376537,8.850578,9.914458,9.782416,8.903395,8.137552,7.884786,8.209232,8.82417,8.582722,8.782671,8.971302,8.873214,8.390318,8.801534,9.242931,9.9257765,10.223814,8.68081,7.0774446,6.971811,7.250985,7.1566696,6.2814207,5.9230213,5.8400235,5.696664,5.3269467,4.745962,4.8025517,4.938366,5.221313,5.6325293,6.058836,5.3609,5.2326307,5.342037,5.5306683,5.855114,6.2927384,7.141579,7.6697464,7.696155,7.6093845,6.971811,6.2361493,5.798525,5.617439,5.194905,5.4438977,5.292993,4.8365054,4.285702,3.953711,4.2517486,4.5799665,4.696918,4.7308717,5.1647234,5.198677,5.1156793,4.949684,4.847823,5.0553174,5.27413,4.9685473,4.7346444,4.772371,4.90064,4.398881,3.682082,3.451952,3.8178966,4.285702,4.45547,5.0968165,5.6476197,5.8626595,5.802297,5.372218,5.666483,6.3455553,7.092535,7.6131573,8.194141,8.809079,9.314611,9.612649,9.665465,9.514561,9.661693,9.97482,10.238904,10.163452,1.6335466,1.8787673,1.8938577,1.9051756,2.033445,2.2862108,2.4597516,2.757789,2.8936033,2.8294687,2.7615614,2.8747404,3.1199608,3.429316,3.832987,4.436607,4.4630156,4.749735,4.9459114,5.0062733,5.2326307,5.1458607,5.323174,5.666483,6.1229706,6.677546,7.2585306,7.424526,7.3981175,7.164215,6.466279,6.1041074,5.8928404,5.8173876,5.9305663,6.3153744,6.221059,6.519096,6.5568223,6.296511,6.326692,7.0887623,7.488661,7.858378,8.307321,8.733627,8.809079,9.114662,9.012801,8.439363,7.937603,7.9941926,8.118689,8.729855,9.676784,10.253995,12.883514,15.758255,17.029629,17.425755,20.270313,20.53817,21.67373,20.477808,17.53139,17.191853,10.684074,8.375228,7.8810134,6.9567204,3.5160866,1.5241405,1.0412445,1.2902378,1.4034165,0.422534,0.23013012,0.09808825,0.026408374,0.003772625,0.0,0.003772625,0.030181,0.03772625,0.018863125,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.041498873,0.094315626,0.0754525,0.23390275,0.41498876,0.4678055,0.34330887,0.124496624,0.060362,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.02263575,0.03772625,0.02263575,0.10940613,0.27540162,0.3169005,0.2867195,0.2565385,0.4376245,0.6828451,0.4640329,1.056335,1.358145,1.2713746,0.9280658,0.7054809,1.3430545,1.7731338,2.0598533,2.1051247,1.6222287,2.5238862,3.8141239,4.4894238,4.376245,4.1272516,3.742444,4.112161,4.666737,5.111907,5.455216,5.8702044,6.1795597,6.673774,7.6848373,9.608876,10.902886,11.431054,11.23865,10.925522,11.653639,12.019584,12.800517,13.27964,13.543724,14.48688,14.215251,13.132507,12.751472,13.204187,13.238141,13.200415,12.951422,12.249713,11.249968,10.49167,11.027383,12.053536,13.04951,13.917213,14.999957,13.924759,12.762791,12.506252,13.158916,13.728582,12.81938,12.151625,12.23085,13.038192,14.015302,14.120935,14.879233,16.407146,18.014284,18.214233,17.14658,17.37671,18.26705,19.266796,19.923233,19.53088,19.353567,19.278114,19.413929,20.100546,20.621168,21.571869,22.315077,22.36412,21.368149,21.353058,21.051247,20.88148,20.89657,20.775846,19.813826,19.817598,20.489126,21.820864,24.103302,26.110338,26.710184,24.967232,21.719002,19.579924,18.761265,19.081938,19.783646,20.98334,23.673222,25.736847,24.861599,22.688566,20.557034,19.48938,18.968758,18.376457,17.844517,17.482344,17.399347,17.210714,16.912678,16.690092,16.603323,16.588232,16.791954,16.72782,16.84477,17.391802,18.421728,17.991648,17.95015,17.908651,17.640795,17.063583,17.139036,17.836971,18.848034,19.915688,20.836208,20.572124,20.028866,18.708447,17.184307,17.127718,18.097282,18.33873,18.568861,18.666948,17.64834,17.033401,16.625957,16.588232,16.788181,16.810818,15.954432,16.26756,17.297485,18.293459,18.184053,16.776863,16.490145,17.384256,18.489635,17.784155,19.855326,20.232588,19.11589,17.595524,17.625704,18.119919,18.176508,14.2077055,7.5490227,4.4818783,4.093298,2.8143783,1.8976303,1.629774,1.3204187,1.2034674,1.5958204,2.5238862,3.7273536,4.6629643,6.175787,8.43559,10.891568,13.132507,14.890551,14.939595,14.464244,13.800262,13.132507,12.510024,13.023102,13.253232,13.328684,13.313594,13.166461,13.634267,13.743673,13.396591,12.694883,11.921495,11.796998,11.604594,11.2801485,10.7557535,9.95973,8.75249,7.5792036,6.670001,6.4511886,7.5301595,8.269594,9.065618,9.688101,10.631257,13.106099,15.671484,15.735619,13.992666,11.170743,8.039464,6.8171334,6.530414,6.2097406,5.828706,6.2814207,5.515578,5.1269975,5.2552667,5.2288585,3.5462675,7.2660756,6.33801,4.7874613,4.5196047,5.3458095,6.417235,9.076936,11.925267,13.958713,14.5283785,12.253486,10.665211,8.473316,6.3531003,6.960493,6.300284,7.1264887,7.586749,7.424526,7.967784,12.14408,13.788944,14.867915,15.784663,15.4074,11.962994,9.001483,6.187105,4.214022,4.8025517,6.2323766,8.031919,9.514561,10.982111,13.758763,11.77059,8.160188,5.20245,3.3123648,1.0450171,0.33953625,0.150905,0.15467763,0.1659955,0.15467763,0.1961765,0.32067314,0.482896,0.6488915,0.76207024,0.80734175,0.9808825,1.0789708,1.0223814,0.8563859,0.98465514,1.2826926,2.0673985,3.218049,4.172523,4.9421387,5.2628117,5.523123,5.8626595,6.1606965,6.145606,5.523123,4.8440504,4.5233774,4.847823,4.5950575,5.27413,5.5268955,4.9459114,4.063117,4.561104,4.4215164,4.4139714,4.459243,3.6179473,3.4142256,3.7914882,4.4931965,5.3156285,6.089017,6.72659,7.322665,7.4999785,7.5075235,8.216777,8.514814,7.877241,7.224577,7.0510364,7.4018903,7.6320205,6.960493,6.4210076,6.3832817,6.5530496,8.326183,8.6581745,7.492433,5.904158,6.1229706,6.670001,6.688864,6.187105,5.6287565,5.9418845,5.349582,4.9232755,4.938366,5.349582,5.7872066,6.8133607,7.4207535,7.3679366,6.858632,6.5455046,7.213259,7.809334,9.186342,10.789707,10.616167,10.178542,9.861642,10.03141,10.653893,11.283921,12.128989,13.626721,14.811326,15.120681,14.396337,13.230596,12.81938,13.245687,14.117163,14.558559,14.479335,14.332202,14.158662,12.585477,6.79827,9.582467,10.11818,10.201178,10.910432,12.577931,14.852824,16.407146,18.025602,19.50447,19.662922,21.311558,21.820864,22.024584,22.326395,22.673477,21.952906,21.134245,19.825144,18.953669,20.8098,18.384,17.33144,16.0827,14.215251,12.445889,17.056038,16.905132,16.761772,15.954432,8.382772,10.816116,11.993175,16.452417,22.432028,21.881226,17.327667,12.083718,10.344538,12.019584,12.736382,11.185833,10.61994,10.997202,11.668729,11.378237,10.310584,8.284684,9.710737,14.237886,16.750456,11.544232,10.842525,12.898605,14.154889,9.246704,7.4396167,8.544995,9.695646,9.665465,8.888305,7.3113475,6.149379,5.8211603,6.1078796,6.1418333,7.118943,7.2962565,6.911449,6.217286,5.4703064,5.323174,5.1345425,4.659192,4.055572,3.893349,3.2369123,2.6597006,2.546522,3.0143273,3.9084394,4.06689,4.168751,4.3649273,4.515832,4.191386,4.4101987,4.52715,4.45547,4.3800178,4.779916,5.5797124,5.4174895,5.4703064,6.017337,6.4474163,6.7039547,7.2472124,7.4282985,7.0472636,6.375736,6.530414,6.485142,6.8058157,7.3490734,7.2924843,7.141579,6.9454026,6.9189944,6.930312,6.507778,6.911449,7.3490734,8.424272,9.778644,10.099318,9.608876,8.729855,7.8395147,7.4018903,7.967784,8.326183,8.669493,8.907167,8.990166,8.918486,8.869441,9.0807085,9.548513,9.582467,7.8131065,6.9982195,7.0359454,7.3792543,7.3981175,6.3832817,6.0286546,5.8437963,5.745708,5.5382137,4.9232755,5.05909,5.168496,5.3986263,5.7004366,5.824933,5.2552667,4.9723196,5.070408,5.4438977,5.7796617,6.255012,7.1793056,7.756517,7.7301087,7.356619,6.8133607,6.119198,5.745708,5.753253,5.7909794,5.847569,5.7004366,5.3156285,4.7006907,3.8895764,3.99521,4.164978,4.244203,4.353609,4.878004,4.859141,4.7874613,4.768598,4.817642,4.847823,4.949684,4.678055,4.534695,4.666737,4.859141,4.4894238,3.942393,3.7160356,3.9122121,4.236658,4.4101987,4.949684,5.534441,5.8928404,5.783434,5.6476197,6.1908774,7.009537,7.7225633,7.967784,8.703445,9.4013815,9.88805,10.084227,10.03141,9.484379,9.714509,10.370946,10.8576145,10.321902,1.690136,2.1466236,2.052308,1.991946,2.1466236,2.282438,2.293756,2.5578396,2.776652,2.8143783,2.7011995,3.127506,3.3274553,3.4896781,3.7235808,4.0895257,4.293247,4.7120085,4.9685473,4.961002,4.8138695,4.4630156,4.6931453,5.2137675,5.7306175,5.945657,6.4021444,6.511551,6.488915,6.25124,5.4174895,5.05909,4.9345937,5.081726,5.43258,5.775889,6.047518,6.571913,6.741681,6.5832305,6.7831798,7.3905725,7.7376537,7.8734684,7.9828744,8.375228,9.21275,9.216523,8.729855,8.22055,8.296002,8.084735,8.103599,8.75249,9.997457,11.389555,13.35132,16.946632,20.440083,24.159891,30.479038,31.24488,30.067822,25.419947,19.655376,18.99894,12.936331,8.918486,6.066381,4.146115,3.5689032,1.2789198,0.362172,0.120724,0.094315626,0.041498873,0.049044125,0.030181,0.018863125,0.02263575,0.026408374,0.060362,0.241448,0.23390275,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.05281675,0.17354076,0.46026024,0.633801,0.47912338,0.120724,0.02263575,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.033953626,0.026408374,0.018863125,0.026408374,0.06790725,0.1358145,0.17354076,0.16222288,0.3470815,0.68661773,0.9242931,0.5885295,0.83752275,1.1393328,1.0487897,0.73566186,0.9808825,1.4562333,1.9994912,2.776652,3.3274553,2.5314314,3.5236318,5.172269,5.8966126,5.251494,3.9273026,4.561104,4.738417,5.0439997,5.7381625,6.730363,6.8737226,7.303802,7.907422,8.937348,10.978339,11.812089,12.155397,12.487389,12.902377,13.124963,13.211733,13.7700815,13.702174,13.041965,12.974057,12.1252165,11.710228,12.091263,13.034419,13.687083,12.393073,11.634775,10.816116,10.020092,9.993684,10.914205,11.785681,12.864652,14.015302,14.728328,14.675511,13.472044,12.683565,12.826925,13.370183,13.430545,12.853333,11.993175,11.849815,14.083209,14.966003,16.350557,17.346529,17.738882,17.99542,18.055782,18.0671,18.644312,19.783646,20.866388,20.23636,19.542198,19.119663,19.281887,20.30804,20.798481,21.27006,21.647322,21.526598,20.179771,20.111864,20.157135,20.4514,20.911661,21.236107,20.032639,19.33093,19.519562,20.545715,21.918951,24.695602,26.136745,24.989868,21.90386,19.4592,18.934805,18.874443,19.168707,20.285404,23.303505,24.903097,25.03514,24.197617,22.89606,21.662413,19.757236,18.414183,17.742655,17.67852,17.961468,18.172735,17.701157,17.142809,16.693865,16.15438,16.358103,16.561823,16.94286,17.508753,18.104828,18.0671,18.146326,18.199142,18.052011,17.463482,17.04472,17.365393,18.104828,19.01403,19.908142,20.108091,20.108091,19.372429,18.259504,18.010511,18.840488,19.17248,19.440336,19.610106,19.15739,17.795471,17.078674,16.991903,17.23335,17.225805,16.603323,16.131744,15.98084,16.16947,16.607096,16.693865,16.690092,17.165443,17.746428,17.078674,18.848034,18.802763,17.742655,16.735365,17.1164,17.014538,18.523588,15.260268,8.329956,6.33801,4.2819295,2.6106565,1.4713237,0.98465514,1.2449663,0.7997965,0.94315624,1.8146327,3.1765501,4.4177437,6.224831,8.428044,10.963248,13.615403,16.026112,15.69412,15.049001,14.298248,13.528633,12.713746,12.940104,12.849561,13.034419,13.539951,13.875714,13.841762,13.860624,13.819125,13.4644985,12.400619,11.793225,11.548005,11.276376,10.763299,9.97482,8.488406,7.2887115,6.6586833,6.719045,7.4282985,8.013056,8.66572,8.967529,9.420244,11.438599,11.887542,12.193124,12.811834,12.393073,7.8017883,6.7643166,8.371455,9.442881,8.948667,7.9753294,6.8774953,6.175787,6.1078796,5.9984736,4.22534,5.8588867,5.0062733,4.4516973,5.0062733,5.5080323,7.7150183,11.661184,14.9358225,16.180788,15.086727,9.955957,8.473316,7.375482,6.138061,7.009537,7.541477,7.3113475,7.115171,7.8961043,10.740664,13.441863,12.838243,11.18206,10.967021,14.894323,11.940358,9.650374,7.537705,5.9984736,6.2851934,7.54525,8.2507305,8.563859,9.22784,11.574413,10.676529,9.020347,6.168242,2.6898816,0.16222288,0.1056335,0.071679875,0.071679875,0.090543,0.08299775,0.090543,0.1358145,0.24899325,0.40367088,0.513077,0.60362,0.95447415,1.1016065,0.95447415,0.784706,0.69039035,0.79602385,1.3732355,2.3692086,3.399135,4.2328854,4.67051,4.8855495,4.9119577,4.6554193,4.9157305,4.8025517,4.255521,3.7160356,4.123479,4.5950575,5.2250857,5.2854476,4.6214657,3.640583,4.247976,4.2706113,4.1197066,3.9386206,3.5990841,2.8521044,3.187868,3.9197574,4.606375,5.062863,5.8173876,6.8737226,7.17176,7.0284004,8.145098,8.062099,7.454707,6.8963585,6.7756343,7.3000293,7.8432875,7.360391,6.8850408,6.6662283,6.1720147,7.5565677,8.371455,7.5263867,5.9607477,6.651138,7.4773426,7.175533,6.368191,5.7117543,5.907931,5.2665844,5.1647234,5.311856,5.4401255,5.281675,6.4021444,7.2396674,7.4509344,6.9944468,6.138061,7.5565677,8.812852,10.084227,11.09529,11.09529,10.514306,9.556059,9.34102,10.061591,10.95193,12.064855,13.920986,14.977322,14.992412,15.01882,14.2944765,13.611631,13.890805,14.924504,15.365902,14.664193,14.053028,14.120935,13.611631,9.446653,9.439108,9.703192,10.11818,11.45369,15.380992,18.119919,19.60256,20.360857,20.545715,19.927006,23.303505,24.608833,23.895807,22.537663,23.216734,22.277351,20.168453,18.33873,18.316093,21.700138,21.081429,21.42851,20.43631,17.18808,12.170488,19.54597,21.779364,21.183289,17.520071,7.9715567,13.053283,13.124963,16.195879,22.858335,26.283878,21.277605,13.830443,9.774872,10.370946,12.30253,11.106608,10.834979,11.502733,12.294985,11.548005,10.812344,8.620448,10.208723,14.766054,15.411173,10.186088,8.948667,10.570895,12.434572,10.457717,6.9680386,8.627994,10.653893,10.774617,9.235386,7.1264887,6.058836,5.9003854,6.187105,6.1078796,7.092535,7.6395655,7.484888,6.7114997,5.7570257,5.6476197,5.3948536,4.406426,3.0520537,2.6634734,2.474842,2.3390274,2.4031622,2.8596497,3.9122121,4.0895257,4.0517993,4.3385186,4.696918,4.0782075,4.38379,4.2819295,4.08198,4.2328854,5.3156285,6.2851934,6.126743,5.80607,5.794752,6.0776987,6.7831798,7.91874,8.028146,6.9982195,6.0814714,6.4926877,6.7944975,7.115171,7.375482,7.2924843,7.8244243,8.028146,7.8131065,7.3377557,6.9793563,7.2057137,7.375482,7.9526935,9.005256,10.223814,9.955957,9.49947,8.382772,7.17176,7.466025,8.00551,8.2507305,8.4544525,8.854351,9.684328,9.250477,9.1976595,9.186342,8.646856,6.7643166,6.4474163,6.752999,7.2396674,7.3905725,6.6322746,6.277648,5.9117036,5.7494807,5.6551647,5.149633,5.0779533,5.0062733,5.0779533,5.2628117,5.3646727,5.311856,5.1835866,5.243949,5.458988,5.50426,5.715527,6.56814,7.24344,7.3188925,6.790725,6.3945994,6.0626082,5.8626595,5.828706,5.96452,5.9003854,5.847569,5.515578,4.749735,3.5538127,3.5953116,3.9461658,4.3611546,4.7308717,5.0779533,4.949684,4.8327327,4.7572803,4.7535076,4.8553686,4.8365054,4.6742826,4.678055,4.8629136,4.979865,4.696918,4.3649273,4.195159,4.2592936,4.485651,4.727099,4.991183,5.4891696,6.006019,5.904158,6.4436436,7.032173,7.575431,7.99042,8.20546,9.439108,10.0465,10.291721,10.374719,10.438853,9.465516,9.673011,10.487898,11.148107,10.676529,1.7391801,1.629774,1.5845025,1.6524098,1.8184053,2.0145817,2.0145817,1.931584,1.9579924,2.1164427,2.2748928,2.8332415,3.059599,3.1237335,3.2218218,3.5387223,3.2972744,3.482133,3.8782585,4.2291126,4.2404304,4.08198,3.92353,3.9688015,4.112161,3.9688015,4.5535583,4.9647746,5.111907,5.1232247,5.3571277,5.379763,5.413717,5.455216,5.485397,5.4476705,6.0701537,6.3531003,6.530414,6.9567204,8.103599,8.360137,7.9941926,7.4811153,7.277394,7.828197,8.390318,7.7716074,7.33021,7.541477,7.9791017,7.5905213,8.122461,9.654147,12.061082,15.015047,14.720782,22.805517,32.052223,37.91111,38.495865,36.485058,30.139502,22.307531,15.848798,13.626721,9.940866,7.1604424,4.878004,2.776652,0.6413463,0.5055317,0.21503963,0.0452715,0.041498873,0.0150905,0.0150905,0.0150905,0.026408374,0.06413463,0.1358145,0.24899325,0.9695646,0.9016574,0.090543,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.17354076,0.38103512,1.1242423,1.0940613,0.663982,0.20372175,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.026408374,0.06790725,0.090543,0.08677038,0.0754525,0.11317875,0.29426476,0.31312788,0.19994913,0.32067314,0.49044126,0.44139713,0.6752999,1.1393328,1.237421,1.5656394,1.7127718,2.0975795,3.2972744,6.058836,5.070408,4.45547,4.3686996,4.6856003,4.991183,4.696918,5.1458607,6.587003,8.695901,10.574668,7.4509344,6.8963585,7.605612,8.963757,11.0613365,13.822898,14.162435,14.083209,14.539697,15.456445,15.543215,15.573396,15.011275,14.060574,13.656902,10.740664,11.072655,11.962994,12.272349,12.404391,11.159425,11.268831,10.823661,9.797507,10.054046,11.276376,12.351574,13.102326,13.347548,12.909923,13.128735,13.494679,13.140053,12.306303,12.344029,13.577678,13.087236,12.272349,12.166716,13.472044,14.705692,16.048746,16.343012,16.177015,17.897333,19.180025,20.130728,20.572124,20.60985,20.658894,19.794964,19.493153,20.032639,20.904116,20.843754,20.1345,19.859098,19.715738,19.164934,17.395575,16.576914,17.23335,18.949896,21.043703,22.567842,20.749437,19.670467,19.146072,19.108345,19.621422,21.636003,23.039421,23.001694,21.632233,19.972277,18.65563,18.214233,18.331184,19.28566,21.971767,21.326649,22.069857,23.590223,24.888006,24.582424,20.760756,18.761265,18.225552,18.51227,18.708447,19.025349,18.059555,17.248442,17.21826,17.7917,16.41092,16.535416,16.607096,16.505234,17.516298,18.372684,18.23687,18.244415,18.61036,18.644312,18.463226,18.417955,18.259504,18.176508,18.79899,19.300749,19.810055,20.16468,20.123182,19.379974,19.915688,20.48158,21.122927,21.454918,20.658894,18.817854,18.135008,17.799244,17.297485,16.418465,16.969267,16.161926,14.7321005,13.664448,14.1926155,14.335975,14.1926155,14.215251,14.441608,14.464244,16.090246,17.237123,16.893814,15.724301,16.06761,16.335466,16.395828,13.087236,8.216777,8.560086,5.2628117,3.7084904,2.4031622,1.2449663,1.5241405,0.86770374,0.65643674,1.3204187,2.7728794,4.395108,6.2021956,8.118689,10.340765,12.672247,14.524607,14.283158,14.037937,13.600313,12.823153,11.627231,11.921495,12.038446,12.472299,13.3626375,14.509516,14.000212,13.302276,12.996693,13.034419,12.740154,11.800771,11.4838705,11.295239,10.7218,9.231613,8.096053,7.5565677,7.6282477,7.7338815,6.6850915,10.578441,10.725573,9.627739,9.190115,10.740664,13.185325,13.483362,13.196642,11.231105,3.8443048,1.9429018,3.9725742,6.6360474,7.4018903,4.5309224,5.142088,5.43258,5.010046,3.9348478,2.7011995,4.06689,3.3123648,2.444661,2.6898816,4.4705606,6.620957,10.38981,11.351829,9.665465,10.054046,10.774617,11.9064045,9.797507,5.6287565,5.4476705,8.096053,10.03141,10.884023,10.970794,11.276376,11.314102,9.831461,8.299775,7.7414265,8.744945,9.74469,9.06939,8.6732645,8.348819,5.7381625,7.3377557,8.82417,8.345046,6.5832305,6.790725,5.9984736,8.98262,7.4207535,1.5430037,0.1358145,0.10186087,0.071679875,0.049044125,0.033953626,0.0452715,0.0452715,0.06413463,0.11317875,0.21881226,0.42630664,0.452715,0.6149379,0.814887,0.88279426,0.56589377,0.44139713,0.4678055,0.59607476,1.0072908,2.1051247,3.2029586,3.8820312,4.2404304,4.3121104,4.044254,3.7386713,3.863168,3.7160356,3.2935016,3.2821836,4.2819295,4.878004,4.9119577,4.349837,3.3123648,3.6179473,3.9499383,3.8103511,3.3764994,3.5236318,2.6219745,2.7879698,3.3689542,4.002755,4.6252384,5.80607,6.379509,6.571913,6.8133607,7.707473,7.194396,7.1378064,7.254758,7.1906233,6.530414,7.3000293,7.281166,7.3679366,7.6395655,7.3717093,7.394345,7.4735703,7.0849895,6.4436436,6.530414,6.7379084,6.6360474,6.7756343,6.934085,6.1041074,5.5306683,5.4212623,5.534441,5.674028,5.723072,5.9532022,6.560595,7.194396,7.2358947,5.783434,7.0170827,8.971302,10.876478,12.1101265,12.208215,11.84227,10.310584,9.495697,9.876732,10.574668,11.747954,13.155144,14.5283785,15.580941,16.022339,15.471535,15.573396,16.72782,17.784155,16.03743,15.354584,15.282904,15.056546,14.283158,12.940104,10.11818,10.148361,11.581959,14.2077055,19.04421,20.628714,20.88148,19.983595,19.047983,20.111864,26.593233,26.29897,22.620659,18.968758,18.79899,18.531134,18.361366,18.063328,18.150099,19.881733,20.836208,23.578907,23.914669,19.859098,11.657412,17.384256,18.923487,20.474035,21.092747,14.709465,16.882498,13.215506,13.947394,19.312067,19.53088,16.822134,14.128481,11.506506,9.895596,11.155652,11.091517,11.378237,11.378237,11.170743,11.536687,11.766817,9.024119,9.676784,13.494679,13.641812,8.367682,6.043745,6.398372,8.529905,10.910432,9.714509,11.427281,13.113645,12.811834,9.552286,7.122716,6.587003,6.6020937,6.587003,6.7454534,7.466025,7.8998766,7.779153,7.0284004,5.783434,5.80607,5.5004873,4.447925,3.0181,2.3956168,2.5314314,2.3993895,2.3201644,2.6182017,3.6330378,4.1310244,4.2102494,4.5233774,4.881777,4.2706113,4.432834,4.719554,4.6818275,4.534695,5.1571784,5.3646727,5.828706,6.221059,6.3342376,6.1041074,6.63982,7.405663,7.454707,6.7039547,5.934339,6.670001,7.2358947,7.564113,7.6697464,7.643338,7.7301087,7.6886096,7.6018395,7.5905213,7.798016,7.5527954,7.6018395,7.748972,7.9791017,8.4544525,9.35611,9.397609,8.7751255,8.00551,7.91874,7.786698,8.035691,8.145098,8.280911,9.291975,9.329701,9.137298,8.98262,8.45068,6.4247804,5.8136153,6.1908774,6.3945994,6.228604,6.485142,6.277648,5.8702044,5.4665337,5.1760416,5.0062733,4.881777,4.659192,4.478106,4.3875628,4.3649273,4.98741,5.251494,5.3986263,5.5306683,5.613666,5.4438977,5.9682927,6.507778,6.6058664,6.058836,5.7909794,5.692891,5.4250345,5.160951,5.5985756,6.1003346,6.089017,5.613666,4.8742313,4.22534,4.191386,4.3083377,4.5535583,4.908185,5.372218,5.2628117,4.859141,4.504514,4.3913355,4.561104,4.610148,4.61392,4.6214657,4.6516466,4.7006907,4.5535583,4.52715,4.776143,5.1458607,5.1571784,5.0477724,5.485397,6.0739264,6.466279,6.3945994,7.3717093,7.8319697,8.137552,8.473316,8.865668,9.510788,9.967276,9.820143,9.374973,9.64283,8.937348,9.107117,9.7220545,10.321902,10.4049,0.8224323,0.8601585,0.9318384,1.0223814,1.1657411,1.4298248,1.6712729,1.7919968,1.7354075,1.6524098,1.8599042,2.0296721,2.2484846,2.4295704,2.5276587,2.565385,2.776652,3.138824,3.308592,3.3312278,3.6066296,3.7009451,3.591539,3.519859,3.531177,3.4896781,3.7952607,3.9801195,4.1536603,4.236658,3.9876647,4.1008434,4.5309224,4.851596,5.0062733,5.311856,5.7117543,6.1795597,6.537959,6.7944975,7.149124,6.6549106,6.511551,6.647365,6.990674,7.462252,8.09228,8.009283,8.424272,9.303293,9.371201,10.269085,12.50248,14.5283785,17.071129,23.118647,25.608578,26.90636,28.788902,29.539654,23.922215,21.470009,19.349794,15.652621,10.853842,7.8508325,5.172269,3.1840954,1.8184053,0.995973,0.6149379,0.56212115,0.4640329,0.2867195,0.10186087,0.124496624,0.663982,0.6149379,0.362172,0.16976812,0.17354076,0.44139713,0.62248313,0.56589377,0.3470815,0.2867195,0.14713238,0.05281675,0.00754525,0.0,0.0,0.0,0.00754525,0.018863125,0.041498873,0.10186087,0.42630664,0.513077,0.38480774,0.14713238,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0452715,0.090543,0.116951376,0.116951376,0.11317875,0.090543,0.30935526,0.3961256,0.35462674,0.56589377,0.5696664,0.362172,0.663982,1.3732355,1.5882751,1.1280149,1.0978339,1.6071383,2.7728794,4.7535076,5.247721,5.247721,5.160951,5.2779026,5.7570257,6.228604,6.4210076,7.5716586,9.537196,10.782163,8.956212,9.597558,9.703192,9.137298,10.661438,11.91395,13.132507,14.50197,15.667711,15.724301,16.376965,17.010767,16.84477,15.916705,15.082954,12.664702,11.966766,11.189606,10.314357,11.076427,12.789199,13.053283,12.513797,11.706455,11.057564,11.476325,12.242168,12.894833,12.958967,11.944131,11.861133,11.785681,11.151879,10.601076,11.966766,12.396846,12.272349,12.121444,12.253486,12.777881,14.030393,15.32063,15.437581,15.230087,17.60684,18.644312,18.561316,18.62545,19.25925,20.051502,20.160908,19.38752,19.240387,19.896824,20.194862,19.859098,18.444365,17.248442,16.65614,16.13929,15.456445,14.652876,14.996184,16.84477,19.651604,19.647831,19.436563,19.647831,20.085455,19.708193,20.530624,21.669958,22.428255,22.39053,21.41342,19.957186,19.266796,19.195116,20.104319,22.839472,21.666185,21.609596,21.934042,22.522572,23.88449,21.236107,20.013775,19.180025,18.534906,18.731083,19.36111,19.010258,18.150099,17.399347,17.523844,17.372938,17.320122,16.810818,16.150608,16.478827,17.901106,19.50447,20.394812,20.37972,19.97605,19.081938,18.184053,18.184053,19.123436,20.16468,20.560806,20.557034,20.8098,21.371922,21.722775,21.624687,21.526598,21.722775,21.937815,21.319103,18.931032,18.082191,17.542706,16.652367,15.343266,15.648849,15.230087,14.426518,13.5663595,12.970284,13.234368,14.022847,14.437836,14.147344,13.392818,14.068119,14.011529,13.083464,12.117672,12.917468,14.709465,15.992157,14.260523,10.4049,8.707218,7.9300575,7.375482,5.5193505,2.6898816,1.086516,0.72811663,0.9695646,1.6033657,2.4559789,3.3576362,5.3986263,7.3792543,9.525878,11.793225,13.890805,13.6682205,13.604086,13.917213,14.27184,13.800262,13.075918,12.479843,12.51757,13.170234,13.8870325,14.34352,14.4152,14.045483,13.400364,12.864652,11.495189,11.231105,11.268831,10.846297,9.231613,8.68081,8.001738,7.865923,8.469543,9.525878,12.543978,11.18206,10.144588,11.487643,14.649103,14.286931,12.121444,11.053791,10.446399,6.126743,3.9008942,5.0175915,7.8961043,10.242677,9.073163,6.3719635,4.606375,3.5047686,2.674791,1.5882751,1.8146327,2.8294687,3.7801702,4.508287,5.5570765,5.1873593,6.0626082,6.224831,5.8437963,7.213259,14.93205,21.134245,21.390783,15.286676,6.4134626,6.549277,7.5490227,8.050782,8.213005,9.737145,8.884532,8.786444,10.33322,11.864905,9.133525,9.25425,7.284939,5.564622,4.8629136,4.357382,6.952948,8.333729,9.110889,9.099571,7.3151197,6.3153744,4.4630156,2.637065,1.8448136,3.2142766,0.8526133,0.15467763,0.08299775,0.06790725,0.02263575,0.011317875,0.06413463,0.124496624,0.1961765,0.35462674,0.44516975,0.52439487,0.65643674,0.7507524,0.5394854,0.6149379,0.5017591,0.543258,0.87902164,1.4600059,2.2069857,2.7879698,3.3010468,3.7575345,4.104616,4.191386,3.942393,3.651901,3.399135,3.0746894,3.7914882,4.134797,4.274384,4.1800685,3.640583,3.350091,3.4594972,3.4330888,3.199186,3.1576872,2.8219235,3.0445085,3.3161373,3.6971724,4.817642,5.0439997,5.515578,5.624984,5.583485,6.436098,7.115171,7.564113,7.5527954,7.232122,7.141579,7.8696957,7.564113,7.356619,7.6622014,8.175279,8.190369,7.937603,7.537705,7.333983,7.8961043,7.039718,5.8966126,5.674028,6.326692,6.541732,5.6778007,5.3269467,5.3609,5.6589375,6.138061,6.319147,6.696409,6.670001,6.2097406,5.8211603,7.383027,8.89585,10.020092,10.552032,10.423763,11.4838705,10.868933,9.978593,10.016319,11.989402,13.026875,13.302276,13.641812,14.445381,15.716756,15.712983,16.641048,18.101055,18.964987,17.354074,16.946632,15.294222,13.679539,12.706201,12.340257,11.853588,13.015556,14.543469,16.052519,18.055782,19.90437,20.066593,20.093,21.654867,26.555508,36.1342,39.156075,35.609806,27.657114,19.60256,16.807045,16.429781,16.84477,17.40689,18.467,19.127209,20.934296,22.213217,20.828663,14.196388,15.792209,16.761772,17.863379,17.014538,9.303293,11.457462,10.608622,10.295494,10.963248,9.97482,10.729345,10.978339,10.608622,10.0276375,10.152134,10.257768,11.246195,11.751727,11.434827,10.948157,10.457717,8.831716,8.416726,9.431562,9.967276,7.779153,6.006019,6.126743,8.00551,9.895596,12.166716,13.298503,13.041965,10.914205,6.221059,5.8136153,6.017337,5.987156,5.692891,5.9494295,7.0246277,8.039464,7.997965,6.900131,5.73439,6.228604,5.330719,4.025391,2.9501927,2.3956168,2.1579416,2.323937,2.674791,3.078462,3.4859054,3.8178966,4.3121104,4.515832,4.3686996,4.187614,4.561104,4.557331,4.6214657,4.772371,4.5950575,4.5497856,5.221313,6.0211096,6.515323,6.40969,6.1833324,6.2323766,6.617184,6.990674,6.5832305,6.485142,6.3531003,6.3417826,6.7077274,7.828197,8.175279,8.179051,8.096053,7.7301087,6.3945994,6.8133607,7.3868,8.137552,8.688355,8.258276,8.439363,9.0543,9.073163,8.420499,8.00551,7.9791017,7.6848373,7.4509344,7.54525,8.171506,8.156415,8.397863,8.60913,8.401636,7.303802,5.824933,5.8173876,6.2097406,6.3229194,5.885295,5.7494807,5.6853456,5.4891696,5.194905,5.1043615,4.825187,4.429062,4.3611546,4.606375,4.719554,5.379763,5.7117543,5.885295,5.9682927,5.956975,6.0211096,6.349328,6.3342376,5.87775,5.3986263,5.168496,4.9534564,4.9232755,5.191132,5.80607,5.8702044,5.59103,5.111907,4.6629643,4.5799665,4.7874613,4.9232755,5.172269,5.4891696,5.59103,5.3458095,5.1269975,4.9421387,4.870459,5.0515447,5.413717,5.5306683,5.3948536,5.081726,4.749735,4.357382,4.357382,4.6629643,5.070408,5.2779026,5.4740787,5.674028,5.8437963,5.9607477,6.013564,7.1378064,7.8131065,8.692128,9.884277,10.978339,10.355856,10.170997,10.174769,10.253995,10.423763,9.405154,9.4013815,9.948412,10.487898,10.355856,0.6413463,0.69039035,0.72811663,0.7394345,0.7696155,0.8978847,1.0487897,1.237421,1.3241913,1.327964,1.4449154,1.5467763,1.7278622,1.8674494,1.9164935,1.9089483,2.2069857,2.5578396,2.7502437,2.7879698,2.9086938,2.8898308,2.9916916,3.1576872,3.2859564,3.2067313,3.4330888,3.610402,3.832987,3.9499383,3.5839937,3.6594462,3.8593953,4.093298,4.3083377,4.5007415,4.7421894,5.300538,5.7192993,5.9192486,6.217286,6.0248823,6.0286546,6.439871,7.1604424,7.816879,8.707218,9.084481,9.789962,10.808571,11.268831,12.6345215,14.973549,16.984358,19.097027,23.443092,22.786655,21.820864,22.522572,22.454664,14.777372,11.7894535,11.5857315,10.676529,8.14887,5.6778007,3.772625,2.4031622,1.4524606,0.97710985,1.20724,1.1619685,0.7997965,0.452715,0.29049212,0.33576363,0.69793564,0.7469798,0.70170826,0.66020936,0.60362,0.69039035,0.7432071,0.7507524,0.6828451,0.4979865,0.24522063,0.08299775,0.00754525,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.011317875,0.1056335,0.16222288,0.14335975,0.06790725,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.030181,0.08299775,0.11317875,0.116951376,0.13204187,0.14713238,0.22258487,0.27917424,0.3169005,0.43385187,0.40367088,0.4376245,0.6149379,0.94692886,1.4034165,0.935611,1.1657411,1.720317,2.3956168,3.199186,3.9763467,4.6026025,5.4363527,6.2399216,6.1720147,6.579458,6.8171334,7.9489207,9.782416,10.861387,10.925522,10.970794,10.144588,9.333474,11.144334,11.98563,13.045737,14.124708,15.086727,15.856343,16.950403,16.803272,15.882751,14.800008,14.317112,11.895086,11.295239,10.827434,10.269085,10.861387,11.887542,12.525115,13.038192,13.302276,12.789199,11.955449,12.434572,13.358865,13.853079,13.023102,13.147598,12.615658,11.69891,11.031156,11.615912,11.744182,11.981857,12.128989,12.208215,12.457208,14.468017,14.894323,14.562332,14.592513,16.414692,17.91997,18.51227,18.580177,18.704676,19.651604,19.628967,19.021576,18.448135,18.323639,18.817854,17.825653,16.143063,15.173498,15.181043,15.264041,15.437581,14.754736,14.649103,15.856343,18.4255,19.17248,19.274342,19.38752,19.583696,19.372429,19.398838,20.013775,20.832436,21.470009,21.537916,20.23636,19.523335,19.481836,20.50799,23.322369,21.224789,18.995167,18.334957,19.564833,21.624687,21.38701,21.002203,19.768555,18.202915,18.025602,18.38023,18.523588,18.65563,18.678267,18.18028,18.534906,18.987621,18.444365,17.237123,17.1164,17.557796,18.61036,19.568605,20.1345,20.383493,19.478064,18.331184,18.052011,18.957441,20.57967,20.794708,20.990885,21.651094,22.56407,22.820608,21.949133,21.360603,21.262514,21.41342,21.107838,19.168707,17.64834,16.444872,15.347038,14.003984,14.015302,13.7851715,13.754991,13.751218,13.004238,13.268322,13.902123,13.9888935,13.430545,12.940104,13.158916,13.532406,12.913695,11.570641,11.204697,13.781399,14.596286,13.102326,10.069136,7.5792036,6.3719635,7.0057645,6.149379,3.3161373,0.86770374,0.6828451,0.7054809,1.1053791,1.8372684,2.6295197,4.5120597,6.3229194,8.190369,10.269085,12.743927,14.215251,14.505743,14.34352,14.222796,14.396337,13.192869,12.276122,12.189351,12.7477,13.026875,14.245432,14.245432,13.513543,12.736382,12.785426,11.710228,11.099063,10.917976,10.604849,9.065618,8.575176,8.088508,8.548768,10.080454,11.970539,13.079691,11.966766,10.174769,9.261794,10.782163,11.359374,8.59404,7.1868505,7.2924843,4.5120597,3.4557245,4.6629643,7.3075747,10.397354,12.781653,8.367682,4.3347464,3.338773,4.715781,4.4705606,3.9612563,6.115425,8.394091,9.529651,9.556059,10.442626,11.940358,11.45369,9.06939,7.5603404,11.45369,16.437326,18.350048,15.282904,7.605612,5.828706,5.692891,5.621211,5.402399,6.221059,7.454707,8.047009,9.099571,10.091772,8.884532,7.8696957,6.549277,6.149379,6.307829,5.0553174,4.7308717,5.1835866,6.8473144,8.586494,7.7112455,5.621211,5.0439997,4.9534564,4.9685473,5.3458095,1.6939086,0.38858038,0.10186087,0.05281675,0.0150905,0.033953626,0.05281675,0.08299775,0.14713238,0.271629,0.34330887,0.3961256,0.452715,0.52062225,0.5696664,0.6488915,0.5055317,0.48666862,0.7054809,1.0412445,1.6863633,2.3163917,2.8822856,3.3123648,3.5349495,3.99521,3.8707132,3.5160866,3.108643,2.6182017,3.3764994,3.8858037,3.9914372,3.7688525,3.531177,3.2369123,3.0822346,3.0181,2.9539654,2.7653341,2.8106055,3.1727777,3.31991,3.4330888,4.398881,4.8440504,5.4250345,5.772116,5.828706,5.836251,6.1003346,6.507778,6.964266,7.375482,7.6584287,7.4207535,7.122716,7.1679873,7.5226145,7.726336,8.141325,8.09228,7.4773426,6.700182,6.673774,6.4021444,5.6023483,5.5457587,6.2097406,6.270103,5.3571277,4.983638,5.1798143,5.764571,6.3417826,6.730363,7.250985,7.352846,7.115171,7.2472124,7.8696957,9.250477,10.650121,11.472552,11.261286,10.933067,11.072655,11.121698,11.155652,11.876224,12.789199,13.015556,13.487134,14.392565,15.181043,15.105591,16.392056,18.135008,19.236614,18.406637,17.384256,14.434063,12.423254,12.298758,13.072145,12.853333,14.603831,16.637276,18.368912,20.315586,23.514772,25.129456,26.638506,30.479038,40.023777,58.973675,70.98194,70.265144,55.55945,30.12441,20.153362,16.124199,14.747191,14.422746,15.245177,16.878725,18.810308,20.8098,20.53817,13.521088,11.242422,12.408164,13.985121,13.151371,7.2924843,8.514814,9.167479,9.110889,8.529905,7.9413757,8.356364,9.288202,9.903141,9.940866,9.737145,9.590013,10.355856,11.034928,11.257513,11.287694,10.593531,9.4127,8.66572,8.699674,9.276885,7.2472124,6.0701537,6.1305156,7.4735703,9.835234,16.195879,16.161926,13.856852,10.823661,6.0286546,6.651138,7.1378064,6.8435416,5.983383,5.6061206,6.5756855,7.6207023,7.816879,7.0585814,6.0776987,6.2135134,5.194905,3.99521,3.1425967,2.7540162,2.2560298,2.2183034,2.584248,3.127506,3.4934506,3.712263,4.2894745,4.4894238,4.2819295,4.3385186,4.8402777,4.3875628,4.2404304,4.568649,4.45547,4.6516466,5.409944,6.043745,6.273875,6.2361493,6.043745,5.8890676,6.4210076,7.3151197,7.273621,7.5037513,6.722818,5.873977,5.8211603,7.3415284,8.114917,8.390318,8.345046,7.8131065,6.25124,6.692637,7.5603404,8.371455,8.918486,9.26934,8.933576,9.42779,9.58624,8.99771,8.009283,8.160188,7.6923823,7.284939,7.364164,8.118689,7.8432875,7.8131065,8.031919,8.228095,7.8508325,6.2814207,5.855114,6.0324273,6.2323766,5.855114,5.915476,5.8400235,5.7079816,5.5985756,5.583485,5.349582,5.0251365,4.9459114,5.1458607,5.3646727,5.515578,5.6325293,5.715527,5.7306175,5.613666,5.772116,6.0286546,6.047518,5.8173876,5.692891,5.2892203,4.9232755,4.7572803,4.8855495,5.3571277,5.6513925,5.553304,5.0666356,4.432834,4.164978,4.266839,4.3649273,4.5460134,4.7572803,4.8138695,4.6856003,4.617693,4.6214657,4.6856003,4.779916,5.036454,5.3344917,5.323174,5.0025005,4.715781,4.466788,4.678055,5.0666356,5.4401255,5.704209,5.855114,5.794752,5.8136153,5.885295,5.692891,6.6247296,7.8244243,9.092027,10.272858,11.257513,10.38981,10.03141,10.20495,10.631257,10.7218,9.857869,9.665465,10.035183,10.638803,10.933067,0.56589377,0.6451189,0.66020936,0.633801,0.6073926,0.6413463,0.663982,0.8186596,0.995973,1.1091517,1.1204696,1.2864652,1.4411428,1.5467763,1.5807298,1.5279131,1.780679,2.0975795,2.2862108,2.293756,2.1994405,2.1277604,2.3692086,2.6710186,2.8785129,2.9313297,3.078462,3.259548,3.4859054,3.5990841,3.270866,3.2972744,3.2482302,3.3651814,3.6783094,3.983892,4.3913355,4.8855495,5.251494,5.4967146,5.832478,6.2135134,6.2927384,6.730363,7.575431,8.269594,9.22784,9.903141,10.638803,11.536687,12.468526,13.36641,14.796235,16.052519,17.316349,19.640285,16.501461,17.05981,19.31584,19.210207,10.612394,7.232122,6.990674,6.952948,5.956975,4.6554193,3.4179983,2.425798,1.6373192,1.2034674,1.4864142,2.161714,1.4977322,0.7130261,0.4074435,0.5998474,0.5093044,0.62625575,0.7432071,0.7696155,0.72811663,0.8563859,1.0450171,1.0487897,0.8224323,0.5357128,0.2678564,0.090543,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.011317875,0.049044125,0.08299775,0.1056335,0.14335975,0.18863125,0.15467763,0.17731337,0.3055826,0.49421388,0.3169005,0.58098423,0.6149379,0.5357128,1.2449663,1.0336993,1.3091009,2.0372176,2.8143783,2.8936033,2.9841464,3.6066296,4.7233267,5.7079816,5.342037,5.5495315,6.387054,7.8319697,9.5032425,10.684074,11.102836,11.057564,10.374719,10.035183,12.181807,12.796744,13.992666,14.509516,14.554788,15.788436,16.478827,15.852571,14.418973,13.030646,12.90615,10.676529,10.661438,11.185833,11.344283,10.989656,11.0613365,11.751727,12.785426,13.59654,13.340002,12.098808,12.506252,13.577678,14.373701,13.973803,13.588995,13.113645,12.340257,11.521597,11.3820095,11.796998,12.083718,12.31762,12.623203,13.219278,15.00373,14.93205,14.456699,14.558559,15.754482,17.123945,18.18028,18.519815,18.4255,18.85558,18.214233,17.89356,17.380484,16.818363,17.010767,15.811071,14.347293,13.830443,14.332202,14.807553,15.675257,15.826162,15.814844,16.195879,17.523844,18.580177,18.912169,18.908396,18.795218,18.640541,18.048239,18.229324,18.919714,19.881733,20.92675,20.06282,19.640285,19.74592,20.598532,22.522572,19.036665,15.607349,15.067864,17.508753,20.258997,21.436056,21.609596,20.277859,18.28214,17.814335,17.787928,18.221779,19.112118,19.923233,19.595015,19.90437,20.043957,19.429018,18.384,18.142553,18.033148,18.127462,18.731083,19.700647,20.46649,19.998686,19.153618,19.029121,20.017548,21.820864,21.83218,21.94536,22.639523,23.58268,23.646814,21.824636,20.606077,20.160908,20.16468,19.772327,18.549997,16.859861,15.267814,14.060574,13.230596,13.113645,12.902377,13.241914,13.834216,13.456953,13.392818,13.385274,13.215506,13.000465,13.215506,13.068373,13.879487,14.094527,13.12119,11.34051,12.698656,13.147598,11.3669195,8.050782,5.885295,4.689373,5.9192486,5.934339,3.7688525,1.1091517,0.6828451,0.41498876,0.55080324,1.0450171,1.6071383,3.2520027,4.991183,6.741681,8.801534,11.853588,14.385019,14.841507,14.369928,13.936077,14.313339,12.966512,11.92904,11.721546,12.155397,12.313848,13.50977,13.313594,12.611885,12.132762,12.464753,11.578186,10.744436,10.220041,9.767326,8.66572,8.194141,8.379,9.125979,10.427535,12.377983,11.917723,12.140307,10.4049,7.5603404,7.960239,10.457717,8.831716,8.069645,8.744945,7.01331,4.647874,5.541986,6.5455046,7.454707,10.993429,7.7716074,4.044254,3.3915899,5.349582,5.406172,4.9987283,7.2962565,9.756008,11.046246,11.057564,13.88326,16.45619,16.056292,12.577931,8.544995,8.582722,10.47658,12.196897,12.306303,9.986138,7.5716586,6.5002327,5.7117543,5.0025005,5.036454,6.934085,7.0472636,6.9152217,7.3188925,8.280911,6.439871,5.6400743,6.79827,8.571404,7.3377557,4.2630663,3.651901,4.745962,6.2663302,6.4247804,6.820906,7.364164,6.6850915,5.5004873,6.6360474,2.0673985,0.44139713,0.07922512,0.02263575,0.00754525,0.030181,0.041498873,0.056589376,0.10186087,0.19240387,0.2263575,0.27917424,0.33576363,0.39989826,0.49044126,0.6073926,0.47535074,0.41121614,0.5470306,0.80734175,1.3505998,1.9429018,2.5389767,2.9841464,3.0143273,3.429316,3.3350005,3.0860074,2.8143783,2.4597516,3.2218218,3.8405323,3.8895764,3.561358,3.6594462,3.500996,3.059599,2.7540162,2.674791,2.5616124,2.8407867,3.1576872,3.169005,3.1199608,3.8895764,4.7308717,5.27413,5.8098426,6.1041074,5.4438977,5.2967653,5.6513925,6.307829,7.009537,7.4282985,6.651138,6.326692,6.670001,7.4584794,8.058327,8.458225,8.439363,7.6584287,6.462507,5.904158,5.8966126,5.696664,5.723072,5.938112,5.8588867,5.1835866,4.6629643,5.081726,6.187105,6.670001,7.4169807,8.084735,8.397863,8.465771,8.816625,8.446907,9.348565,11.00852,12.449662,12.23085,11.219787,11.631002,12.279895,12.528888,12.261031,12.536433,12.653384,13.422999,14.566105,14.7321005,14.898096,16.018566,17.497435,18.55377,18.225552,17.395575,14.724555,12.751472,12.359119,12.759018,13.577678,15.482853,18.240643,21.07011,22.639523,26.023567,29.158619,32.138992,37.254673,48.972446,74.52066,96.00199,97.86189,76.16175,38.62036,23.337458,16.746683,14.0983,13.030646,13.5663595,15.531898,17.644567,19.583696,19.15739,12.313848,8.182823,7.877241,8.959985,9.295748,7.0284004,7.911195,8.737399,9.024119,8.83926,8.790216,8.60913,9.567377,10.487898,10.774617,10.435081,9.937095,9.80128,10.170997,10.684074,10.484125,10.657665,10.087999,9.280658,8.703445,8.782671,6.6549106,6.349328,6.466279,6.6850915,7.748972,15.490398,16.324148,13.819125,10.280403,6.752999,7.33021,7.779153,7.4735703,6.5756855,6.0512905,6.375736,6.903904,7.062354,6.7680893,6.40969,6.4511886,5.3986263,4.2630663,3.5462675,3.2520027,2.7804246,2.4899325,2.5427492,2.938875,3.519859,3.6179473,4.168751,4.515832,4.5309224,4.640329,4.7874613,4.025391,3.8367596,4.4403796,4.779916,5.2590394,5.8626595,6.2097406,6.228604,6.1644692,6.085244,5.9796104,6.4247804,7.2094865,7.3415284,7.7225633,7.066127,6.221059,6.009792,7.213259,7.6508837,7.854605,7.9225125,7.6923823,6.749226,7.2472124,8.122461,8.756263,9.114662,9.759781,9.771099,10.110635,10.208723,9.691874,8.405409,8.186596,7.6320205,7.1604424,7.0585814,7.4773426,7.7112455,7.647111,7.7037,7.9828744,8.280911,7.0472636,6.217286,6.009792,6.1720147,5.9720654,5.983383,5.904158,5.828706,5.798525,5.798525,5.511805,5.323174,5.342037,5.511805,5.6023483,5.455216,5.383536,5.3609,5.3910813,5.515578,5.6589375,5.855114,5.945657,5.926794,5.9494295,5.413717,4.979865,4.678055,4.5912848,4.8629136,5.409944,5.5985756,5.1798143,4.4215164,4.08198,3.9499383,3.983892,4.074435,4.187614,4.3686996,4.346064,4.3686996,4.4441524,4.534695,4.5460134,4.666737,4.9685473,5.0025005,4.7610526,4.659192,4.7006907,5.0175915,5.4438977,5.9305663,6.537959,6.519096,6.0362,5.772116,5.7909794,5.534441,6.3531003,8.145098,9.725827,10.672756,11.306557,10.412445,10.038955,10.099318,10.378491,10.536942,9.95973,9.756008,10.114408,10.819888,11.231105,0.422534,0.52439487,0.56212115,0.56212115,0.5696664,0.63002837,0.62625575,0.69793564,0.8299775,0.94692886,0.91674787,1.1280149,1.2713746,1.3958713,1.4600059,1.3468271,1.5543215,1.8448136,1.9353566,1.7919968,1.6184561,1.5807298,1.7919968,2.022127,2.2069857,2.4559789,2.4899325,2.6106565,2.8143783,2.9728284,2.8445592,2.837014,2.806833,2.969056,3.399135,4.0517993,4.779916,5.1760416,5.481624,5.7909794,6.0324273,6.673774,6.790725,7.2094865,8.00551,8.477088,9.318384,10.125726,10.86516,11.615912,12.540206,12.777881,13.128735,13.45318,14.083209,15.841252,13.087236,16.686321,20.500444,19.515789,9.850324,6.2436943,5.093044,4.696918,4.2894745,4.0178456,3.2067313,2.3578906,1.6260014,1.2185578,1.388326,3.0407357,2.263575,1.0035182,0.39989826,0.7922512,0.3470815,0.392353,0.47157812,0.43385187,0.44516975,0.7884786,1.1280149,1.0676528,0.66020936,0.38858038,0.20749438,0.0754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.030181,0.00754525,0.018863125,0.049044125,0.094315626,0.150905,0.21503963,0.1961765,0.21881226,0.35839936,0.66020936,0.36594462,0.6413463,0.633801,0.44894236,1.1732863,1.327964,1.3770081,2.335255,3.7688525,3.8065786,3.0860074,2.9086938,3.1652324,3.5160866,3.3840446,3.7952607,5.4967146,7.2094865,8.507269,9.789962,9.310839,10.016319,10.676529,11.317875,13.245687,13.460726,14.8339615,15.290449,14.992412,16.31283,15.328176,15.026365,13.860624,12.162943,12.132762,10.18986,10.665211,11.857361,12.408164,11.268831,11.314102,11.5857315,12.147853,12.725064,12.702429,12.272349,12.728837,13.517315,14.1058445,13.9888935,12.815607,12.540206,12.068627,11.351829,11.378237,12.185578,12.23085,12.528888,13.385274,14.392565,15.169725,15.430037,15.241405,15.056546,15.712983,16.278877,17.006994,17.512526,17.621931,17.38803,16.403374,16.018566,15.660167,15.199906,14.973549,14.400109,13.585222,13.479589,14.094527,14.494425,15.32063,16.263786,16.708956,16.663685,16.780636,17.803017,18.168962,18.1086,17.82188,17.48989,16.524097,16.497688,17.093763,18.184053,19.859098,19.523335,19.4592,19.57615,19.862871,20.387266,16.222288,13.170234,13.705947,17.240896,20.145817,21.092747,21.651094,20.843754,19.123436,18.402864,18.251959,18.806536,19.727057,20.594759,20.900343,21.009748,20.270313,19.523335,19.149845,19.059301,18.949896,18.632996,18.94235,19.938324,20.915434,20.990885,20.775846,21.262514,22.582933,24.042938,23.669449,23.265778,23.567589,24.412657,24.718239,22.21699,20.26277,19.217752,18.749947,17.803017,17.048492,15.848798,14.396337,13.196642,13.068373,13.011784,12.766563,12.97783,13.539951,13.58145,13.396591,12.845788,12.600568,12.917468,13.664448,13.494679,14.483108,15.509261,15.513034,13.50977,12.0233555,12.291212,10.182315,6.0362,4.6516466,5.3910813,6.126743,5.794752,4.142342,1.720317,0.724344,0.32444575,0.271629,0.36971724,0.4640329,1.7580433,3.4934506,5.4250345,7.696155,10.853842,13.2607765,13.826671,13.690856,13.547497,13.619176,12.366665,11.472552,11.212241,11.465008,11.721546,12.261031,12.272349,12.113899,11.981857,11.883769,11.042474,10.303039,9.601331,8.850578,7.9451485,7.91874,8.805306,9.2995205,9.374973,10.295494,9.431562,10.4049,9.390063,6.971811,8.137552,11.291467,12.325166,13.355092,14.143571,12.083718,7.0963078,8.345046,8.20546,5.5570765,5.8098426,5.3080835,4.2894745,3.9876647,4.293247,3.7273536,3.92353,5.481624,7.0963078,8.194141,8.922258,11.691365,14.48688,14.762281,12.279895,9.14107,9.695646,8.880759,8.922258,10.416218,12.355347,10.223814,8.922258,7.779153,6.832224,6.8435416,7.2057137,6.096562,5.4665337,6.138061,7.77538,6.198423,5.5080323,6.8774953,9.21275,9.159933,5.8702044,5.191132,4.9232755,4.3385186,4.2064767,9.348565,9.216523,6.017337,3.5839937,7.383027,2.0145817,0.29803738,0.030181,0.0,0.0,0.0,0.030181,0.056589376,0.0754525,0.124496624,0.150905,0.1961765,0.30181,0.3961256,0.32821837,0.48666862,0.40367088,0.33953625,0.42630664,0.6790725,1.0601076,1.4977322,2.0900342,2.6710186,2.8143783,2.8936033,2.6408374,2.5540671,2.686109,2.6710186,3.2670932,3.7575345,3.7575345,3.5274043,3.983892,4.0103,3.3689542,2.6974268,2.372981,2.5125682,2.987919,3.0671442,2.8747404,2.8106055,3.5349495,4.538468,4.881777,5.3986263,5.8890676,5.111907,5.0062733,5.4778514,5.934339,6.1833324,6.4134626,6.085244,5.9305663,6.4474163,7.647111,9.0543,9.009028,8.6732645,7.877241,6.934085,6.598321,6.1418333,6.0814714,5.8664317,5.5570765,5.824933,5.406172,4.5912848,5.0138187,6.515323,7.149124,8.235641,8.873214,9.291975,9.593785,9.733373,8.9788475,9.107117,10.423763,12.064855,12.027128,11.827179,12.483616,13.407909,13.913441,13.226823,12.842015,12.604341,13.287186,14.437836,14.381247,15.275358,16.188334,17.199398,17.874697,17.274849,17.482344,16.580687,14.890551,13.0646,12.0724,14.524607,16.105335,19.130981,22.854563,23.48459,25.378448,29.652832,33.900806,38.75995,47.904793,70.91026,93.74219,94.87775,71.08757,37.443302,23.333685,17.308804,14.822643,13.6833105,14.04171,15.467763,17.380484,18.384,17.108854,12.234623,8.605357,5.8513412,5.2552667,6.40969,7.2094865,8.379,8.737399,9.084481,9.5183325,9.420244,9.827688,10.842525,11.781908,12.162943,11.676274,10.884023,9.737145,10.642575,12.479843,10.601076,10.386037,10.11818,9.691874,9.14107,8.639311,6.990674,6.9944468,6.7944975,5.828706,4.798779,10.133271,13.192869,12.396846,9.001483,7.069899,7.032173,7.2623034,7.284939,7.1038527,7.194396,6.651138,6.356873,6.126743,6.039973,6.439871,6.9227667,6.0248823,4.9459114,4.266839,3.9574835,3.6028569,3.1954134,2.806833,2.7313805,3.4934506,3.4783602,4.014073,4.5309224,4.8025517,4.938366,4.45547,3.7348988,3.7688525,4.5837393,5.240176,5.8211603,6.2889657,6.6586833,6.85486,6.700182,6.3417826,6.175787,6.3116016,6.617184,6.749226,6.7567716,6.8661776,6.9152217,6.937857,7.164215,6.9982195,6.937857,7.0774446,7.3075747,7.3075747,7.9451485,8.541223,8.926031,9.144843,9.431562,10.314357,10.608622,10.484125,9.982366,9.031664,8.182823,7.575431,7.0963078,6.6850915,6.326692,7.537705,7.748972,7.635793,7.7414265,8.477088,7.748972,6.779407,6.3153744,6.330465,6.0248823,5.6589375,5.7117543,5.7683434,5.7117543,5.7004366,5.3080835,5.119452,5.2665844,5.5268955,5.3344917,5.3646727,5.251494,5.1458607,5.2250857,5.6815734,5.832478,5.938112,5.938112,5.8588867,5.775889,5.2250857,4.8968673,4.644101,4.4743333,4.564876,5.062863,5.3948536,5.2062225,4.678055,4.5120597,4.1800685,4.1310244,4.1574326,4.22534,4.45547,4.4441524,4.425289,4.3686996,4.3007927,4.3121104,4.45547,4.644101,4.6327834,4.4705606,4.5309224,4.979865,5.2326307,5.5080323,6.017337,6.9567204,6.8963585,6.1041074,5.572167,5.572167,5.6363015,6.4926877,8.612903,10.291721,11.019837,11.46878,10.612394,10.382264,10.155907,9.899368,10.148361,9.782416,9.805053,10.359629,11.0613365,11.004747,0.45648763,0.44516975,0.41498876,0.422534,0.48666862,0.59607476,0.6187105,0.6526641,0.70170826,0.7582976,0.7922512,0.9280658,1.0525624,1.1506506,1.2110126,1.237421,1.4562333,1.629774,1.6222287,1.4713237,1.3732355,1.0940613,1.1317875,1.3505998,1.5656394,1.5430037,1.5543215,1.6109109,1.8674494,2.3088465,2.746471,2.6597006,2.9049213,3.289729,3.7462165,4.3347464,4.8968673,5.4740787,5.915476,6.1795597,6.3644185,6.5455046,6.7643166,7.4018903,8.22055,8.394091,9.333474,10.163452,11.0613365,11.808316,11.793225,12.796744,13.000465,13.585222,14.939595,16.648594,14.939595,19.327158,22.665932,20.240133,9.767326,5.934339,4.7912335,4.8025517,4.9345937,4.6554193,3.6669915,2.7879698,2.0673985,1.6335466,1.6939086,2.916239,2.2296214,1.0601076,0.3734899,0.7167987,0.35085413,0.13204187,0.15467763,0.31312788,0.27540162,0.32444575,0.47157812,0.44894236,0.25276586,0.1659955,0.1056335,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.041498873,0.090543,0.030181,0.02263575,0.056589376,0.1056335,0.150905,0.32444575,0.41121614,0.41876137,0.34330887,0.18485862,0.32821837,0.43007925,0.5281675,0.6375736,0.7469798,1.5543215,1.6825907,2.5917933,4.0970707,4.3800178,4.195159,2.7389257,1.539231,1.1996948,1.418507,2.848332,4.8063245,5.9607477,6.349328,7.3868,7.484888,8.122461,10.18986,12.864652,13.611631,13.475817,13.215506,14.166207,16.471281,19.059301,15.01882,15.16218,14.758509,13.000465,13.000465,10.559577,10.93684,11.736636,11.978085,12.098808,12.027128,11.661184,11.54046,11.921495,12.785426,13.81158,14.068119,14.007756,13.856852,13.611631,13.502225,12.283667,11.295239,11.148107,11.732863,12.00072,11.84227,12.449662,13.660675,13.917213,15.07541,16.244923,16.422237,15.652621,15.030138,15.309312,15.682802,15.596032,15.192361,15.290449,15.203679,13.936077,12.815607,12.46098,12.800517,12.996693,13.502225,14.32843,14.8339615,13.747445,13.539951,14.577423,15.83748,16.758,17.255987,17.429527,16.976812,16.233604,15.660167,15.852571,15.120681,15.0376835,15.467763,16.463736,18.297232,18.233097,18.025602,17.557796,17.176762,17.716248,15.9695215,13.728582,15.079182,19.032892,19.54597,19.54597,20.873934,21.45869,20.63626,19.134754,19.40261,20.055275,20.587215,20.73812,20.50799,20.911661,20.73812,20.326904,20.02132,20.157135,18.874443,18.693357,19.379974,20.723028,22.49239,22.80929,23.163918,23.876944,24.899324,25.800982,24.457928,23.7864,24.084438,25.12191,26.121656,24.107073,21.719002,19.63274,17.999193,16.448645,15.596032,14.841507,13.856852,12.898605,12.785426,12.800517,12.672247,12.611885,12.664702,12.725064,13.898351,13.43809,12.743927,12.577931,13.075918,14.139798,16.124199,17.191853,17.195625,17.686066,13.717264,12.370438,10.03141,6.5568223,5.247721,9.386291,8.345046,5.934339,3.9688015,2.2598023,0.8299775,0.30935526,0.23013012,0.2565385,0.18485862,0.5998474,2.022127,4.346064,6.858632,8.239413,10.570895,11.8045435,12.2119875,12.057309,11.581959,10.631257,10.453944,10.597303,10.7557535,10.819888,10.929295,11.872451,12.385528,11.993175,11.016065,10.8576145,10.370946,9.910686,9.107117,6.8359966,8.118689,8.6581745,9.042982,8.805306,6.4247804,6.6549106,5.0666356,3.5575855,3.6330378,6.379509,7.220804,12.079946,15.841252,15.184815,8.605357,5.9682927,11.793225,15.777118,13.43809,6.1041074,5.7872066,6.7680893,6.907676,5.6551647,4.044254,4.2517486,4.779916,5.406172,5.956975,6.2851934,4.749735,7.375482,8.028146,6.771862,9.87296,13.27964,10.257768,8.986393,11.038701,11.3669195,8.99771,8.820397,8.616675,8.054554,8.650629,8.114917,6.368191,5.794752,6.8359966,7.9941926,8.75249,9.2995205,8.7751255,7.484888,6.911449,6.5832305,8.431817,8.424272,6.013564,4.1197066,9.186342,9.544742,7.0246277,4.9421387,8.103599,2.1692593,0.27540162,0.0,0.0,0.0,0.0,0.0,0.030181,0.0754525,0.0754525,0.150905,0.15845025,0.20749438,0.29049212,0.29049212,0.21503963,0.27917424,0.3169005,0.33953625,0.5357128,0.814887,1.1695137,1.6222287,2.1654868,2.776652,2.9237845,2.674791,2.546522,2.6823363,2.8521044,3.1954134,3.4557245,3.350091,3.169005,3.7537618,4.266839,3.7273536,2.7615614,2.0485353,2.305074,3.169005,3.048281,2.7011995,2.6785638,3.3274553,4.398881,4.678055,5.093044,5.564622,4.991183,4.708236,5.2892203,5.726845,5.6287565,5.20245,6.058836,7.039718,7.798016,8.224322,8.469543,8.345046,7.7037,7.0057645,6.8058157,7.7225633,7.2924843,6.609639,5.975838,5.802297,6.6058664,5.9230213,4.9459114,4.7648253,5.73439,7.492433,8.66572,9.103344,9.865415,10.627484,9.673011,9.224068,9.046755,9.314611,9.9257765,10.514306,10.684074,12.804289,15.052773,15.656394,12.909923,13.373956,13.268322,13.392818,13.807808,13.856852,15.358356,17.05981,18.591496,19.1423,17.471025,17.923742,18.787672,17.833199,15.467763,14.709465,16.222288,16.791954,18.459454,21.202152,22.948877,22.888515,28.521046,34.040394,36.80573,37.36785,45.01119,49.02149,43.007923,30.120638,23.028103,19.338476,16.539188,14.434063,13.430545,14.543469,16.007248,17.463482,17.052265,15.067864,13.932304,12.049765,9.695646,7.6923823,6.6360474,6.8661776,7.5490227,8.152642,8.744945,9.016574,8.284684,9.774872,10.650121,11.529142,12.238396,11.812089,10.785934,9.4127,14.50197,22.171717,17.852062,10.759526,8.695901,9.914458,12.019584,11.947904,10.34831,8.209232,6.3644185,5.5306683,6.2851934,6.6058664,9.291975,10.306811,8.68081,6.5455046,6.4474163,6.379509,6.8133607,7.707473,8.514814,7.598067,6.692637,5.9607477,5.6325293,6.013564,6.9152217,6.9491754,6.3644185,5.5797124,5.20245,4.496969,4.0517993,3.3764994,2.7879698,3.4330888,3.410453,3.9348478,4.349837,4.561104,5.036454,4.436607,4.2064767,4.4177437,4.8855495,5.142088,5.6551647,6.6247296,7.7225633,8.484633,8.299775,6.983129,6.2135134,5.885295,5.885295,6.1041074,5.836251,6.379509,6.971811,6.9189944,5.5985756,6.4926877,6.832224,6.752999,6.700182,7.432071,7.6886096,7.7225633,7.828197,8.296002,9.446653,10.386037,10.336992,9.6051035,8.850578,9.0957985,8.544995,8.088508,7.605612,7.0585814,6.485142,7.5603404,7.564113,7.435844,7.6093845,8.024373,7.756517,7.4169807,7.164215,6.85486,6.013564,5.168496,5.3344917,5.6513925,5.772116,5.8588867,5.6513925,5.1156793,5.040227,5.3458095,5.0666356,5.5193505,5.4212623,5.2364035,5.1835866,5.2175403,5.621211,5.6589375,5.5306683,5.3986263,5.3873086,4.825187,4.878004,4.82896,4.515832,4.3347464,4.466788,4.666737,4.927048,5.0741806,4.745962,4.293247,4.134797,4.1762958,4.2592936,4.1498876,4.1498876,3.8480775,3.3840446,3.029418,3.187868,3.5047686,3.85185,4.002755,4.006528,4.164978,5.3269467,5.515578,5.240176,4.979865,5.1873593,5.50426,5.2175403,5.1156793,5.4778514,6.089017,6.8435416,8.616675,9.797507,10.148361,10.834979,10.612394,10.944386,10.789707,10.163452,10.103089,9.782416,10.227587,10.970794,11.3820095,10.650121,0.52062225,0.47912338,0.44516975,0.45648763,0.5357128,0.7054809,0.6790725,0.70170826,0.7205714,0.7507524,0.86770374,0.8639311,0.90543,0.98842776,1.056335,1.0035182,1.3317367,1.3619176,1.297783,1.237421,1.1883769,1.1431054,1.2336484,1.3317367,1.3845534,1.418507,1.4298248,1.4901869,1.6637276,1.9881734,2.4672968,2.6634734,2.8898308,3.0633714,3.199186,3.3953626,4.014073,4.8440504,5.6287565,6.319147,7.0585814,7.4094353,7.967784,8.639311,9.507015,10.868933,12.140307,12.396846,13.200415,14.317112,13.698401,14.11339,14.441608,14.151116,14.007756,16.097792,15.611122,15.83748,15.901614,14.117163,7.960239,6.432326,5.907931,5.8400235,5.7570257,5.300538,4.3611546,3.5160866,2.8558772,2.3465726,1.8523588,2.203213,1.7354075,0.9507015,0.38858038,0.6451189,0.33576363,0.116951376,0.049044125,0.08299775,0.06790725,0.09808825,0.16222288,0.1659955,0.10940613,0.08299775,0.049044125,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.049044125,0.07922512,0.094315626,0.071679875,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.02263575,0.07922512,0.18485862,0.26408374,0.181086,0.12826926,0.11317875,0.38858038,1.4222796,1.3091009,0.8865669,0.56589377,0.452715,0.35462674,0.52062225,0.6828451,0.87902164,1.2525115,2.0673985,1.720317,1.931584,2.5087957,3.5839937,5.613666,5.5759397,4.821415,3.610402,2.2975287,1.3468271,2.372981,3.7650797,4.61392,4.8968673,5.4438977,6.907676,8.20546,9.439108,10.665211,11.891314,13.70972,13.705947,13.936077,14.841507,15.260268,12.306303,15.39231,17.003222,15.354584,14.43029,13.970031,14.169979,13.543724,12.347801,12.577931,12.37421,11.947904,12.54775,13.7851715,13.615403,14.800008,14.675511,14.283158,14.290704,15.015047,13.860624,12.687338,11.830952,11.551778,12.049765,12.894833,12.928786,12.743927,12.785426,13.355092,14.3095665,15.264041,15.690348,14.984866,12.479843,12.181807,13.532406,14.569878,14.517061,13.762536,13.8719425,13.732355,13.336229,12.830698,12.498707,12.400619,12.804289,13.788944,15.007503,15.690348,15.509261,15.252723,15.414946,15.841252,15.70921,16.052519,15.901614,15.441354,14.939595,14.754736,15.01882,14.996184,15.158407,15.554533,15.792209,15.811071,16.946632,17.64834,17.523844,17.335213,15.316857,14.509516,15.430037,16.912678,16.116653,21.94536,21.624687,21.107838,21.813318,20.62494,20.560806,21.130472,21.82841,22.137764,21.545462,20.296722,20.560806,20.98334,21.058792,21.145563,20.040184,19.198889,19.210207,20.043957,21.062565,23.499681,24.654104,24.695602,23.963715,22.982832,24.012758,24.495655,24.091984,23.186554,22.888515,22.8357,22.315077,21.258741,19.670467,17.621931,15.546988,13.966258,12.619431,11.706455,11.921495,11.853588,11.92904,12.030901,12.053536,11.921495,12.272349,12.113899,11.706455,11.559323,12.4307995,13.675766,15.32063,16.343012,16.939087,18.549997,14.837734,12.381755,10.057818,7.835742,6.7643166,7.5527954,6.175787,4.315883,2.8558772,1.8787673,0.6752999,0.241448,0.271629,0.44516975,0.392353,0.6790725,1.841041,3.4745877,5.1458607,6.398372,8.141325,9.608876,10.269085,10.257768,10.397354,10.216269,9.993684,9.537196,9.035437,9.035437,10.484125,11.16697,11.408418,11.438599,11.419736,11.223559,11.351829,10.529396,8.661947,6.858632,10.299266,9.220296,7.454707,6.515323,5.583485,8.99771,10.612394,9.352338,6.5455046,5.9003854,8.4544525,7.364164,5.1798143,3.3350005,2.1353056,7.7225633,12.355347,11.77059,7.6131573,7.435844,11.84227,14.856597,13.053283,7.4094353,3.2859564,4.002755,6.092789,9.4013815,11.993175,10.144588,5.8702044,6.1908774,6.7756343,6.462507,7.2585306,7.960239,7.2585306,6.507778,6.1116524,5.534441,3.7801702,5.138315,6.85486,7.6697464,7.798016,10.110635,10.4049,9.288202,7.99042,8.348819,12.396846,11.898859,9.397609,7.0812173,6.790725,5.511805,6.1606965,7.9413757,9.771099,10.272858,8.209232,7.533932,6.4247804,5.0741806,5.6853456,5.873977,2.3993895,0.030181,0.0,0.0,0.0,0.0,0.026408374,0.06413463,0.06413463,0.08677038,0.1056335,0.13204187,0.181086,0.27917424,0.18485862,0.19240387,0.2678564,0.36594462,0.422534,0.65643674,0.8526133,1.1846043,1.7731338,2.655928,3.0746894,3.1539145,3.1916409,3.1916409,2.867195,2.8445592,2.8332415,2.9049213,3.127506,3.5575855,3.7990334,3.8782585,3.1614597,1.991946,1.6825907,2.4220252,2.6031113,2.5238862,2.5201135,2.9728284,3.2369123,3.4368613,3.9273026,4.534695,4.52715,4.859141,5.251494,5.511805,5.402399,4.5912848,5.4288073,6.5455046,7.7376537,8.262049,6.8435416,7.141579,7.5792036,7.424526,6.9265394,7.3075747,6.5568223,5.8966126,5.455216,5.2628117,5.240176,5.406172,5.028909,5.194905,6.221059,7.6886096,8.782671,9.024119,9.544742,10.223814,9.710737,10.412445,10.582213,10.487898,10.4049,10.612394,12.079946,13.106099,14.27184,15.154634,14.313339,14.784918,14.049255,13.792717,14.015302,12.989148,14.460471,16.807045,18.16519,17.912424,16.678776,17.157898,18.829172,19.40261,18.704676,18.640541,18.131235,18.082191,19.191343,21.605824,24.903097,25.174726,29.716967,32.59925,31.486328,27.653341,26.70264,24.60506,20.907888,16.939087,15.811071,15.045229,15.531898,16.614641,17.214487,15.833707,15.856343,15.863888,15.452672,14.471789,13.053283,11.955449,11.989402,10.49167,7.805561,7.3075747,8.213005,8.375228,8.575176,9.061845,9.529651,12.66093,15.147089,14.264296,10.585986,8.001738,9.593785,15.679029,18.116146,16.739138,19.33093,12.128989,9.435335,9.631512,10.616167,9.797507,9.167479,8.213005,7.435844,8.726082,15.39231,9.782416,9.597558,8.07719,5.1760416,7.5603404,7.118943,7.1981683,7.383027,7.5603404,7.914967,7.7716074,7.0359454,6.375736,6.039973,5.855114,6.228604,6.8774953,7.2094865,6.790725,5.349582,4.5912848,4.3083377,3.7575345,3.1840954,3.8103511,4.4516973,4.7610526,4.738417,4.5799665,4.6931453,5.119452,5.138315,4.817642,4.5007415,4.776143,5.172269,5.855114,6.8171334,7.6886096,7.752744,6.541732,5.9682927,6.1418333,6.609639,6.360646,5.8664317,6.436098,6.9189944,6.802043,6.2361493,6.541732,5.8928404,5.6023483,6.2361493,7.6131573,7.3905725,7.2887115,7.4697976,8.031919,8.993938,9.103344,8.907167,8.13378,7.405663,8.228095,8.929804,8.710991,8.258276,7.7942433,7.0963078,6.6058664,6.7114997,7.2962565,7.9791017,8.111144,7.8923316,7.1378064,6.7341356,6.719045,6.270103,5.50426,5.2552667,5.1232247,5.0439997,5.2854476,5.692891,5.304311,5.0477724,5.1269975,4.991183,5.4740787,5.696664,5.534441,5.168496,5.0968165,4.825187,5.0515447,5.3948536,5.6551647,5.836251,4.9723196,4.708236,4.346064,3.8254418,3.712263,4.3611546,4.7874613,4.991183,4.908185,4.3913355,4.183841,4.349837,4.3196554,3.9876647,3.712263,3.682082,3.6066296,3.4557245,3.31991,3.410453,3.6594462,3.942393,4.0706625,4.085753,4.274384,4.859141,5.292993,5.3344917,5.1156793,5.1269975,4.7421894,4.6742826,5.372218,6.537959,7.149124,7.3981175,7.8432875,8.122461,8.669493,10.699164,11.4838705,11.223559,10.280403,9.382519,9.623966,9.786189,10.544487,10.725573,10.246449,10.137043,0.6073926,0.52062225,0.51684964,0.513077,0.5357128,0.694163,0.6526641,0.6752999,0.694163,0.7054809,0.77338815,0.7696155,0.8337501,0.9016574,0.9620194,1.056335,1.2411937,1.2525115,1.1581959,1.0374719,0.9695646,1.0110635,1.0223814,1.1016065,1.237421,1.3241913,1.4109617,1.4713237,1.5845025,1.7957695,2.093807,2.2296214,2.4899325,2.8143783,3.1539145,3.4783602,4.1008434,4.7006907,5.3458095,6.058836,6.820906,7.696155,8.75249,9.691874,10.631257,12.121444,12.619431,12.808062,13.743673,14.886778,14.075664,14.656648,14.969776,15.441354,16.524097,18.689585,16.939087,13.588995,11.276376,10.321902,8.75249,7.911195,7.647111,7.4773426,7.1793056,6.828451,5.6589375,4.727099,4.002755,3.3878171,2.7238352,2.1692593,1.659955,1.0902886,0.6111652,0.6149379,0.30935526,0.1056335,0.02263575,0.018863125,0.00754525,0.02263575,0.05281675,0.056589376,0.041498873,0.041498873,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.041498873,0.08299775,0.14713238,0.17354076,0.0754525,0.03772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.018863125,0.06413463,0.14335975,0.21503963,0.20749438,0.32067314,0.60362,1.0223814,1.4449154,0.9393836,0.72811663,0.5281675,0.35085413,0.5055317,0.94692886,0.79602385,0.724344,1.0223814,1.5731846,2.5917933,2.8822856,3.6141748,5.1571784,7.1000805,6.375736,5.6891184,4.7912335,3.712263,2.7728794,2.9766011,3.5424948,3.8820312,4.055572,4.768598,6.25124,7.5188417,8.66572,9.767326,10.884023,12.098808,12.860879,13.490907,13.905896,13.645585,12.283667,14.188843,15.192361,14.317112,13.743673,14.290704,14.019074,13.558814,13.283413,13.328684,13.174006,13.347548,14.27184,15.282904,14.6302395,15.426264,15.082954,14.388792,14.045483,14.652876,14.471789,13.619176,12.7477,12.2270775,12.102581,13.034419,12.709973,12.185578,12.068627,12.555296,13.034419,13.2607765,13.804035,14.264296,13.27964,12.479843,13.641812,15.086727,15.679029,14.837734,15.245177,15.086727,14.222796,12.951422,11.989402,11.8045435,11.959221,12.555296,13.472044,14.351066,15.347038,15.422491,15.354584,15.252723,14.588741,14.588741,14.517061,14.196388,13.807808,13.849306,14.222796,14.388792,14.720782,15.226315,15.543215,15.584714,16.380737,17.18808,17.618158,17.618158,16.659912,15.792209,16.188334,17.463482,17.701157,21.100292,20.670212,19.715738,19.636513,19.915688,21.088974,21.560553,22.115128,22.854563,23.205416,22.481071,22.00195,21.813318,21.862362,21.986858,21.081429,20.417446,20.391039,21.062565,22.160398,23.171463,24.608833,24.963459,23.812809,21.820864,23.605314,24.586197,24.080666,22.496162,21.337967,21.375692,21.247423,20.4514,18.848034,16.659912,14.954685,13.947394,12.936331,12.030901,12.1252165,12.457208,12.306303,12.053536,11.951676,12.15917,12.464753,11.834724,11.34051,11.619685,12.898605,13.9888935,13.777626,14.124708,15.633758,17.640795,15.46399,13.306048,11.642321,10.31813,8.552541,7.647111,6.1078796,4.534695,3.1048703,1.5920477,0.6451189,0.32067314,0.30181,0.44516975,0.7997965,0.8941121,1.7014539,3.270866,4.9345937,5.311856,6.56814,8.145098,9.118435,9.5183325,10.329447,10.978339,10.612394,10.095545,9.971047,10.450171,11.189606,11.133017,11.00852,11.148107,11.4838705,10.933067,10.627484,9.782416,8.27714,6.673774,10.186088,9.982366,7.647111,4.851596,3.338773,7.805561,11.148107,11.54046,9.495697,7.888559,7.424526,4.9949555,3.380272,3.802806,5.956975,5.587258,6.009792,6.0814714,7.066127,12.608112,15.592259,14.705692,10.8576145,6.5643673,5.945657,6.971811,7.009537,8.160188,10.499215,12.061082,7.1038527,5.4212623,4.8440504,4.3875628,4.2630663,5.7306175,6.485142,5.975838,4.8402777,4.908185,5.696664,6.387054,7.5565677,8.488406,7.1793056,9.261794,10.499215,11.3971,11.69891,10.370946,10.933067,12.54775,12.510024,10.79348,10.0465,7.2887115,6.0512905,6.356873,7.2887115,6.9944468,6.4511886,5.8928404,4.927048,3.942393,4.1008434,4.22534,1.7240896,0.018863125,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.071679875,0.05281675,0.08299775,0.1056335,0.13958712,0.28294688,0.19994913,0.17731337,0.23013012,0.331991,0.41498876,0.5319401,0.60362,0.97333723,1.7089992,2.5804756,2.927557,3.0671442,3.229367,3.2746384,2.7238352,2.686109,2.704972,2.7389257,2.8445592,3.169005,3.289729,3.4179983,3.0030096,2.1579416,1.6524098,2.1277604,2.3993895,2.3956168,2.372981,2.9313297,3.1312788,3.3274553,3.4783602,3.62172,3.8782585,4.425289,4.5799665,4.772371,4.983638,4.7346444,5.5570765,6.511551,7.515069,7.9451485,6.63982,6.349328,6.971811,7.5188417,7.6395655,7.643338,6.8850408,6.119198,5.9796104,6.0626082,4.9534564,4.9345937,4.8327327,5.1232247,6.013564,7.443389,8.473316,8.707218,9.26934,10.106862,10.005001,10.246449,10.27663,10.023865,9.7296,9.948412,11.529142,12.898605,14.056801,14.8339615,14.894323,14.894323,14.449154,14.479335,14.750964,13.860624,14.694374,16.761772,18.33873,18.602814,17.640795,19.681786,20.130728,19.557287,18.848034,19.183798,18.565088,19.681786,20.458946,21.794455,27.570343,27.506208,26.412148,24.322113,21.824636,20.051502,18.92726,17.437073,15.7657995,14.18507,13.038192,15.490398,15.773345,16.090246,16.761772,16.222288,16.429781,14.3095665,12.989148,13.498452,14.792462,14.445381,12.506252,10.231359,8.590267,8.258276,7.4207535,6.9793563,7.4584794,8.865668,10.702937,11.876224,15.841252,17.380484,14.898096,10.419991,11.3669195,15.513034,16.437326,14.011529,14.369928,10.733118,9.42779,10.306811,11.962994,11.725319,8.933576,7.5829763,7.175533,10.012547,21.183289,24.880463,23.190327,15.46399,6.964266,8.884532,7.2170315,7.4094353,7.6207023,7.3490734,7.4471617,7.8621507,7.745199,7.3415284,6.9680386,7.001992,6.8435416,6.960493,7.066127,6.7869525,5.6325293,4.738417,4.938366,4.908185,4.3913355,4.1989317,4.938366,4.8100967,4.564876,4.5196047,4.5724216,5.0062733,5.2364035,5.142088,4.927048,5.142088,5.2099953,5.481624,6.0512905,6.7077274,6.9454026,6.7341356,6.537959,6.7454534,7.1981683,7.175533,6.7039547,6.8359966,6.964266,6.7680893,6.1908774,6.3644185,5.904158,5.9682927,6.670001,7.066127,7.383027,7.564113,7.8432875,8.303548,8.880759,8.254503,7.575431,6.900131,6.7077274,7.8998766,8.473316,8.465771,7.986647,7.3717093,7.164215,6.375736,6.3945994,7.073672,7.937603,8.160188,8.031919,7.2057137,6.5756855,6.300284,5.802297,5.4438977,5.1571784,4.9459114,4.908185,5.2250857,5.4476705,5.2854476,5.100589,5.0213637,4.9459114,4.90064,5.089271,5.251494,5.2137675,4.8742313,4.851596,5.2854476,5.8626595,6.277648,6.217286,5.5457587,5.0779533,4.5724216,4.146115,4.2706113,4.5233774,4.459243,4.266839,4.074435,3.9386206,3.942393,4.1083884,4.063117,3.8141239,3.7386713,3.8858037,3.7348988,3.4972234,3.3651814,3.519859,3.5538127,3.7348988,3.832987,3.9122121,4.3121104,4.919503,5.379763,5.6551647,5.745708,5.6891184,4.90064,4.8100967,5.43258,6.405917,6.9944468,7.0510364,7.360391,7.8810134,8.816625,10.627484,11.234878,10.804798,10.072908,9.64283,9.97482,10.7218,11.348056,11.2801485,10.680302,10.450171,0.6073926,0.55080324,0.56589377,0.5470306,0.52062225,0.6413463,0.5772116,0.60362,0.633801,0.6413463,0.6413463,0.7167987,0.8224323,0.88279426,0.9242931,1.0638802,1.1091517,1.1506506,1.1053791,0.995973,0.95824677,0.965792,0.9393836,1.0601076,1.2789198,1.3241913,1.3958713,1.4600059,1.50905,1.5807298,1.750498,1.8825399,2.2711203,2.7917426,3.3236825,3.7613072,4.3007927,4.6629643,5.292993,6.228604,7.115171,8.284684,9.442881,10.427535,11.291467,12.306303,12.23085,12.936331,14.019074,14.909414,14.890551,16.188334,16.957949,18.995167,21.737865,22.266033,20.081682,15.135772,11.374464,10.253995,10.748209,10.1294985,9.937095,9.563604,8.854351,8.088508,6.858632,5.926794,5.142088,4.349837,3.410453,2.3088465,1.7429527,1.2713746,0.7997965,0.58475685,0.36971724,0.23767537,0.14713238,0.07922512,0.018863125,0.0150905,0.03772625,0.041498873,0.030181,0.03772625,0.033953626,0.033953626,0.018863125,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.03772625,0.06790725,0.14335975,0.21881226,0.211267,0.13204187,0.056589376,0.0150905,0.0150905,0.018863125,0.018863125,0.0150905,0.011317875,0.00754525,0.00754525,0.00754525,0.011317875,0.05281675,0.10940613,0.116951376,0.32444575,0.76207024,0.995973,0.9318384,0.8186596,0.36594462,0.43007925,0.38858038,0.21503963,0.48666862,0.9205205,0.8601585,0.7582976,0.88279426,1.3166461,3.1652324,3.4255435,3.9801195,5.172269,5.824933,5.353355,5.221313,4.9949555,4.4894238,3.7877154,3.9650288,4.0178456,3.9650288,4.0895257,4.927048,6.1720147,6.9793563,7.8244243,8.790216,9.582467,10.035183,11.9064045,13.490907,14.007756,13.600313,13.253232,13.340002,13.245687,12.872196,12.626976,13.023102,12.498707,12.566614,13.502225,14.347293,14.362384,14.483108,15.067864,15.705438,15.192361,15.196134,15.015047,14.403882,13.758763,14.11339,15.116908,14.84528,13.81158,12.709973,12.415709,12.740154,12.559069,12.208215,12.012038,12.261031,12.042219,11.921495,12.298758,13.030646,13.422999,13.211733,14.456699,15.826162,16.573141,16.516552,16.852316,16.395828,15.245177,13.6682205,12.128989,11.868678,11.714001,11.627231,11.608367,11.710228,13.415455,14.505743,15.154634,15.271586,14.50197,14.200161,13.72481,13.102326,12.694883,13.189097,13.630494,14.034165,14.705692,15.414946,15.403628,15.475307,15.833707,16.422237,17.105082,17.670975,17.852062,16.98813,16.976812,18.361366,20.36463,21.277605,20.99843,19.591242,18.116146,18.614132,20.628714,21.519053,22.258488,23.288414,24.537153,24.544699,23.435547,22.22076,21.632233,22.111355,22.122673,21.843498,21.82841,22.409393,23.707176,23.507227,24.039167,24.061802,23.16769,21.813318,22.997923,23.737356,23.575134,22.57916,21.345512,20.394812,19.496925,18.52736,17.267305,15.4074,14.48688,14.283158,13.830443,13.124963,13.12119,13.404137,12.838243,12.219532,12.049765,12.543978,13.117417,12.166716,11.348056,11.446144,12.400619,13.008011,12.585477,13.268322,14.962231,15.365902,15.467763,13.687083,12.128989,11.272603,9.955957,8.729855,7.0472636,5.0553174,3.0369632,1.4034165,0.62625575,0.34330887,0.271629,0.422534,1.0978339,1.026154,1.7278622,3.308592,4.8402777,4.3800178,5.96452,7.4396167,8.409182,9.110889,10.416218,11.661184,11.548005,11.302785,11.555551,12.359119,12.106354,11.759273,11.676274,11.857361,11.940358,11.234878,10.597303,9.835234,9.1825695,9.310839,10.435081,9.473062,6.888813,3.7462165,1.7014539,4.6214657,7.756517,9.989911,10.623712,9.382519,7.8961043,5.764571,4.606375,5.0968165,6.952948,3.1840954,3.127506,5.2288585,8.575176,12.902377,12.0724,9.348565,7.066127,7.062354,10.691619,11.385782,8.20546,6.971811,9.544742,13.792717,9.465516,5.907931,4.315883,4.0216184,2.4861598,4.1197066,5.3759904,5.198677,4.2291126,4.798779,7.1981683,6.9755836,7.2094865,8.0206,6.587003,7.33021,8.692128,11.174516,13.215506,11.193378,8.756263,12.600568,15.509261,15.214996,14.426518,8.941121,6.304056,6.0022464,6.156924,3.5349495,5.798525,6.1720147,5.2967653,4.0178456,3.3689542,2.5276587,1.2449663,0.3169005,0.0,0.0,0.0,0.0,0.0,0.011317875,0.05281675,0.10186087,0.10940613,0.10186087,0.12826926,0.27917424,0.23013012,0.1961765,0.20749438,0.271629,0.392353,0.4678055,0.49044126,0.8601585,1.6260014,2.5012503,2.927557,3.0030096,3.1010978,3.097325,2.3616633,2.41448,2.5616124,2.546522,2.444661,2.6710186,2.6823363,2.7238352,2.5125682,2.082489,1.7655885,2.0749438,2.323937,2.3277097,2.3088465,2.8822856,3.169005,3.5387223,3.6669915,3.5764484,3.6594462,3.953711,3.9801195,4.247976,4.7308717,4.8553686,5.7796617,6.4964604,7.111398,7.3717093,6.63982,6.2399216,6.677546,7.3000293,7.699928,7.707473,7.062354,6.485142,6.273875,6.126743,5.149633,4.6516466,4.745962,5.2628117,6.0701537,7.0585814,7.854605,8.171506,8.756263,9.540969,9.661693,9.65792,9.691874,9.507015,9.337247,9.899368,11.129244,12.608112,13.8719425,14.68683,15.033911,15.049001,15.060319,15.199906,15.237633,14.611377,15.516807,17.463482,19.391293,20.455173,20.010002,21.851044,21.258741,19.94964,18.953669,18.629223,19.146072,21.05502,21.394556,21.4436,26.710184,25.944342,22.07363,18.078419,16.060064,17.255987,16.633503,16.475054,15.724301,14.694374,15.064092,18.02183,17.810562,16.150608,14.260523,12.872196,14.505743,12.332711,11.23865,12.875969,15.663939,17.135263,12.872196,9.699419,9.718282,10.306811,8.050782,7.798016,8.280911,9.276885,11.623458,10.631257,15.871433,19.957186,19.229069,13.762536,11.732863,13.019329,13.166461,11.117926,9.208978,8.635539,8.597813,10.846297,14.083209,13.970031,9.35611,7.9451485,7.7942433,10.7557535,22.484844,34.8251,32.493618,21.439827,10.091772,9.367428,7.352846,7.7942433,8.288457,7.9489207,7.4207535,7.9338303,8.231868,8.16396,7.9036493,7.967784,7.4584794,6.9454026,6.6586833,6.439871,5.7683434,5.0854983,5.617439,5.9003854,5.413717,4.61392,5.1081343,4.666737,4.3649273,4.534695,4.7535076,5.0779533,5.451443,5.7192993,5.8664317,6.0211096,5.9796104,5.87775,5.9532022,6.2625575,6.696409,7.4018903,7.443389,7.4018903,7.54525,7.84706,7.605612,7.3453007,7.1868505,6.971811,6.258785,6.198423,6.1644692,6.700182,7.4697976,7.2585306,7.7904706,8.0206,8.265821,8.560086,8.654402,7.654656,6.952948,6.620957,6.7831798,7.6282477,8.186596,7.9489207,7.424526,7.0548086,7.194396,6.4549613,6.5002327,7.0849895,7.786698,8.009283,8.009283,7.4207535,6.609639,5.783434,5.0138187,5.1760416,5.010046,4.825187,4.8553686,5.2779026,5.6363015,5.311856,4.8855495,4.6516466,4.6290107,4.357382,4.447925,4.745962,4.949684,4.5761943,5.119452,5.6778007,5.9984736,6.0362,5.9305663,5.7381625,5.330719,4.8440504,4.4818783,4.5309224,4.466788,4.063117,3.6179473,3.380272,3.5462675,3.651901,3.742444,3.7273536,3.6669915,3.7914882,4.032936,3.874486,3.5387223,3.2670932,3.3161373,3.3312278,3.3764994,3.3915899,3.5462675,4.221567,5.0251365,5.4288073,5.7872066,6.0739264,5.9003854,5.160951,5.0515447,5.3986263,6.017337,6.688864,6.8171334,7.273621,8.001738,8.929804,9.97482,10.155907,10.1294985,10.33322,10.801025,11.151879,11.374464,11.446144,11.3669195,11.133017,10.736891,0.55080324,0.58475685,0.59607476,0.56589377,0.5357128,0.6187105,0.5281675,0.5470306,0.59230214,0.6073926,0.55080324,0.7054809,0.80734175,0.8639311,0.8978847,0.91674787,0.935611,1.0223814,1.0714256,1.0676528,1.0751982,1.0336993,1.0487897,1.1959221,1.3958713,1.3920987,1.3392819,1.3996439,1.4034165,1.3619176,1.4939595,1.7165444,2.2447119,2.8219235,3.308592,3.6971724,4.2630663,4.644101,5.572167,7.0170827,8.190369,9.22784,9.982366,10.725573,11.529142,12.245941,12.31762,13.88326,15.045229,15.62244,17.180534,19.198889,20.474035,23.322369,26.529099,25.348267,25.276588,20.73812,15.62244,12.396846,12.08749,12.027128,11.917723,11.295239,10.084227,8.590267,7.4584794,6.579458,5.7117543,4.6856003,3.4217708,2.3503454,1.8448136,1.4071891,0.9205205,0.6451189,0.5583485,0.4640329,0.331991,0.17354076,0.05281675,0.026408374,0.041498873,0.05281675,0.0452715,0.0452715,0.060362,0.06413463,0.056589376,0.03772625,0.0150905,0.003772625,0.0,0.0,0.003772625,0.011317875,0.0452715,0.0754525,0.124496624,0.21503963,0.35839936,0.26408374,0.12826926,0.0452715,0.030181,0.03772625,0.041498873,0.033953626,0.026408374,0.02263575,0.02263575,0.030181,0.026408374,0.06790725,0.116951376,0.056589376,0.482896,1.0525624,0.9016574,0.20372175,0.15845025,0.21881226,0.38103512,0.33953625,0.20372175,0.48666862,0.754525,0.98842776,1.0299267,1.0978339,1.7693611,2.9539654,3.108643,3.1237335,3.1840954,2.7653341,3.308592,3.8858037,4.1574326,4.0291634,3.6481283,4.515832,4.5535583,4.395108,4.478106,5.0666356,6.2889657,6.692637,7.1868505,7.960239,8.446907,8.6581745,10.929295,13.075918,14.015302,13.800262,13.977575,13.241914,12.577931,12.37421,12.415709,12.015811,11.559323,11.778135,13.030646,15.30554,15.230087,15.00373,15.041456,15.343266,15.501716,14.735873,14.950912,14.852824,14.317112,14.392565,15.712983,16.007248,14.962231,13.407909,13.309821,12.600568,12.823153,12.849561,12.506252,12.562841,11.774363,11.936585,12.136535,12.189351,12.657157,13.321139,14.826416,15.852571,16.331694,17.4333,17.267305,16.920223,16.290195,15.241405,13.63804,13.087236,12.46098,11.638548,10.687846,9.869187,11.389555,13.174006,14.739646,15.55076,15.026365,14.728328,13.822898,12.770335,12.2270775,13.034419,13.573905,14.264296,15.184815,15.79598,14.973549,15.241405,15.611122,16.105335,16.758,17.625704,18.429274,17.972786,17.255987,17.686066,21.085201,22.382984,22.379211,20.772074,18.531134,17.908651,19.568605,21.05502,22.337713,23.526089,24.85028,25.182272,24.333431,22.741383,21.503962,22.382984,23.4695,23.329912,22.956423,23.107328,24.333431,24.340977,23.54118,22.60557,22.03213,22.167944,22.26226,22.31885,22.548979,22.714975,22.160398,20.394812,18.372684,16.97304,16.143063,14.905642,14.547242,14.811326,14.875461,14.634012,14.679284,14.241659,13.20796,12.408164,12.238396,12.66093,13.343775,12.543978,11.593277,11.170743,11.287694,11.517824,12.510024,13.792717,14.320885,12.487389,14.664193,13.181552,11.45369,10.872705,10.79348,9.680555,8.069645,5.402399,2.4295704,1.2034674,0.5696664,0.41121614,0.35462674,0.41876137,0.98465514,0.965792,1.780679,3.1425967,4.22534,3.6745367,5.904158,7.066127,7.91874,8.98262,10.54826,12.162943,12.679792,12.736382,12.872196,13.551269,12.940104,12.804289,12.917468,12.97783,12.608112,12.091263,11.491416,10.774617,10.695392,12.774108,11.2801485,7.8621507,5.032682,3.3312278,1.327964,2.7540162,4.610148,7.5226145,10.178542,9.307066,9.0957985,7.273621,4.927048,3.1048703,2.8181508,2.8596497,4.919503,7.1378064,8.167733,7.17176,3.983892,3.5085413,5.221313,8.733627,13.792717,13.400364,8.469543,7.1000805,10.917976,15.094273,12.064855,7.6584287,5.5495315,5.3344917,2.5578396,2.7200627,3.6028569,3.7575345,3.259548,3.7198083,5.9418845,5.492942,5.13077,5.696664,6.1342883,6.043745,6.937857,9.216523,11.563096,10.93684,8.182823,12.170488,15.543215,15.82239,15.399856,8.612903,6.2021956,7.0812173,8.126234,4.191386,6.1531515,7.0887623,6.4926877,4.817642,3.4557245,2.9501927,1.8297231,0.69793564,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.19994913,0.16222288,0.1056335,0.1358145,0.27540162,0.2678564,0.23390275,0.211267,0.23390275,0.33953625,0.452715,0.49421388,0.7922512,1.4637785,2.4107075,3.2105038,3.199186,3.0822346,2.9049213,2.0560806,2.0673985,2.2258487,2.233394,2.1051247,2.1768045,2.0258996,2.082489,1.9957186,1.7882242,1.8259505,2.082489,2.305074,2.3805263,2.4220252,2.7728794,3.0256453,3.561358,3.9914372,4.1197066,3.9310753,3.783943,3.7386713,4.1197066,4.749735,4.957229,5.9720654,6.466279,6.7039547,6.72659,6.356873,6.5002327,6.6360474,6.771862,6.960493,7.3188925,6.8435416,6.6586833,6.066381,5.270357,5.3609,4.610148,4.9421387,5.87775,6.8397694,7.1566696,7.484888,7.7829256,8.201687,8.669493,8.903395,9.125979,9.533423,9.593785,9.525878,10.344538,11.234878,12.117672,13.332457,14.649103,15.294222,15.777118,16.01102,15.848798,15.388537,14.962231,16.418465,18.274595,20.157135,21.688822,22.488617,22.33394,21.956678,21.100292,19.651604,17.644567,19.670467,21.651094,21.677504,20.730574,22.665932,20.843754,18.406637,16.558052,16.24115,18.127462,16.923996,16.078928,14.86037,14.694374,19.164934,19.440336,20.22127,18.678267,14.060574,7.7037,11.019837,10.729345,10.668983,12.3893,15.17727,19.466745,14.241659,10.416218,11.3669195,12.917468,11.046246,10.887795,10.4049,9.884277,11.925267,10.26154,14.754736,19.99114,21.802,17.30503,10.61994,10.47658,10.306811,8.299775,7.4018903,7.4584794,7.6622014,10.887795,15.218769,13.917213,10.023865,9.733373,10.220041,12.2119875,19.979822,32.806747,30.237589,20.485353,11.0613365,8.75249,7.6923823,8.461998,9.193887,8.971302,7.816879,8.013056,8.265821,8.443134,8.43559,8.137552,7.496206,6.7039547,6.2851934,6.2021956,5.836251,5.6551647,6.1418333,6.307829,5.824933,5.0213637,4.983638,4.496969,4.3196554,4.647874,5.1043615,5.492942,5.885295,6.3417826,6.790725,7.039718,7.164215,6.802043,6.470052,6.507778,7.0849895,8.20546,8.318638,8.00551,7.786698,8.118689,8.213005,7.828197,7.5565677,7.3868,6.6662283,6.307829,6.405917,7.149124,8.152642,8.43559,8.356364,8.390318,8.52236,8.586494,8.299775,7.322665,7.0057645,7.0170827,7.152897,7.33021,8.243186,7.5829763,7.1793056,7.4735703,7.5188417,6.888813,6.990674,7.33021,7.598067,7.673519,7.8395147,7.707473,6.952948,5.6778007,4.395108,4.7912335,4.8100967,4.7421894,4.8365054,5.292993,6.1041074,5.4438977,4.5460134,4.08198,4.134797,4.187614,4.3309736,4.508287,4.617693,4.504514,5.243949,5.6551647,5.462761,4.991183,5.172269,5.4174895,5.2854476,4.919503,4.478106,4.1197066,3.9989824,3.651901,3.2784111,3.0746894,3.2331395,3.308592,3.3727267,3.4029078,3.4594972,3.6443558,3.8405323,3.8178966,3.5236318,3.1010978,2.916239,3.059599,2.9841464,2.8936033,3.0822346,3.9461658,4.881777,5.281675,5.594803,5.8211603,5.5004873,5.194905,5.1458607,5.3646727,5.855114,6.617184,6.990674,7.4471617,7.99042,8.541223,8.937348,8.952439,9.57115,10.653893,11.740409,12.053536,11.068882,10.544487,10.567122,10.77839,10.382264,0.6111652,0.6828451,0.65643674,0.6187105,0.63002837,0.7167987,0.59607476,0.5998474,0.663982,0.68661773,0.56589377,0.6488915,0.6526641,0.70170826,0.7809334,0.73188925,0.7809334,0.91297525,1.0148361,1.026154,0.91674787,1.0148361,1.0374719,1.0940613,1.2223305,1.4034165,1.2336484,1.2826926,1.3355093,1.3241913,1.3128735,1.3845534,1.8787673,2.323937,2.6219745,3.0369632,4.123479,4.851596,6.1644692,7.960239,9.0957985,9.7296,9.914458,10.469034,11.710228,13.441863,14.0907545,16.28265,17.542706,18.119919,21.02484,22.918697,23.280869,23.922215,25.419947,27.128946,31.852272,28.373913,20.281631,12.332711,10.453944,11.710228,11.951676,11.204697,9.8239155,8.469543,7.149124,6.115425,4.9685473,3.7009451,2.7011995,2.2862108,1.9806281,1.5731846,1.1355602,1.0374719,0.8299775,0.5772116,0.331991,0.150905,0.0754525,0.041498873,0.041498873,0.0452715,0.0452715,0.0452715,0.071679875,0.0754525,0.13204187,0.18485862,0.0754525,0.026408374,0.00754525,0.0,0.0,0.0,0.060362,0.150905,0.211267,0.24899325,0.33576363,0.33576363,0.18863125,0.060362,0.011317875,0.0,0.02263575,0.030181,0.03772625,0.0452715,0.0452715,0.094315626,0.071679875,0.05281675,0.056589376,0.030181,0.35839936,0.23013012,0.09808825,0.10940613,0.120724,0.6111652,0.8526133,0.6752999,0.4376245,1.0374719,1.780679,1.3015556,0.9507015,1.2449663,1.8297231,1.9881734,2.1315331,1.9844007,1.9089483,2.897376,3.0822346,2.7238352,2.2296214,2.0749438,2.806833,3.663219,4.0216184,4.0291634,3.893349,3.904667,5.1873593,5.956975,7.3679366,9.107117,9.397609,8.83926,8.888305,9.842778,11.299012,12.178034,13.690856,12.887287,12.113899,12.528888,14.11339,13.468271,13.102326,12.83447,13.215506,15.546988,14.437836,15.580941,16.007248,15.501716,16.603323,15.79598,16.090246,16.697638,16.87118,15.8676605,16.320375,16.588232,16.320375,15.592259,14.909414,13.468271,12.83447,12.721292,12.842015,12.879742,12.31762,12.981603,13.679539,14.022847,14.449154,13.679539,14.019074,14.588741,15.294222,16.84477,16.11288,16.761772,17.36162,17.36162,17.105082,15.811071,14.260523,12.879742,11.846043,11.076427,12.2270775,13.355092,14.445381,15.135772,14.709465,14.68683,14.479335,13.837989,13.230596,13.837989,13.804035,14.928277,15.735619,15.7657995,15.596032,16.497688,16.81459,17.50498,18.478317,18.599041,19.60256,19.093256,16.331694,13.920986,17.77661,19.960958,21.368149,21.02484,19.43279,18.55377,19.055529,20.096773,21.73032,23.360094,23.726038,24.703148,25.269043,25.05023,24.540926,25.114365,25.56708,25.103046,23.759993,22.541435,23.405365,23.676994,23.29596,22.469755,21.70391,21.790682,21.764273,21.394556,21.405874,21.918951,22.432028,21.696367,19.519562,17.448391,16.150608,15.380992,15.245177,15.697892,16.222288,16.546734,16.633503,15.275358,13.758763,12.830698,12.611885,12.58925,12.736382,12.257258,12.098808,12.37421,12.37421,13.132507,13.962485,13.023102,10.804798,10.133271,12.815607,12.574159,12.14408,12.208215,11.3669195,9.171251,8.439363,6.1606965,2.4974778,0.76207024,0.482896,0.9507015,0.9507015,0.362172,0.16976812,0.7054809,1.4147344,2.2899833,3.2105038,3.9688015,5.406172,6.1531515,7.575431,9.756008,11.491416,13.551269,14.524607,14.532151,14.124708,14.283158,14.060574,13.79649,13.241914,12.570387,12.37421,12.193124,11.359374,10.612394,10.235131,10.038955,10.529396,6.971811,4.5120597,3.904667,1.50905,7.273621,8.99771,9.918231,10.502988,8.4544525,5.7306175,3.9688015,2.293756,1.0978339,2.0749438,5.7004366,3.410453,1.146878,1.1280149,1.8636768,1.690136,3.5877664,5.66271,7.284939,9.0807085,7.0774446,4.719554,5.775889,10.114408,13.702174,12.079946,9.876732,7.1868505,4.779916,4.1197066,3.180323,3.0897799,3.0256453,2.9011486,3.4029078,4.7950063,4.7044635,3.4444065,2.8521044,6.255012,7.122716,7.1302614,7.6848373,9.522105,12.694883,9.473062,10.114408,9.522105,6.9755836,6.1342883,5.5495315,6.1229706,7.6810646,9.099571,8.329956,5.4363527,4.5233774,3.6745367,2.9313297,4.2894745,4.5309224,2.2220762,0.38480774,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.211267,0.1659955,0.120724,0.17731337,0.33576363,0.3470815,0.3055826,0.26408374,0.26408374,0.35085413,0.4376245,0.48666862,0.77716076,1.4222796,2.3503454,3.6066296,3.572676,3.2821836,3.0331905,2.4107075,2.022127,1.8297231,1.9164935,2.0787163,1.8448136,1.4939595,1.7165444,1.8561316,1.7882242,1.9240388,1.9957186,2.323937,2.6483827,2.8219235,2.8219235,2.957738,3.1916409,3.5387223,3.9310753,4.2102494,4.063117,3.7273536,3.99521,4.919503,5.798525,6.530414,6.8133607,6.6624556,6.270103,6.0286546,6.198423,5.938112,5.907931,6.3531003,7.111398,6.937857,6.779407,6.089017,5.191132,5.2628117,4.776143,5.349582,6.760544,8.280911,8.68081,8.36391,8.239413,8.280911,8.526133,9.061845,8.646856,9.661693,9.997457,9.442881,9.673011,10.469034,10.774617,12.174261,14.611377,16.418465,16.77309,16.954176,16.490145,15.803526,16.218515,16.965494,17.38803,18.010511,19.534653,22.843245,22.111355,23.133736,22.398075,19.123436,15.290449,18.097282,20.930523,21.553007,20.357084,20.372175,16.878725,15.358356,16.301512,18.23687,17.701157,19.055529,16.014793,13.219278,13.830443,19.53088,16.026112,19.628967,24.17121,22.68102,7.3868,11.083972,11.578186,10.631257,10.880251,15.82239,22.733839,17.282394,12.638294,13.162688,14.418973,15.418718,12.559069,9.676784,8.98262,11.046246,10.242677,8.375228,14.373701,25.008732,24.888006,12.264804,8.322411,8.152642,8.918486,9.857869,8.379,8.103599,10.819888,13.856852,10.072908,10.38981,12.15917,14.109617,15.513034,16.218515,22.288668,19.466745,12.593022,6.8359966,7.6923823,7.960239,8.831716,9.175024,8.7600355,8.269594,8.073418,7.9451485,8.07719,8.246958,7.7829256,7.122716,6.205968,5.828706,6.066381,6.2851934,6.360646,6.4436436,6.228604,5.7419353,5.3269467,4.3611546,4.036709,4.2328854,4.738417,5.2628117,5.583485,5.798525,6.25124,6.9680386,7.673519,7.8961043,7.3905725,6.9755836,7.0246277,7.4773426,8.624221,8.892077,8.646856,8.27714,8.179051,8.5563135,8.2507305,7.9791017,7.8017883,7.0963078,6.9982195,6.779407,7.164215,8.265821,9.582467,8.397863,8.68081,8.8618965,8.495952,8.239413,7.5075235,7.0585814,6.820906,6.85486,7.356619,8.013056,7.6207023,7.8206515,8.605357,8.299775,8.167733,7.8961043,7.515069,7.220804,7.356619,7.745199,8.107371,7.9300575,6.8246784,4.515832,4.29702,4.5724216,4.9685473,5.2590394,5.3571277,5.832478,5.5570765,4.696918,3.8292143,3.953711,4.5007415,4.9949555,5.160951,5.089271,5.247721,5.040227,4.768598,4.5309224,4.5007415,4.927048,5.1232247,5.2364035,4.9987283,4.4139714,3.7537618,3.1916409,2.9426475,2.8634224,2.8521044,2.8521044,2.8521044,2.916239,2.9841464,3.0709167,3.2670932,3.4594972,3.5274043,3.31991,2.938875,2.7313805,2.7313805,2.6483827,2.5276587,2.625747,3.4330888,4.398881,4.961002,5.240176,5.2552667,4.9119577,5.1571784,5.1647234,5.402399,5.945657,6.470052,7.1302614,7.5226145,7.937603,8.375228,8.560086,8.729855,9.431562,10.061591,10.370946,10.469034,9.688101,9.235386,9.295748,9.514561,9.001483,0.84129536,0.94315624,0.8941121,0.875249,0.91297525,0.9016574,0.83752275,0.7394345,0.69793564,0.73188925,0.79602385,0.8903395,0.8903395,0.8978847,0.90543,0.7696155,0.84884065,0.8526133,0.8941121,0.94315624,0.84129536,1.026154,1.2298758,1.2298758,1.1280149,1.3317367,1.1317875,1.2600567,1.3694628,1.3770081,1.4713237,1.3505998,1.7429527,2.1579416,2.5201135,3.1576872,3.904667,5.353355,6.7152724,7.567886,7.8734684,8.692128,9.359882,10.03141,11.246195,13.905896,13.958713,15.667711,17.520071,19.059301,20.88148,19.15739,20.873934,22.394302,23.107328,25.419947,34.15735,31.535372,21.55678,10.963248,9.231613,12.276122,11.940358,10.265312,8.518587,7.175533,5.4665337,3.953711,2.7313805,1.8561316,1.3355093,1.1129243,0.95447415,0.7432071,0.59230214,0.8186596,1.3807807,0.9242931,0.4074435,0.20372175,0.10186087,0.08299775,0.0754525,0.056589376,0.041498873,0.08299775,0.06790725,0.049044125,0.07922512,0.12826926,0.08677038,0.041498873,0.011317875,0.0,0.003772625,0.02263575,0.094315626,0.15845025,0.17354076,0.16222288,0.18863125,0.16976812,0.150905,0.10186087,0.03772625,0.03772625,0.05281675,0.049044125,0.0452715,0.056589376,0.094315626,0.06413463,0.06413463,0.05281675,0.02263575,0.018863125,0.08299775,0.05281675,0.030181,0.071679875,0.18485862,0.7394345,0.47157812,0.43007925,1.0412445,2.1013522,1.2336484,0.8111144,1.0035182,1.4562333,1.2713746,1.4675511,1.8221779,2.1994405,2.2975287,1.6675003,2.0636258,2.1654868,2.1466236,2.3163917,3.0897799,4.293247,3.8782585,3.8254418,4.478106,4.52715,5.3609,7.1981683,8.892077,9.748463,9.533423,8.337502,8.348819,8.89585,10.269085,13.713491,14.9358225,14.456699,14.290704,14.750964,14.445381,14.215251,12.830698,12.189351,12.830698,13.913441,13.7700815,15.377219,16.0827,15.494171,15.490398,16.697638,17.572887,18.033148,17.889788,16.856089,17.135263,16.961721,16.580687,16.195879,15.98084,13.35132,11.815862,11.77059,12.657157,12.97783,13.166461,13.36641,13.819125,14.400109,14.634012,13.894578,13.924759,14.237886,14.596286,15.00373,15.324403,16.244923,16.882498,16.999449,16.995676,15.984612,14.554788,13.234368,12.14408,11.004747,12.238396,13.332457,14.396337,15.377219,16.052519,16.03743,16.607096,16.935314,16.675003,15.988385,15.471535,16.290195,17.37671,17.95015,17.486116,17.286167,17.21826,17.63325,18.4255,19.029121,20.066593,19.327158,17.255987,14.916959,13.981348,17.191853,20.002459,20.647577,19.455427,18.859352,20.055275,21.34174,22.7527,24.031622,24.642786,24.963459,25.25018,25.32186,25.468992,26.434784,25.92925,25.042685,23.695858,22.398075,22.24717,22.058538,21.53037,21.307787,21.390783,21.14179,21.420965,21.439827,21.23988,21.171972,21.869907,22.111355,21.371922,19.621422,17.286167,15.260268,15.241405,15.701665,16.248695,16.603323,16.569368,15.245177,13.536179,12.366665,12.083718,12.4307995,12.419481,11.978085,12.00072,12.551523,12.864652,14.381247,15.124454,13.20796,9.869187,9.473062,11.427281,11.966766,11.099063,9.420244,8.107371,8.850578,8.763808,6.1116524,2.0975795,0.8601585,0.65643674,0.73566186,0.6526641,0.41121614,0.44894236,0.8978847,1.7995421,2.546522,3.0709167,3.8556228,5.142088,6.1833324,7.8696957,10.133271,11.955449,12.755245,13.04951,12.347801,11.925267,14.807553,14.471789,13.736128,12.585477,11.355601,10.740664,10.899114,10.1294985,10.242677,11.11038,10.661438,8.612903,5.1798143,2.6031113,1.4826416,0.7922512,2.2371666,2.9916916,4.3083377,5.5495315,4.195159,1.9693103,1.5618668,1.9240388,3.5123138,8.288457,9.314611,6.8774953,4.0517993,2.3616633,1.7769064,2.5804756,3.8292143,4.195159,3.8292143,4.353609,5.4665337,4.979865,5.4891696,7.54525,9.650374,6.560595,5.847569,4.90064,3.3576362,3.1199608,2.5691576,4.425289,5.5759397,4.9534564,3.500996,4.044254,5.1647234,5.5797124,5.379763,6.0626082,6.2927384,5.2099953,4.285702,4.459243,6.126743,5.6098933,5.9532022,6.33801,7.277394,10.612394,8.152642,7.6320205,7.3717093,6.587003,5.3759904,3.470815,2.3126192,2.3654358,3.1576872,3.2633207,2.033445,0.77338815,0.10940613,0.049044125,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.14335975,0.13204187,0.1659955,0.29049212,0.4074435,0.38103512,0.30181,0.23767537,0.24899325,0.362172,0.33953625,0.4074435,0.6752999,1.2600567,2.263575,3.3764994,3.2482302,3.0935526,3.2746384,3.2784111,2.7200627,2.1956677,2.0636258,2.1353056,1.6863633,1.2864652,1.3128735,1.4826416,1.6410918,1.7655885,1.8561316,2.1692593,2.6446102,3.029418,2.8822856,3.6330378,3.8593953,4.236658,4.659192,4.236658,4.002755,3.5877664,3.8178966,4.8629136,6.25124,6.085244,5.674028,5.7306175,6.255012,6.5266414,5.847569,5.670255,5.6853456,5.8136153,6.205968,5.451443,5.5683947,5.855114,5.9984736,6.0701537,5.6287565,5.836251,6.9755836,8.386545,8.439363,8.903395,8.75249,8.820397,9.122208,8.869441,8.209232,8.89585,9.314611,9.397609,10.612394,11.740409,11.793225,12.887287,15.052773,16.233604,16.637276,16.72782,16.87118,16.863634,15.950659,16.109108,16.13929,15.871433,16.26756,19.398838,21.058792,22.009495,21.013521,18.19537,15.056546,16.644821,18.69713,20.243906,20.866388,20.711712,17.818108,16.897587,16.437326,16.007248,16.260014,17.84829,15.584714,15.433809,16.94286,13.268322,11.133017,17.73511,23.19787,20.52308,5.59103,8.605357,10.710483,10.578441,10.702937,17.372938,20.474035,17.87847,14.324657,11.510279,8.122461,8.624221,8.280911,8.171506,8.7600355,9.876732,10.231359,9.850324,17.554024,31.471237,39.03535,17.16167,8.733627,7.1038527,8.126234,10.148361,7.5188417,6.617184,9.110889,12.208215,8.68081,6.3417826,6.5945487,7.6320205,8.533678,9.250477,10.767072,10.906659,9.265567,7.6622014,10.155907,9.778644,9.2844305,8.9788475,8.850578,8.526133,8.243186,8.179051,7.84706,7.333983,7.2698483,7.333983,6.356873,5.7494807,6.039973,6.8850408,6.930312,6.983129,6.48137,5.583485,5.1798143,4.5460134,4.247976,4.6516466,5.406172,5.4212623,5.975838,6.1342883,6.458734,6.9869013,7.2358947,7.2396674,7.4018903,7.432071,7.375482,7.6093845,8.699674,9.450426,9.676784,9.446653,9.107117,8.75249,8.458225,8.175279,7.748972,6.911449,7.1868505,7.567886,8.137552,8.899622,9.789962,8.311093,8.235641,8.345046,8.209232,8.179051,7.6810646,6.937857,6.541732,6.7379084,7.466025,8.22055,8.797762,9.167479,9.295748,9.118435,9.14107,8.386545,7.7037,7.360391,7.0849895,7.533932,8.058327,7.877241,6.749226,4.979865,3.9876647,4.496969,4.983638,4.983638,5.0515447,5.2628117,4.5196047,3.8820312,3.85185,4.353609,4.2592936,4.496969,4.610148,4.5799665,4.847823,4.217795,4.2517486,4.4743333,4.817642,5.624984,5.372218,4.90064,4.436607,4.0480266,3.682082,3.6443558,3.5424948,3.2670932,2.927557,2.8407867,2.8709676,2.7653341,2.6144292,2.5389767,2.704972,2.7540162,2.7917426,2.674791,2.425798,2.2183034,2.2107582,2.1541688,2.1843498,2.41448,2.957738,3.610402,4.2894745,4.7610526,4.9949555,5.1835866,5.3571277,5.323174,5.4665337,5.8513412,6.25124,6.937857,7.3113475,7.432071,7.4509344,7.594294,8.654402,9.669238,10.38981,10.582213,10.016319,9.431562,9.963503,10.201178,9.639057,8.695901,0.87147635,0.90920264,0.875249,0.8941121,0.9695646,0.9808825,1.0148361,0.8865669,0.8299775,0.8865669,0.90920264,0.935611,0.91297525,0.9280658,0.95447415,0.87147635,0.91297525,1.0072908,1.116697,1.1657411,1.0525624,1.0412445,1.1355602,1.1129243,1.0035182,1.0940613,1.1204696,1.1959221,1.3920987,1.6184561,1.629774,1.569412,1.8485862,2.1503963,2.4371157,2.9803739,3.953711,5.5457587,6.587003,6.8737226,7.175533,8.201687,9.235386,10.442626,11.947904,13.822898,14.464244,16.750456,18.365139,18.776354,19.251705,17.987877,19.327158,20.575897,21.38701,23.75622,33.28587,31.72023,22.598024,12.3289385,10.197406,11.491416,10.555805,8.820397,7.1340337,5.7607985,3.8971217,2.3993895,1.3656902,0.8299775,0.72811663,0.73188925,0.66020936,0.5055317,0.43007925,0.76207024,1.2789198,0.83752275,0.3470815,0.16222288,0.09808825,0.12826926,0.13958712,0.116951376,0.08299775,0.08299775,0.049044125,0.02263575,0.030181,0.05281675,0.03772625,0.018863125,0.003772625,0.0,0.003772625,0.011317875,0.041498873,0.124496624,0.16976812,0.15845025,0.1358145,0.10940613,0.14335975,0.116951376,0.0452715,0.071679875,0.049044125,0.03772625,0.041498873,0.049044125,0.060362,0.026408374,0.030181,0.026408374,0.00754525,0.00754525,0.00754525,0.003772625,0.011317875,0.049044125,0.116951376,0.36594462,0.19240387,0.31312788,0.8299775,1.2110126,1.297783,1.2713746,1.5467763,1.8033148,0.9997456,1.3392819,1.9730829,2.4597516,2.4974778,1.9353566,2.2975287,2.2447119,2.022127,2.0145817,2.727608,3.9914372,4.2706113,4.6629643,5.240176,5.05909,5.243949,5.9607477,6.651138,7.224577,8.084735,7.375482,7.424526,8.088508,9.273112,10.933067,12.868423,13.766309,13.804035,13.513543,13.758763,13.600313,12.913695,12.623203,13.0646,13.981348,13.947394,16.59955,17.440845,15.83748,15.030138,16.233604,17.80679,18.889534,19.040438,18.229324,18.119919,17.248442,15.901614,14.867915,15.445127,13.890805,12.4307995,11.736636,11.940358,12.615658,13.483362,13.585222,13.604086,13.721037,13.58145,14.203933,14.656648,14.679284,14.600059,15.328176,15.23386,15.848798,16.358103,16.58446,17.003222,16.422237,14.822643,13.151371,11.834724,10.774617,11.638548,12.645839,13.502225,14.305794,15.528125,16.4826,17.976559,18.542452,17.942604,17.191853,16.867407,17.18808,18.082191,18.976303,18.772581,18.53868,18.599041,18.689585,18.787672,19.134754,20.689075,18.444365,16.490145,15.411173,12.31762,16.324148,19.36111,20.66644,20.225042,18.772581,19.429018,20.68153,22.567842,24.601288,25.778347,25.891525,25.948114,25.71044,25.506718,26.223516,25.00496,23.695858,22.567842,21.820864,21.564325,20.723028,20.345766,20.628714,21.38701,22.050993,22.367893,22.33394,22.005722,21.820864,22.590479,23.031876,22.805517,21.65864,19.595015,16.886269,15.958203,16.086473,16.403374,16.35433,15.686575,14.603831,13.181552,11.951676,11.348056,11.721546,11.891314,11.732863,12.053536,12.815607,13.140053,15.056546,14.954685,12.936331,10.521852,10.661438,12.453435,12.913695,11.136789,8.348819,7.914967,9.310839,8.13378,5.1232247,2.3277097,3.1010978,4.1272516,2.746471,1.1581959,0.66020936,1.6448646,1.4071891,1.871222,2.5767028,3.3576362,4.3347464,5.198677,6.428553,7.594294,8.314865,8.2507305,8.578949,9.148616,9.276885,9.480607,11.46878,11.446144,10.842525,10.884023,11.578186,11.68382,10.148361,10.306811,10.035183,8.778898,7.5301595,5.292993,3.1765501,1.7467253,1.0223814,0.44516975,0.94315624,1.1996948,1.871222,2.7917426,2.9539654,3.5877664,3.5500402,2.848332,2.927557,6.647365,8.782671,8.627994,6.809588,4.3385186,2.625747,2.9841464,3.682082,3.5990841,2.927557,3.1539145,5.1571784,5.66271,5.089271,4.3121104,4.6554193,5.13077,5.73439,4.6327834,2.4823873,2.4295704,2.1956677,3.3689542,4.7120085,5.3080835,4.5233774,4.889322,5.1798143,5.836251,6.6020937,6.507778,5.3948536,3.8405323,3.783943,4.7535076,3.863168,3.531177,3.8480775,4.561104,5.764571,7.8998766,7.1868505,7.7904706,7.5565677,5.9305663,3.9612563,2.8936033,1.7844516,1.9542197,2.9803739,2.686109,4.112161,2.5314314,0.8224323,0.15467763,0.0,0.0,0.071679875,0.124496624,0.120724,0.056589376,0.1056335,0.1056335,0.15845025,0.271629,0.34330887,0.38103512,0.3961256,0.3470815,0.28294688,0.33953625,0.3470815,0.3961256,0.543258,0.9393836,1.8033148,2.916239,2.776652,2.5880208,2.7125173,2.6898816,2.3465726,2.1051247,2.0560806,2.003264,1.4750963,1.2185578,1.2713746,1.4901869,1.690136,1.659955,1.5882751,1.9655377,2.4484336,2.7691069,2.7238352,3.3048196,3.6254926,4.29702,5.0515447,4.745962,4.3724723,4.1612053,4.1574326,4.5497856,5.6778007,5.402399,5.1798143,5.4212623,6.0701537,6.598321,6.571913,6.1116524,5.553304,5.243949,5.541986,5.2628117,5.1760416,5.191132,5.2892203,5.5382137,5.7796617,6.3719635,7.224577,8.0206,8.213005,8.790216,8.597813,8.624221,9.084481,9.431562,9.239159,9.578695,9.718282,9.812597,10.902886,11.740409,11.898859,13.011784,14.969776,15.950659,16.309057,16.278877,16.637276,17.025856,15.958203,15.558306,15.731846,15.128226,14.698147,17.697384,20.590988,21.590733,20.458946,17.886015,15.482853,14.554788,15.411173,17.025856,18.45568,18.840488,17.840744,17.56157,17.123945,16.678776,17.365393,15.577168,13.287186,14.200161,16.735365,14.019074,14.407655,17.72002,20.225042,18.059555,7.220804,9.507015,10.269085,10.020092,10.887795,16.607096,17.395575,15.916705,13.626721,11.2650585,8.843033,8.379,8.484633,8.869441,9.250477,9.344792,10.702937,10.797253,15.30554,23.45441,28.02683,12.234623,6.9454026,6.9944468,9.756008,15.147089,11.570641,7.9489207,7.2698483,8.409182,6.115425,5.2590394,5.745708,6.119198,6.096562,6.5455046,6.9982195,7.424526,7.8395147,8.597813,10.38981,10.487898,9.842778,9.352338,9.092027,8.296002,7.6848373,7.7640624,7.6697464,7.213259,6.8850408,6.477597,6.1342883,6.0211096,6.296511,7.1340337,7.092535,6.9454026,6.319147,5.402399,4.98741,4.504514,4.5724216,5.1873593,5.824933,5.4438977,5.907931,6.2399216,6.4549613,6.5756855,6.620957,6.8133607,7.333983,7.7301087,7.9262853,8.201687,8.98262,9.74469,10.155907,9.914458,8.733627,7.997965,7.8131065,7.854605,7.8432875,7.5263867,7.9300575,8.420499,8.707218,8.869441,9.35611,8.677037,8.243186,8.013056,7.9451485,8.009283,7.8017883,7.073672,6.571913,6.6850915,7.435844,7.4773426,8.397863,9.099571,9.265567,9.359882,9.669238,8.990166,8.262049,7.7301087,6.9567204,7.360391,7.5188417,6.7379084,5.323174,4.610148,4.247976,4.776143,5.089271,4.9685473,5.0741806,5.292993,4.6931453,4.183841,4.0895257,4.1536603,4.1008434,3.9801195,4.002755,4.2706113,4.7912335,4.534695,4.2291126,4.164978,4.406426,4.817642,4.2630663,4.195159,4.104616,3.7575345,3.187868,3.0860074,3.138824,3.0520537,2.8332415,2.8106055,2.8822856,2.757789,2.584248,2.463524,2.463524,2.3578906,2.2484846,2.1466236,2.0560806,1.9806281,1.8863125,1.9391292,2.0372176,2.173032,2.4371157,2.8407867,3.5160866,4.1272516,4.5535583,4.8553686,5.372218,5.6325293,5.666483,5.624984,5.7909794,6.149379,6.587003,6.862405,6.9567204,7.0510364,8.246958,9.061845,9.386291,9.258021,8.8769865,9.001483,9.895596,10.231359,9.537196,8.209232,0.935611,0.9620194,0.9808825,1.026154,1.0940613,1.1431054,1.177059,1.0487897,0.98465514,1.0035182,0.9280658,0.98465514,0.9808825,0.97710985,0.98842776,0.98465514,1.0035182,1.0751982,1.1581959,1.1959221,1.1129243,1.0374719,1.0374719,1.0374719,1.0223814,1.056335,1.1808317,1.1544232,1.3355093,1.6712729,1.7014539,1.7542707,1.9768555,2.2673476,2.6182017,3.1048703,4.146115,5.194905,5.9494295,6.5002327,7.375482,8.262049,9.544742,10.842525,12.079946,13.487134,15.188588,17.557796,18.931032,19.017803,18.900852,19.455427,20.168453,20.934296,22.201899,24.971004,31.599506,29.517017,22.077402,14.086982,11.793225,10.650121,9.035437,7.484888,6.1720147,4.927048,3.0218725,1.6561824,0.8337501,0.52439487,0.6451189,0.69039035,0.633801,0.46026024,0.331991,0.58098423,0.7884786,0.4979865,0.20749438,0.1056335,0.071679875,0.12826926,0.1659955,0.15467763,0.1056335,0.094315626,0.056589376,0.03772625,0.026408374,0.018863125,0.00754525,0.00754525,0.003772625,0.00754525,0.018863125,0.018863125,0.0150905,0.07922512,0.14713238,0.1659955,0.09808825,0.07922512,0.150905,0.14713238,0.060362,0.056589376,0.026408374,0.018863125,0.02263575,0.026408374,0.018863125,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.056589376,0.08299775,0.071679875,0.2565385,0.5470306,0.5093044,1.3920987,1.4071891,1.3845534,1.4562333,1.0450171,1.4600059,2.0372176,2.584248,2.8521044,2.5389767,2.6182017,2.3428001,2.082489,2.2711203,3.4179983,3.783943,4.323428,4.825187,5.0515447,4.749735,4.515832,4.561104,4.6742826,5.081726,6.477597,6.326692,6.507778,7.0170827,7.6018395,7.7640624,9.861642,11.815862,12.54775,12.393073,13.079691,12.83447,12.494934,12.7477,13.490907,13.807808,13.547497,16.029884,17.380484,16.705183,16.086473,16.561823,18.365139,19.73083,20.213724,20.69662,19.564833,17.142809,15.00373,14.056801,14.554788,14.260523,12.917468,11.676274,11.2650585,11.993175,12.672247,13.174006,13.373956,13.249459,12.872196,14.407655,15.101818,14.796235,14.211478,14.958458,14.886778,15.30554,15.63753,15.784663,16.13929,15.912932,15.143317,14.003984,12.645839,11.197151,11.551778,12.057309,12.434572,12.958967,14.471789,16.501461,18.331184,18.94235,18.516043,18.444365,18.063328,17.523844,17.784155,18.723537,19.123436,19.006485,19.327158,19.40261,19.202662,19.353567,20.598532,16.890041,14.120935,13.781399,12.974057,16.697638,18.670721,19.881733,20.53817,20.07791,19.621422,20.519308,22.330168,24.412657,25.92925,26.136745,26.366877,26.178246,25.616123,25.186045,23.888262,22.77911,22.020813,21.53037,20.972023,20.206179,20.032639,20.477808,21.402102,22.522572,23.099783,22.99415,22.499935,22.156626,22.767792,23.386503,23.55627,22.873425,21.187061,18.62545,17.139036,16.690092,16.546734,16.078928,14.747191,14.132254,13.332457,12.30253,11.438599,11.593277,11.604594,11.751727,12.566614,13.72481,14.079436,15.497944,14.7736,13.392818,12.377983,12.298758,14.456699,13.185325,10.419991,8.329956,9.314611,9.533423,6.8133607,4.425289,4.236658,6.700182,8.0206,5.1156793,1.9994912,1.026154,2.9011486,1.9881734,2.2409391,2.8822856,3.651901,4.8025517,5.511805,7.115171,8.130007,7.6886096,5.5495315,5.541986,6.5040054,7.541477,8.367682,9.2844305,10.220041,8.688355,8.627994,10.427535,10.910432,9.654147,8.975075,7.956466,6.2814207,4.2592936,2.6898816,1.6825907,1.5807298,1.8599042,1.1053791,1.2261031,1.1280149,1.539231,2.463524,3.1727777,6.360646,5.956975,4.8402777,4.696918,6.013564,8.854351,9.352338,8.231868,6.7643166,6.7567716,6.2625575,4.6818275,3.6896272,3.6669915,3.6858547,5.3948536,5.3910813,4.5233774,3.3350005,2.0673985,5.775889,6.8473144,5.089271,2.463524,3.0558262,2.8030603,3.6254926,4.640329,5.142088,4.606375,4.5988297,4.5837393,5.2326307,6.300284,6.651138,4.851596,3.6971724,3.85185,4.8327327,5.028909,6.1229706,6.5832305,6.205968,5.2552667,4.4818783,5.379763,6.7454534,7.2094865,6.092789,3.3953626,2.5691576,1.8523588,1.81086,2.173032,1.8184053,3.904667,3.2218218,1.6184561,0.38858038,0.2867195,0.38103512,0.4376245,0.5055317,0.5093044,0.271629,0.14335975,0.1056335,0.13958712,0.20749438,0.26408374,0.31312788,0.36971724,0.35462674,0.29049212,0.30181,0.35462674,0.36594462,0.4376245,0.7205714,1.418507,2.3654358,2.3126192,2.1541688,2.1390784,1.871222,1.901403,1.9127209,1.8900851,1.720317,1.2110126,1.1129243,1.2902378,1.5807298,1.8033148,1.7580433,1.5203679,1.7882242,2.1956677,2.4861598,2.5238862,3.1539145,3.591539,4.2064767,4.8025517,4.6554193,4.2706113,4.1762958,4.1008434,4.1800685,4.949684,5.010046,5.240176,5.492942,5.798525,6.379509,6.620957,6.1305156,5.5570765,5.2628117,5.3156285,5.406172,5.172269,4.9345937,4.9459114,5.3873086,6.043745,6.828451,7.5527954,8.062099,8.213005,8.137552,8.0206,8.314865,9.0957985,10.050273,10.736891,10.785934,10.54826,10.457717,11.038701,11.7026825,11.883769,13.068373,15.049001,15.901614,16.233604,15.98084,15.890297,16.071383,15.961976,15.16218,15.399856,15.17727,14.890551,16.840998,19.519562,21.247423,20.904116,18.75372,16.448645,14.139798,14.079436,15.007503,15.882751,15.886524,16.74291,16.965494,17.184307,17.520071,17.56157,13.641812,12.540206,13.407909,16.724047,24.265524,26.974268,25.235088,20.75321,14.656648,7.496206,9.344792,9.733373,9.782416,10.736891,13.985121,13.577678,12.483616,11.604594,11.144334,10.582213,9.714509,9.26934,8.809079,8.356364,8.397863,10.419991,11.212241,12.438345,13.853079,13.298503,7.2472124,5.7872066,6.9567204,11.378237,22.235851,19.595015,11.959221,7.4471617,7.254758,5.6287565,5.564622,6.2663302,6.2814207,5.753253,6.3945994,6.4247804,6.7680893,7.9036493,9.329701,9.57115,10.280403,9.737145,9.216523,8.926031,8.00551,7.3868,7.3113475,7.4094353,7.3188925,6.677546,6.043745,6.175787,6.3455553,6.477597,7.145352,6.858632,6.5530496,6.1003346,5.5193505,4.979865,4.9157305,5.070408,5.5080323,5.8966126,5.492942,5.824933,6.247467,6.3945994,6.300284,6.40969,6.688864,7.2283497,7.647111,7.9300575,8.416726,8.76758,9.559832,10.001229,9.695646,8.6732645,7.7225633,7.33021,7.3981175,7.745199,8.111144,8.812852,8.975075,8.959985,8.98262,9.107117,8.59404,8.031919,7.7602897,7.865923,8.186596,7.594294,6.8435416,6.477597,6.647365,7.0963078,7.2698483,8.050782,8.616675,8.790216,9.031664,9.510788,9.0807085,8.533678,8.190369,7.8961043,7.2698483,6.5455046,5.2326307,3.8480775,3.9197574,4.255521,4.689373,5.0062733,5.1043615,5.0213637,5.062863,4.727099,4.3800178,4.104616,3.6971724,3.5802212,3.6254926,4.0404816,4.7120085,5.1571784,4.644101,3.9612563,3.7009451,3.9008942,4.074435,3.4783602,3.4444065,3.338773,2.957738,2.5314314,2.4559789,2.5427492,2.5917933,2.5616124,2.584248,2.6483827,2.5314314,2.3956168,2.305074,2.2183034,1.9881734,1.7769064,1.6788181,1.6863633,1.7014539,1.6071383,1.720317,1.8146327,1.8448136,1.9768555,2.252257,2.7917426,3.451952,4.08198,4.5196047,5.1534057,5.5268955,5.5683947,5.4476705,5.541986,5.6325293,5.9682927,6.3531003,6.688864,6.990674,7.7414265,8.065872,7.9828744,7.7338815,7.7716074,8.782671,9.812597,9.967276,9.0957985,7.77538,1.086516,1.177059,1.2525115,1.3015556,1.3392819,1.3996439,1.3241913,1.1921495,1.0978339,1.0336993,0.91674787,1.0638802,1.0676528,1.0186088,0.98842776,1.0525624,1.086516,1.0035182,0.9695646,1.0035182,0.9507015,1.0072908,1.0450171,1.086516,1.1431054,1.2110126,1.297783,1.2147852,1.3053282,1.5882751,1.7957695,1.871222,2.0749438,2.4295704,2.9237845,3.4670424,4.3422914,4.644101,5.353355,6.7039547,8.194141,8.646856,9.955957,10.774617,11.314102,13.343775,15.701665,17.738882,19.65915,20.98334,20.549488,21.896315,22.696112,23.75622,25.676485,28.853037,30.263998,26.012249,19.91946,14.841507,12.664702,10.038955,7.914967,6.590776,5.7872066,4.659192,2.795515,1.50905,0.8111144,0.6111652,0.7167987,0.67152727,0.59607476,0.42630664,0.271629,0.40367088,0.3055826,0.16222288,0.08299775,0.071679875,0.0452715,0.08299775,0.12826926,0.124496624,0.08677038,0.10186087,0.07922512,0.07922512,0.06413463,0.030181,0.0150905,0.011317875,0.003772625,0.018863125,0.0452715,0.0452715,0.060362,0.0754525,0.11317875,0.13958712,0.056589376,0.05281675,0.150905,0.17354076,0.08677038,0.00754525,0.003772625,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.011317875,0.030181,0.0452715,0.06413463,0.0754525,0.20749438,0.44139713,0.6149379,1.4034165,1.1732863,0.87147635,0.97710985,1.50905,1.659955,1.8485862,2.565385,3.3312278,2.6710186,2.8181508,2.4371157,2.4371157,3.199186,4.568649,3.8782585,3.953711,4.014073,3.8254418,3.6783094,3.240685,3.7009451,4.0178456,4.2328854,5.451443,5.413717,5.621211,5.715527,5.7117543,5.994701,7.533932,9.737145,11.517824,12.510024,13.057055,12.630749,11.947904,12.528888,13.758763,12.90615,12.562841,13.539951,15.165953,16.603323,16.837225,16.807045,18.504726,19.640285,20.093,21.937815,20.643805,17.41821,15.4074,15.07541,14.237886,14.079436,12.823153,11.714001,11.329193,11.570641,11.487643,12.494934,13.287186,13.377728,13.098554,14.339747,14.675511,14.02662,13.072145,13.215506,13.86817,14.347293,14.667966,14.803781,14.66042,14.483108,15.116908,15.335721,14.520834,12.67602,12.51757,12.30253,12.061082,12.196897,13.50977,15.977067,17.542706,18.28214,18.606586,19.270569,18.636768,17.440845,17.105082,17.80679,18.49718,18.26705,18.791445,19.293203,19.496925,19.61765,19.640285,15.663939,12.076173,11.449917,14.543469,17.014538,17.629477,18.48209,20.274086,22.288668,21.03993,21.481327,22.401848,23.409138,24.910643,25.484081,26.061293,26.31406,25.804754,23.982576,23.133736,22.782883,22.413166,21.726547,20.65135,20.496672,20.492899,20.847527,21.519053,22.224533,23.043194,23.1941,22.714975,22.10381,22.326395,23.29596,23.84299,23.41291,21.96045,19.942095,18.644312,17.550251,16.795727,16.0412,14.456699,14.25675,14.04171,13.290957,12.291212,12.1101265,11.717773,12.162943,13.45318,14.977322,15.509261,15.848798,14.943368,14.437836,14.460471,13.626721,16.286423,12.713746,9.318384,8.918486,10.7218,9.088254,5.4363527,4.025391,6.0022464,9.382519,10.593531,6.7680893,2.9011486,1.6825907,3.5160866,2.5314314,2.9728284,3.5387223,4.0178456,5.292993,6.3719635,8.552541,9.922004,9.178797,5.6363015,5.413717,6.2927384,7.356619,8.243186,9.156161,11.189606,8.303548,6.858632,8.069645,7.99042,8.748717,5.8890676,4.304565,4.432834,2.2711203,1.4901869,1.2261031,2.1164427,3.289729,2.3465726,1.8259505,1.5845025,2.1353056,3.1124156,3.2633207,7.062354,6.560595,6.6322746,8.201687,8.213005,10.140816,9.461743,8.465771,8.7600355,11.2650585,9.884277,5.9003854,3.9008942,4.515832,4.432834,5.6023483,4.1574326,3.6971724,4.2517486,2.2786655,6.145606,6.9227667,5.2137675,3.2557755,4.90064,4.244203,5.402399,6.0324273,5.3458095,4.0895257,3.5689032,4.0895257,4.817642,5.4891696,6.405917,4.3724723,3.983892,3.4255435,3.3651814,6.9491754,11.219787,12.121444,10.374719,7.1038527,3.8367596,4.3007927,5.040227,5.8928404,5.9117036,3.3538637,2.173032,1.961765,1.81086,1.3392819,0.724344,0.814887,1.8259505,1.6939086,0.5394854,0.663982,0.8978847,0.9242931,1.0148361,1.0789708,0.70170826,0.3055826,0.16976812,0.14335975,0.15845025,0.23013012,0.21503963,0.2263575,0.24899325,0.271629,0.27917424,0.32067314,0.30181,0.35839936,0.6149379,1.1581959,1.780679,1.931584,1.9579924,1.8976303,1.478869,1.7844516,1.750498,1.599593,1.3996439,1.0940613,1.0487897,1.3053282,1.6410918,1.9164935,2.0862615,1.6863633,1.6410918,1.9089483,2.2560298,2.263575,3.3274553,3.8707132,4.055572,4.006528,3.821669,3.7273536,3.5274043,3.5462675,3.9310753,4.647874,5.0439997,5.553304,5.764571,5.8098426,6.375736,6.0626082,5.6853456,5.666483,5.847569,5.4740787,5.4212623,5.1534057,5.05909,5.292993,5.80607,6.7039547,7.2962565,7.9791017,8.620448,8.563859,7.567886,7.635793,8.375228,9.454198,10.612394,11.9064045,11.664956,11.144334,11.046246,11.502733,12.264804,12.147853,13.124963,15.052773,15.701665,16.097792,15.928022,15.241405,14.781145,15.999702,15.16218,15.098045,15.335721,15.663939,16.120426,17.610613,20.311813,21.296469,19.772327,17.052265,15.286676,14.867915,14.815099,14.460471,13.4644985,14.905642,15.441354,16.388283,17.271078,15.818617,12.653384,13.29473,13.389046,17.067356,36.960407,41.197063,36.00216,24.405111,11.910177,6.485142,7.443389,8.643084,9.42779,9.805053,10.4049,9.952185,9.1976595,9.382519,10.306811,10.291721,9.820143,8.846806,7.5792036,6.790725,7.835742,10.080454,11.461235,11.133017,9.125979,6.3153744,6.047518,6.6850915,8.013056,12.521342,25.389767,24.959686,15.513034,9.303293,8.888305,7.141579,6.1418333,6.541732,6.5643673,6.2097406,7.250985,6.5530496,7.069899,8.326183,9.363655,8.75249,9.6201935,9.020347,8.511042,8.431817,7.937603,7.5603404,7.020855,6.930312,7.118943,6.651138,6.3719635,6.4549613,6.477597,6.458734,6.8359966,6.156924,5.87775,5.873977,5.8173876,5.1835866,5.7909794,5.6513925,5.560849,5.7192993,5.7419353,5.8513412,6.0701537,6.145606,6.156924,6.507778,6.651138,7.066127,7.1981683,7.213259,8.009283,8.084735,9.099571,9.556059,9.276885,9.4013815,8.337502,7.496206,7.2094865,7.5792036,8.443134,9.495697,9.103344,8.922258,9.25425,9.050528,7.997965,7.665974,7.756517,8.054554,8.439363,7.092535,6.349328,6.25124,6.530414,6.6134114,7.786698,8.2507305,8.273367,8.152642,8.213005,8.918486,8.899622,8.620448,8.567632,9.22784,7.224577,5.4703064,3.9499383,3.006782,3.3123648,3.8895764,4.2328854,4.6554193,4.9949555,4.606375,4.406426,4.3385186,4.2819295,4.0404816,3.3123648,2.8558772,3.3953626,4.353609,5.1534057,5.2137675,4.1083884,3.451952,3.2633207,3.410453,3.6330378,3.3915899,3.006782,2.4823873,2.0183544,2.0183544,2.1541688,2.1541688,2.1579416,2.1843498,2.1466236,2.142851,2.0636258,1.991946,1.9466745,1.8674494,1.569412,1.388326,1.3317367,1.358145,1.3656902,1.3505998,1.4562333,1.5316857,1.5618668,1.6750455,1.8863125,2.2220762,2.8294687,3.6179473,4.304565,4.7836885,5.032682,5.1647234,5.281675,5.4703064,5.6287565,5.80607,6.1305156,6.609639,7.1264887,7.224577,7.0585814,6.802043,6.651138,6.7944975,8.405409,9.488152,9.393836,8.356364,7.4697976,1.2223305,1.3317367,1.3656902,1.4222796,1.5241405,1.6335466,1.388326,1.2185578,1.1016065,1.0299267,0.9922004,0.9808825,0.86770374,0.80734175,0.8563859,0.9922004,1.0638802,0.9808825,0.9695646,1.0110635,0.83752275,0.935611,1.116697,1.1544232,1.0789708,1.1732863,1.4562333,1.4901869,1.5882751,1.8561316,2.1956677,2.1466236,2.2748928,2.5012503,2.8181508,3.2972744,4.406426,4.8025517,5.7306175,7.3377557,8.68081,8.903395,9.797507,10.182315,10.729345,13.977575,15.562078,18.587723,22.57916,25.32186,22.858335,21.93027,23.967487,27.144037,30.135729,32.15031,29.234072,22.80929,17.30503,14.128481,11.6875925,8.952439,7.0170827,6.1795597,5.794752,4.255521,2.5616124,1.3204187,0.6790725,0.5093044,0.41121614,0.48666862,0.45648763,0.41498876,0.47535074,0.7922512,0.35462674,0.16222288,0.10186087,0.08299775,0.0452715,0.033953626,0.041498873,0.0452715,0.041498873,0.0150905,0.05281675,0.09808825,0.090543,0.041498873,0.0150905,0.003772625,0.0,0.018863125,0.0452715,0.0452715,0.1659955,0.181086,0.13204187,0.071679875,0.0452715,0.071679875,0.13204187,0.14335975,0.090543,0.030181,0.018863125,0.05281675,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.00754525,0.00754525,0.0452715,0.08299775,0.10186087,0.13204187,0.26031113,0.62625575,1.6863633,1.7618159,1.8900851,2.3390274,2.595566,1.7391801,1.6184561,2.5767028,3.5123138,1.8787673,3.6481283,3.0897799,3.0671442,3.8858037,3.3123648,3.6669915,3.8556228,3.3350005,2.516341,2.7615614,1.8938577,2.474842,2.7728794,2.9464202,5.036454,4.7044635,4.432834,4.6818275,5.247721,5.247721,6.749226,8.820397,10.838752,12.5326605,13.962485,13.192869,12.909923,13.29473,13.615403,12.223305,12.404391,12.095036,12.027128,12.381755,12.770335,13.0646,15.150862,16.324148,16.177015,16.618414,19.413929,19.900597,19.398838,18.104828,15.0905,13.430545,12.970284,13.041965,12.974057,12.083718,12.049765,12.717519,13.309821,13.585222,13.853079,13.856852,13.287186,12.355347,11.544232,11.642321,12.30253,12.694883,13.483362,14.366156,14.0983,13.415455,13.8870325,14.867915,15.607349,15.226315,14.471789,14.079436,13.45318,12.679792,12.559069,14.2077055,15.626213,16.576914,17.14658,17.731337,17.644567,17.350302,17.369165,17.569115,17.165443,16.750456,17.4333,18.678267,19.678013,19.349794,18.395319,16.335466,14.11339,12.883514,14.007756,15.373446,16.38451,18.052011,20.43631,22.643295,22.058538,22.416937,22.367893,22.141537,23.544952,24.838963,25.133228,25.306768,25.114365,23.22428,22.748928,22.967741,22.828154,22.092491,21.345512,21.05502,21.236107,21.696367,22.198126,22.49239,22.590479,23.548725,23.835445,23.254461,22.948877,24.084438,24.348522,24.257978,23.593996,21.409647,20.48158,18.919714,17.527617,16.505234,15.456445,15.052773,14.781145,13.936077,12.73261,12.268577,12.121444,13.000465,14.245432,15.399856,16.203424,16.044973,14.86037,14.607604,15.199906,14.539697,17.105082,13.615403,10.419991,9.891823,10.453944,8.156415,4.9760923,2.6785638,2.9501927,7.3717093,11.216014,7.405663,3.7877154,3.0897799,2.9313297,3.0407357,3.5802212,4.2064767,5.0025005,6.4549613,8.420499,11.117926,12.472299,11.227332,6.94163,7.1981683,7.2094865,6.934085,6.8359966,7.8734684,9.948412,8.171506,7.175533,7.6584287,6.379509,6.4134626,3.4859054,1.7354075,1.7957695,0.7922512,0.9393836,2.1315331,3.7348988,4.5309224,2.7011995,2.3956168,2.674791,2.384299,1.5882751,1.6033657,3.470815,4.870459,5.9192486,6.858632,8.043237,9.092027,9.107117,8.990166,8.846806,7.9791017,5.4288073,3.92353,3.2444575,3.3123648,4.164978,5.3759904,3.3236825,2.4861598,3.4142256,2.7313805,3.561358,4.134797,4.191386,4.4743333,6.7454534,5.511805,5.406172,6.0211096,6.4926877,5.492942,5.3344917,5.247721,5.692891,6.428553,6.515323,2.938875,2.4220252,2.7087448,3.2369123,5.142088,11.61214,13.59654,13.2607765,11.197151,6.4247804,4.349837,3.610402,3.7575345,4.134797,3.8895764,2.1805773,2.11267,2.3428001,1.9202662,0.26031113,0.51684964,0.58098423,0.36594462,0.12826926,0.45648763,0.69039035,0.965792,1.2864652,1.4826416,1.2525115,0.63002837,0.33576363,0.20749438,0.1659955,0.23013012,0.21503963,0.1961765,0.23767537,0.3169005,0.3055826,0.2678564,0.24899325,0.27540162,0.38858038,0.65643674,1.1431054,1.6410918,1.9164935,1.8825399,1.6033657,1.7957695,1.5354583,1.2525115,1.2185578,1.50905,1.3770081,1.5165952,1.750498,2.052308,2.5616124,1.8184053,1.4411428,1.50905,1.7882242,1.7391801,2.9464202,3.5877664,3.5575855,3.150142,3.0520537,3.712263,3.2444575,3.1652324,3.953711,5.0515447,5.270357,5.583485,6.1003346,6.790725,7.462252,6.779407,5.836251,5.802297,6.3531003,5.7079816,5.342037,4.7535076,4.6554193,5.0968165,5.462761,7.4773426,8.080963,8.488406,9.061845,9.307066,8.246958,8.458225,9.14107,10.076681,11.627231,12.178034,11.434827,10.842525,11.219787,12.770335,13.468271,12.725064,12.762791,13.834216,14.237886,14.811326,15.950659,15.799753,14.939595,16.403374,16.218515,15.497944,14.815099,14.569878,14.984866,15.607349,18.059555,19.353567,18.323639,15.626213,15.441354,15.067864,14.57365,14.064346,13.671993,13.306048,14.019074,15.460217,16.158154,13.536179,12.411936,12.049765,10.925522,14.562332,35.507946,40.683987,35.779575,24.888006,13.626721,9.110889,6.9227667,6.6247296,7.2924843,7.8810134,7.232122,8.280911,8.186596,8.152642,8.337502,7.8734684,8.058327,7.533932,7.2962565,8.069645,10.314357,12.306303,12.279895,10.944386,9.2844305,8.575176,6.549277,9.676784,13.072145,14.66042,15.199906,15.331948,12.483616,10.020092,8.82417,7.2623034,6.3229194,6.692637,7.149124,7.3377557,7.752744,6.9454026,6.8359966,7.2585306,8.009283,8.850578,9.22784,8.544995,8.160188,8.341274,8.254503,7.6320205,6.688864,6.085244,6.126743,6.760544,6.6360474,6.304056,6.2323766,6.3229194,5.9192486,4.821415,4.8402777,5.353355,5.7419353,5.402399,6.439871,6.085244,5.553304,5.572167,6.379509,5.7909794,5.3986263,5.3194013,5.59103,6.1644692,6.2021956,6.7869525,6.6662283,6.187105,7.322665,7.7150183,8.975075,9.623966,9.597558,10.269085,9.242931,8.265821,7.745199,7.9300575,8.89585,9.703192,8.903395,8.537451,8.869441,8.394091,7.6584287,7.9526935,8.4544525,8.537451,7.7829256,6.6586833,6.4247804,6.319147,6.198423,6.515323,7.9451485,8.345046,8.145098,7.6508837,7.066127,8.639311,9.556059,9.390063,8.631766,8.66572,7.1038527,4.90064,3.338773,2.8634224,3.0822346,3.7047176,4.0970707,4.164978,3.9612563,3.6934,3.863168,4.3196554,4.727099,4.606375,3.3274553,2.6898816,3.0558262,3.482133,3.5689032,3.4330888,3.410453,3.4594972,3.1237335,2.5314314,2.4107075,3.059599,3.2557755,2.9086938,2.2748928,1.9693103,2.0183544,1.9730829,1.9127209,1.8297231,1.6335466,1.5731846,1.6675003,1.7580433,1.7316349,1.5241405,1.2562841,1.237421,1.2789198,1.2940104,1.2826926,1.2449663,1.3468271,1.5052774,1.6260014,1.6033657,1.6750455,1.8787673,2.3578906,3.0935526,3.874486,4.4743333,4.798779,4.870459,4.8629136,5.081726,5.775889,6.187105,6.541732,6.832224,6.820906,6.6360474,6.3644185,6.1606965,5.9532022,5.4174895,6.722818,7.699928,7.91874,7.5188417,7.201941,1.1242423,1.2411937,1.4298248,1.4864142,1.4335974,1.4864142,1.4071891,1.1393328,0.9507015,0.9016574,0.845068,0.754525,0.76207024,0.784706,0.7997965,0.845068,1.0374719,1.0110635,0.9808825,1.0110635,1.0336993,1.0940613,1.2713746,1.3505998,1.2902378,1.2223305,1.3694628,1.5731846,1.7127718,1.8863125,2.4031622,2.2673476,2.5012503,3.0558262,3.6896272,3.9801195,4.983638,6.319147,8.043237,9.318384,8.424272,8.83926,10.914205,12.298758,13.226823,16.490145,18.663176,23.495909,28.1551,29.52079,24.224026,28.415411,31.452375,31.361832,29.313295,29.64906,25.208681,20.394812,16.55428,13.619176,10.114408,7.164215,5.3194013,4.5460134,4.3309736,3.6707642,2.4333432,1.3958713,0.8337501,0.69793564,0.6187105,0.62625575,0.69793564,0.66020936,0.52439487,0.5017591,0.20749438,0.08677038,0.056589376,0.049044125,0.02263575,0.030181,0.026408374,0.0150905,0.00754525,0.003772625,0.041498873,0.08677038,0.0754525,0.018863125,0.0150905,0.003772625,0.00754525,0.026408374,0.041498873,0.033953626,0.07922512,0.1056335,0.08677038,0.041498873,0.0452715,0.14713238,0.3470815,0.362172,0.19240387,0.090543,0.049044125,0.0452715,0.030181,0.003772625,0.011317875,0.030181,0.030181,0.02263575,0.02263575,0.02263575,0.1358145,0.16976812,0.15467763,0.24899325,0.754525,1.1506506,1.6788181,2.2409391,2.6408374,2.5804756,2.1843498,1.5958204,1.629774,2.1805773,2.203213,2.1390784,2.3314822,2.8181508,3.0671442,1.9994912,2.6446102,1.991946,2.1051247,3.0369632,2.8332415,3.4632697,4.217795,4.1989317,3.3878171,2.6634734,1.750498,2.0673985,2.3654358,2.7879698,4.878004,4.4215164,4.4139714,4.878004,5.4703064,5.4703064,6.971811,7.7225633,9.718282,12.528888,13.302276,12.1252165,11.796998,11.834724,11.910177,11.857361,11.627231,11.529142,11.532914,11.514051,11.268831,11.1631975,12.577931,13.287186,13.27964,14.7736,14.969776,16.840998,18.470772,18.606586,16.618414,15.697892,15.267814,15.313085,15.16218,13.502225,12.996693,12.925014,13.13628,13.762536,15.222542,14.460471,13.36641,12.061082,10.646348,9.201432,9.7220545,11.065109,12.223305,13.162688,14.807553,14.739646,14.211478,14.532151,15.679029,16.32792,16.203424,16.18456,16.244923,16.026112,14.841507,15.188588,16.437326,17.45971,17.772837,17.56157,16.320375,15.358356,15.105591,15.62244,16.569368,16.769318,17.165443,18.459454,19.964731,19.606333,18.33873,18.429274,18.12369,16.086473,11.359374,11.7894535,13.664448,16.505234,19.368656,20.82489,21.304014,22.7527,23.507227,23.209188,22.8357,22.081175,22.22076,22.594252,22.556524,21.503962,21.145563,21.598278,21.805773,21.560553,21.53037,22.183035,22.50748,22.658386,22.941332,23.820354,24.69183,25.966978,26.597006,26.261242,25.378448,25.548216,25.159636,25.099274,24.793692,22.239624,21.05502,19.470518,18.044466,17.093763,16.678776,16.471281,15.701665,14.366156,12.97783,12.562841,12.989148,13.7700815,15.120681,16.565596,16.961721,16.13929,13.754991,13.113645,14.505743,15.211224,16.33924,13.781399,10.770844,9.005256,8.669493,8.016829,5.5080323,3.1124156,2.4220252,4.636556,8.744945,8.035691,6.1418333,4.247976,1.0638802,2.5276587,3.240685,4.2404304,6.0022464,8.431817,11.283921,12.955194,11.823407,8.929804,7.956466,8.428044,7.6923823,7.17176,7.1566696,6.79827,7.967784,6.6549106,5.6815734,5.458988,4.0216184,2.3616633,2.6597006,2.5880208,1.7542707,1.720317,1.1846043,1.3920987,2.252257,3.169005,3.0181,2.848332,2.4182527,2.9501927,4.0782075,3.8367596,2.7238352,2.5993385,4.4743333,7.6282477,9.6051035,9.940866,8.948667,8.273367,8.035691,6.8435416,9.009028,10.763299,9.940866,6.9793563,4.8855495,6.006019,4.6214657,3.9273026,4.7610526,5.5985756,4.006528,3.5651307,3.7537618,4.104616,4.2064767,5.0251365,5.372218,4.7912335,4.006528,4.919503,4.3007927,3.9914372,4.2517486,4.52715,3.451952,2.082489,1.7844516,2.2296214,3.4066803,5.643847,7.77538,10.163452,11.589504,11.321648,9.0957985,5.5080323,3.7462165,3.0445085,3.5877664,6.5266414,7.5037513,6.296511,4.3422914,2.6144292,1.6373192,1.3392819,0.91297525,0.41876137,0.0452715,0.090543,0.18863125,0.29803738,0.69039035,1.177059,1.1431054,0.73188925,0.59607476,0.43385187,0.21503963,0.1659955,0.26408374,0.23767537,0.20749438,0.21503963,0.23013012,0.25276586,0.24899325,0.27540162,0.362172,0.5357128,0.935611,1.7014539,2.0447628,1.8674494,1.7731338,1.9202662,1.6976813,1.2826926,1.0110635,1.3505998,1.267602,1.4411428,1.7693611,2.1315331,2.3805263,1.8976303,1.5958204,1.599593,1.9127209,2.4107075,3.1010978,3.429316,3.3350005,2.938875,2.5389767,3.4896781,3.308592,3.3727267,4.247976,5.696664,6.013564,6.5568223,6.651138,6.368191,6.5228686,6.677546,6.198423,5.9607477,6.205968,6.537959,5.292993,4.7874613,5.1269975,5.670255,5.010046,6.507778,7.0057645,7.643338,8.507269,8.624221,8.537451,9.148616,9.937095,10.604849,11.042474,11.423509,11.623458,11.608367,11.593277,12.038446,12.189351,11.846043,12.170488,13.166461,13.675766,13.43809,14.252977,14.445381,14.015302,14.622695,14.173752,12.857106,12.427027,13.324911,14.667966,14.928277,16.750456,18.384,18.94235,18.384,17.508753,15.690348,14.5132885,14.166207,13.45318,12.510024,13.298503,13.958713,14.260523,15.611122,14.720782,10.804798,13.204187,21.869907,27.389257,27.517527,22.515026,18.52736,15.467763,7.0359454,5.240176,5.7796617,7.0548086,7.9036493,7.598067,7.8395147,7.5716586,7.488661,7.6093845,7.2623034,7.9941926,7.3453007,7.1981683,8.597813,11.729091,13.27964,11.212241,9.612649,10.457717,13.615403,12.781653,15.007503,19.859098,23.235598,17.346529,13.407909,11.23865,9.805053,8.544995,7.3717093,6.628502,7.062354,7.7678347,8.299775,8.66572,7.937603,7.488661,7.5226145,7.967784,8.495952,8.152642,7.9413757,8.00551,8.190369,8.035691,7.2170315,6.2399216,5.6325293,5.5004873,5.5382137,5.7306175,5.783434,5.670255,5.4250345,5.138315,4.244203,4.1310244,5.0439997,6.405917,6.8171334,7.073672,6.700182,6.066381,5.764571,6.609639,5.7683434,4.961002,5.0025005,5.7192993,5.934339,6.2323766,6.8246784,7.062354,6.934085,7.092535,7.462252,8.703445,9.318384,9.367428,10.47658,9.899368,8.873214,8.52236,8.956212,9.224068,9.865415,9.574923,9.307066,9.031664,7.745199,7.8810134,8.793989,9.152389,8.601585,7.756517,7.2283497,6.8435416,6.6020937,6.628502,7.164215,7.4282985,7.122716,7.224577,7.8621507,8.311093,8.722309,9.092027,8.8618965,8.228095,8.118689,6.828451,5.3948536,4.2102494,3.4896781,3.289729,3.6481283,3.6971724,3.6254926,3.4594972,3.0822346,3.5274043,3.8971217,4.123479,4.0178456,3.2520027,2.6068838,2.6483827,2.8822856,3.1048703,3.361409,3.3538637,3.108643,2.7841973,2.5087957,2.3880715,2.7502437,2.7917426,2.5087957,2.0900342,1.8825399,1.8523588,1.8938577,1.8184053,1.6260014,1.4977322,1.5656394,1.7655885,1.7542707,1.5015048,1.2940104,1.0940613,1.1242423,1.2864652,1.448688,1.4637785,1.4675511,1.5920477,1.6712729,1.6561824,1.6033657,1.7919968,2.022127,2.3654358,2.7992878,3.229367,3.9914372,4.357382,4.4177437,4.38379,4.5912848,5.3873086,5.9117036,6.168242,6.3229194,6.7114997,6.907676,6.8737226,6.670001,6.4926877,6.700182,7.0849895,7.1604424,6.9152217,6.5832305,6.628502,1.0525624,1.0374719,1.1808317,1.3204187,1.3694628,1.3015556,1.3091009,1.1657411,1.0223814,0.94315624,0.8903395,0.8903395,0.8337501,0.814887,0.8526133,0.8903395,1.0374719,1.1053791,1.0601076,0.98842776,1.0940613,1.2525115,1.388326,1.4298248,1.327964,1.0714256,1.1506506,1.3543724,1.6524098,2.0447628,2.5389767,2.5502944,2.6332922,3.1614597,4.0706625,4.8629136,5.8400235,7.7150183,9.261794,9.842778,9.4127,10.091772,12.079946,13.905896,15.531898,18.357594,20.417446,25.717985,29.192572,28.913399,26.076384,33.406593,34.83642,30.897799,25.751938,27.19308,24.046711,19.65915,15.169725,11.129244,7.496206,4.9685473,3.4481792,2.7351532,2.5087957,2.335255,1.8259505,1.3958713,1.1959221,1.3128735,1.7618159,1.0223814,0.77338815,0.6488915,0.5696664,0.72811663,0.27540162,0.090543,0.03772625,0.026408374,0.0150905,0.018863125,0.018863125,0.00754525,0.0,0.00754525,0.0452715,0.090543,0.0754525,0.0150905,0.00754525,0.0,0.041498873,0.06413463,0.05281675,0.041498873,0.033953626,0.0452715,0.03772625,0.02263575,0.056589376,0.15467763,0.3470815,0.38103512,0.2263575,0.08677038,0.041498873,0.033953626,0.049044125,0.09808825,0.23390275,0.45648763,0.35085413,0.150905,0.026408374,0.0754525,0.2678564,0.38858038,1.2826926,2.7426984,3.4745877,2.637065,3.2859564,3.9159849,4.085753,4.38379,2.8445592,3.0558262,3.531177,3.4670424,2.7540162,2.5767028,2.987919,3.1539145,2.6597006,1.5241405,2.4710693,2.022127,2.1277604,2.7351532,1.7919968,2.8445592,3.772625,3.6330378,2.6785638,2.3390274,2.3163917,2.3880715,2.1164427,2.0485353,3.682082,3.7650797,4.191386,4.568649,4.927048,5.6891184,6.5530496,7.6320205,9.903141,12.449662,12.449662,11.646093,10.861387,10.736891,11.355601,12.23085,11.932813,11.393328,10.740664,10.284176,10.518079,11.016065,11.532914,11.9064045,12.215759,12.792972,12.898605,15.154634,17.689838,19.040438,18.168962,17.350302,16.697638,16.263786,15.882751,15.192361,14.086982,13.5663595,13.3626375,13.690856,15.245177,14.483108,13.604086,12.615658,11.231105,8.865668,8.737399,9.431562,11.23865,13.585222,15.022593,15.735619,15.799753,15.743164,15.90916,16.444872,16.856089,17.523844,17.976559,17.7502,16.361876,16.060064,17.421982,18.670721,18.79899,17.599297,15.422491,13.7700815,13.128735,13.721037,15.482853,16.995676,17.569115,18.334957,19.138527,18.523588,18.565088,19.417702,19.059301,17.13149,14.9358225,12.030901,13.079691,15.731846,18.4255,20.360857,21.24365,22.839472,24.340977,24.74842,22.869654,20.956932,20.55326,21.088974,21.594505,20.689075,19.398838,19.678013,20.413673,21.05502,21.60205,22.714975,23.431774,23.477045,23.16769,23.420456,24.865372,26.910133,27.970242,27.845745,27.706158,27.170444,25.78212,24.869144,24.125937,21.594505,20.621168,19.436563,18.406637,17.655886,17.056038,16.867407,16.343012,15.422491,14.351066,13.6682205,13.70972,14.226569,15.614895,16.957949,16.033657,15.07541,13.792717,14.237886,15.852571,15.482853,15.988385,13.091009,9.869187,8.043237,7.9941926,6.571913,4.927048,3.9348478,4.164978,5.847569,8.688355,8.326183,5.926794,2.9313297,1.0601076,2.6634734,3.5462675,4.708236,6.4964604,8.597813,11.212241,12.219532,11.593277,9.820143,7.914967,7.232122,6.1229706,5.802297,6.2135134,6.0626082,6.126743,5.7004366,5.247721,4.3611546,1.7844516,1.1317875,1.3543724,1.4260522,1.4147344,2.4672968,3.9197574,3.127506,2.142851,2.0258996,2.8521044,4.5761943,3.8443048,2.9011486,2.6332922,2.5540671,2.9992368,3.482133,5.2590394,7.6018395,7.798016,7.496206,7.84706,7.9489207,7.8621507,8.582722,10.457717,12.683565,12.31762,9.469289,7.281166,8.013056,5.4401255,3.9197574,4.6252384,5.5306683,4.2027044,4.29702,5.1534057,5.7796617,4.8440504,3.983892,4.4403796,6.651138,8.458225,5.1043615,4.115934,3.1576872,3.7009451,4.6856003,2.5201135,2.0749438,1.8523588,4.2064767,8.179051,9.5032425,7.5565677,7.069899,7.5263867,8.382772,9.0807085,6.40969,4.3913355,2.9539654,2.969056,6.2361493,7.567886,6.0512905,3.7084904,1.9881734,1.7919968,1.931584,1.50905,0.7582976,0.06790725,0.0,0.1056335,0.14335975,0.331991,0.62248313,0.70170826,0.60362,0.6073926,0.5055317,0.28294688,0.150905,0.20749438,0.19994913,0.19240387,0.211267,0.26031113,0.3169005,0.2867195,0.26031113,0.29426476,0.3772625,0.67152727,1.3204187,1.8485862,2.0447628,1.9429018,1.7052265,1.6712729,1.4864142,1.1846043,1.1921495,1.1355602,1.1883769,1.4826416,1.9240388,2.2258487,1.9504471,1.7089992,1.6184561,1.9278114,3.0181,3.1463692,3.0746894,3.0105548,2.8596497,2.2371666,3.1954134,3.169005,3.4594972,4.5007415,5.8400235,5.6325293,5.9607477,6.3455553,6.462507,6.156924,6.304056,6.398372,6.039973,5.4740787,5.6098933,4.9345937,4.8968673,5.402399,5.9720654,5.7306175,6.255012,6.458734,6.79827,7.462252,8.397863,8.409182,9.26934,10.042727,10.336992,10.280403,10.827434,11.050018,11.41219,11.800771,11.52537,11.627231,11.631002,11.993175,12.7477,13.498452,13.430545,13.083464,13.358865,14.324657,15.181043,13.528633,12.838243,12.725064,12.913695,13.241914,13.449409,14.796235,16.614641,18.187824,18.761265,18.270823,16.407146,14.962231,14.339747,13.562587,13.011784,13.781399,13.924759,13.479589,14.498198,11.631002,14.581196,26.265015,37.514984,27.09122,23.054512,19.263023,14.916959,9.922004,4.9119577,4.5497856,5.9532022,7.2698483,7.752744,7.7716074,7.1264887,7.1076255,7.33021,7.7640624,8.710991,8.371455,7.322665,6.971811,8.016829,10.438853,12.257258,12.823153,15.316857,19.983595,24.133482,19.595015,14.02662,13.7851715,16.678776,11.959221,10.152134,9.820143,9.178797,8.0206,7.7301087,8.126234,8.016829,8.458225,9.322156,9.318384,8.624221,8.209232,8.280911,8.552541,8.231868,7.3792543,7.6584287,7.960239,7.8810134,7.7338815,7.5905213,6.356873,5.6325293,5.5382137,4.738417,4.7308717,5.270357,5.3986263,4.9534564,4.587512,4.104616,3.9310753,4.7120085,6.145606,6.971811,6.349328,6.168242,6.126743,6.1531515,6.428553,5.8211603,5.485397,5.726845,6.247467,6.156924,6.4964604,6.620957,6.9227667,7.3113475,7.2170315,7.5188417,8.461998,8.975075,9.065618,9.831461,10.121953,9.469289,9.058073,9.0543,8.601585,9.903141,10.487898,10.378491,9.695646,8.68081,8.582722,9.065618,9.261794,8.903395,8.299775,7.4094353,6.6662283,6.40969,6.7039547,7.3415284,7.5603404,7.2472124,7.488661,8.235641,8.329956,8.326183,8.296002,8.326183,8.273367,7.7716074,6.651138,5.772116,5.1760416,4.610148,3.5538127,3.0558262,2.9237845,3.1237335,3.3764994,3.1954134,3.62172,3.9084394,3.8895764,3.5123138,2.8332415,2.384299,2.3880715,2.5616124,2.7313805,2.8558772,2.7540162,2.3692086,2.2484846,2.384299,2.233394,2.3201644,2.191895,1.8900851,1.599593,1.6410918,1.7240896,1.7580433,1.6675003,1.5015048,1.4298248,1.3996439,1.4637785,1.4222796,1.2713746,1.1883769,1.1619685,1.1959221,1.2826926,1.3807807,1.418507,1.327964,1.3845534,1.4260522,1.3958713,1.327964,1.5920477,1.9240388,2.305074,2.7351532,3.2331395,3.8178966,4.044254,4.1083884,4.214022,4.5912848,5.304311,5.975838,6.2889657,6.2399216,6.1342883,6.3908267,6.628502,6.749226,6.8397694,7.1566696,6.9869013,7.164215,7.3377557,7.462252,7.8017883,1.0450171,0.9922004,1.1053791,1.2902378,1.4034165,1.2713746,1.2940104,1.2713746,1.2261031,1.1732863,1.1091517,1.116697,1.0487897,0.995973,0.9922004,1.026154,1.1506506,1.1996948,1.1393328,1.0450171,1.0751982,1.2638294,1.4373702,1.478869,1.3543724,1.1129243,1.1242423,1.3241913,1.7542707,2.2447119,2.4295704,2.8936033,3.097325,3.5953116,4.5724216,5.8664317,7.6848373,9.386291,10.227587,10.56335,11.823407,12.404391,14.079436,15.935568,17.63325,19.436563,20.85507,26.781864,30.335678,30.188545,30.580898,37.86961,35.379677,28.487091,23.190327,26.091475,24.265524,19.21398,13.253232,8.111144,4.9459114,3.3840446,2.4069347,1.8259505,1.5543215,1.6146835,1.388326,1.2487389,1.1883769,1.3204187,1.8900851,1.1280149,0.77338815,0.573439,0.49044126,0.69793564,0.2678564,0.08677038,0.026408374,0.00754525,0.00754525,0.030181,0.026408374,0.011317875,0.0,0.00754525,0.030181,0.06413463,0.05281675,0.011317875,0.0,0.003772625,0.049044125,0.06413463,0.0452715,0.033953626,0.041498873,0.049044125,0.060362,0.0754525,0.07922512,0.331991,0.3734899,0.29049212,0.16976812,0.06413463,0.049044125,0.06413463,0.120724,0.211267,0.32067314,0.482896,0.3470815,0.14713238,0.060362,0.19994913,0.4640329,0.6375736,2.0673985,4.1083884,4.0970707,3.3161373,3.640583,3.92353,3.8292143,3.8178966,2.7615614,3.1463692,3.429316,3.0030096,2.1768045,2.4484336,3.1916409,3.2255943,2.5767028,2.4899325,2.7426984,2.4333432,2.4974778,2.6597006,1.4298248,2.3767538,2.897376,2.9766011,2.7917426,2.704972,2.8106055,3.0558262,2.9954643,2.8596497,3.5387223,4.055572,4.7421894,4.7572803,4.5007415,5.6098933,5.945657,7.6923823,9.759781,11.11038,10.7557535,11.159425,10.555805,10.574668,11.563096,12.596795,12.566614,11.668729,10.967021,10.868933,11.148107,11.102836,11.072655,11.408418,11.864905,11.608367,11.951676,14.045483,16.94286,19.28566,19.300749,18.576405,17.554024,16.592005,15.999702,16.022339,14.909414,14.2077055,13.951167,14.203933,15.041456,14.245432,14.245432,13.924759,12.887287,11.457462,10.668983,10.578441,11.932813,14.075664,14.966003,15.992157,17.139036,17.252214,16.588232,16.7995,17.301258,18.074646,18.225552,17.637022,16.94286,16.588232,17.60684,18.640541,18.859352,17.927513,15.754482,14.139798,13.313594,13.483362,14.800008,16.84477,17.554024,17.916197,18.040693,17.16167,17.795471,18.87067,18.504726,16.758,15.629986,13.615403,14.539697,16.094019,17.399347,19.017803,20.296722,21.869907,23.741129,24.680513,22.205671,20.319359,19.425245,19.772327,20.82489,21.24365,19.572378,18.938578,19.534653,20.677757,20.817345,21.843498,22.99415,23.488363,23.148827,22.409393,23.145054,25.616123,27.506208,28.09851,28.279596,27.24967,25.608578,23.816582,21.971767,19.806282,19.33093,18.51227,18.199142,18.251959,17.538933,16.912678,16.693865,16.29774,15.62244,15.060319,14.664193,14.784918,15.784663,16.659912,15.033911,14.34352,14.2077055,15.199906,16.852316,17.689838,17.795471,14.354838,10.314357,7.5527954,6.8963585,4.7572803,3.500996,3.361409,4.485651,6.937857,8.695901,8.167733,6.0626082,3.5839937,2.3918443,3.199186,4.5120597,6.198423,7.9791017,9.450426,11.102836,12.121444,12.619431,11.695138,7.4282985,6.379509,5.2628117,5.028909,5.5570765,5.66271,5.2665844,5.5570765,5.836251,4.8553686,0.814887,0.90920264,0.86770374,1.2185578,2.0447628,2.9728284,5.5759397,5.4174895,4.398881,3.519859,2.9124665,4.5120597,3.953711,2.6106565,1.5845025,1.7052265,2.5804756,3.097325,4.5724216,6.6058664,7.0887623,6.9680386,8.386545,9.0807085,8.952439,10.110635,10.612394,12.400619,12.808062,10.974566,7.865923,8.386545,4.9534564,3.6179473,5.062863,4.6252384,4.3422914,4.8327327,5.349582,5.409944,4.798779,4.5799665,4.0291634,6.4436436,9.510788,5.3382645,4.191386,2.9237845,3.410453,4.8440504,3.7462165,2.4107075,2.233394,5.0515447,9.469289,10.876478,8.458225,6.398372,5.6551647,6.379509,7.907422,6.609639,4.7572803,3.5802212,3.8820312,6.0776987,6.700182,5.1232247,3.4972234,2.6823363,2.2258487,2.282438,1.5656394,0.6752999,0.060362,0.0,0.16976812,0.14713238,0.15845025,0.24899325,0.2867195,0.38103512,0.47157812,0.47912338,0.38480774,0.2565385,0.19994913,0.23767537,0.2565385,0.2565385,0.331991,0.4678055,0.3734899,0.27540162,0.26408374,0.29426476,0.52062225,0.9242931,1.448688,1.9164935,2.0372176,1.5618668,1.5203679,1.448688,1.2261031,1.0450171,0.9922004,1.0525624,1.3128735,1.7089992,2.0372176,1.871222,1.7957695,1.7014539,1.9542197,3.3764994,3.2444575,2.8294687,2.625747,2.584248,2.071171,2.9426475,2.9992368,3.470815,4.5535583,5.4212623,5.251494,5.5457587,6.0362,6.4021444,6.2851934,5.885295,6.1908774,6.138061,5.560849,5.1760416,5.1647234,5.111907,5.2892203,5.66271,5.8966126,5.7796617,5.934339,6.205968,6.72659,7.914967,8.254503,9.220296,9.831461,9.835234,9.714509,10.469034,10.465261,10.861387,11.717773,11.989402,11.981857,12.08749,12.196897,12.506252,13.517315,14.000212,12.868423,12.702429,13.86817,14.48688,13.174006,14.32843,14.743419,13.536179,12.166716,12.736382,14.2077055,16.03743,17.674747,18.572634,19.047983,17.882242,16.26756,15.071637,14.84528,14.109617,14.762281,15.697892,17.603067,22.918697,17.882242,25.19359,39.325844,47.91611,31.803228,19.715738,15.78089,11.812089,6.511551,5.462761,5.873977,6.8774953,10.967021,16.052519,15.445127,8.631766,6.930312,7.466025,9.156161,12.672247,10.061591,8.480861,7.533932,7.273621,8.239413,10.653893,13.147598,18.749947,27.136492,34.64779,25.174726,14.007756,8.89585,9.914458,9.431562,9.903141,9.884277,9.061845,7.967784,7.986647,9.623966,9.533423,9.514561,9.850324,9.322156,8.639311,8.386545,8.544995,8.726082,8.171506,7.073672,7.356619,7.6018395,7.352846,7.1302614,7.537705,6.149379,5.462761,5.6853456,4.719554,4.4177437,5.1081343,5.4212623,4.957229,4.3007927,4.323428,4.3121104,4.7120085,5.5457587,6.398372,5.462761,5.485397,5.881522,6.1606965,5.9305663,5.7872066,5.873977,6.145606,6.417235,6.360646,6.417235,6.277648,6.6586833,7.454707,7.7376537,7.745199,8.27714,8.846806,9.224068,9.442881,9.737145,9.480607,9.288202,9.216523,8.748717,10.0465,10.676529,10.61994,10.084227,9.537196,9.25425,9.454198,9.325929,8.7600355,8.356364,7.4584794,6.6624556,6.48137,6.9680386,7.696155,7.7338815,7.7640624,8.024373,8.288457,7.858378,7.960239,7.6886096,7.6508837,7.7904706,7.3792543,6.3719635,5.7494807,5.3080835,4.696918,3.410453,2.7728794,2.6634734,2.8558772,3.1539145,3.3727267,3.451952,3.519859,3.4066803,3.059599,2.5314314,2.323937,2.3390274,2.4597516,2.565385,2.5578396,2.4069347,1.9994912,1.8976303,2.1202152,2.1466236,2.372981,2.1466236,1.7354075,1.4260522,1.5316857,1.6637276,1.6071383,1.5015048,1.4411428,1.4637785,1.3543724,1.3355093,1.2638294,1.1393328,1.0789708,1.1846043,1.2487389,1.2713746,1.2789198,1.3091009,1.1393328,1.1431054,1.1657411,1.1506506,1.1242423,1.3770081,1.7014539,2.0749438,2.5276587,3.1576872,3.7009451,3.783943,3.8782585,4.168751,4.564876,5.100589,5.5797124,5.881522,6.0211096,6.1418333,6.224831,6.5643673,6.930312,7.194396,7.322665,7.092535,7.322665,7.6395655,7.911195,8.262049,1.2411937,1.2789198,1.3958713,1.5241405,1.5769572,1.4298248,1.4071891,1.4034165,1.418507,1.4222796,1.3166461,1.2261031,1.2110126,1.177059,1.1129243,1.1091517,1.2147852,1.177059,1.1355602,1.116697,1.0374719,1.1657411,1.4222796,1.5052774,1.4071891,1.4260522,1.358145,1.6524098,2.1805773,2.6295197,2.4823873,3.3350005,3.9122121,4.534695,5.492942,7.0510364,9.87296,10.834979,11.140562,11.959221,14.434063,15.011275,16.539188,18.157644,19.48561,20.640032,22.371666,28.97376,33.508453,34.72324,37.058495,41.36306,34.39125,26.431011,23.133736,25.518036,24.12971,18.214233,11.219787,5.670255,3.1652324,2.6332922,2.173032,1.7467253,1.4411428,1.4977322,1.1355602,0.91674787,0.7469798,0.67152727,0.87902164,0.8262049,0.67152727,0.4640329,0.3055826,0.33953625,0.16976812,0.06790725,0.018863125,0.0,0.0,0.03772625,0.03772625,0.0150905,0.0,0.003772625,0.00754525,0.011317875,0.011317875,0.011317875,0.0,0.011317875,0.02263575,0.026408374,0.02263575,0.011317875,0.06413463,0.09808825,0.150905,0.19240387,0.1358145,0.51684964,0.38103512,0.16976812,0.071679875,0.0452715,0.08299775,0.120724,0.18863125,0.24899325,0.211267,0.094315626,0.026408374,0.02263575,0.1056335,0.29049212,0.55457586,0.69793564,1.901403,3.4066803,2.546522,3.127506,3.2369123,3.1614597,2.8521044,1.9466745,2.0787163,1.6976813,1.2940104,1.0751982,0.98465514,1.9429018,2.7389257,2.8256962,2.6823363,3.821669,2.7426984,2.5993385,2.7615614,2.674791,1.841041,2.203213,2.214531,2.9351022,4.063117,3.9310753,3.2218218,3.5349495,4.025391,4.274384,4.2781568,4.9044123,5.7607985,5.66271,4.949684,5.5004873,5.9305663,7.5829763,8.692128,8.797762,8.756263,10.31813,10.642575,11.068882,11.974312,12.759018,12.698656,11.676274,11.472552,12.208215,12.362892,10.948157,10.842525,11.2801485,11.672502,11.634775,11.819634,13.204187,15.78089,18.504726,19.304522,19.24416,18.19537,16.999449,16.165699,15.8676605,15.230087,14.728328,14.769827,15.184815,15.218769,14.158662,14.909414,15.222542,14.78869,15.23386,14.351066,14.071891,14.102073,14.2944765,14.649103,15.460217,17.308804,18.03692,17.512526,17.60684,17.897333,18.12369,17.572887,16.625957,16.739138,16.735365,16.984358,17.38803,17.77661,17.927513,16.720274,15.79598,15.143317,14.871688,15.214996,16.509007,17.037174,17.342756,17.414436,16.693865,16.795727,17.799244,17.663431,15.746937,12.808062,15.079182,16.648594,16.939087,16.524097,17.139036,18.663176,20.258997,21.900087,22.598024,20.424992,19.538425,18.568861,18.52736,19.859098,22.443346,21.537916,19.942095,19.768555,20.662666,19.80251,20.175999,21.375692,22.545206,22.903606,21.722775,20.847527,22.888515,25.404858,26.955406,27.087448,25.43881,24.20139,22.107582,19.383747,17.746428,17.787928,17.169216,17.57666,18.689585,18.184053,16.791954,16.731592,16.690092,16.346785,16.335466,15.739391,15.373446,15.641303,15.946886,14.698147,14.422746,14.637785,15.301767,16.735365,19.625195,19.99114,16.399601,11.419736,7.122716,5.089271,3.2670932,1.9278114,1.5430037,2.6634734,5.934339,7.877241,7.877241,7.2472124,6.2663302,4.187614,3.9273026,5.583485,7.798016,9.771099,11.287694,11.646093,12.947649,14.015302,12.951422,7.145352,6.85486,5.9305663,5.8513412,6.387054,5.5985756,5.1760416,5.4250345,6.1003346,5.6891184,1.4109617,0.88279426,1.1129243,2.0447628,3.0935526,3.138824,4.9232755,6.4021444,7.17176,6.511551,3.399135,2.6785638,2.3616633,2.0485353,1.750498,1.9127209,1.3053282,0.9997456,2.2371666,4.9949555,7.967784,8.635539,10.106862,10.676529,10.087999,9.552286,10.008774,12.064855,12.83447,10.872705,6.198423,6.458734,3.953711,3.8669407,5.8400235,3.9650288,4.538468,4.8025517,4.093298,2.9992368,3.3651814,6.0626082,4.5724216,4.244203,5.783434,5.240176,4.2328854,3.1350515,3.1463692,4.2819295,5.383536,2.625747,2.6483827,4.142342,6.19465,8.27714,8.096053,7.1566696,6.4926877,6.477597,6.8435416,6.2814207,4.8629136,4.557331,5.5759397,6.3908267,6.277648,4.8138695,4.093298,4.1498876,2.9728284,2.2711203,1.0601076,0.22258487,0.00754525,0.0,0.17731337,0.14335975,0.15845025,0.21881226,0.094315626,0.18485862,0.30181,0.41876137,0.47535074,0.392353,0.26031113,0.32067314,0.33576363,0.28294688,0.3734899,0.5998474,0.47535074,0.32067314,0.27917424,0.3055826,0.47157812,0.6828451,1.0072908,1.4600059,1.9957186,1.6486372,1.4147344,1.2487389,1.1091517,0.97333723,0.91674787,1.1016065,1.3996439,1.7127718,1.9957186,1.7995421,1.9089483,1.9127209,2.0787163,3.3840446,3.270866,2.704972,2.293756,2.173032,2.0183544,2.757789,2.8634224,3.4179983,4.406426,4.727099,5.1798143,5.80607,6.096562,6.092789,6.3719635,5.553304,5.6589375,6.1305156,6.33801,5.5985756,5.7306175,5.3609,5.0779533,5.1156793,5.330719,5.2099953,5.515578,5.975838,6.537959,7.352846,8.284684,9.390063,9.854096,9.748463,10.008774,10.691619,10.453944,10.616167,11.653639,13.20796,13.245687,13.234368,12.853333,12.540206,13.475817,14.188843,13.102326,12.415709,12.626976,12.540206,13.038192,15.509261,16.263786,14.509516,12.351574,13.098554,14.966003,16.678776,17.80679,18.742401,20.100546,19.60256,18.101055,16.81459,17.342756,15.735619,16.837225,19.87796,25.997158,38.224236,30.84121,34.6742,42.890972,45.765713,30.663897,14.162435,10.133271,9.159933,7.677292,7.9791017,7.865923,7.865923,16.475054,28.747402,26.310287,11.336739,6.964266,7.8131065,11.2650585,17.463482,12.709973,10.050273,8.29223,7.092535,6.952948,9.291975,11.302785,16.180788,25.031366,36.900043,25.702894,15.041456,9.016574,8.616675,11.714001,11.993175,11.080199,9.861642,8.888305,8.360137,10.31813,10.823661,10.442626,9.661693,8.846806,8.356364,8.197914,8.22055,8.311093,8.375228,7.224577,7.1264887,7.1378064,6.8473144,6.3945994,6.6813188,5.583485,5.20245,5.696664,5.2779026,4.6252384,5.0213637,5.3609,5.142088,4.4630156,4.8968673,5.0138187,4.957229,5.0025005,5.560849,5.0439997,5.2665844,5.7004366,5.881522,5.413717,5.5457587,5.6778007,5.8513412,6.0626082,6.273875,6.0512905,6.058836,6.5455046,7.383027,8.062099,7.888559,8.13378,8.899622,9.782416,9.846551,9.42779,9.310839,9.480607,9.771099,9.831461,10.246449,10.020092,9.857869,9.891823,9.684328,9.661693,9.948412,9.390063,8.20546,7.964011,7.6395655,7.1000805,6.9869013,7.4735703,8.265821,7.8319697,8.194141,8.484633,8.296002,7.673519,7.7942433,7.3905725,6.9793563,6.820906,6.888813,5.975838,5.383536,4.689373,3.8103511,3.0030096,3.006782,3.048281,2.9464202,2.8822856,3.399135,3.1199608,2.927557,2.8785129,2.848332,2.5314314,2.4333432,2.384299,2.4107075,2.4672968,2.4182527,2.3126192,2.0145817,1.8221779,1.9051756,2.2748928,2.8445592,2.6144292,2.161714,1.8221779,1.7052265,1.6976813,1.5769572,1.4901869,1.4901869,1.5618668,1.4713237,1.4939595,1.3920987,1.1657411,1.0374719,1.1280149,1.2185578,1.237421,1.2034674,1.2147852,1.0601076,1.0450171,1.0412445,1.0186088,1.0450171,1.2600567,1.5052774,1.7316349,2.0372176,2.674791,3.3538637,3.4481792,3.6745367,4.142342,4.353609,4.5950575,4.7610526,5.119452,5.7683434,6.598321,6.507778,6.7379084,7.032173,7.213259,7.1981683,7.33021,7.383027,7.3868,7.4169807,7.5792036,1.8749946,1.961765,1.9278114,1.9240388,1.9051756,1.6486372,1.5505489,1.478869,1.4260522,1.3392819,1.1431054,1.0940613,0.97333723,0.9620194,1.0374719,0.97710985,0.80734175,0.8639311,0.9507015,0.98842776,1.0374719,1.1959221,1.3996439,1.418507,1.3770081,1.7542707,1.6675003,2.1692593,2.916239,3.5462675,3.6934,4.032936,4.659192,5.5495315,6.8058157,8.635539,10.393582,10.650121,11.517824,13.324911,14.618922,16.618414,17.889788,19.164934,21.032385,23.925987,29.73583,35.315544,37.92243,38.56,41.993088,42.015724,33.251915,26.63096,24.872917,22.49239,21.651094,16.376965,9.820143,4.5309224,2.4559789,2.1390784,1.6750455,1.2411937,0.9016574,0.59607476,0.4376245,0.3772625,0.33576363,0.3169005,0.42630664,0.4640329,0.34330887,0.211267,0.1659955,0.29049212,0.23013012,0.1056335,0.018863125,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0150905,0.041498873,0.018863125,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.011317875,0.0,0.02263575,0.094315626,0.20372175,0.29426476,0.24522063,0.15845025,0.08299775,0.06413463,0.08299775,0.0452715,0.094315626,0.09808825,0.08677038,0.08677038,0.1358145,0.05281675,0.011317875,0.018863125,0.056589376,0.1056335,0.15467763,0.15845025,0.8903395,2.1579416,2.7917426,3.2067313,4.3347464,4.6554193,3.9122121,3.1425967,1.9957186,1.3958713,1.2034674,1.4373702,2.305074,2.0108092,1.6184561,1.9051756,2.3918443,1.3430545,1.4298248,1.9994912,2.6446102,2.8407867,1.9391292,2.0485353,2.595566,3.610402,4.772371,5.43258,4.3196554,3.127506,2.293756,2.263575,3.5085413,4.2404304,5.66271,6.730363,6.9152217,6.19465,7.6093845,7.533932,7.175533,7.2924843,8.194141,9.024119,10.174769,11.121698,11.891314,13.075918,11.404645,10.054046,9.465516,10.008774,11.947904,11.117926,11.065109,11.242422,11.634775,12.770335,13.102326,12.853333,13.426772,15.143317,17.240896,18.889534,19.04421,18.16519,16.810818,15.626213,14.977322,15.339493,15.618668,15.584714,15.852571,14.694374,14.588741,15.082954,15.686575,15.8676605,16.13929,16.248695,15.939341,15.113135,13.856852,14.452927,15.977067,17.301258,17.95015,18.097282,18.474545,18.26705,17.621931,16.810818,16.252468,16.618414,16.535416,16.497688,16.550507,16.28265,16.293968,15.8676605,15.701665,16.15438,17.240896,16.961721,16.927769,17.28994,17.912424,18.402864,18.376457,18.644312,17.335213,14.93205,14.298248,15.98084,16.697638,16.610868,16.478827,17.640795,18.323639,19.636513,20.315586,19.779873,18.142553,18.485863,18.13878,18.150099,19.353567,22.367893,22.967741,22.062311,21.439827,21.364376,20.583443,19.715738,19.930779,21.005976,22.17549,22.126446,20.575897,21.092747,22.552752,24.220253,25.75571,22.790428,21.288923,19.828917,18.085964,16.82968,17.037174,16.659912,17.274849,18.534906,18.157644,16.24115,16.41092,16.803272,16.837225,17.225805,16.29774,15.418718,15.143317,15.282904,14.894323,14.781145,15.113135,15.943113,16.365646,14.5132885,17.271078,14.04171,9.208978,5.406172,3.5387223,2.5767028,1.327964,0.5696664,0.94315624,2.9464202,6.790725,8.216777,7.91874,6.651138,5.247721,4.6742826,5.6476197,7.115171,8.993938,12.193124,11.299012,12.083718,13.170234,12.58925,7.7678347,7.888559,7.020855,8.039464,9.552286,5.8890676,4.5724216,3.4444065,3.3727267,3.85185,3.0218725,1.2638294,0.6149379,1.1016065,2.1956677,2.806833,3.0520537,4.274384,5.772116,6.2814207,3.9989824,2.191895,1.2902378,0.76584285,0.4376245,0.47157812,0.5583485,0.7167987,1.6146835,3.6481283,6.94163,7.835742,9.465516,9.718282,8.197914,6.255012,8.880759,13.245687,12.811834,7.7376537,4.8666863,3.9159849,4.859141,5.243949,4.429062,3.5839937,4.8440504,4.9647746,3.9273026,2.6446102,2.9766011,4.745962,5.534441,5.406172,4.847823,4.776143,4.2404304,3.3161373,3.097325,3.6254926,3.904667,2.3201644,2.9200118,3.8292143,4.274384,4.5761943,4.2102494,5.292993,6.458734,7.001992,6.8661776,6.205968,5.511805,5.0779533,4.927048,4.7912335,4.719554,4.002755,3.2029586,2.6785638,2.595566,1.6788181,0.76207024,0.19994913,0.03772625,0.0,0.0,0.1358145,0.34330887,0.44894236,0.1659955,0.13204187,0.23013012,0.392353,0.47535074,0.3055826,0.27917424,0.23767537,0.21503963,0.2263575,0.27540162,0.482896,0.47157812,0.35839936,0.2678564,0.3055826,0.35462674,0.48666862,0.724344,1.1280149,1.7995421,1.8749946,1.6712729,1.4411428,1.267602,1.0827434,1.0336993,1.1883769,1.5731846,2.093807,2.5314314,2.082489,2.1503963,2.2560298,2.384299,3.006782,2.8219235,2.4371157,2.1654868,2.0900342,2.0900342,2.565385,2.704972,3.2972744,4.214022,4.4101987,4.9232755,5.994701,6.4511886,6.043745,5.43258,5.3344917,5.2628117,5.6853456,6.156924,5.342037,5.2326307,5.451443,5.534441,5.4174895,5.4174895,5.73439,5.87775,6.066381,6.587003,7.7829256,8.526133,10.140816,10.834979,10.789707,12.14408,12.098808,11.427281,11.378237,12.366665,13.977575,15.184815,15.094273,14.147344,13.109872,13.060828,12.853333,12.344029,12.204442,12.551523,12.955194,14.079436,13.826671,13.792717,14.241659,14.143571,13.59654,15.033911,16.595778,17.753973,19.31584,20.63626,19.893051,19.48561,20.017548,20.30804,18.429274,21.915178,27.317577,33.644268,42.374123,30.520536,25.242634,28.751175,30.018778,4.7610526,7.3113475,8.729855,9.107117,8.782671,8.329956,6.7944975,7.828197,17.399347,29.079393,24.061802,10.7218,6.9567204,8.420499,12.691111,19.270569,14.743419,9.465516,7.164215,7.964011,8.394091,8.416726,9.484379,9.450426,10.631257,19.821371,15.354584,10.042727,7.7301087,9.224068,12.313848,10.774617,11.031156,11.442371,11.057564,9.64283,9.81637,10.325675,9.944639,8.846806,8.590267,8.873214,8.575176,8.111144,7.997965,8.865668,7.643338,7.484888,7.413208,6.94163,6.089017,5.4778514,5.5193505,5.6400743,5.6287565,5.6287565,4.2404304,4.112161,4.4403796,4.8553686,5.4174895,5.8702044,5.4401255,4.9157305,4.7044635,4.851596,5.1458607,5.7306175,6.145606,6.085244,5.402399,4.98741,5.0854983,5.3571277,5.6287565,5.8588867,6.066381,6.3945994,6.752999,7.01331,6.9869013,7.575431,7.960239,8.82417,10.11818,11.031156,10.740664,10.344538,10.227587,10.393582,10.469034,10.186088,9.246704,8.873214,9.25425,9.537196,9.81637,9.805053,9.024119,8.001738,8.269594,8.197914,7.7301087,7.5112963,7.8017883,8.484633,8.228095,8.537451,9.061845,9.295748,8.575176,7.673519,7.1340337,6.730363,6.436098,6.4247804,5.617439,5.070408,4.402653,3.6141748,3.0520537,3.308592,3.4745877,3.429316,3.3123648,3.5085413,3.519859,3.350091,3.3010468,3.2633207,2.7011995,2.4182527,2.2484846,2.1390784,2.003264,1.7089992,1.6712729,1.690136,1.8448136,2.1768045,2.7011995,3.0181,2.8407867,2.7200627,2.6710186,2.1805773,1.8523588,1.9089483,1.9240388,1.7693611,1.5882751,1.5731846,1.6071383,1.5467763,1.4034165,1.3430545,1.20724,1.1846043,1.1355602,1.0676528,1.1280149,1.0940613,1.0110635,0.935611,0.8865669,0.83752275,1.1808317,1.4864142,1.4864142,1.3807807,1.8297231,2.4408884,2.8521044,3.4481792,4.0970707,4.1197066,3.874486,4.398881,5.3759904,6.2436943,6.19465,6.2814207,6.330465,6.175787,5.9909286,6.270103,6.881268,7.1981683,7.2472124,7.201941,7.3868,1.7052265,1.7995421,1.7844516,1.8146327,1.8599042,1.720317,1.5241405,1.3958713,1.3317367,1.3053282,1.267602,1.0902886,0.9507015,0.86770374,0.8337501,0.84129536,0.8865669,0.9393836,1.0299267,1.1506506,1.2562841,1.297783,1.6146835,1.8033148,1.7731338,1.7429527,2.1051247,2.7426984,3.519859,4.3611546,5.2288585,5.1232247,5.455216,6.360646,7.756517,9.344792,9.616421,10.86516,12.377983,13.800262,15.143317,18.161417,18.848034,19.466745,21.564325,25.989614,31.456148,35.636215,36.798183,36.198338,38.07333,35.86257,27.577888,21.156881,18.478317,15.373446,13.166461,10.084227,6.4549613,3.1727777,1.7240896,1.1921495,0.814887,0.68661773,0.6790725,0.41121614,0.28294688,0.24522063,0.20749438,0.211267,0.4376245,0.4376245,0.34330887,0.2263575,0.15467763,0.21503963,0.23390275,0.18863125,0.1056335,0.033953626,0.02263575,0.003772625,0.00754525,0.0150905,0.011317875,0.0150905,0.030181,0.0150905,0.0,0.0,0.0,0.011317875,0.0150905,0.011317875,0.003772625,0.0,0.13204187,0.13204187,0.124496624,0.16222288,0.23013012,0.12826926,0.06790725,0.05281675,0.06413463,0.056589376,0.21503963,0.2867195,0.25276586,0.150905,0.10186087,0.05281675,0.06790725,0.12826926,0.19240387,0.19240387,0.19240387,0.18485862,0.56589377,1.0827434,0.83752275,2.0749438,3.0369632,2.8634224,2.142851,2.886058,1.4939595,1.2034674,1.5505489,1.9466745,1.6825907,1.0186088,0.88279426,1.026154,1.1393328,0.84129536,2.003264,2.305074,2.3616633,2.2447119,1.4864142,2.173032,3.531177,3.9008942,3.5123138,4.504514,4.6516466,3.9499383,3.6141748,3.9084394,4.168751,6.013564,7.1566696,7.3453007,7.073672,7.575431,7.496206,7.6622014,7.99042,8.707218,10.355856,10.853842,11.970539,13.370183,14.332202,13.758763,12.498707,13.011784,12.894833,12.400619,14.449154,15.426264,14.641558,13.04951,11.808316,12.272349,13.411682,13.287186,13.2607765,14.071891,15.852571,16.882498,18.7839,20.032639,19.97605,18.810308,18.153872,17.003222,16.29774,16.365646,16.91645,15.901614,16.199652,16.429781,16.218515,16.188334,17.14658,17.889788,17.784155,16.803272,15.528125,15.618668,16.301512,17.120173,17.844517,18.485863,17.644567,17.836971,17.554024,16.686321,16.493916,16.791954,17.410664,17.82188,17.836971,17.599297,16.859861,15.871433,15.543215,15.829934,15.716756,15.70921,15.882751,16.459963,17.380484,18.316093,17.520071,18.43682,18.557543,17.20317,15.554533,16.06761,16.444872,16.486372,16.414692,16.87118,17.799244,18.323639,18.644312,18.670721,18.02183,19.466745,19.757236,19.821371,20.353312,21.794455,22.745155,22.171717,21.02484,20.206179,20.545715,20.617395,19.851553,20.11941,21.568098,22.613113,21.805773,21.21347,21.711456,23.073374,23.98635,21.722775,19.908142,18.531134,17.327667,15.769572,16.524097,17.071129,17.761518,18.293459,17.72002,16.535416,16.222288,16.21097,16.41092,17.191853,16.078928,15.516807,15.16218,14.84528,14.551015,15.4074,16.350557,16.648594,15.282904,10.948157,12.14408,10.4049,7.281166,4.6931453,4.957229,2.6068838,1.1996948,0.66775465,0.98842776,2.1881225,3.6707642,5.7607985,7.4282985,7.986647,7.092535,4.485651,3.7650797,4.357382,5.9192486,8.345046,9.869187,10.616167,10.695392,10.27663,9.635284,8.194141,7.039718,6.8359966,6.8473144,4.9119577,5.028909,4.293247,3.5877664,3.2935016,3.2670932,1.8674494,1.0525624,0.84884065,1.1996948,1.9655377,3.4972234,4.0103,4.1612053,3.9725742,2.8521044,1.659955,1.0299267,0.7130261,0.56212115,0.52062225,0.6187105,1.9278114,3.078462,4.7610526,9.725827,8.273367,9.986138,12.472299,14.196388,14.483108,14.841507,13.234368,10.495442,8.084735,8.07719,4.0291634,4.0517993,5.3948536,6.156924,5.292993,3.4972234,3.1614597,3.5236318,4.236658,5.3571277,5.7306175,4.112161,3.4217708,4.5422406,6.326692,4.274384,3.289729,2.6898816,2.6936543,4.432834,5.4401255,4.927048,4.22534,4.085753,4.6629643,4.715781,5.9305663,7.17176,7.6584287,6.9869013,6.4549613,6.436098,6.3832817,5.9682927,5.070408,5.1835866,4.3121104,2.8558772,1.6146835,1.7655885,2.3428001,1.20724,0.21503963,0.00754525,0.0,0.0,0.026408374,0.124496624,0.21503963,0.13204187,0.19240387,0.2678564,0.41498876,0.5281675,0.32821837,0.29426476,0.23013012,0.21881226,0.271629,0.29803738,0.573439,0.62248313,0.5319401,0.422534,0.4376245,0.31312788,0.3772625,0.7394345,1.2411937,1.4826416,1.841041,1.7467253,1.5769572,1.4675511,1.3015556,1.3619176,1.4977322,1.8674494,2.5729303,3.6669915,2.886058,2.746471,2.9237845,3.1161883,3.0558262,2.71629,2.2711203,2.1654868,2.3088465,2.0673985,2.335255,2.5616124,2.9992368,3.6481283,4.2630663,4.432834,5.5457587,6.115425,5.7381625,5.089271,4.9534564,4.7950063,5.028909,5.4740787,5.3269467,5.1798143,5.3156285,5.6061206,5.9230213,6.149379,6.2135134,6.1305156,6.247467,6.779407,7.8319697,8.009283,8.941121,9.937095,10.736891,11.487643,11.2801485,11.370691,11.634775,11.978085,12.3289385,13.615403,13.622949,13.200415,12.940104,13.196642,13.309821,12.925014,12.238396,11.774363,12.393073,14.962231,14.596286,14.324657,14.792462,14.268067,12.664702,14.569878,16.214743,17.086218,19.927006,21.013521,20.956932,21.190834,21.432283,19.723284,18.0671,20.692848,25.959433,31.482555,34.14603,26.219744,18.976303,14.50197,12.740154,11.487643,11.283921,10.231359,9.405154,8.937348,8.024373,8.062099,7.854605,9.865415,12.615658,10.672756,8.843033,8.439363,10.450171,12.947649,11.068882,8.707218,7.1264887,8.643084,11.668729,10.699164,10.178542,11.8045435,12.792972,12.30253,11.434827,6.428553,5.028909,6.722818,9.295748,8.809079,11.774363,15.007503,14.581196,11.140562,9.899368,9.593785,10.035183,9.88805,9.0807085,8.7751255,8.809079,8.337502,7.707473,7.352846,7.7904706,6.862405,6.952948,7.281166,7.284939,6.6247296,6.326692,6.255012,6.255012,6.0739264,5.349582,4.447925,4.2064767,4.568649,5.353355,6.247467,5.8588867,5.704209,5.2099953,4.6026025,4.927048,4.9760923,5.5268955,6.149379,6.439871,6.0626082,4.8742313,4.961002,5.1798143,5.119452,5.1269975,5.6287565,6.2323766,6.730363,6.8133607,6.096562,7.201941,7.9338303,8.639311,9.337247,9.725827,10.33322,10.197406,9.835234,9.7296,10.355856,9.95973,9.092027,8.401636,8.273367,8.816625,10.250222,10.680302,9.922004,8.6581745,8.428044,8.854351,8.473316,8.035691,8.009283,8.59404,8.375228,8.616675,9.175024,9.65792,9.416472,8.201687,7.2283497,6.5756855,6.3531003,6.692637,5.6513925,4.61392,4.044254,3.92353,3.7235808,3.7273536,3.9725742,3.8367596,3.410453,3.4972234,3.4217708,3.682082,3.8103511,3.5274043,2.7615614,2.6672459,2.5502944,2.4408884,2.3503454,2.282438,2.0598533,2.0258996,2.123988,2.2484846,2.2258487,2.71629,2.5201135,2.3390274,2.4333432,2.6106565,2.4069347,2.3993895,2.1466236,1.6675003,1.4147344,1.3958713,1.4034165,1.448688,1.4750963,1.3543724,1.2789198,1.3807807,1.3543724,1.1808317,1.1053791,1.1959221,1.1581959,1.1204696,1.0638802,0.83752275,1.0525624,1.3430545,1.4637785,1.539231,2.0372176,2.3088465,2.6068838,3.0407357,3.5802212,4.08198,4.425289,4.957229,5.80607,6.6020937,6.477597,6.4926877,6.5040054,6.48137,6.6020937,7.2358947,7.33021,7.4282985,7.605612,7.884786,8.2507305,1.7542707,1.8523588,1.9278114,2.003264,2.033445,1.8863125,1.6524098,1.5128226,1.418507,1.327964,1.1959221,1.026154,1.0223814,1.0186088,0.95824677,0.90920264,1.0374719,1.0827434,1.1280149,1.2261031,1.4222796,1.4411428,1.7316349,1.9655377,2.0560806,2.142851,2.8143783,3.4972234,4.172523,4.878004,5.670255,5.832478,6.428553,7.1906233,8.0206,9.027891,9.382519,10.7218,12.042219,13.321139,15.539442,17.323895,17.64834,19.406384,23.209188,27.411894,32.188038,37.27731,39.5522,38.808994,37.771523,30.475266,22.21699,16.550507,13.622949,10.163452,7.5075235,5.764571,4.1083884,2.4220252,1.267602,0.7092535,0.43007925,0.40367088,0.4640329,0.30181,0.56212115,0.44516975,0.2678564,0.2565385,0.543258,0.331991,0.2867195,0.2263575,0.150905,0.23390275,0.30181,0.26031113,0.18863125,0.124496624,0.06790725,0.02263575,0.011317875,0.011317875,0.011317875,0.02263575,0.0150905,0.003772625,0.0,0.0,0.00754525,0.124496624,0.08299775,0.02263575,0.00754525,0.00754525,0.181086,0.24899325,0.2263575,0.21503963,0.392353,0.59230214,0.46026024,0.29803738,0.20749438,0.09808825,0.18485862,0.2263575,0.56212115,1.1355602,1.4750963,0.38103512,0.124496624,0.1358145,0.14335975,0.15845025,0.18485862,0.35085413,1.1016065,1.9164935,1.3128735,1.8599042,2.516341,2.9313297,3.1312788,3.5387223,1.9164935,1.3920987,1.5845025,1.8938577,1.5241405,0.724344,1.0487897,1.0450171,0.6526641,1.2034674,2.3314822,2.1805773,1.720317,1.569412,2.0145817,2.493705,3.0897799,3.1652324,2.938875,3.4934506,3.0558262,3.4179983,4.08198,4.617693,4.636556,5.1571784,5.6815734,6.881268,8.552541,9.65792,9.220296,8.631766,9.216523,10.906659,12.23085,13.758763,13.766309,13.555041,13.389046,12.494934,12.038446,12.804289,13.238141,13.257004,14.27184,14.754736,14.498198,13.981348,13.615403,13.739901,14.781145,15.347038,15.690348,16.003475,16.418465,16.705183,17.297485,18.372684,19.662922,20.4514,20.070366,18.99894,18.214233,18.025602,18.070873,17.7502,17.946377,17.874697,17.312576,16.569368,17.48989,18.68204,18.889534,17.953922,16.788181,16.260014,16.94286,18.225552,19.074392,18.03692,18.346275,19.349794,19.379974,18.45568,18.323639,17.738882,18.251959,19.247932,19.76101,18.451908,17.297485,16.199652,15.663939,15.505488,14.841507,15.362129,15.105591,14.977322,15.513034,16.886269,16.505234,17.369165,18.13878,17.984104,16.592005,16.071383,16.497688,16.501461,16.090246,16.648594,17.852062,19.108345,19.685556,19.47429,18.961214,19.274342,20.375948,22.028357,23.09601,21.560553,21.58696,21.371922,20.304268,19.047983,19.523335,20.334448,20.462717,20.877707,21.779364,22.60557,22.17549,20.715485,20.477808,21.817091,23.186554,21.349285,19.753464,18.244415,16.833452,15.69412,16.350557,16.716501,17.052265,17.297485,17.078674,16.803272,16.286423,15.79598,15.626213,16.109108,16.018566,15.984612,15.565851,14.928277,14.849052,14.958458,14.856597,15.513034,15.543215,11.18206,11.634775,8.99771,6.1116524,4.881777,6.2625575,3.6292653,1.6750455,1.1016065,1.6373192,2.0447628,3.097325,5.4703064,7.8206515,9.058073,8.341274,5.036454,3.7084904,3.7084904,4.644101,6.349328,8.695901,9.774872,9.6201935,9.050528,9.680555,8.07719,7.2358947,6.4738245,5.458988,4.221567,4.6742826,4.636556,3.983892,3.2067313,3.4255435,2.5087957,1.9089483,1.5128226,1.4750963,2.2220762,4.515832,4.1989317,3.1840954,2.372981,1.6373192,1.0714256,0.76207024,1.0789708,1.5128226,0.69039035,0.9922004,3.9159849,6.092789,7.7338815,12.664702,9.880505,12.645839,16.395828,18.651857,19.002712,17.746428,12.947649,9.914458,9.789962,9.529651,3.8443048,2.9200118,4.191386,5.4967146,5.089271,3.048281,2.987919,3.8103511,4.9044123,6.1418333,6.356873,4.7308717,3.9197574,4.82896,6.6134114,3.9273026,3.270866,3.4972234,3.8820312,4.112161,4.961002,5.379763,5.3458095,5.119452,5.2628117,5.66271,6.3455553,6.94163,7.149124,6.72659,6.006019,5.9305663,5.915476,5.5495315,4.610148,4.5799665,3.8103511,2.8256962,2.1503963,2.3428001,2.674791,1.3053282,0.2263575,0.0452715,0.00754525,0.0,0.0,0.0452715,0.11317875,0.11317875,0.16976812,0.22258487,0.3169005,0.41121614,0.362172,0.20372175,0.17354076,0.19994913,0.23390275,0.26031113,0.44139713,0.62248313,0.6451189,0.513077,0.3734899,0.29049212,0.32821837,0.6187105,1.1204696,1.6033657,1.9429018,1.8825399,1.7731338,1.6788181,1.358145,1.6712729,2.033445,2.41448,3.0407357,4.4101987,3.3727267,3.1199608,3.2105038,3.2972744,3.138824,2.746471,2.3163917,2.2711203,2.4786146,2.214531,2.5389767,2.8558772,3.1048703,3.4632697,4.346064,4.255521,4.5196047,5.0175915,5.2364035,4.2630663,4.315883,4.085753,4.0480266,4.3083377,4.6026025,4.847823,5.3382645,5.96452,6.5002327,6.587003,6.530414,6.515323,6.6020937,6.9227667,7.677292,7.9036493,8.465771,9.133525,9.854096,10.736891,10.940613,11.41219,12.1252165,12.759018,12.687338,13.12119,12.759018,12.2270775,12.132762,13.102326,13.830443,13.543724,12.815607,12.2119875,12.291212,13.645585,14.901869,15.309312,14.879233,14.362384,12.51757,13.472044,14.962231,16.59955,19.908142,21.153109,20.892797,20.63626,20.69662,20.172226,19.927006,20.655123,21.87368,23.948624,28.106056,27.355305,24.197617,23.111101,26.66114,35.496628,32.584164,20.209951,11.472552,9.612649,8.031919,8.224322,7.3981175,7.092535,7.854605,9.239159,15.4074,17.923742,17.674747,14.400109,6.7114997,6.722818,6.3417826,8.737399,11.978085,9.042982,7.2396674,8.903395,11.680047,13.407909,12.121444,8.00551,7.8508325,8.858124,9.0957985,7.496206,14.230342,16.912678,14.766054,10.095545,8.296002,8.91094,8.692128,8.360137,8.22055,8.197914,7.61693,7.492433,7.333983,7.149124,7.4584794,7.01331,6.900131,6.9227667,6.937857,6.8774953,7.194396,6.952948,6.4738245,5.8928404,5.149633,4.8025517,4.7836885,5.1043615,5.692891,6.398372,6.349328,5.832478,5.100589,4.5233774,4.568649,4.689373,5.2175403,6.0626082,6.7341356,6.3644185,5.349582,5.1081343,5.010046,4.9987283,5.594803,5.8513412,6.058836,6.628502,7.2170315,6.7077274,7.250985,7.8508325,8.13378,8.047009,7.8696957,8.6581745,9.050528,9.107117,9.250477,10.284176,9.673011,8.692128,8.224322,8.262049,7.9036493,9.763554,10.352083,9.880505,8.963757,8.597813,8.869441,8.7600355,8.60913,8.582722,8.66572,9.178797,9.525878,9.665465,9.6201935,9.491924,8.284684,7.1566696,6.5002327,6.3153744,6.2021956,5.3080835,4.315883,3.7688525,3.7235808,3.7462165,3.4330888,3.5085413,3.380272,3.0822346,3.2821836,3.3161373,3.6858547,3.7801702,3.3727267,2.6219745,2.674791,2.5314314,2.293756,2.0787163,2.0145817,1.8033148,1.8976303,1.8900851,1.7542707,1.8221779,2.293756,2.1881225,2.1013522,2.2899833,2.6521554,2.6332922,2.384299,2.0296721,1.6675003,1.3543724,1.2223305,1.2110126,1.2600567,1.297783,1.2562841,1.2826926,1.2600567,1.1431054,1.0299267,1.1619685,1.2562841,1.2713746,1.2261031,1.1053791,0.9016574,0.9922004,1.2185578,1.4713237,1.7165444,2.0183544,2.3013012,2.505023,2.8106055,3.2331395,3.6066296,4.036709,4.617693,5.353355,6.006019,6.089017,6.439871,6.692637,6.881268,7.1038527,7.5301595,7.4811153,7.4018903,7.3113475,7.303802,7.533932,1.7316349,1.8561316,2.022127,2.1277604,2.1277604,2.0145817,1.7844516,1.6524098,1.5354583,1.3996439,1.2713746,1.0676528,1.1280149,1.1732863,1.1053791,1.0186088,1.2185578,1.1581959,1.1242423,1.2261031,1.3958713,1.4939595,1.6335466,1.8372684,2.0975795,2.3692086,3.3727267,4.08198,4.689373,5.2590394,5.7306175,6.458734,7.284939,7.665974,7.779153,8.503497,9.005256,10.163452,11.461235,13.113645,16.044973,17.56157,18.48209,21.424738,26.34424,30.528082,35.432495,40.540627,41.79314,38.477,33.233055,24.159891,17.372938,13.12119,10.412445,7.0057645,4.6742826,3.7009451,3.2067313,2.505023,1.1317875,0.5357128,0.32067314,0.29049212,0.30181,0.26031113,0.7582976,0.73566186,0.58098423,0.51684964,0.6149379,0.35462674,0.23767537,0.17354076,0.150905,0.23390275,0.30181,0.26408374,0.211267,0.16222288,0.06790725,0.030181,0.03772625,0.033953626,0.02263575,0.03772625,0.011317875,0.00754525,0.003772625,0.003772625,0.02263575,0.15467763,0.090543,0.018863125,0.00754525,0.00754525,0.124496624,0.26031113,0.27917424,0.23390275,0.35839936,0.633801,0.52439487,0.33576363,0.211267,0.10940613,0.13958712,0.97710985,1.5958204,1.6561824,1.5279131,0.482896,0.3055826,0.30935526,0.2867195,0.49421388,0.35839936,1.2562841,2.4899325,3.338773,3.0558262,2.3126192,2.7879698,3.2444575,3.451952,4.1762958,2.5238862,1.8523588,1.5731846,1.4034165,1.3807807,0.88279426,1.267602,1.3015556,0.98842776,1.569412,2.2409391,2.1654868,1.8485862,1.7278622,2.173032,2.5201135,2.6672459,2.71629,2.7917426,3.059599,2.463524,3.0181,3.9122121,4.5422406,4.508287,4.4743333,4.938366,6.752999,9.265567,10.325675,9.846551,9.288202,9.8239155,11.159425,11.555551,13.498452,13.113645,11.872451,10.876478,10.868933,11.299012,12.178034,12.777881,13.155144,14.147344,14.143571,14.377474,14.762281,15.022593,14.671739,15.184815,16.275105,17.120173,17.20317,16.346785,16.686321,16.550507,16.840998,17.803017,19.051756,19.293203,19.462973,19.47429,19.31584,19.059301,18.964987,18.829172,18.666948,18.28214,17.282394,17.384256,17.904879,18.146326,17.87847,17.342756,16.939087,17.57666,19.28566,20.621168,18.68204,19.938324,20.847527,20.806026,20.30804,20.930523,19.568605,19.164934,19.613878,20.025093,18.700903,17.467255,16.505234,15.875206,15.384765,14.584969,15.618668,15.222542,14.34352,13.86817,14.607604,15.0376835,15.660167,16.429781,16.897587,16.18456,15.535669,16.380737,16.569368,15.905387,16.13929,17.21826,19.01403,20.334448,20.700394,20.353312,19.63274,20.756983,22.696112,23.850534,22.066084,21.104065,20.715485,19.779873,18.58395,18.832945,20.232588,21.394556,22.21699,22.63575,22.594252,22.024584,20.11941,19.436563,20.617395,22.382984,20.99843,19.866644,18.289686,16.55428,15.931795,15.690348,15.928022,16.290195,16.501461,16.33924,16.595778,16.33924,15.848798,15.365902,15.116908,15.675257,16.188334,15.852571,15.226315,16.233604,14.358611,13.70972,14.592513,15.214996,11.6875925,11.038701,7.756517,4.9987283,4.3800178,5.945657,4.5912848,2.4182527,1.6335466,2.2220762,1.9579924,3.4179983,5.572167,8.013056,9.714509,9.035437,5.726845,4.7346444,4.7044635,5.1835866,6.6360474,7.907422,8.552541,8.182823,7.3679366,7.647111,7.1076255,6.688864,5.9532022,4.8742313,3.8405323,4.266839,4.727099,4.640329,4.2404304,4.568649,4.074435,3.7650797,3.6179473,3.270866,2.033445,4.8553686,4.666737,3.591539,2.7426984,2.1805773,1.6825907,1.2600567,1.4298248,1.7919968,1.0374719,1.2298758,3.9876647,6.5756855,8.643084,12.238396,10.502988,12.095036,14.188843,15.384765,15.728074,15.562078,11.3820095,8.582722,8.345046,7.6207023,3.31991,2.5993385,3.31991,4.0291634,3.942393,3.2633207,3.6179473,4.3913355,5.1835866,5.824933,5.798525,4.798779,4.0970707,4.221567,4.991183,5.0439997,5.0666356,4.9987283,4.647874,3.682082,3.6896272,5.6589375,6.1606965,5.0138187,5.2967653,5.9532022,6.205968,6.058836,5.7607985,5.8211603,5.194905,5.20245,5.5985756,5.904158,5.3986263,4.6629643,3.663219,2.9049213,2.5616124,2.4597516,2.7728794,1.2600567,0.14713238,0.060362,0.00754525,0.0,0.018863125,0.07922512,0.15845025,0.1659955,0.16976812,0.20372175,0.2565385,0.30935526,0.34330887,0.150905,0.13204187,0.16222288,0.18863125,0.23013012,0.3055826,0.52439487,0.6111652,0.4979865,0.3169005,0.2867195,0.331991,0.5583485,1.0035182,1.6410918,2.1088974,2.082489,2.0145817,2.033445,1.9391292,2.293756,2.7615614,3.127506,3.591539,4.7648253,3.6594462,3.5462675,3.6330378,3.440634,2.8294687,2.6295197,2.3314822,2.263575,2.3880715,2.3088465,2.7992878,3.1350515,3.1350515,3.1425967,4.0103,4.285702,4.1989317,4.3913355,4.6629643,3.9574835,4.014073,3.7613072,3.7877154,4.1310244,4.3083377,4.67051,5.413717,6.145606,6.6020937,6.6360474,6.477597,6.752999,7.0812173,7.356619,7.77538,7.911195,8.216777,8.597813,9.1976595,10.423763,10.948157,11.385782,12.095036,12.97783,13.460726,13.630494,13.155144,12.370438,11.955449,12.943876,14.053028,13.698401,13.29473,13.358865,13.50977,14.003984,15.856343,16.286423,15.271586,15.546988,12.925014,12.5326605,13.328684,15.0905,18.440592,20.62494,20.613623,19.840235,19.470518,20.387266,23.020557,22.726294,21.179516,20.598532,23.748674,24.552244,27.785383,32.15031,37.91111,46.901276,39.25039,23.160145,11.868678,9.359882,10.355856,8.661947,8.903395,9.884277,10.891568,11.680047,17.395575,21.73032,20.69662,14.011529,5.0741806,5.8702044,7.3981175,9.325929,10.457717,8.748717,4.5988297,5.1760416,9.49947,14.196388,13.505998,10.212496,10.295494,9.963503,8.050782,5.987156,14.928277,19.153618,17.21826,11.257513,6.990674,8.5563135,7.91874,7.4207535,7.673519,7.564113,6.277648,6.5341864,6.7944975,6.771862,7.4169807,7.175533,7.1566696,7.122716,7.1264887,7.4999785,8.412953,7.7037,6.688864,5.8626595,4.8968673,5.1232247,5.4703064,5.6589375,5.8211603,6.5266414,6.33801,5.4438977,4.6516466,4.255521,4.0480266,4.745962,5.1043615,5.824933,6.6322746,6.300284,5.6023483,5.2175403,4.9232755,4.82896,5.379763,5.80607,5.9682927,6.4021444,7.0585814,7.2924843,7.5792036,7.5565677,7.2094865,6.696409,6.33801,7.2924843,7.960239,8.243186,8.52236,9.699419,9.646602,9.073163,8.635539,8.243186,7.066127,8.714764,9.4127,9.5032425,9.190115,8.578949,8.718536,8.937348,9.107117,9.167479,9.159933,10.18986,10.514306,10.20495,9.684328,9.740918,8.643084,7.3075747,6.541732,6.304056,5.7192993,4.7044635,3.92353,3.5538127,3.5349495,3.5802212,3.2369123,3.2859564,3.2369123,3.097325,3.380272,3.4783602,3.399135,3.218049,2.916239,2.3578906,2.6974268,2.4107075,2.0145817,1.7542707,1.6109109,1.4147344,1.4826416,1.4713237,1.3920987,1.6071383,1.8636768,1.901403,1.9164935,2.04099,2.3767538,2.4597516,2.1277604,1.8033148,1.6146835,1.3845534,1.1619685,1.1544232,1.1808317,1.1619685,1.1280149,1.2110126,1.0978339,1.0223814,1.0751982,1.2185578,1.2336484,1.2336484,1.1657411,1.0299267,0.8865669,0.97710985,1.1732863,1.4335974,1.720317,2.0183544,2.5427492,2.7426984,2.8747404,3.097325,3.4557245,3.6858547,4.1197066,4.6742826,5.240176,5.66271,6.326692,6.888813,7.24344,7.4471617,7.756517,7.745199,7.635793,7.375482,7.0812173,7.0284004,1.569412,1.7240896,1.9127209,2.022127,2.0145817,1.961765,1.81086,1.7052265,1.5920477,1.4939595,1.4713237,1.2336484,1.2185578,1.2185578,1.177059,1.1732863,1.3732355,1.177059,1.086516,1.2110126,1.2789198,1.4826416,1.4524606,1.5958204,2.003264,2.4069347,3.6443558,4.323428,4.878004,5.3948536,5.6287565,6.851087,7.756517,7.9036493,7.726336,8.552541,8.892077,9.97482,11.680047,14.030393,17.214487,19.859098,22.009495,25.416174,30.256453,35.119366,40.823574,43.73227,40.763214,32.704887,24.205162,17.814335,13.792717,11.083972,8.714764,5.798525,4.074435,3.4142256,3.289729,2.9086938,1.2147852,0.5998474,0.42630664,0.33953625,0.2263575,0.23767537,0.62248313,0.784706,0.7922512,0.69793564,0.5357128,0.44516975,0.21881226,0.1056335,0.15845025,0.211267,0.23013012,0.20749438,0.181086,0.150905,0.056589376,0.041498873,0.0754525,0.08299775,0.05281675,0.049044125,0.02263575,0.0150905,0.00754525,0.00754525,0.030181,0.0754525,0.033953626,0.0,0.003772625,0.0,0.0150905,0.17354076,0.25276586,0.20749438,0.16222288,0.1961765,0.19994913,0.14335975,0.06790725,0.08677038,0.120724,1.8146327,2.3918443,1.3128735,0.31312788,0.7130261,0.8601585,0.98842776,1.1808317,1.358145,1.0072908,2.4408884,3.7047176,4.134797,4.3611546,2.8709676,3.2520027,3.1954134,2.8219235,4.6818275,3.270866,2.4031622,1.5920477,0.90920264,0.98842776,1.026154,1.1808317,1.3996439,1.5920477,1.6373192,1.7919968,2.2484846,2.5276587,2.4069347,1.8938577,2.1994405,2.6068838,2.7728794,2.8143783,3.3048196,3.31991,3.108643,3.399135,4.006528,3.8593953,4.61392,5.4212623,6.7643166,8.379,9.288202,8.907167,9.220296,9.476834,9.442881,9.405154,10.593531,10.699164,9.752235,8.797762,9.910686,10.8576145,12.121444,12.815607,13.287186,15.116908,15.045229,15.256495,15.46399,15.335721,14.490653,14.618922,15.746937,16.648594,16.569368,15.237633,15.973294,16.403374,16.31283,15.894069,15.75071,16.463736,17.870924,18.931032,19.319613,19.40261,19.025349,18.606586,18.387774,18.248188,17.72002,16.746683,16.060064,16.090246,16.72782,17.301258,17.7502,18.221779,19.870417,21.681276,20.455173,21.462463,21.488873,21.183289,21.349285,22.918697,21.749184,20.398582,19.462973,18.968758,18.372684,17.4333,16.822134,16.124199,15.264041,14.524607,15.754482,15.762027,14.720782,13.29473,12.672247,13.528633,14.0983,14.641558,15.086727,15.026365,14.958458,16.161926,16.678776,16.086473,15.516807,15.886524,17.482344,19.625195,21.383238,21.579414,20.77962,21.27006,21.96045,22.398075,22.786655,21.55678,20.673985,19.768555,18.99894,19.059301,20.843754,22.401848,23.348776,23.537407,23.054512,21.677504,19.68933,18.829172,19.534653,20.934296,20.22127,19.60256,18.233097,16.486372,15.958203,14.754736,15.165953,15.916705,16.214743,15.720529,15.943113,16.150608,16.086473,15.626213,14.781145,15.335721,16.143063,16.029884,15.784663,18.161417,14.388792,13.93985,14.222796,13.426772,10.521852,8.571404,5.847569,3.8141239,3.270866,4.38379,4.776143,2.8822856,1.8599042,2.1956677,1.6939086,3.4179983,5.028909,7.3113475,9.488152,9.216523,6.9265394,6.368191,6.4964604,6.934085,7.937603,7.2924843,6.8737226,6.198423,5.3269467,4.8629136,5.7079816,5.5985756,5.2250857,4.7233267,3.6971724,4.0782075,4.738417,5.372218,5.8211603,6.066381,6.1116524,5.9720654,5.9418845,5.1232247,1.4260522,3.9197574,4.4630156,4.266839,3.983892,3.6971724,2.9124665,2.1541688,1.6524098,1.4864142,1.5845025,1.50905,2.335255,4.3611546,7.141579,9.514561,9.922004,9.329701,8.59404,8.167733,8.107371,9.778644,8.635539,6.4134626,4.6252384,4.564876,2.795515,2.9652832,3.259548,3.0218725,2.7615614,3.5349495,4.353609,4.9647746,5.149633,4.7346444,4.327201,4.2102494,3.9989824,3.5538127,2.9652832,7.073672,7.8432875,6.5455046,4.644101,3.7914882,3.2821836,5.783434,6.1305156,4.2819295,5.349582,5.836251,5.926794,5.349582,4.5422406,4.67051,4.4177437,4.715781,5.624984,6.609639,6.5530496,5.6551647,4.6252384,3.6141748,2.7125173,1.9730829,2.6106565,1.1204696,0.026408374,0.030181,0.0,0.00754525,0.041498873,0.12826926,0.23013012,0.24522063,0.21881226,0.23390275,0.26408374,0.28294688,0.271629,0.16976812,0.120724,0.124496624,0.17354076,0.24899325,0.271629,0.41876137,0.49421388,0.44139713,0.34330887,0.29426476,0.35462674,0.6111652,1.056335,1.5769572,2.2484846,2.2447119,2.2107582,2.4371157,2.837014,3.1199608,3.451952,3.7386713,4.063117,4.6554193,3.7348988,4.002755,4.1989317,3.6669915,2.3503454,2.354118,2.2447119,2.142851,2.1503963,2.3465726,2.9615107,3.2218218,2.9992368,2.7238352,3.361409,4.2781568,4.606375,4.5007415,4.2404304,4.255521,4.0404816,3.7877154,4.093298,4.745962,4.719554,4.859141,5.492942,5.926794,6.047518,6.33801,6.2927384,6.730363,7.281166,7.748972,8.058327,7.798016,7.9526935,8.3525915,9.0543,10.325675,11.09529,11.34051,11.536687,12.136535,13.58145,14.2944765,14.305794,13.50977,12.525115,12.672247,14.109617,13.932304,13.962485,14.709465,15.354584,16.003475,17.176762,17.180534,16.539188,18.002966,14.4152,13.200415,13.091009,13.93985,16.697638,19.742147,20.489126,20.06282,19.670467,20.590988,25.008732,24.703148,22.990377,21.519053,20.289177,17.908651,25.804754,31.946589,33.595226,37.292397,25.868889,16.403374,10.86516,10.378491,15.203679,10.933067,12.815607,15.056546,15.0376835,13.290957,12.449662,16.580687,17.006994,11.657412,5.05909,5.8400235,9.5183325,10.740664,9.382519,10.589758,4.327201,4.115934,8.499724,13.264549,11.446144,8.865668,9.016574,8.529905,6.4549613,4.255521,13.192869,21.353058,21.319103,13.543724,6.360646,8.175279,7.643338,7.2660756,7.605612,7.2585306,5.666483,6.0776987,6.375736,6.2814207,7.322665,7.0510364,7.326438,7.575431,7.752744,8.326183,9.344792,8.130007,6.8925858,6.1795597,4.847823,5.4401255,6.039973,6.092789,5.9305663,6.779407,5.6589375,4.6742826,4.134797,3.9801195,3.7914882,5.1760416,5.2175403,5.50426,6.1908774,5.9909286,5.300538,5.0062733,4.798779,4.5837393,4.4818783,5.3156285,5.9607477,6.1342883,6.2021956,7.164215,7.752744,7.0887623,6.1720147,5.6023483,5.617439,6.696409,7.360391,7.54525,7.707473,8.83926,9.65792,9.7069645,9.009028,7.8206515,6.6134114,7.816879,8.424272,8.903395,9.148616,8.473316,8.688355,9.152389,9.473062,9.627739,9.989911,11.046246,11.136789,10.465261,9.74469,10.227587,9.246704,7.673519,6.571913,6.0739264,5.3910813,4.164978,3.5538127,3.4368613,3.5387223,3.4368613,3.2255943,3.410453,3.4557245,3.3274553,3.500996,3.6368105,2.9916916,2.546522,2.4786146,2.1654868,2.5993385,2.1164427,1.6335466,1.4562333,1.2864652,1.0751982,0.965792,1.0186088,1.1959221,1.3656902,1.388326,1.5241405,1.5580941,1.5354583,1.750498,1.841041,1.6750455,1.50905,1.448688,1.448688,1.2261031,1.2147852,1.2336484,1.1808317,1.0148361,1.0638802,0.9922004,1.0714256,1.2638294,1.2223305,1.1732863,1.1506506,1.086516,0.9808825,0.8865669,1.146878,1.3355093,1.4600059,1.6373192,2.1051247,2.8181508,3.0822346,3.0671442,3.0860074,3.5953116,3.6292653,3.8367596,4.2064767,4.7308717,5.3910813,6.1644692,6.900131,7.2698483,7.375482,7.7716074,7.8734684,7.888559,7.7414265,7.4697976,7.1981683,1.4335974,1.5203679,1.6410918,1.7391801,1.7429527,1.5731846,1.6448646,1.6071383,1.5731846,1.5430037,1.4335974,1.3732355,1.2487389,1.1808317,1.2600567,1.539231,1.4071891,1.3166461,1.2826926,1.3015556,1.388326,1.5845025,1.5430037,1.6637276,2.1164427,2.8219235,3.7763977,4.214022,4.5422406,4.8855495,5.081726,6.398372,7.643338,8.492179,9.061845,9.918231,10.552032,11.819634,13.815352,16.542961,19.911915,22.733839,25.35204,28.720995,33.165146,38.390232,44.117077,43.177692,35.35704,24.41643,18.0671,14.916959,12.774108,10.582213,8.152642,6.1644692,4.52715,3.6330378,3.0369632,2.3503454,1.2525115,0.90920264,0.84129536,0.6149379,0.23767537,0.150905,0.17731337,0.14713238,0.1358145,0.15467763,0.1659955,0.30181,0.19994913,0.13204187,0.18485862,0.26031113,0.211267,0.16222288,0.16222288,0.18863125,0.150905,0.090543,0.11317875,0.120724,0.08677038,0.060362,0.02263575,0.00754525,0.0,0.00754525,0.030181,0.00754525,0.0,0.00754525,0.011317875,0.0,0.02263575,0.18485862,0.32067314,0.34330887,0.26031113,0.08677038,0.10186087,0.1056335,0.06413463,0.0754525,0.08677038,0.21881226,0.482896,0.72811663,0.6413463,2.3503454,2.173032,2.5804756,3.5538127,2.5804756,2.4823873,2.372981,2.6898816,3.187868,2.9464202,2.674791,2.7087448,3.1539145,4.1197066,5.7079816,4.8138695,2.806833,1.50905,1.1355602,0.3055826,0.48666862,0.935611,1.1996948,1.2864652,1.6637276,1.2600567,1.8561316,2.1843498,2.0673985,2.3956168,1.9202662,2.1768045,2.4672968,2.7804246,3.7688525,3.5990841,2.9237845,2.9237845,3.4934506,3.2520027,4.032936,4.447925,5.100589,6.307829,8.103599,8.394091,8.75249,8.544995,8.405409,10.223814,10.344538,10.303039,9.812597,9.333474,10.054046,10.593531,11.879996,13.6682205,15.456445,16.493916,15.309312,15.354584,15.494171,15.196134,14.524607,15.124454,15.886524,16.090246,15.603577,14.909414,14.543469,14.607604,14.879233,14.969776,14.298248,14.298248,15.056546,16.218515,17.437073,18.402864,18.168962,17.772837,16.969267,16.15438,16.388283,15.192361,14.864142,14.93205,15.482853,17.165443,18.33873,19.217752,20.462717,21.688822,21.470009,21.62846,21.58696,21.503962,21.636003,22.307531,23.103556,22.337713,21.02484,19.542198,17.640795,17.4333,17.56157,16.4826,14.509516,13.837989,14.622695,15.154634,14.916959,13.966258,12.940104,13.072145,14.049255,14.837734,15.211224,15.746937,15.79598,16.459963,16.886269,16.697638,15.992157,15.113135,16.365646,18.75372,21.088974,22.01704,21.481327,21.915178,22.164171,22.03213,22.26226,21.87368,21.122927,20.37972,19.938324,20.036411,21.839725,23.371412,23.733583,23.446865,24.457928,21.420965,19.43279,18.55377,18.48209,18.55377,18.787672,18.632996,17.889788,16.667458,15.396083,14.811326,15.022593,15.660167,16.124199,15.546988,15.339493,15.501716,15.641303,15.539442,15.135772,16.052519,16.546734,16.637276,17.025856,19.089483,15.70921,14.505743,13.015556,10.374719,7.322665,5.383536,3.682082,2.9954643,3.31991,3.8443048,3.8103511,2.2975287,1.2185578,1.1431054,1.327964,2.3277097,3.531177,5.406172,7.594294,8.91094,9.95973,8.382772,7.8961043,8.6581745,7.277394,6.2889657,5.613666,5.093044,4.640329,4.22534,5.13077,5.300538,5.1835866,4.768598,3.5839937,3.8782585,4.768598,5.692891,6.1418333,5.613666,6.8133607,6.617184,5.492942,3.8405323,1.9994912,1.780679,1.871222,2.2296214,2.6597006,2.806833,2.3428001,1.9429018,1.9504471,2.2560298,2.305074,2.6597006,2.04099,3.1727777,6.488915,10.163452,9.846551,11.6875925,12.427027,10.7218,7.1566696,5.4476705,5.8890676,5.692891,4.908185,6.40969,2.9766011,2.6597006,3.2784111,3.410453,2.3956168,2.897376,4.606375,5.311856,4.4403796,3.0369632,3.3538637,5.3269467,6.5228686,5.9796104,4.2102494,7.0812173,8.118689,7.3377557,5.6853456,5.0515447,4.244203,4.4177437,5.194905,6.3153744,7.643338,6.900131,6.63982,6.187105,5.3269467,4.304565,4.1197066,4.2027044,4.4403796,4.5988297,4.3196554,6.2361493,7.0812173,6.187105,4.08198,2.4710693,2.0070364,0.77338815,0.018863125,0.0,0.0,0.03772625,0.018863125,0.018863125,0.071679875,0.18485862,0.24522063,0.2678564,0.2678564,0.24899325,0.19994913,0.17354076,0.13204187,0.124496624,0.18863125,0.33576363,0.3470815,0.44139713,0.52062225,0.51684964,0.38103512,0.28294688,0.31312788,0.69793564,1.358145,1.9089483,2.2748928,2.173032,2.2107582,2.5578396,2.9615107,3.5839937,3.6934,3.821669,4.032936,3.9386206,3.4859054,4.168751,4.4139714,3.7047176,2.595566,2.1654868,2.1315331,2.1390784,2.1768045,2.5804756,3.0671442,3.2067313,3.006782,2.8030603,3.2670932,3.8405323,4.5233774,4.644101,4.2894745,4.304565,3.7650797,3.4859054,3.6481283,4.2781568,5.2175403,5.3910813,5.5683947,5.311856,5.0062733,5.873977,6.6813188,6.470052,6.458734,7.069899,7.9489207,7.424526,7.696155,8.280911,8.899622,9.461743,11.0613365,11.54046,11.200924,10.982111,12.483616,13.456953,14.554788,14.27184,12.804289,12.0233555,14.637785,15.848798,16.056292,15.754482,15.546988,15.682802,17.172989,18.30855,19.040438,20.979568,18.28214,17.580433,17.312576,17.112627,17.82188,19.557287,20.326904,21.817091,23.4695,22.50748,22.17549,21.251196,19.421474,17.346529,16.663685,17.029629,23.537407,25.608578,21.790682,19.7761,13.585222,10.072908,12.415709,18.51227,20.964478,16.803272,17.572887,15.414946,10.838752,12.740154,8.873214,9.616421,10.978339,10.163452,5.583485,8.941121,10.880251,11.778135,11.774363,10.770844,5.583485,8.307321,9.767326,7.5527954,6.0286546,5.4778514,5.5495315,5.6778007,5.455216,4.6252384,10.861387,20.349539,20.598532,11.438599,5.0062733,6.273875,6.115425,6.221059,6.952948,7.352846,6.537959,6.8435416,6.832224,6.432326,6.9567204,6.9567204,6.802043,6.881268,7.3981175,8.360137,8.386545,7.3679366,6.6850915,6.485142,5.692891,6.009792,6.40969,6.5228686,6.458734,6.790725,4.9949555,4.146115,4.032936,4.293247,4.3800178,5.5759397,5.3080835,5.3080835,5.832478,5.66271,4.5988297,4.214022,4.323428,4.640329,4.776143,4.983638,5.9418845,6.058836,5.5495315,6.4549613,7.0510364,6.6813188,5.696664,4.957229,5.8136153,6.228604,7.0548086,7.435844,7.5716586,8.744945,8.975075,8.503497,7.77538,7.149124,6.881268,8.16396,7.888559,7.7301087,8.201687,8.66572,8.873214,9.329701,9.725827,10.038955,10.514306,11.45369,11.231105,10.084227,9.0807085,10.11818,9.310839,7.854605,6.330465,5.1835866,4.7308717,4.217795,3.712263,3.5424948,3.5839937,3.2670932,2.8030603,2.8785129,2.927557,2.7540162,2.546522,2.987919,2.776652,2.595566,2.5804756,2.3503454,1.8749946,1.2864652,0.8978847,0.77338815,0.76207024,0.63002837,0.5319401,0.5017591,0.52062225,0.5357128,0.65643674,0.7054809,0.68661773,0.6413463,0.6413463,0.7884786,0.87902164,1.0072908,1.20724,1.448688,1.3015556,1.237421,1.2713746,1.2562841,0.91674787,0.86770374,0.8903395,0.94692886,1.026154,1.1581959,1.20724,1.358145,1.3656902,1.237421,1.2525115,1.7769064,1.9089483,1.841041,1.8259505,2.1654868,2.6068838,2.8521044,2.9501927,3.0105548,3.2029586,3.4255435,3.772625,4.1612053,4.5724216,5.036454,5.7796617,6.3417826,6.4926877,6.4134626,6.6850915,6.964266,7.152897,7.3075747,7.3717093,7.1868505,1.3241913,1.3694628,1.3958713,1.5580941,1.8184053,1.9504471,1.8674494,1.8485862,1.7919968,1.7052265,1.7014539,1.5430037,1.5467763,1.5543215,1.50905,1.4675511,1.4713237,1.4901869,1.4977322,1.5052774,1.5731846,1.9730829,2.0749438,2.2748928,2.6446102,2.9313297,3.6292653,4.06689,4.425289,4.9119577,5.7419353,7.1264887,8.088508,9.0807085,10.269085,11.555551,12.755245,14.418973,15.814844,17.814335,22.892288,25.868889,28.517273,32.131447,36.91136,41.977997,44.93951,41.800686,33.14251,22.767792,17.689838,14.694374,11.879996,9.416472,7.360391,5.66271,3.9801195,2.8898308,2.1353056,1.5656394,1.1280149,1.3430545,1.0638802,0.62248313,0.28294688,0.2263575,0.3470815,0.44516975,0.362172,0.181086,0.19240387,0.3734899,0.26031113,0.16222288,0.16976812,0.17354076,0.116951376,0.1659955,0.24899325,0.30935526,0.31312788,0.241448,0.21503963,0.17354076,0.10186087,0.03772625,0.018863125,0.0150905,0.00754525,0.00754525,0.030181,0.0150905,0.026408374,0.06413463,0.08677038,0.02263575,0.03772625,0.124496624,0.16976812,0.17731337,0.24899325,0.28294688,0.24899325,0.21503963,0.29803738,0.663982,0.43007925,0.86770374,1.3920987,1.8938577,2.71629,3.8971217,3.663219,3.1916409,2.8747404,2.2975287,2.1805773,2.191895,2.6031113,3.0633714,2.6031113,3.097325,3.6934,4.4630156,4.821415,3.5462675,3.983892,2.5125682,1.4939595,1.5128226,1.3656902,1.2562841,1.539231,1.569412,1.3920987,1.7127718,1.6109109,2.252257,2.5276587,2.3088465,2.4333432,2.3163917,2.1013522,2.1164427,2.2975287,2.1805773,2.6446102,2.7011995,3.1312788,3.6594462,2.957738,4.538468,5.0062733,5.7909794,7.066127,7.7376537,7.2283497,7.2623034,7.0887623,7.0774446,8.722309,9.186342,10.310584,10.714255,10.529396,11.434827,13.155144,13.792717,14.769827,16.06761,16.22606,15.912932,15.79598,15.663939,15.505488,15.528125,14.943368,14.468017,14.037937,13.7700815,13.943622,12.845788,12.528888,12.423254,12.272349,12.147853,12.951422,13.434318,14.226569,15.448899,16.705183,16.063837,15.607349,15.154634,14.64533,14.154889,13.924759,14.520834,14.890551,14.890551,15.286676,16.91645,17.814335,18.251959,18.599041,19.357338,18.75372,20.013775,21.375692,22.235851,23.163918,23.654358,23.028103,21.688822,19.806282,17.297485,16.437326,16.350557,15.83748,14.815099,14.32843,13.977575,14.037937,14.053028,13.834216,13.45318,12.736382,13.060828,14.109617,15.064092,14.622695,14.739646,15.75071,16.286423,15.973294,15.430037,14.581196,15.241405,16.927769,18.97253,20.515535,21.462463,22.33394,22.677248,22.481071,22.17549,21.843498,21.51528,20.922977,20.4099,20.938068,22.186808,23.4695,24.789919,25.744392,25.544443,22.703657,20.545715,19.18757,18.429274,17.761518,17.874697,18.26705,18.184053,17.41821,16.275105,15.777118,16.222288,16.712729,16.697638,15.977067,15.573396,15.456445,15.607349,15.924251,16.233604,16.478827,17.082445,17.557796,17.976559,18.964987,16.863634,15.218769,12.464753,9.171251,8.031919,6.247467,4.032936,2.5012503,2.1503963,2.867195,2.6483827,1.7693611,1.1506506,1.0751982,1.2185578,2.11267,2.9200118,4.014073,5.458988,7.032173,10.023865,10.03141,8.59404,7.043491,6.485142,7.3113475,6.760544,6.273875,5.9418845,4.4705606,5.0138187,6.096562,5.8966126,4.398881,3.3915899,3.7499893,4.7006907,6.2625575,7.1906233,4.9685473,4.2894745,4.8402777,4.4705606,2.8822856,1.6448646,1.4750963,1.9164935,2.776652,3.591539,3.6028569,2.444661,2.04099,2.2560298,2.6031113,2.2447119,3.3878171,3.187868,3.150142,5.1534057,11.442371,13.588995,13.732355,12.6345215,10.850069,8.729855,7.3453007,5.66271,5.032682,5.3873086,5.2364035,2.3918443,1.780679,1.7844516,1.81086,2.323937,4.395108,6.198423,6.126743,4.5007415,3.5236318,3.4594972,5.5759397,7.0774446,6.7152724,4.7610526,6.730363,6.8058157,5.666483,4.2630663,3.8065786,4.4177437,5.27413,5.9984736,6.488915,6.900131,7.2283497,9.5032425,11.02361,10.729345,9.186342,6.94163,5.983383,5.915476,5.624984,3.2444575,4.447925,4.8742313,4.4894238,4.014073,4.9119577,2.0749438,0.6375736,0.090543,0.0,0.0,0.018863125,0.03772625,0.03772625,0.0452715,0.14713238,0.18863125,0.2678564,0.29049212,0.24522063,0.18485862,0.16222288,0.120724,0.1358145,0.20749438,0.23767537,0.32821837,0.42630664,0.452715,0.39989826,0.331991,0.30181,0.32067314,0.62248313,1.2298758,1.9429018,1.9579924,2.11267,2.5578396,2.9803739,2.6295197,3.1539145,3.3010468,3.3953626,3.4670424,3.2520027,3.289729,3.610402,3.5689032,3.1161883,2.8256962,2.1353056,2.233394,2.3277097,2.3126192,2.7728794,3.006782,2.9464202,3.0218725,3.338773,3.6556737,4.5120597,4.8138695,4.821415,4.821415,5.0968165,4.4818783,4.327201,3.99521,3.8782585,5.413717,5.4665337,5.462761,5.2665844,5.0515447,5.311856,6.217286,6.3531003,6.4474163,6.8699503,7.6207023,7.145352,7.6320205,8.529905,9.0957985,8.397863,10.533169,11.604594,11.732863,11.555551,12.2270775,12.098808,13.498452,13.95494,13.011784,12.23085,14.766054,15.746937,15.878979,15.173498,12.936331,14.351066,16.01102,16.976812,17.440845,18.746174,17.904879,18.346275,18.104828,17.757746,20.458946,20.911661,20.82489,22.04722,23.609087,21.677504,21.952906,22.14531,21.632233,20.043957,17.25976,21.65864,24.17498,21.417192,15.720529,15.16218,18.45568,17.916197,18.063328,18.451908,13.679539,15.237633,16.641048,14.226569,9.718282,10.227587,7.8621507,9.099571,11.895086,13.234368,9.125979,10.001229,12.0082655,12.50248,10.536942,6.8435416,5.1798143,5.670255,5.379763,4.06689,4.172523,4.568649,4.7610526,4.779916,4.659192,4.4516973,6.560595,10.480352,10.355856,6.530414,5.553304,6.677546,6.8246784,6.85486,7.1264887,7.488661,7.443389,7.2924843,6.809588,6.4511886,7.3490734,7.9451485,7.6810646,7.364164,7.4396167,7.9941926,8.567632,7.333983,6.296511,6.089017,5.9607477,6.326692,6.3644185,5.904158,5.2967653,5.409944,4.817642,4.538468,4.5007415,4.6290107,4.8440504,5.9230213,5.704209,5.541986,5.7570257,5.6363015,4.7421894,4.45547,4.5837393,4.821415,4.738417,5.111907,5.704209,5.824933,5.6023483,5.9796104,6.0701537,5.9003854,5.6589375,5.6853456,6.4738245,7.3377557,7.462252,7.3717093,7.3377557,7.375482,6.8661776,6.8737226,6.673774,6.2436943,6.247467,7.001992,7.0057645,7.149124,7.7187905,8.386545,9.092027,9.627739,9.937095,10.125726,10.465261,10.895341,10.540714,9.748463,9.016574,8.98262,8.907167,7.956466,6.398372,4.6516466,3.289729,3.470815,3.470815,3.451952,3.3840446,3.0445085,2.8143783,2.7691069,2.7125173,2.6106565,2.5616124,2.9200118,3.029418,2.9426475,2.595566,1.7882242,1.0601076,0.77338815,0.663982,0.56589377,0.45648763,0.4979865,0.49044126,0.47912338,0.48666862,0.4979865,0.49421388,0.46026024,0.42630664,0.39989826,0.35839936,0.39989826,0.47912338,0.59607476,0.7432071,0.9016574,1.1053791,1.1280149,1.1581959,1.2713746,1.4147344,1.3166461,1.1695137,1.0978339,1.1506506,1.2940104,1.4977322,1.6373192,1.6410918,1.5165952,1.3241913,1.6637276,1.8523588,1.8372684,1.7618159,1.9466745,2.463524,2.9803739,3.350091,3.5689032,3.7537618,3.4745877,3.712263,3.9084394,4.036709,4.606375,5.304311,5.9909286,6.3644185,6.356873,6.145606,6.1833324,6.4436436,6.8850408,7.322665,7.432071,1.2525115,1.3317367,1.4147344,1.6146835,1.8976303,2.0900342,1.9466745,1.9127209,1.8749946,1.7957695,1.7240896,1.5769572,1.5015048,1.4939595,1.5467763,1.659955,1.7995421,1.8334957,1.8334957,1.8523588,1.9202662,2.142851,2.3918443,2.5767028,2.7200627,2.9615107,3.8141239,4.515832,5.13077,5.723072,6.3455553,7.3905725,8.488406,9.948412,11.5857315,12.721292,13.800262,15.082954,16.644821,19.470518,25.431265,28.041922,30.977024,34.760967,39.269253,43.766224,46.60701,42.977745,33.949852,23.443092,18.199142,14.70192,11.981857,9.97482,8.288457,6.1795597,3.85185,2.4522061,1.6109109,1.1242423,0.9507015,1.3732355,1.1695137,0.69039035,0.25276586,0.150905,0.39989826,0.5319401,0.44894236,0.26408374,0.29049212,0.331991,0.25276586,0.16222288,0.10940613,0.08677038,0.181086,0.1961765,0.22258487,0.2678564,0.26031113,0.20749438,0.20372175,0.15845025,0.06790725,0.030181,0.06790725,0.05281675,0.030181,0.026408374,0.02263575,0.02263575,0.049044125,0.06413463,0.056589376,0.02263575,0.018863125,0.071679875,0.1659955,0.30935526,0.5357128,0.66775465,0.5394854,0.62625575,0.91297525,0.90920264,1.2600567,1.7580433,2.6898816,3.6971724,3.7650797,5.0062733,4.485651,3.7499893,3.8820312,5.485397,5.311856,4.5196047,4.4177437,5.0741806,5.300538,6.356873,6.3531003,6.2814207,6.058836,4.5422406,4.689373,3.3689542,2.4333432,2.305074,1.961765,1.6637276,1.6109109,1.690136,1.7995421,1.8599042,1.3317367,1.5279131,1.8259505,1.9240388,1.8636768,1.8900851,1.81086,1.7580433,1.8938577,2.3805263,2.535204,2.71629,3.108643,3.5462675,3.5047686,5.304311,5.515578,6.3908267,8.09228,8.688355,7.9300575,8.058327,8.707218,9.906913,12.091263,10.510533,10.8576145,11.796998,12.313848,11.69891,14.713238,15.588487,15.792209,15.943113,15.792209,15.916705,15.848798,15.331948,14.667966,14.762281,13.773854,12.736382,12.019584,11.9064045,12.604341,12.370438,12.31762,12.23085,12.102581,12.151625,12.038446,12.291212,12.838243,13.856852,15.758255,15.565851,15.758255,15.362129,14.366156,13.72481,14.139798,15.026365,15.396083,15.147089,15.071637,15.720529,15.82239,15.660167,15.603577,16.094019,16.33924,17.674747,19.059301,20.142044,21.262514,22.847017,23.043194,21.983086,19.91946,17.229578,15.814844,15.528125,15.313085,15.033911,15.456445,14.901869,14.34352,14.181297,14.535924,15.237633,14.124708,13.396591,13.626721,14.234114,13.502225,13.128735,14.037937,14.6302395,14.437836,14.136025,13.694629,13.879487,14.999957,16.97304,19.346022,20.8098,21.907633,22.862108,23.314823,22.349031,22.058538,22.126446,21.78691,21.224789,21.55678,22.288668,23.824127,25.204908,25.959433,26.102793,23.8279,21.541689,19.48938,18.006739,17.527617,17.320122,17.77661,18.233097,18.384,18.270823,18.199142,18.580177,18.923487,18.802763,17.87847,17.16167,17.120173,17.301258,17.425755,17.369165,17.369165,17.935059,18.976303,19.836462,19.274342,18.51227,16.335466,12.691111,8.83926,7.375482,5.8211603,3.9461658,2.5427492,2.0900342,2.7426984,2.4522061,1.7127718,1.1808317,1.0676528,1.1355602,2.2786655,2.9351022,3.5953116,4.447925,5.379763,8.397863,8.975075,7.7037,5.8966126,5.6098933,7.8810134,7.8017883,7.0170827,6.1606965,4.889322,5.1269975,6.168242,6.1229706,4.821415,3.7990334,3.2633207,3.5764484,4.7648253,5.975838,5.4665337,3.3350005,4.168751,4.3422914,3.0143273,2.1315331,3.62172,4.425289,4.749735,4.425289,2.8822856,3.5538127,3.5160866,4.0291634,5.3759904,6.858632,4.659192,3.8858037,4.0970707,4.961002,6.255012,7.9225125,8.620448,8.590267,7.624475,5.070408,5.1534057,4.123479,3.9159849,4.587512,4.3121104,2.2748928,1.780679,1.8033148,2.0070364,2.7804246,5.0062733,6.7567716,6.4210076,4.5497856,3.8556228,3.8669407,4.6252384,5.8400235,6.5832305,5.292993,5.9305663,5.6589375,5.1345425,4.5799665,3.7763977,3.92353,4.82896,5.80607,6.730363,8.039464,8.243186,10.672756,12.67602,13.890805,16.237377,10.469034,7.039718,6.115425,6.0286546,3.2784111,3.3878171,4.957229,5.010046,3.531177,3.4557245,1.327964,0.362172,0.0452715,0.0,0.0,0.003772625,0.02263575,0.026408374,0.033953626,0.10940613,0.20372175,0.35085413,0.34330887,0.20372175,0.1659955,0.15467763,0.13958712,0.15845025,0.211267,0.241448,0.35085413,0.43007925,0.45648763,0.41876137,0.32067314,0.30935526,0.32821837,0.55080324,1.0223814,1.6788181,1.4524606,1.7655885,2.5767028,3.2557755,2.6031113,2.9652832,2.867195,2.8445592,2.9426475,2.7351532,3.187868,3.4745877,3.2935016,2.867195,2.957738,2.0975795,2.033445,2.1843498,2.3880715,2.8785129,2.969056,2.957738,3.2105038,3.6556737,3.7801702,4.825187,5.2137675,5.3646727,5.4778514,5.541986,4.8855495,4.719554,4.2781568,3.9461658,5.243949,5.1043615,5.142088,5.2137675,5.311856,5.5759397,5.8890676,5.8626595,5.9230213,6.307829,7.069899,7.1264887,7.4999785,8.311093,9.084481,8.744945,9.597558,10.876478,11.514051,11.672502,12.728837,11.7026825,12.883514,13.894578,13.977575,13.985121,15.70921,15.70921,14.954685,13.736128,11.668729,12.853333,14.109617,15.241405,16.014793,16.165699,16.724047,18.233097,18.417955,17.45971,17.969013,16.931541,16.893814,18.663176,20.885252,20.070366,20.16468,19.470518,19.47429,19.38752,16.13929,16.45619,20.655123,20.421219,17.139036,21.881226,17.912424,13.721037,11.106608,10.352083,10.208723,13.000465,13.460726,11.774363,9.484379,9.488152,8.084735,7.3717093,9.348565,12.340257,10.997202,10.7218,11.423509,10.091772,6.9265394,5.3458095,5.511805,5.564622,4.745962,3.6745367,4.349837,5.138315,5.2628117,5.111907,4.9685473,4.9760923,5.7004366,6.6058664,6.4021444,5.6363015,6.6813188,6.673774,6.937857,7.326438,7.654656,7.677292,7.9791017,7.8131065,7.443389,7.281166,7.858378,7.854605,7.5829763,7.4169807,7.6018395,8.2507305,8.6581745,7.61693,6.5455046,6.2663302,6.960493,6.5040054,6.2097406,5.624984,4.8063245,4.3347464,4.7006907,4.9157305,5.0025005,4.9232755,4.5761943,5.726845,5.6400743,5.194905,4.9723196,5.2628117,4.8855495,4.8440504,5.13077,5.3986263,4.9421387,5.100589,5.093044,5.081726,5.142088,5.281675,5.2326307,5.3458095,5.59103,5.938112,6.3644185,7.383027,7.405663,7.0170827,6.590776,6.300284,5.8928404,5.9305663,5.8588867,5.6287565,5.7419353,6.5040054,6.6813188,6.8699503,7.375482,8.231868,8.89585,9.676784,10.076681,10.125726,10.378491,10.487898,10.140816,9.465516,8.91094,9.22784,8.869441,7.7640624,6.398372,5.0025005,3.5236318,3.3576362,3.350091,3.3576362,3.3350005,3.3010468,2.8445592,2.71629,2.637065,2.584248,2.7917426,2.8181508,2.957738,2.6106565,1.7882242,1.1431054,0.7092535,0.5470306,0.47535074,0.39989826,0.3169005,0.35839936,0.392353,0.4074435,0.4074435,0.4074435,0.362172,0.29049212,0.23013012,0.1961765,0.16976812,0.18485862,0.23013012,0.32067314,0.44139713,0.55080324,0.76584285,0.9393836,1.0223814,1.0487897,1.1091517,1.1619685,1.146878,1.146878,1.2034674,1.327964,1.4977322,1.5430037,1.5316857,1.4864142,1.388326,1.9240388,2.1805773,2.1466236,2.0145817,2.1654868,2.6068838,3.1614597,3.6783094,3.9801195,3.863168,3.4745877,3.7877154,4.183841,4.504514,5.0515447,5.292993,5.6853456,6.066381,6.2625575,6.085244,6.0814714,6.217286,6.387054,6.590776,6.94163,1.4222796,1.478869,1.6524098,1.8297231,1.9542197,2.052308,1.9278114,1.8448136,1.7769064,1.690136,1.5430037,1.5015048,1.4864142,1.5203679,1.6637276,1.9957186,1.991946,2.0485353,2.0749438,2.0975795,2.2484846,2.3654358,2.7389257,2.8785129,2.8596497,3.3312278,4.0291634,4.8327327,5.7570257,6.719045,7.5527954,8.492179,9.64283,11.223559,12.868423,13.63804,14.339747,15.4074,17.512526,21.311558,27.430756,30.214954,33.764996,36.967953,40.638718,47.531303,49.176167,44.98478,35.84371,25.314314,19.625195,16.275105,13.834216,11.480098,8.846806,6.009792,3.6330378,2.203213,1.358145,1.0186088,1.3656902,1.4977322,1.1921495,0.7582976,0.3961256,0.18863125,0.35462674,0.56212115,0.5093044,0.29803738,0.41121614,0.27917424,0.21881226,0.2263575,0.2263575,0.071679875,0.17731337,0.15845025,0.15467763,0.18863125,0.15467763,0.13204187,0.14335975,0.120724,0.060362,0.041498873,0.090543,0.06790725,0.049044125,0.049044125,0.0150905,0.033953626,0.049044125,0.0452715,0.026408374,0.0150905,0.00754525,0.033953626,0.124496624,0.31312788,0.6451189,0.8186596,0.59607476,0.66775465,1.0035182,0.8224323,1.3619176,2.1805773,3.4255435,4.3875628,3.5047686,4.5233774,4.191386,3.7348988,4.0706625,5.7872066,6.63982,6.722818,6.9755836,7.5490227,7.809334,8.499724,7.911195,7.2962565,6.673774,4.8365054,5.485397,4.719554,3.5424948,2.6106565,2.1994405,2.0862615,1.6109109,1.629774,2.0673985,1.9089483,1.1129243,1.056335,1.327964,1.5203679,1.2411937,1.6976813,1.9278114,1.8938577,1.8825399,2.4786146,2.6823363,2.7728794,3.3727267,4.5460134,5.80607,7.0963078,6.56814,7.0246277,8.827943,9.891823,10.042727,10.227587,11.272603,13.358865,16.022339,13.43809,11.883769,11.815862,12.393073,11.491416,14.045483,14.928277,14.803781,14.637785,15.690348,16.0412,15.735619,14.705692,13.490907,13.241914,12.81938,11.808316,10.925522,10.585986,10.914205,11.664956,12.653384,13.158916,13.223051,13.641812,12.67602,12.559069,12.823153,13.43809,14.830189,15.154634,15.746937,15.871433,15.331948,14.475562,14.675511,15.565851,16.06761,15.977067,15.961976,15.377219,14.999957,14.7321005,14.566105,14.588741,15.294222,15.90916,16.580687,17.380484,18.289686,20.50799,21.353058,20.462717,18.5085,17.191853,15.682802,15.430037,15.565851,15.803526,16.463736,15.999702,14.950912,14.313339,14.517061,15.422491,14.950912,14.275613,14.094527,14.203933,13.517315,12.377983,12.7477,13.321139,13.45318,13.189097,13.132507,13.321139,14.317112,16.078928,17.972786,19.519562,20.77962,21.87368,22.39053,21.394556,21.711456,22.171717,22.213217,22.07363,22.760246,22.948877,24.008986,24.752193,24.963459,25.39354,23.997667,21.820864,19.527107,17.784155,17.282394,17.05981,17.444618,18.372684,19.610106,20.73812,21.277605,21.519053,21.915178,22.194353,21.35683,20.225042,20.07791,20.010002,19.681786,19.300749,19.229069,19.670467,20.911661,22.326395,22.382984,20.46649,17.112627,13.290957,9.763554,7.0887623,5.191132,3.7348988,2.848332,2.5125682,2.5804756,2.282438,1.6373192,1.1695137,1.0299267,0.995973,2.2296214,2.7389257,3.6028569,4.9534564,5.983383,9.005256,8.526133,7.2170315,6.2814207,5.4250345,7.492433,8.567632,8.043237,6.466279,5.553304,5.9117036,5.5570765,4.798779,3.8782585,2.987919,3.0030096,6.579458,7.7037,5.6325293,4.9044123,2.1843498,2.4333432,2.674791,2.0108092,1.6373192,3.6254926,5.6815734,6.828451,6.2135134,3.108643,4.4818783,4.1989317,4.8930945,7.567886,11.59705,6.428553,4.768598,4.3007927,3.8480775,3.3538637,3.4745877,4.991183,6.096562,6.0701537,5.27413,4.459243,3.6028569,3.651901,4.1536603,3.2670932,2.7615614,2.8256962,2.7502437,2.5804756,3.1350515,4.5422406,6.149379,6.255012,4.9647746,4.1989317,4.478106,4.6629643,5.142088,5.5985756,5.0251365,5.311856,5.3948536,6.039973,6.488915,4.4743333,4.8063245,5.7192993,6.19465,6.198423,6.651138,7.194396,9.186342,11.736636,14.3095665,16.72782,10.272858,6.6322746,5.353355,4.991183,3.1199608,2.9200118,4.919503,4.991183,2.9615107,2.6068838,0.80734175,0.14335975,0.0,0.0,0.0,0.0,0.018863125,0.041498873,0.056589376,0.056589376,0.29049212,0.38103512,0.33576363,0.22258487,0.13958712,0.124496624,0.14713238,0.1961765,0.2565385,0.29426476,0.3470815,0.36594462,0.40367088,0.422534,0.31312788,0.33576363,0.35839936,0.5017591,0.83752275,1.4034165,1.1883769,1.6222287,2.3918443,2.9539654,2.546522,2.7691069,2.5238862,2.4408884,2.5540671,2.282438,2.9237845,3.2821836,3.138824,2.8747404,3.482133,2.3880715,1.9844007,1.9994912,2.2862108,2.8030603,2.7502437,2.7804246,3.289729,4.025391,4.093298,5.3080835,5.541986,5.6287565,5.80607,5.7079816,5.070408,4.7874613,4.4441524,4.255521,5.05909,4.8440504,4.708236,4.7836885,5.194905,6.058836,6.092789,5.8437963,5.794752,6.0248823,6.221059,7.2585306,7.598067,7.986647,8.495952,8.503497,8.726082,10.103089,11.065109,11.570641,13.102326,12.238396,12.826925,13.981348,14.830189,14.535924,15.992157,15.897841,14.652876,12.657157,10.303039,11.114153,11.706455,12.902377,14.362384,14.603831,15.660167,17.357847,17.448391,15.818617,14.494425,13.45318,13.992666,15.977067,18.485863,19.798737,19.708193,16.840998,15.414946,15.731846,14.1926155,11.8045435,17.048492,19.783646,18.700903,21.319103,13.298503,9.303293,6.832224,5.8400235,8.748717,10.838752,10.86516,10.057818,9.344792,9.367428,8.367682,6.530414,6.8359966,8.903395,9.009028,8.416726,8.420499,7.141579,5.323174,6.3116016,6.907676,6.7379084,5.80607,4.9421387,5.794752,6.911449,7.194396,7.0057645,6.530414,5.7909794,5.7494807,5.5382137,5.560849,6.058836,7.1000805,6.541732,7.183078,7.8998766,8.228095,8.345046,8.379,8.156415,8.0206,8.084735,8.216777,7.8319697,7.598067,7.4735703,7.541477,8.050782,8.503497,8.099826,7.224577,6.643593,7.4811153,6.802043,6.156924,5.617439,5.119452,4.4630156,5.010046,4.9044123,4.821415,4.859141,4.538468,5.2854476,5.541986,5.270357,4.8365054,5.0138187,5.142088,5.402399,5.6363015,5.666483,5.2590394,5.0062733,4.6214657,4.459243,4.5724216,4.715781,4.5799665,4.9119577,5.2552667,5.50426,5.885295,6.688864,6.722818,6.304056,5.8098426,5.6778007,5.4740787,5.379763,5.3269467,5.3986263,5.8211603,6.0550632,6.138061,6.3531003,6.881268,7.7942433,8.816625,9.7296,9.982366,9.763554,9.989911,10.291721,9.759781,8.8618965,8.262049,8.820397,8.66572,7.435844,6.156924,5.1760416,4.1612053,3.6368105,3.7198083,3.7273536,3.5274043,3.5575855,2.9200118,2.7313805,2.637065,2.5880208,2.867195,2.848332,2.704972,2.022127,1.0336993,0.6149379,0.48666862,0.40367088,0.35462674,0.31312788,0.27540162,0.26408374,0.2678564,0.271629,0.2678564,0.26408374,0.241448,0.181086,0.124496624,0.09808825,0.08677038,0.09808825,0.10940613,0.150905,0.2263575,0.32067314,0.44894236,0.6451189,0.80734175,0.875249,0.8186596,0.965792,1.116697,1.2864652,1.448688,1.4977322,1.4750963,1.3958713,1.327964,1.3091009,1.3656902,1.8976303,2.2069857,2.1994405,2.0636258,2.2447119,2.6936543,3.108643,3.440634,3.6443558,3.6971724,3.6330378,4.08198,4.640329,5.111907,5.4967146,5.5759397,5.7872066,6.0512905,6.277648,6.3908267,6.255012,6.1418333,6.006019,6.017337,6.5341864,1.6033657,1.5769572,1.8221779,1.9542197,1.9164935,1.9504471,1.9278114,1.7844516,1.6448646,1.539231,1.388326,1.4373702,1.6033657,1.7089992,1.7957695,2.1466236,1.9164935,1.9881734,2.093807,2.2069857,2.5125682,2.686109,3.0218725,3.1199608,3.1576872,3.9159849,4.2630663,4.9647746,6.0776987,7.4811153,8.899622,10.329447,11.551778,12.811834,13.996439,14.637785,15.101818,16.592005,19.40261,23.548725,28.74363,32.414394,36.783092,39.069305,41.60828,51.88491,51.488785,45.863804,36.790638,27.400576,22.133991,18.983849,16.063837,12.438345,8.288457,4.927048,3.2935016,2.203213,1.5958204,1.5618668,2.3692086,1.9466745,1.4147344,1.0374719,0.80356914,0.44894236,0.32444575,0.56212115,0.5357128,0.28294688,0.5017591,0.32821837,0.23767537,0.33576363,0.452715,0.14713238,0.11317875,0.08677038,0.10186087,0.1358145,0.1056335,0.1056335,0.120724,0.120724,0.09808825,0.060362,0.06413463,0.05281675,0.060362,0.06790725,0.02263575,0.041498873,0.03772625,0.033953626,0.033953626,0.02263575,0.026408374,0.018863125,0.026408374,0.13204187,0.482896,0.67152727,0.39989826,0.4074435,0.7130261,0.6111652,1.0676528,2.505023,3.9801195,4.5724216,3.3651814,3.380272,3.410453,3.2444575,2.9539654,2.897376,4.98741,6.779407,7.8961043,8.280911,8.190369,7.8923316,7.3792543,6.9227667,6.058836,3.5877664,5.379763,5.541986,4.2064767,2.4559789,2.3088465,2.625747,1.9164935,1.6675003,2.0183544,1.7693611,1.2826926,1.3053282,1.4147344,1.3166461,0.8563859,1.8372684,2.3163917,2.4069347,2.2711203,2.123988,2.867195,3.0445085,4.104616,6.273875,8.571404,9.325929,8.367682,8.065872,9.088254,10.419991,12.3893,13.034419,13.800262,15.297995,17.30503,15.264041,12.268577,10.638803,10.710483,10.834979,11.510279,11.970539,11.974312,12.419481,15.339493,15.75071,15.049001,13.705947,12.377983,11.895086,12.14408,11.491416,10.725573,10.148361,9.574923,10.646348,12.468526,13.641812,14.102073,15.098045,14.320885,14.200161,14.313339,14.456699,14.622695,14.977322,15.286676,15.901614,16.380737,15.505488,15.596032,16.161926,16.70141,16.969267,16.97304,15.999702,15.807299,15.641303,15.324403,15.241405,15.467763,15.271586,15.199906,15.358356,15.422491,17.048492,17.938831,17.176762,15.803526,16.833452,16.524097,16.708956,16.94286,17.040947,17.097536,16.923996,15.924251,14.792462,14.04171,13.992666,14.637785,14.947141,15.01882,14.830189,14.230342,12.559069,12.37421,13.057055,13.713491,13.162688,13.117417,13.630494,14.743419,15.992157,16.403374,17.972786,19.4592,20.22127,20.123182,19.527107,20.673985,21.394556,21.866135,22.541435,24.156118,23.910898,24.088211,24.269297,24.227798,23.914669,22.967741,21.21347,19.410156,18.006739,17.120173,17.029629,17.399347,18.757492,20.934296,23.073374,24.205162,24.529608,25.186045,26.057522,25.729303,24.224026,23.639269,23.05074,22.31885,22.077402,21.97554,22.273579,23.156372,24.710693,26.913906,21.809546,16.818363,13.170234,10.627484,7.466025,5.100589,3.8367596,3.3312278,3.0369632,2.233394,1.9202662,1.4713237,1.1317875,0.9620194,0.8526133,1.8146327,2.2183034,3.731126,6.405917,8.710991,11.932813,10.140816,8.469543,8.167733,6.5756855,6.749226,8.956212,9.246704,7.2962565,6.4436436,6.5756855,4.4101987,2.5578396,1.8146327,1.177059,2.71629,10.382264,11.725319,5.7381625,2.8558772,0.69039035,0.08677038,0.11317875,0.2565385,0.44516975,1.9353566,4.8742313,7.3453007,7.816879,5.1269975,6.119198,5.4288073,5.666483,8.194141,13.143826,7.828197,5.5495315,3.5877664,2.0862615,4.032936,3.3840446,5.138315,6.620957,7.4471617,9.514561,6.2399216,4.45547,4.146115,4.266839,2.7313805,3.5575855,4.123479,3.8178966,3.1312788,3.682082,4.032936,5.2590394,6.0739264,5.8626595,4.6856003,5.0062733,5.6098933,5.481624,4.7874613,4.8666863,5.7909794,7.4169807,9.65792,10.691619,6.9680386,7.7640624,8.080963,7.4094353,5.9532022,4.61392,5.5004873,6.900131,9.710737,12.510024,11.555551,7.443389,5.3910813,4.1197066,3.1312788,2.674791,2.9313297,3.9763467,3.802806,2.6182017,2.8521044,0.65643674,0.0452715,0.0,0.003772625,0.02263575,0.003772625,0.030181,0.06790725,0.08677038,0.041498873,0.35839936,0.34330887,0.3055826,0.30935526,0.15467763,0.09808825,0.150905,0.241448,0.32067314,0.33953625,0.3470815,0.29803738,0.30935526,0.36594462,0.29426476,0.36971724,0.40367088,0.513077,0.7696155,1.177059,1.1657411,1.7391801,2.2069857,2.354118,2.4484336,2.637065,2.5389767,2.4522061,2.3993895,2.1315331,2.6785638,3.0369632,3.0671442,3.150142,4.1762958,2.9916916,2.2673476,1.9957186,2.161714,2.7540162,2.4786146,2.4484336,3.2142766,4.3724723,4.5912848,5.7192993,5.534441,5.3571277,5.564622,5.560849,5.243949,4.8402777,4.538468,4.5120597,4.9119577,4.8063245,4.508287,4.3875628,4.847823,6.349328,6.6624556,6.2889657,6.0286546,5.934339,5.2854476,7.0963078,7.7112455,7.726336,7.598067,7.6395655,8.375228,9.688101,10.559577,11.125471,12.653384,12.740154,12.845788,13.898351,15.045229,13.622949,15.335721,16.124199,15.297995,12.853333,9.450426,10.050273,10.186088,11.076427,12.792972,14.268067,15.011275,15.916705,15.365902,13.52486,12.344029,12.306303,13.622949,15.230087,17.08999,20.160908,20.277859,15.422491,12.215759,12.868423,15.154634,12.189351,14.8339615,18.059555,18.28214,13.370183,8.710991,8.831716,8.495952,6.960493,7.9715567,9.076936,9.5183325,9.42779,9.175024,9.382519,8.59404,7.54525,6.598321,5.847569,5.1458607,4.8365054,5.149633,5.696664,6.5341864,8.152642,8.511042,8.2507305,7.5490227,7.0472636,7.8508325,8.892077,9.367428,9.325929,8.526133,6.439871,5.73439,5.5759397,5.945657,6.587003,7.01331,6.9265394,7.8810134,8.480861,8.5563135,9.144843,8.744945,8.3525915,8.299775,8.503497,8.458225,8.29223,8.22055,8.096053,7.956466,8.016829,8.643084,8.688355,8.0206,7.1906233,7.4584794,7.3490734,6.628502,6.085244,5.8890676,5.572167,5.6098933,4.8440504,4.376245,4.52715,4.8025517,4.9044123,5.3986263,5.6098933,5.3873086,5.111907,5.560849,5.915476,5.7909794,5.342037,5.292993,4.776143,4.4215164,4.247976,4.2706113,4.515832,4.195159,4.5120597,4.666737,4.666737,5.292993,5.745708,5.73439,5.50426,5.3156285,5.4476705,5.2892203,5.111907,5.1232247,5.50426,6.4134626,5.66271,5.413717,5.666483,6.3417826,7.2924843,8.854351,9.635284,9.590013,9.171251,9.325929,9.97482,9.152389,7.9941926,7.3453007,7.748972,8.265821,7.201941,5.907931,5.0515447,4.5950575,4.063117,4.2517486,4.2291126,3.7952607,3.4670424,2.897376,2.7238352,2.595566,2.4710693,2.595566,2.6785638,2.1503963,1.3543724,0.63002837,0.32444575,0.2867195,0.27917424,0.29426476,0.3055826,0.27917424,0.23013012,0.181086,0.14713238,0.1358145,0.14713238,0.15467763,0.1358145,0.124496624,0.120724,0.10940613,0.120724,0.13958712,0.12826926,0.10940613,0.16222288,0.23390275,0.30935526,0.49421388,0.7130261,0.7092535,0.8262049,1.086516,1.4298248,1.7089992,1.7014539,1.5354583,1.4147344,1.3204187,1.2940104,1.4147344,1.6524098,1.9164935,1.9768555,1.9353566,2.2220762,2.625747,2.8332415,2.8445592,2.897376,3.4745877,3.9801195,4.5912848,5.070408,5.3156285,5.3910813,5.7192993,6.0512905,6.221059,6.3116016,6.6850915,6.398372,6.0701537,5.881522,5.9796104,6.458734,1.1129243,1.0902886,1.3770081,1.5845025,1.6675003,1.9391292,2.1202152,1.9466745,1.7957695,1.7655885,1.6939086,1.5958204,1.690136,1.6712729,1.5354583,1.5731846,1.7052265,1.6373192,1.8334957,2.3390274,2.7917426,2.927557,2.8219235,2.8596497,3.2444575,4.014073,4.7836885,5.5495315,6.5643673,7.7640624,8.790216,11.400873,13.419228,14.418973,14.879233,16.173243,16.893814,19.429018,23.088465,26.815819,29.158619,33.738586,38.81654,41.325333,42.9702,50.247593,51.16434,43.40782,34.68174,28.86058,26.016022,20.60985,15.165953,10.627484,7.17176,4.1800685,3.289729,2.7087448,2.8634224,3.4179983,3.2972744,2.6483827,2.3767538,1.9994912,1.4147344,0.9016574,0.52062225,0.44516975,0.392353,0.32821837,0.48666862,0.6111652,0.43007925,0.35839936,0.42630664,0.3055826,0.24522063,0.17354076,0.124496624,0.120724,0.1659955,0.1659955,0.23013012,0.23013012,0.14713238,0.060362,0.03772625,0.041498873,0.06413463,0.08299775,0.0452715,0.056589376,0.041498873,0.041498873,0.056589376,0.0452715,0.071679875,0.041498873,0.02263575,0.090543,0.33576363,0.5055317,0.30181,0.63002837,1.2336484,0.67152727,2.282438,4.2064767,6.092789,7.224577,6.515323,4.587512,3.874486,3.0143273,2.082489,2.595566,3.2670932,3.2670932,3.5877664,4.5422406,5.798525,5.2364035,5.583485,5.3269467,4.1612053,2.9916916,3.8443048,4.4516973,3.9574835,2.7841973,2.625747,3.0897799,2.867195,2.2975287,1.720317,1.4637785,1.8070874,1.8448136,1.5845025,1.1393328,0.7469798,1.4562333,2.1013522,2.5767028,2.757789,2.5012503,3.2331395,4.0782075,5.168496,6.5832305,8.314865,10.038955,10.70671,10.114408,9.092027,9.507015,13.045737,15.935568,16.471281,14.984866,13.822898,11.431054,9.808825,9.276885,9.431562,9.125979,9.088254,9.4013815,9.590013,10.26154,13.106099,13.253232,12.751472,11.944131,11.332966,11.566868,10.661438,10.299266,10.469034,10.684074,9.963503,10.585986,10.933067,11.68382,12.925014,14.143571,14.803781,16.214743,16.837225,16.67123,17.255987,16.840998,16.29774,15.633758,15.188588,15.641303,18.191597,17.70493,17.274849,17.546478,16.693865,17.191853,17.384256,16.712729,15.690348,15.897841,15.618668,15.539442,15.422491,14.875461,13.336229,13.505998,13.807808,13.649357,13.660675,15.686575,19.225298,20.323132,19.47429,17.916197,17.625704,18.406637,18.5085,17.274849,15.17727,13.807808,14.358611,14.679284,14.698147,14.351066,13.59654,12.423254,12.479843,13.845533,15.260268,14.11339,13.456953,13.920986,14.652876,15.131999,15.181043,16.927769,18.836716,19.772327,19.466745,18.53868,19.478064,20.100546,20.843754,22.081175,24.091984,23.850534,24.612606,25.672712,25.831163,23.375185,21.032385,19.960958,19.308294,18.61036,17.7917,17.14658,17.63325,19.36111,21.986858,24.73333,26.151836,27.174217,28.12492,29.011486,29.524563,27.962696,26.812046,25.75571,24.955914,25.054003,24.933279,25.129456,25.276588,25.767029,27.755201,20.89657,14.720782,10.529396,8.431817,7.3717093,5.9305663,4.7836885,4.0970707,3.5538127,2.3201644,1.8787673,1.5580941,1.2487389,0.97333723,0.9016574,1.3656902,1.9730829,3.8895764,7.2698483,11.261286,13.422999,13.43809,12.121444,10.446399,9.567377,7.3453007,8.952439,9.684328,8.386545,7.4471617,5.1156793,2.9652832,1.7316349,1.2864652,0.6413463,1.3015556,3.1124156,3.6028569,2.282438,0.67152727,0.34330887,0.20372175,0.3734899,0.7394345,0.94692886,4.0480266,4.0970707,4.304565,5.907931,8.179051,11.427281,12.064855,10.359629,8.273367,9.446653,7.1378064,5.0251365,3.3312278,2.2862108,2.0900342,3.2972744,5.010046,7.3000293,9.258021,9.001483,6.888813,5.081726,3.9273026,3.6481283,4.3196554,3.904667,3.9273026,3.9763467,4.2706113,5.66271,5.696664,5.9909286,6.7152724,7.1000805,5.4174895,4.9760923,5.0968165,5.50426,6.198423,7.432071,8.578949,13.800262,18.23687,18.746174,13.898351,12.117672,9.548513,8.3525915,8.971302,10.133271,8.75249,8.473316,9.001483,10.038955,11.261286,8.586494,5.311856,3.0897799,2.505023,3.0671442,3.3236825,2.9766011,2.957738,2.8030603,0.6413463,0.12826926,0.0,0.0,0.02263575,0.1056335,0.02263575,0.0,0.0,0.041498873,0.21503963,0.23767537,0.34330887,0.4074435,0.3734899,0.29049212,0.15467763,0.18485862,0.26031113,0.30181,0.29049212,0.47157812,0.4074435,0.32821837,0.30935526,0.26031113,0.331991,0.422534,0.66775465,0.935611,0.8224323,0.95824677,1.7165444,2.293756,2.4710693,2.595566,2.9464202,3.338773,3.1312788,2.5804756,2.837014,3.0331905,3.2029586,3.4594972,3.7952607,4.0895257,3.5538127,2.8030603,2.3390274,2.4484336,3.2029586,2.6068838,2.4823873,3.150142,4.2630663,4.8365054,5.0553174,4.8553686,4.6856003,4.7421894,4.9760923,5.7419353,5.3571277,4.7044635,4.349837,4.5309224,4.689373,5.142088,5.2137675,5.1760416,6.224831,6.8737226,6.33801,5.66271,5.2250857,4.7610526,5.8588867,7.0774446,7.4735703,7.322665,8.103599,8.956212,9.673011,9.839006,9.846551,10.895341,11.332966,11.857361,13.151371,14.441608,13.487134,14.671739,15.856343,16.15438,14.93205,11.793225,11.563096,12.053536,12.189351,12.313848,14.2077055,14.460471,14.169979,13.340002,12.355347,11.978085,11.306557,13.328684,14.558559,14.898096,17.610613,18.402864,13.905896,12.913695,18.02183,25.604805,16.203424,12.913695,15.214996,18.97253,16.433554,11.012292,8.797762,7.3151197,6.1644692,7.020855,7.61693,7.8961043,8.560086,9.491924,9.733373,9.699419,10.27663,9.635284,7.586749,5.583485,6.1342883,6.620957,7.2358947,7.786698,7.673519,8.2507305,9.473062,10.016319,9.789962,9.948412,9.352338,9.25425,9.510788,9.159933,6.439871,6.2323766,6.4926877,6.9680386,7.515069,8.088508,8.880759,8.933576,8.590267,8.375228,8.986393,9.035437,8.710991,8.526133,8.650629,8.89585,8.956212,9.329701,9.97482,10.567122,10.484125,10.34831,9.318384,8.503497,8.228095,7.9941926,8.130007,8.246958,7.496206,6.2927384,6.3153744,5.87775,5.7570257,5.2137675,4.436607,4.5460134,4.9119577,4.776143,4.8742313,5.3080835,5.5382137,6.126743,5.9494295,5.292993,4.5724216,4.3649273,4.2291126,4.2706113,4.398881,4.5761943,4.821415,4.1989317,4.08198,4.08198,4.172523,4.6856003,5.221313,5.2628117,5.2137675,5.251494,5.3269467,5.2628117,5.2288585,5.3344917,5.7909794,6.9265394,5.9494295,5.3684454,5.458988,6.2663302,7.5829763,8.461998,8.846806,8.944894,8.888305,8.729855,8.801534,8.107371,7.3717093,7.1981683,8.043237,8.137552,7.356619,6.3153744,5.4250345,4.9119577,4.398881,3.8971217,3.7613072,3.712263,2.806833,2.4522061,2.493705,2.354118,2.0070364,1.9844007,1.4826416,0.95447415,0.5357128,0.31312788,0.33576363,0.24899325,0.23767537,0.27917424,0.32821837,0.3055826,0.2565385,0.23390275,0.211267,0.18485862,0.18485862,0.18485862,0.18485862,0.21503963,0.2565385,0.24522063,0.2565385,0.3961256,0.36594462,0.16222288,0.0754525,0.10186087,0.09808825,0.116951376,0.18485862,0.3055826,0.36594462,0.7922512,1.1846043,1.3807807,1.478869,1.6260014,1.7089992,1.7882242,1.8787673,1.9542197,1.9655377,1.9579924,1.9881734,2.1843498,2.746471,2.5767028,2.6521554,2.8030603,3.0218725,3.4481792,4.376245,5.240176,5.3986263,4.90064,4.485651,5.05909,5.613666,5.915476,6.0286546,6.3342376,6.307829,6.043745,6.089017,6.40969,6.40969,1.418507,1.539231,1.8938577,2.1654868,2.282438,2.41448,2.5767028,2.516341,2.3767538,2.252257,2.1692593,2.0145817,1.8674494,1.7354075,1.6222287,1.5241405,1.5807298,1.6373192,1.7354075,1.9579924,2.4371157,2.4559789,2.584248,2.897376,3.4142256,4.123479,4.647874,5.5457587,6.6624556,8.062099,10.0465,12.355347,13.917213,14.901869,15.818617,17.50498,19.768555,22.33394,25.650078,30.00746,35.55699,42.12513,50.25891,54.718155,56.057434,60.644947,56.619556,47.74257,39.974735,34.428974,27.34776,20.006231,14.011529,10.167224,7.816879,4.878004,3.2633207,3.6368105,4.738417,5.4212623,4.6629643,3.380272,3.097325,2.8030603,2.0787163,1.1091517,0.79602385,0.8639311,0.8224323,0.6187105,0.6111652,0.5093044,0.40367088,0.41876137,0.48666862,0.35462674,0.39989826,0.34330887,0.30181,0.32821837,0.3734899,0.3169005,0.35085413,0.34330887,0.2565385,0.16976812,0.1659955,0.181086,0.27917424,0.3470815,0.1056335,0.090543,0.06790725,0.06790725,0.0754525,0.033953626,0.018863125,0.00754525,0.049044125,0.19994913,0.543258,0.6149379,0.43007925,1.1581959,2.1692593,1.0487897,1.8221779,2.4861598,2.9049213,2.916239,2.354118,1.5165952,1.3166461,1.1619685,1.1846043,2.214531,2.0749438,1.9504471,2.1353056,2.7087448,3.5274043,2.595566,3.1765501,3.218049,2.7087448,3.6745367,4.0103,3.4557245,3.1954134,3.4444065,3.440634,3.429316,2.625747,2.0900342,2.1051247,2.173032,2.7200627,2.2258487,1.8749946,1.9730829,1.9429018,2.282438,1.9768555,2.1692593,2.916239,3.199186,3.832987,4.8402777,5.9418845,7.1264887,8.631766,10.042727,11.974312,12.66093,12.038446,11.740409,13.347548,15.645076,16.81459,15.988385,13.226823,11.408418,9.608876,8.941121,9.125979,8.488406,8.952439,9.688101,9.084481,7.960239,9.556059,8.639311,8.643084,8.420499,7.805561,7.647111,8.197914,9.416472,10.54826,11.23865,11.514051,11.521597,11.480098,11.815862,12.774108,14.4152,14.973549,15.577168,16.116653,16.588232,17.086218,17.697384,17.50498,17.093763,16.931541,17.372938,19.48561,21.507734,21.262514,19.051756,17.670975,18.119919,18.576405,18.03692,16.675003,15.826162,15.848798,15.648849,15.154634,14.162435,12.310076,11.936585,11.9064045,11.910177,12.151625,13.36641,17.708702,20.598532,20.972023,19.296976,17.599297,18.274595,19.191343,19.357338,18.327412,16.237377,15.799753,15.471535,15.369675,15.24895,14.524607,13.555041,13.815352,15.260268,17.006994,17.323895,16.52787,16.15438,16.31283,16.74291,16.82968,16.690092,16.893814,17.425755,17.927513,17.686066,18.459454,19.346022,20.621168,22.17549,23.495909,24.031622,24.639013,25.32186,25.604805,24.537153,21.409647,19.828917,19.153618,18.89708,18.731083,18.387774,19.149845,20.587215,22.469755,24.759737,26.555508,27.857063,29.041668,29.939552,29.818829,29.241617,28.264507,27.208172,26.51778,26.751684,26.834682,28.015512,28.766266,28.871899,29.426476,27.547709,20.862616,14.373701,10.069136,6.907676,7.888559,7.3075747,5.5797124,3.4972234,2.2447119,1.991946,1.599593,1.1242423,0.784706,0.98465514,1.3505998,1.7240896,3.0030096,6.047518,11.6875925,19.708193,23.782627,21.934042,15.562078,9.457971,8.59404,9.167479,8.09228,5.9003854,6.72659,3.8103511,1.871222,0.8111144,0.41498876,0.38480774,1.1883769,1.478869,1.3770081,1.1657411,1.2940104,4.1008434,4.429062,3.0445085,1.2902378,1.116697,2.263575,1.9542197,2.1654868,3.6028569,5.6891184,9.393836,14.173752,16.120426,14.807553,13.302276,11.465008,7.575431,3.7914882,1.6109109,1.8938577,2.8596497,2.6068838,3.078462,4.8063245,6.903904,5.564622,4.496969,3.712263,3.5575855,4.708236,3.92353,3.3727267,3.097325,3.7877154,6.771862,6.964266,6.9227667,6.458734,6.0286546,6.749226,6.952948,8.4544525,9.4013815,8.880759,6.930312,7.8923316,19.04421,32.19181,38.009197,26.034885,17.180534,12.691111,9.261794,6.48137,6.8133607,9.103344,8.956212,8.52236,8.582722,8.563859,7.8734684,6.277648,4.104616,2.5917933,3.8971217,3.361409,3.218049,3.1539145,2.4823873,0.17731337,0.033953626,0.0,0.0,0.0150905,0.08299775,0.42630664,0.20372175,0.0,0.060362,0.29803738,0.23390275,0.17354076,0.23013012,0.41121614,0.6073926,0.3169005,0.2867195,0.30935526,0.32067314,0.3734899,0.422534,0.42630664,0.362172,0.29049212,0.36971724,0.3734899,0.38103512,0.5696664,0.8299775,0.7997965,0.9922004,1.9542197,2.776652,3.0218725,2.71629,3.1199608,3.5274043,3.1539145,2.3654358,2.6785638,2.8143783,3.3123648,3.8178966,4.146115,4.285702,4.1083884,3.3840446,2.7200627,2.5125682,2.9464202,3.0520537,3.048281,3.3236825,3.9159849,4.5196047,4.9044123,4.7308717,4.776143,4.9345937,4.217795,4.4894238,4.689373,4.8138695,4.9044123,5.0553174,4.5988297,4.957229,5.4703064,5.7192993,5.5306683,6.488915,6.3832817,6.096562,5.9607477,5.7494807,6.5643673,7.4169807,7.748972,7.696155,8.126234,8.843033,9.710737,9.876732,9.5032425,9.771099,10.876478,11.766817,13.392818,14.996184,14.124708,14.351066,15.660167,16.177015,15.147089,12.966512,11.981857,11.838497,12.045992,12.434572,13.155144,13.502225,13.140053,12.604341,12.102581,11.54046,10.280403,13.20796,15.116908,14.818871,15.165953,13.079691,10.623712,19.987368,35.5004,33.64804,24.639013,18.23687,16.180788,16.769318,14.84528,18.52736,13.381501,8.695901,7.4396167,6.2625575,9.944639,9.537196,10.638803,13.430545,12.687338,11.117926,11.400873,11.400873,10.306811,8.646856,7.8206515,6.900131,6.7454534,7.1076255,6.6360474,6.9265394,8.299775,8.937348,8.899622,10.133271,10.940613,10.910432,10.714255,10.038955,7.598067,7.4509344,7.3490734,7.3717093,7.515069,7.696155,7.964011,8.080963,8.360137,8.8769865,9.488152,8.854351,8.635539,8.646856,8.605357,8.126234,8.635539,8.771353,9.016574,9.424017,9.6051035,10.386037,9.820143,8.99771,8.469543,8.228095,8.216777,7.7904706,7.1264887,6.560595,6.571913,6.428553,5.8890676,5.4250345,5.2590394,5.3910813,5.775889,5.541986,5.081726,4.851596,5.3684454,5.1835866,5.1458607,4.768598,4.104616,3.731126,4.1800685,4.346064,4.515832,4.7912335,5.0553174,4.715781,4.2064767,4.032936,4.146115,3.9159849,4.38379,4.659192,4.8402777,4.9157305,4.7648253,4.9647746,5.3571277,5.7004366,6.096562,6.9755836,6.2323766,5.5570765,5.251494,5.5759397,6.730363,7.254758,7.8621507,8.624221,9.295748,9.303293,9.307066,8.805306,8.016829,7.4207535,7.786698,7.326438,6.470052,5.764571,5.292993,4.6818275,4.568649,4.115934,3.5651307,3.0520537,2.5880208,2.0183544,1.931584,1.9579924,1.9240388,1.8599042,1.4977322,0.91674787,0.4640329,0.2678564,0.21503963,0.2565385,0.27540162,0.2867195,0.28294688,0.21881226,0.211267,0.20749438,0.1961765,0.18485862,0.1961765,0.25276586,0.32067314,0.3734899,0.41498876,0.452715,0.4640329,0.5885295,0.6526641,0.5696664,0.35839936,0.20749438,0.150905,0.13958712,0.14335975,0.15845025,0.21881226,0.47157812,0.7884786,1.0525624,1.1506506,1.2562841,1.388326,1.6335466,1.8976303,1.8938577,1.7693611,1.7429527,1.81086,1.9957186,2.3428001,2.3767538,2.6446102,3.0445085,3.5764484,4.327201,4.8629136,5.353355,5.624984,5.6891184,5.7419353,5.8966126,6.1644692,6.224831,6.0324273,5.8211603,5.7872066,5.798525,6.126743,6.628502,6.7756343,1.8523588,2.071171,2.3163917,2.4861598,2.5201135,2.4031622,2.5691576,2.7351532,2.8181508,2.727608,2.372981,2.0258996,1.8561316,1.7278622,1.5958204,1.5203679,1.5580941,1.5543215,1.7052265,2.0070364,2.2748928,2.6144292,2.927557,3.2821836,3.731126,4.2894745,4.870459,5.73439,6.8246784,8.311093,10.597303,12.804289,13.7851715,14.762281,16.214743,17.912424,21.183289,24.348522,28.558771,34.6742,43.260693,51.647236,60.196003,62.787796,60.071507,59.45657,54.548386,47.35399,39.937008,32.606796,23.907125,15.147089,9.839006,7.1679873,5.80607,3.9159849,3.2633207,3.8103511,4.6629643,5.0779533,4.45547,3.440634,3.3425457,3.2142766,2.5540671,1.3053282,1.0789708,0.87902164,0.70170826,0.66020936,0.9620194,0.7582976,0.56212115,0.543258,0.6187105,0.47535074,0.543258,0.43007925,0.35839936,0.38480774,0.42630664,0.41121614,0.44894236,0.43007925,0.33953625,0.25276586,0.26031113,0.241448,0.23390275,0.211267,0.08677038,0.11317875,0.124496624,0.10940613,0.07922512,0.06790725,0.041498873,0.018863125,0.05281675,0.25276586,0.7884786,0.7394345,0.5055317,0.995973,1.7542707,0.94315624,0.9242931,1.0940613,1.0601076,0.83752275,0.845068,0.59230214,1.2034674,1.5354583,1.3091009,1.1053791,0.9620194,1.1355602,1.5731846,2.1692593,2.795515,2.8256962,3.229367,2.8294687,2.1202152,3.2670932,3.2067313,2.7200627,2.757789,3.1614597,2.686109,2.8143783,2.8256962,2.6898816,2.6597006,3.2821836,2.444661,1.991946,2.2484846,2.8521044,2.7389257,2.7841973,2.3993895,2.4672968,3.1237335,3.7575345,5.2326307,5.772116,6.515323,7.7376537,8.858124,10.453944,12.106354,12.743927,12.245941,11.457462,12.310076,14.203933,15.611122,15.543215,13.562587,10.570895,9.1825695,8.669493,8.337502,7.5075235,7.6923823,8.228095,8.062099,7.5037513,8.235641,7.183078,7.413208,7.488661,7.0246277,6.651138,7.61693,9.016574,9.88805,10.114408,10.419991,10.910432,11.083972,11.2801485,11.962994,13.728582,14.268067,14.871688,15.32063,15.686575,16.33924,16.920223,17.614386,18.150099,18.467,18.693357,19.74592,21.70391,22.77911,21.881226,18.617905,18.648085,19.304522,18.821627,17.078674,15.580941,15.509261,15.558306,15.331948,14.524607,12.932558,11.732863,11.498961,11.46878,11.461235,11.879996,15.580941,18.387774,19.927006,20.138271,19.25925,19.38752,20.258997,21.202152,21.27006,19.236614,18.199142,17.693611,17.557796,17.429527,16.731592,15.788436,15.818617,16.908905,18.885761,21.304014,20.568352,19.960958,19.538425,19.127209,18.331184,17.003222,16.433554,16.490145,16.852316,17.003222,17.493662,18.376457,19.91946,21.790682,23.069601,24.812555,25.838709,26.121656,25.680258,24.578651,22.862108,21.28515,20.096773,19.542198,19.862871,19.859098,20.33822,20.941841,21.847271,23.748674,25.325632,27.325123,29.049213,29.988596,29.818829,29.452883,28.61536,27.770292,27.32135,27.596752,28.404093,30.992115,33.01424,33.361324,32.180492,33.678223,29.094484,21.53037,14.019074,9.5183325,11.046246,9.397609,7.092535,5.1760416,3.2067313,2.704972,1.8221779,1.0751982,0.77716076,1.0525624,1.358145,1.690136,2.3503454,4.3724723,9.533423,23.809036,37.52253,40.906574,31.24488,12.879742,9.537196,9.318384,8.397863,6.2323766,5.5759397,3.0671442,1.5769572,0.68661773,0.21503963,0.23013012,0.62625575,0.6451189,0.7582976,1.2789198,2.372981,6.571913,12.434572,15.294222,13.434318,8.088508,4.851596,2.9200118,2.5691576,3.3727267,4.187614,6.6549106,12.751472,17.067356,17.41821,14.879233,11.642321,8.544995,5.73439,3.651901,2.9992368,3.712263,3.4142256,3.4217708,4.036709,4.5460134,4.432834,4.0216184,3.4330888,3.1840954,4.2102494,3.9348478,3.6896272,3.4934506,3.6368105,4.696918,5.5306683,6.7341356,6.5945487,5.4703064,5.80607,5.9607477,8.130007,9.752235,9.533423,7.435844,7.745199,16.403374,28.057013,35.489082,29.626425,18.89708,13.324911,9.854096,7.6508837,8.13378,8.356364,7.8621507,7.2472124,6.7756343,6.387054,7.1302614,5.168496,3.4066803,2.9049213,2.886058,2.6974268,2.505023,2.142851,1.4109617,0.07922512,0.02263575,0.003772625,0.00754525,0.02263575,0.041498873,0.45648763,0.27917424,0.17354076,0.3055826,0.35839936,0.13958712,0.21881226,0.34330887,0.41876137,0.5017591,0.47535074,0.38858038,0.33953625,0.34330887,0.35085413,0.35462674,0.392353,0.362172,0.29049212,0.31312788,0.32444575,0.331991,0.5357128,0.8186596,0.7922512,1.0525624,1.841041,2.8898308,3.6179473,3.1576872,3.5500402,3.7688525,3.2482302,2.4031622,2.6295197,2.8634224,3.2444575,3.7650797,4.244203,4.3422914,4.104616,3.561358,2.9652832,2.565385,2.625747,2.7917426,3.259548,3.6368105,3.9084394,4.432834,4.9232755,4.5912848,4.7346444,5.2628117,4.7044635,4.5724216,4.8855495,5.2137675,5.2967653,5.032682,4.7006907,4.7950063,5.2137675,5.6513925,5.621211,6.1229706,6.1908774,6.2135134,6.277648,6.1606965,6.8699503,7.4018903,7.484888,7.284939,7.435844,8.412953,9.861642,10.461489,10.11818,9.948412,11.219787,11.819634,12.823153,14.011529,13.8870325,14.864142,15.154634,15.086727,14.592513,13.185325,12.257258,11.872451,11.921495,12.344029,13.132507,12.479843,12.442118,12.347801,11.868678,11.00852,10.63503,12.242168,12.996693,12.351574,12.057309,10.152134,12.355347,23.812809,35.753166,25.499172,18.69713,16.127972,15.686575,15.841252,15.675257,25.706667,21.662413,14.196388,9.220296,7.8961043,10.601076,9.820143,11.080199,14.215251,13.373956,12.487389,13.29473,13.264549,12.491161,13.671993,14.302021,14.086982,12.31762,9.703192,8.401636,8.239413,8.907167,8.518587,7.6697464,9.42779,10.419991,10.736891,10.925522,10.770844,9.318384,8.699674,8.492179,8.646856,9.076936,9.669238,9.216523,8.75249,8.83926,9.405154,9.759781,9.027891,8.771353,8.552541,8.073418,7.164215,7.699928,7.7829256,8.084735,8.729855,9.310839,10.469034,10.529396,9.767326,8.710991,8.137552,8.390318,7.7678347,7.118943,6.8435416,6.8925858,6.439871,6.115425,6.2361493,6.530414,6.1305156,6.2663302,5.926794,5.956975,6.4549613,6.752999,5.3646727,4.90064,4.459243,3.8707132,3.6896272,3.9197574,3.9386206,4.0970707,4.4743333,4.8365054,4.7006907,4.3309736,4.036709,3.8820312,3.6858547,3.9612563,4.025391,4.0593443,4.1197066,4.146115,4.3875628,5.251494,5.832478,6.0739264,6.7680893,6.2097406,5.583485,5.1345425,5.1798143,6.085244,6.7680893,7.4018903,8.039464,8.578949,8.805306,9.167479,8.75249,7.8734684,7.0510364,7.0170827,6.541732,5.9192486,5.5570765,5.3571277,4.7233267,4.2517486,3.5839937,2.8407867,2.2258487,2.003264,1.8184053,1.720317,1.7278622,1.7618159,1.6750455,1.2713746,0.8639311,0.5394854,0.33953625,0.23013012,0.24522063,0.2678564,0.26408374,0.2263575,0.19994913,0.19240387,0.17731337,0.16976812,0.16976812,0.18863125,0.241448,0.3055826,0.35839936,0.42630664,0.5772116,0.69039035,0.80734175,0.8978847,0.91297525,0.7469798,0.60362,0.51684964,0.4376245,0.3734899,0.36971724,0.4376245,0.6375736,0.87147635,1.0487897,1.0601076,1.1506506,1.3015556,1.6109109,1.9693103,2.0673985,1.7655885,1.780679,1.9353566,2.1051247,2.214531,2.161714,2.474842,3.138824,3.9725742,4.6214657,4.949684,5.2779026,5.4174895,5.458988,5.783434,5.8966126,6.2323766,6.3531003,6.205968,6.085244,6.2323766,6.25124,6.3832817,6.63982,6.7944975,2.2296214,2.282438,2.4672968,2.6408374,2.6823363,2.5012503,2.6332922,2.8106055,2.8747404,2.7125173,2.2560298,1.9994912,1.841041,1.7354075,1.6637276,1.6109109,1.6788181,1.6637276,1.8448136,2.1843498,2.3503454,2.886058,3.2935016,3.6669915,4.112161,4.7572803,5.4401255,6.2323766,7.0170827,8.228095,10.819888,13.174006,14.400109,15.901614,18.104828,20.447628,24.340977,27.841972,32.5238,39.646515,50.17214,57.25713,62.9387,62.323765,55.90653,49.587383,46.184475,42.000633,35.040142,25.95566,18.03692,10.280403,6.2135134,4.4215164,3.6368105,2.7426984,2.6823363,3.1652324,3.62172,3.7348988,3.4594972,2.8898308,2.8143783,2.8181508,2.505023,1.5015048,1.0751982,0.7696155,0.5885295,0.6111652,1.0223814,0.76207024,0.5319401,0.48666862,0.60362,0.694163,0.5583485,0.4376245,0.38103512,0.392353,0.43385187,0.44894236,0.49421388,0.48666862,0.4074435,0.32821837,0.27540162,0.23390275,0.17354076,0.10186087,0.071679875,0.14335975,0.1659955,0.14713238,0.1056335,0.060362,0.056589376,0.033953626,0.041498873,0.21503963,0.7997965,0.663982,0.40367088,0.51684964,0.8563859,0.6149379,0.38103512,0.72811663,1.1657411,1.5543215,2.1164427,1.871222,1.8636768,1.6788181,1.1883769,0.55080324,0.41498876,0.65643674,1.056335,1.4750963,1.8448136,2.2786655,2.6672459,2.463524,1.8900851,1.9240388,1.7014539,1.5807298,1.9240388,2.4069347,1.9957186,2.8521044,3.2670932,3.108643,2.9351022,3.9688015,2.6710186,2.5389767,2.9766011,3.3727267,3.1161883,3.5047686,3.3236825,3.4972234,4.191386,4.8063245,6.802043,6.9567204,7.7187905,9.34102,9.903141,10.974566,11.385782,11.593277,11.774363,11.834724,11.747954,12.615658,14.354838,15.679029,14.068119,9.95973,8.843033,8.224322,7.2396674,6.651138,6.7341356,7.3415284,7.635793,7.5263867,7.6923823,6.903904,7.1566696,7.496206,7.484888,7.1981683,7.6622014,8.59404,9.163706,9.178797,9.0957985,9.552286,10.038955,10.4049,11.083972,13.094781,13.29473,13.747445,14.626467,15.592259,15.807299,16.358103,17.384256,18.206688,18.636768,18.976303,19.312067,20.274086,21.470009,21.719002,19.021576,19.221525,19.353567,18.595268,16.961721,15.279131,14.969776,15.113135,15.222542,14.939595,14.060574,12.178034,11.849815,11.819634,11.664956,11.808316,14.11339,15.950659,17.629477,18.851807,18.715992,18.893307,20.040184,21.884998,23.1941,21.78691,20.511763,19.953413,19.647831,19.255478,18.565088,17.942604,17.686066,18.168962,19.711966,22.586706,23.160145,23.375185,22.669704,21.073883,19.229069,17.746428,16.957949,16.45619,16.263786,16.825907,16.939087,17.580433,19.066847,21.09652,22.748928,24.608833,26.008476,26.34424,25.61235,24.420202,24.084438,22.620659,21.1267,20.455173,21.183289,20.904116,20.730574,20.647577,20.866388,21.851044,23.22428,25.46522,27.728794,29.237844,29.283115,28.619133,27.796701,27.151583,27.015768,27.702385,29.426476,32.893517,36.009705,37.292397,35.86257,37.763977,36.92268,31.799456,23.605314,16.293968,14.483108,12.2119875,9.725827,7.175533,4.610148,3.591539,2.2296214,1.3166461,1.0789708,1.1393328,1.448688,1.7731338,2.11267,3.180323,6.432326,21.869907,44.030308,56.540333,50.73426,25.68403,13.52486,8.993938,7.6395655,6.8435416,5.832478,3.5990841,2.0485353,0.9393836,0.24899325,0.1659955,0.21503963,0.32821837,0.98465514,2.2673476,3.863168,7.7225633,16.659912,25.54067,29.743376,25.140774,15.328176,7.888559,4.3686996,4.217795,4.8100967,7.2057137,12.30253,15.264041,14.339747,10.884023,9.0957985,7.8508325,6.741681,5.3609,3.3123648,3.482133,3.7009451,4.025391,4.315883,4.2404304,5.1760416,5.010046,4.055572,3.1312788,3.5651307,3.9876647,3.9688015,4.1989317,4.402653,3.3538637,4.0895257,5.8702044,6.1342883,4.8666863,4.6252384,4.4743333,6.7039547,8.827943,9.348565,7.748972,7.854605,12.751472,19.715738,24.910643,23.371412,15.712983,11.578186,9.099571,7.6320205,7.798016,7.4999785,7.443389,7.2887115,6.881268,6.2663302,5.379763,3.6141748,2.9124665,3.2482302,2.5880208,3.169005,2.757789,1.659955,0.46026024,0.056589376,0.026408374,0.030181,0.033953626,0.060362,0.181086,0.38103512,0.43385187,0.3772625,0.331991,0.48666862,0.24899325,0.29426476,0.38103512,0.3772625,0.28294688,0.44139713,0.38103512,0.32444575,0.32821837,0.29426476,0.35462674,0.422534,0.43007925,0.36594462,0.29049212,0.2565385,0.331991,0.59230214,0.87902164,0.7884786,0.9695646,1.5807298,2.5880208,3.5500402,3.6330378,4.214022,4.085753,3.2784111,2.3578906,2.4295704,2.7728794,3.138824,3.62172,4.104616,4.2706113,3.893349,3.4179983,2.9803739,2.686109,2.584248,2.5276587,3.1425967,3.5500402,3.6443558,4.0895257,4.719554,4.315883,4.3121104,4.9119577,5.0779533,4.6931453,4.9949555,5.2628117,5.149633,4.6856003,4.7950063,4.851596,5.010046,5.304311,5.6287565,5.5495315,5.534441,5.6325293,5.7683434,5.726845,6.48137,7.001992,7.069899,6.9869013,7.594294,8.590267,9.997457,10.95193,11.283921,11.54046,11.970539,12.298758,12.766563,13.226823,13.170234,14.807553,14.452927,14.030393,13.72481,11.996947,11.891314,11.898859,11.668729,11.615912,12.955194,11.566868,11.781908,12.261031,12.15917,11.099063,11.812089,11.827179,11.09529,10.144588,10.050273,9.778644,14.532151,22.379211,26.498919,15.188588,11.717773,16.109108,20.700394,22.228306,21.851044,25.435038,20.157135,13.50977,9.789962,10.121953,10.861387,10.235131,11.314102,13.781399,13.947394,14.203933,15.758255,16.867407,18.270823,23.156372,34.760967,35.636215,29.128437,20.255224,15.705438,14.094527,12.717519,10.808571,9.005256,9.352338,9.627739,9.993684,10.70671,11.41219,11.140562,10.065364,9.80128,9.808825,10.069136,11.083972,10.589758,9.850324,9.635284,9.880505,9.718282,9.291975,8.801534,8.375228,7.91874,7.092535,7.364164,7.7112455,7.986647,8.318638,9.103344,10.310584,10.631257,10.008774,8.922258,8.375228,8.356364,7.8206515,7.4018903,7.2094865,6.832224,6.326692,6.432326,7.062354,7.624475,7.0170827,6.598321,6.066381,6.304056,7.1340337,7.333983,5.541986,4.938366,4.4215164,3.8480775,4.014073,3.832987,3.682082,3.8141239,4.236658,4.696918,4.644101,4.4516973,4.0970707,3.7198083,3.6066296,3.6443558,3.4330888,3.2935016,3.3576362,3.5538127,3.7160356,4.6214657,5.3646727,5.715527,6.145606,5.881522,5.198677,4.7874613,5.032682,6.013564,6.6058664,7.0548086,7.413208,7.7150183,7.997965,8.514814,8.216777,7.5792036,6.9567204,6.5455046,6.228604,5.775889,5.4476705,5.20245,4.7006907,4.1612053,3.4029078,2.5314314,1.7919968,1.5580941,1.7542707,1.6788181,1.599593,1.5920477,1.5279131,1.086516,0.875249,0.67152727,0.43007925,0.26408374,0.2263575,0.23767537,0.22258487,0.17731337,0.1659955,0.17354076,0.17731337,0.18863125,0.1961765,0.17731337,0.20372175,0.29049212,0.3961256,0.52062225,0.6790725,0.83752275,0.97333723,1.0487897,1.056335,1.0148361,0.95824677,0.8601585,0.72811663,0.6187105,0.6375736,0.69039035,0.8639311,1.0827434,1.237421,1.1619685,1.1808317,1.2789198,1.569412,1.901403,1.8485862,1.5882751,1.7089992,1.9353566,2.1353056,2.3428001,2.11267,2.3428001,3.108643,4.063117,4.425289,4.715781,5.0062733,5.119452,5.20245,5.745708,6.1795597,6.6322746,6.7152724,6.4511886,6.2851934,6.2625575,6.2021956,6.2625575,6.4210076,6.477597,2.3956168,2.1843498,2.3880715,2.6219745,2.71629,2.7087448,2.8143783,2.7804246,2.595566,2.3013012,1.9693103,2.0108092,1.8674494,1.8259505,1.9051756,1.841041,1.9730829,2.052308,2.2258487,2.5012503,2.7426984,3.1425967,3.519859,3.942393,4.5233774,5.4174895,6.1229706,7.0284004,7.5792036,8.43559,11.431054,14.302021,16.358103,18.565088,21.360603,24.657877,28.690813,31.625916,35.71167,42.362804,52.164085,56.84214,59.426388,56.861004,48.885674,38.03938,35.783348,33.138737,26.419693,17.263533,12.653384,7.4207535,4.534695,3.1199608,2.493705,2.161714,1.8561316,2.214531,2.4823873,2.4333432,2.3390274,2.052308,1.8976303,2.0485353,2.2711203,1.9240388,1.1431054,0.7696155,0.573439,0.5055317,0.7130261,0.45648763,0.32067314,0.30181,0.4376245,0.84129536,0.46026024,0.44139713,0.45648763,0.41498876,0.45648763,0.4376245,0.452715,0.44516975,0.4074435,0.38480774,0.2565385,0.25276586,0.23013012,0.15845025,0.10186087,0.19240387,0.21503963,0.19240387,0.13958712,0.030181,0.049044125,0.0452715,0.030181,0.124496624,0.5319401,0.40367088,0.18863125,0.08677038,0.15845025,0.32067314,0.32821837,0.98465514,2.1654868,3.3840446,3.8178966,3.4896781,2.0447628,0.9205205,0.6375736,0.7507524,0.43007925,0.41876137,0.47157812,0.49421388,0.55080324,0.5357128,1.0186088,1.4977322,1.478869,0.44139713,0.30181,0.46026024,1.0223814,1.6561824,1.599593,3.2067313,3.3953626,3.127506,3.138824,3.9273026,3.3010468,3.4557245,3.640583,3.591539,3.5500402,4.5460134,4.395108,4.659192,5.617439,6.277648,8.001738,8.062099,9.065618,11.034928,11.404645,11.212241,10.499215,10.438853,11.491416,13.400364,12.1252165,12.064855,13.826671,15.671484,13.498452,10.11818,8.918486,7.8734684,6.620957,6.4474163,6.688864,7.492433,7.8206515,7.5112963,7.284939,6.990674,7.333983,7.835742,8.182823,8.231868,7.9941926,8.299775,8.722309,8.89585,8.507269,8.514814,9.076936,9.7069645,10.555805,12.385528,12.234623,12.31762,13.853079,15.931795,15.543215,16.120426,16.720274,17.048492,17.278622,18.029375,18.45568,18.931032,19.059301,18.863125,18.814081,19.723284,19.051756,17.833199,16.535416,15.033911,14.520834,14.369928,14.607604,14.992412,15.007503,13.102326,12.73261,12.626976,12.423254,12.649611,13.6833105,14.532151,15.501716,16.335466,16.237377,16.84477,18.48209,21.062565,23.352549,22.960196,21.669958,20.832436,20.111864,19.447882,19.04421,18.840488,18.48209,18.648085,19.60256,21.187061,23.378958,25.031366,24.699375,22.4773,20.010002,18.62545,17.87847,17.074902,16.471281,17.301258,17.086218,17.308804,18.41041,20.277859,22.26226,23.36764,24.786146,25.499172,25.272816,24.684286,24.578651,23.126192,21.798227,21.447372,22.296213,21.190834,20.398582,20.070366,20.025093,19.742147,20.877707,22.613113,25.054003,27.423212,28.05324,26.985586,26.182018,25.789665,26.004704,27.094994,29.5472,33.036877,36.817047,39.544655,39.295662,38.60527,41.385696,42.381668,39.159847,32.127674,21.35683,16.592005,12.875969,8.699674,6.013564,4.561104,2.8936033,1.871222,1.5731846,1.2864652,1.6184561,2.0108092,2.2711203,2.674791,3.9348478,15.01882,38.89199,59.0944,63.602684,44.837646,21.847271,9.608876,5.6325293,6.3342376,7.073672,5.3873086,3.059599,1.2185578,0.33576363,0.2263575,0.41876137,0.46026024,1.4411428,3.2784111,4.727099,7.111398,14.252977,26.66114,39.73706,43.769997,32.976517,19.715738,10.020092,6.25124,7.0887623,10.63503,13.456953,12.800517,9.092027,5.9003854,8.009283,7.7338815,6.7077274,5.2779026,2.5012503,2.505023,2.8936033,3.482133,4.323428,5.6815734,7.3453007,7.224577,5.80607,4.0782075,3.5047686,4.266839,4.1536603,4.564876,5.138315,3.7273536,3.9348478,4.930821,5.1043615,4.406426,4.3686996,3.6783094,5.5495315,7.7414265,8.6732645,7.3905725,7.8961043,10.944386,14.362384,15.807299,12.808062,9.710737,8.360137,7.250985,6.0211096,5.4401255,6.7680893,7.284939,7.7112455,7.835742,6.511551,3.0520537,2.5880208,2.886058,2.938875,2.9652832,4.357382,3.5689032,1.7052265,0.03772625,0.0,0.018863125,0.05281675,0.06413463,0.124496624,0.3961256,0.3734899,0.65643674,0.5357128,0.17354076,0.58475685,0.4640329,0.33576363,0.31312788,0.3470815,0.21503963,0.31312788,0.39989826,0.38103512,0.27917424,0.241448,0.43007925,0.5017591,0.49421388,0.4376245,0.35462674,0.23013012,0.362172,0.6752999,0.95824677,0.84884065,0.8941121,1.4977322,2.3126192,3.1576872,4.014073,4.851596,4.395108,3.31991,2.3277097,2.1466236,2.5201135,3.059599,3.4972234,3.783943,4.0970707,3.6745367,3.2142766,2.9501927,2.8822856,2.795515,2.4786146,2.8445592,3.1539145,3.259548,3.5877664,4.4101987,4.1272516,3.8443048,4.085753,4.798779,4.432834,4.7572803,4.98741,4.821415,4.4516973,4.870459,5.0025005,4.8742313,4.7874613,5.311856,4.9459114,4.8063245,4.768598,4.7648253,4.798779,5.66271,6.519096,6.9227667,7.1906233,8.397863,9.22784,9.88805,10.921749,12.276122,13.283413,12.917468,13.230596,13.415455,13.189097,12.785426,14.18507,13.690856,13.196642,12.691111,10.250222,11.148107,11.623458,11.072655,10.412445,12.098808,10.819888,11.219787,12.2119875,12.917468,12.626976,13.290957,12.306303,10.816116,9.87296,10.435081,12.626976,16.954176,19.40261,17.501207,10.325675,10.020092,19.862871,28.377686,30.39604,27.061039,17.591751,10.220041,7.5829763,9.25425,11.740409,11.472552,11.415963,11.627231,12.347801,14.02662,15.792209,18.18028,21.21347,25.533127,32.384212,57.151497,59.19626,47.765205,32.486073,23.356321,19.930779,16.818363,14.022847,11.6875925,10.076681,9.684328,9.861642,10.823661,12.079946,12.423254,11.506506,11.144334,10.646348,10.223814,10.970794,11.072655,10.536942,10.174769,10.061591,9.540969,9.540969,8.812852,8.348819,8.254503,7.756517,7.6395655,8.375228,8.541223,8.156415,8.695901,9.567377,9.940866,9.771099,9.329701,9.186342,8.488406,8.031919,7.8508325,7.665974,6.8737226,6.5568223,6.8473144,7.488661,7.956466,7.4509344,6.7944975,6.1795597,6.0211096,6.3153744,6.628502,5.2552667,4.859141,4.406426,3.9273026,4.5007415,4.1762958,3.8405323,3.832987,4.2064767,4.7308717,4.6554193,4.376245,3.9914372,3.6368105,3.4934506,3.3048196,2.9728284,2.7841973,2.8294687,3.0143273,3.0897799,3.7009451,4.4818783,5.1081343,5.2779026,5.3080835,4.647874,4.4139714,5.0138187,6.1720147,6.537959,6.779407,7.020855,7.2660756,7.4018903,7.7602897,7.5716586,7.3188925,7.073672,6.4964604,6.168242,5.726845,5.270357,4.870459,4.5761943,4.2781568,3.5990841,2.6597006,1.780679,1.4901869,1.7882242,1.6675003,1.5165952,1.4750963,1.448688,1.0374719,0.9242931,0.754525,0.47535074,0.31312788,0.24522063,0.241448,0.23013012,0.18863125,0.15467763,0.18485862,0.20372175,0.2263575,0.23767537,0.1659955,0.20749438,0.36594462,0.56589377,0.72811663,0.7582976,0.8639311,1.0072908,1.0450171,0.9922004,1.0450171,1.0714256,1.0223814,0.9280658,0.86770374,0.9620194,0.97333723,1.0714256,1.2638294,1.4335974,1.327964,1.2562841,1.2638294,1.4750963,1.6863633,1.3694628,1.327964,1.4939595,1.7240896,2.0108092,2.5012503,2.1654868,2.263575,3.0143273,4.025391,4.285702,4.568649,4.859141,5.0477724,5.2628117,5.8626595,6.6624556,7.1076255,7.0472636,6.620957,6.270103,5.9305663,5.8136153,5.907931,6.0324273,5.8626595,2.2107582,2.1768045,2.3126192,2.3126192,2.2220762,2.4408884,2.674791,2.5314314,2.323937,2.1390784,1.8448136,1.8221779,1.8448136,2.0258996,2.2673476,2.2447119,2.463524,2.6106565,2.897376,3.3048196,3.5839937,3.682082,3.7990334,4.22534,4.9760923,5.783434,6.4436436,7.997965,9.224068,10.442626,13.517315,17.425755,19.493153,21.322876,23.692085,26.551735,29.920689,30.94307,33.74613,38.835403,43.106014,51.213383,57.211857,56.7101,48.768723,35.90407,30.618624,23.922215,15.860115,9.563604,11.261286,6.3417826,4.032936,2.8709676,2.233394,2.3201644,2.0749438,2.052308,2.033445,1.901403,1.6335466,1.50905,1.6524098,2.1843498,2.8521044,3.0218725,2.3013012,1.0487897,0.27540162,0.2263575,0.3961256,0.33576363,0.32821837,0.3169005,0.34330887,0.55080324,0.40367088,0.59607476,0.6488915,0.5017591,0.5017591,0.41876137,0.27917424,0.18485862,0.21503963,0.3961256,0.3470815,0.4640329,0.42630664,0.22258487,0.1358145,0.26031113,0.35462674,0.27540162,0.090543,0.090543,0.090543,0.071679875,0.056589376,0.06790725,0.150905,0.19994913,0.1056335,0.056589376,0.1358145,0.32067314,0.26031113,0.33576363,1.3241913,2.4031622,1.1431054,1.6561824,0.8865669,0.362172,0.543258,0.8224323,0.49421388,0.422534,0.4074435,0.392353,0.42630664,0.41498876,0.41121614,0.3772625,0.30935526,0.26031113,0.331991,0.88279426,1.3958713,1.3656902,0.3055826,1.599593,2.323937,3.289729,4.146115,3.4029078,2.474842,2.5087957,3.1312788,4.036709,4.991183,5.5759397,4.979865,4.7308717,5.5570765,7.4018903,8.36391,8.322411,8.744945,10.072908,11.732863,10.684074,10.521852,10.484125,11.068882,14.022847,12.5326605,13.917213,14.064346,12.045992,10.11818,11.091517,9.733373,8.397863,7.888559,7.462252,7.3377557,7.2924843,7.541477,7.786698,7.1868505,7.8206515,8.741172,8.948667,8.601585,9.001483,9.175024,8.914713,8.560086,8.299775,8.179051,9.144843,9.35611,9.880505,10.627484,10.344538,10.808571,11.144334,12.464753,14.347293,14.84528,14.554788,14.637785,14.849052,15.23386,16.11288,17.357847,19.123436,19.338476,18.240643,18.387774,19.47429,19.270569,17.969013,16.180788,14.924504,14.362384,13.600313,13.788944,14.86037,15.531898,14.886778,14.4152,13.728582,12.97783,12.83447,13.758763,14.339747,15.098045,15.958203,16.252468,16.203424,17.13149,19.006485,21.077656,21.896315,20.590988,18.889534,17.53516,17.082445,17.897333,17.312576,17.13149,18.184053,19.968504,20.613623,21.809546,24.152346,25.269043,24.34475,22.111355,19.180025,18.53868,18.350048,18.055782,18.387774,18.191597,17.886015,18.28214,19.542198,21.164427,22.57916,23.639269,24.31834,24.842735,25.695349,24.646559,23.103556,22.228306,22.24717,22.432028,20.70794,19.930779,19.734602,19.557287,18.629223,18.791445,19.572378,21.409647,23.948624,26.061293,25.02382,24.582424,24.827644,25.450129,25.74062,28.26828,31.24488,35.564537,39.82383,40.29918,35.33063,39.042896,47.8482,58.030518,65.730446,38.925945,23.08092,14.260523,9.567377,7.1264887,5.8702044,3.9688015,2.546522,1.9089483,1.5430037,1.7844516,2.5502944,2.625747,2.323937,3.4934506,9.367428,23.89958,41.600735,55.751854,58.426643,33.74236,14.434063,4.961002,4.436607,6.620957,7.707473,4.1989317,1.2449663,0.56589377,0.45648763,1.5203679,1.1996948,1.6561824,2.9313297,2.9464202,3.8858037,7.0585814,15.977067,29.8641,43.671906,52.862022,43.238056,25.616123,10.676529,8.956212,12.095036,12.943876,11.800771,10.499215,12.404391,15.335721,12.717519,7.858378,3.5387223,1.9994912,3.8405323,3.5877664,3.289729,4.032936,5.9494295,8.356364,8.83926,8.152642,6.752999,4.776143,5.070408,5.040227,4.2781568,3.361409,3.8593953,4.9459114,4.678055,4.561104,5.0138187,5.3571277,3.4745877,4.82896,6.4511886,6.9755836,6.620957,7.4773426,9.831461,12.47607,13.505998,10.329447,6.6058664,5.3646727,5.855114,6.8435416,6.6360474,5.613666,4.293247,4.5460134,5.2326307,2.2296214,1.9730829,2.4031622,1.9127209,0.8299775,1.4034165,3.5764484,2.1692593,0.5696664,0.09808825,0.0,0.0,0.0,0.060362,0.17731337,0.27540162,0.5055317,0.7092535,0.62625575,0.35462674,0.36594462,0.29426476,0.36594462,0.43385187,0.45648763,0.52062225,0.47157812,0.8224323,0.7507524,0.25276586,0.1659955,0.52062225,0.47157812,0.33953625,0.3055826,0.42630664,0.29426476,0.34330887,0.62248313,0.995973,1.1280149,1.3128735,2.0372176,2.9615107,3.8065786,4.3196554,4.991183,4.508287,3.6481283,2.8407867,2.1805773,2.4522061,2.9841464,3.289729,3.399135,3.874486,3.4745877,3.410453,3.3312278,3.1124156,2.867195,2.3692086,2.6182017,3.169005,3.6141748,3.6028569,4.6252384,4.606375,4.2404304,4.002755,4.1498876,4.2706113,4.5950575,5.0854983,5.4174895,4.991183,5.0741806,4.7950063,4.255521,4.0178456,5.0666356,4.908185,5.0213637,4.82896,4.3686996,4.3347464,5.247721,6.587003,7.5075235,7.8017883,7.8734684,9.0957985,9.1976595,10.197406,12.027128,12.528888,14.015302,14.362384,13.822898,13.234368,13.992666,14.407655,13.000465,11.853588,11.336739,10.11818,11.031156,10.691619,9.861642,9.488152,10.695392,10.208723,11.185833,12.253486,13.505998,16.509007,14.603831,12.985375,12.049765,12.242168,14.022847,19.859098,23.816582,24.363613,20.564579,12.068627,12.887287,21.23988,26.049976,23.23937,15.731846,9.065618,8.043237,8.650629,9.567377,12.128989,12.642066,13.12119,11.140562,8.397863,10.680302,15.905387,19.538425,22.673477,25.92548,29.40384,48.168877,52.590393,44.200073,29.139755,18.202915,14.70192,13.936077,12.543978,10.359629,10.4049,10.978339,11.434827,12.223305,12.936331,12.313848,12.864652,12.396846,11.744182,11.155652,10.299266,10.702937,10.235131,9.7220545,9.552286,9.673011,9.820143,9.2995205,8.809079,8.465771,7.7829256,7.33021,8.088508,8.567632,8.341274,8.009283,7.8395147,8.89585,9.95973,10.442626,10.4049,9.857869,8.922258,8.288457,8.190369,8.424272,7.677292,7.3905725,7.281166,6.9755836,6.013564,6.670001,6.560595,6.1229706,5.798525,6.043745,4.7006907,4.1272516,3.8443048,3.9273026,4.991183,5.0741806,4.3007927,3.8254418,4.0480266,4.606375,4.4743333,3.7348988,3.2482302,3.2520027,3.3727267,3.006782,2.776652,2.5880208,2.4522061,2.5012503,2.5767028,3.218049,3.9386206,4.447925,4.67051,4.6214657,4.6818275,4.7421894,4.9157305,5.5382137,6.477597,6.9152217,7.194396,7.3868,7.277394,7.5603404,7.3000293,6.8171334,6.398372,6.300284,5.485397,5.05909,4.927048,4.878004,4.6252384,3.8178966,3.1312788,2.3390274,1.659955,1.7693611,1.9542197,1.6033657,1.4034165,1.4750963,1.388326,1.0336993,0.8563859,0.6526641,0.44516975,0.45648763,0.3734899,0.3772625,0.38480774,0.35085413,0.29049212,0.29049212,0.23390275,0.18485862,0.1659955,0.1659955,0.32821837,0.5772116,0.79602385,0.88279426,0.7469798,0.784706,0.8299775,0.83752275,0.814887,0.83752275,0.8639311,0.9997456,1.1619685,1.3505998,1.6335466,1.5958204,1.5128226,1.4524606,1.4147344,1.327964,1.3166461,1.3317367,1.4109617,1.5165952,1.5430037,1.5165952,1.418507,1.5656394,1.9504471,2.2447119,1.9994912,2.0673985,2.9615107,4.38379,5.1873593,5.247721,5.4740787,5.485397,5.3269467,5.4476705,6.0814714,6.3342376,6.4436436,6.5228686,6.560595,6.719045,6.6134114,6.217286,5.617439,5.0213637,1.991946,1.9164935,1.9730829,1.991946,2.0296721,2.3692086,2.8634224,2.8143783,2.6634734,2.5578396,2.372981,2.082489,2.0749438,2.0862615,2.0183544,1.9240388,2.2220762,2.4408884,2.7502437,3.2067313,3.7198083,3.7009451,3.7499893,4.1272516,4.7610526,5.2326307,6.19465,7.907422,9.691874,11.680047,14.811326,17.244669,18.606586,19.859098,21.405874,23.058285,26.019794,26.83091,30.101774,35.809757,39.310753,42.649525,47.233265,45.018734,34.964687,23.028103,19.57615,15.275358,10.521852,6.9944468,7.647111,5.511805,4.08198,3.361409,2.9539654,2.0636258,2.1692593,2.0787163,1.9844007,1.8448136,1.3996439,1.5618668,1.7014539,1.9994912,2.3692086,2.4710693,1.8485862,0.995973,0.513077,0.52439487,0.6790725,0.56589377,0.543258,0.5093044,0.4640329,0.47535074,0.42630664,0.513077,0.59230214,0.58475685,0.4678055,0.392353,0.35462674,0.44894236,0.573439,0.44516975,0.63002837,0.84884065,0.7054809,0.29049212,0.17354076,0.2867195,0.29049212,0.22258487,0.12826926,0.07922512,0.06790725,0.1659955,0.1659955,0.06413463,0.041498873,0.08299775,0.056589376,0.041498873,0.0754525,0.150905,0.15845025,0.15467763,0.32821837,0.5696664,0.47157812,0.7922512,0.73566186,0.73566186,0.8299775,0.6526641,0.47157812,0.482896,0.58475685,0.70170826,0.80734175,0.9205205,0.8262049,0.68661773,0.58475685,0.51684964,0.49044126,0.5093044,0.663982,0.84884065,0.7809334,1.6561824,1.9693103,2.5389767,2.987919,1.7542707,1.9994912,2.2220762,2.5729303,3.0407357,3.4632697,3.6707642,4.4931965,5.221313,5.983383,7.7678347,9.435335,9.14107,9.088254,10.035183,11.295239,9.669238,9.597558,10.287949,11.189606,11.98563,12.359119,13.290957,13.747445,13.479589,12.996693,15.252723,14.611377,12.668475,10.853842,10.427535,9.359882,8.677037,8.473316,8.416726,7.7602897,7.907422,8.533678,9.005256,9.0807085,8.918486,9.382519,9.612649,9.2844305,8.616675,8.386545,9.163706,9.318384,9.42779,9.661693,9.771099,10.967021,12.019584,12.755245,13.181552,13.517315,13.781399,14.535924,14.671739,14.362384,15.07541,16.70141,17.912424,18.03692,17.523844,17.923742,19.11589,19.84778,19.274342,17.550251,15.814844,15.358356,14.713238,14.64533,14.962231,14.471789,14.2944765,14.539697,14.566105,13.996439,12.698656,12.96274,13.479589,13.913441,14.11339,14.102073,14.796235,15.546988,17.078674,19.081938,20.213724,19.998686,18.402864,16.592005,15.860115,17.655886,18.629223,18.399092,18.376457,18.991394,19.685556,20.756983,22.243397,23.26955,23.360094,22.46221,20.06282,19.010258,18.591496,18.342503,18.055782,18.49718,18.568861,19.063074,20.33822,22.322622,23.458181,23.616632,24.133482,25.144547,25.597261,24.363613,23.107328,23.069601,23.790173,23.114874,19.662922,18.357594,18.085964,18.048239,17.765291,18.38023,19.425245,20.455173,21.473782,22.911152,23.212961,23.265778,24.163664,25.661396,26.166927,28.090965,30.39604,32.17672,33.146282,33.632954,31.459919,33.27455,40.608536,50.15328,53.786316,37.662117,25.401085,17.150352,11.940358,7.6622014,5.8211603,4.3309736,3.1237335,2.2069857,1.6750455,1.8334957,2.335255,2.3126192,2.1277604,3.3463185,8.016829,17.818108,29.505701,40.800938,50.406044,36.983044,19.610106,7.964011,4.817642,6.0362,6.205968,3.7688525,1.6448646,0.845068,0.482896,1.0450171,0.90920264,0.84884065,1.0978339,1.3355093,1.2487389,3.1539145,8.869441,18.433046,30.120638,35.79844,32.180492,21.470009,9.507015,5.794752,6.3153744,8.993938,11.038701,12.268577,15.0905,16.388283,13.585222,9.144843,5.1345425,3.2067313,4.7572803,4.738417,4.557331,4.779916,5.1345425,6.8171334,7.914967,7.356619,5.670255,4.9723196,5.3609,4.881777,4.3724723,4.044254,3.470815,3.9122121,4.2064767,4.6856003,5.1571784,4.8930945,4.115934,3.7801702,5.485397,8.488406,9.699419,7.54525,9.608876,11.080199,10.231359,8.412953,6.828451,5.0251365,4.6629643,5.8966126,7.3717093,5.4363527,4.168751,3.380272,3.2067313,4.1197066,4.1574326,3.7462165,2.867195,2.203213,3.138824,3.240685,1.8146327,0.5696664,0.12826926,0.0,0.0,0.0,0.17731337,0.41498876,0.29803738,0.29803738,0.4074435,0.422534,0.3169005,0.23013012,0.46026024,0.49421388,0.58098423,0.70170826,0.56589377,0.43007925,0.5583485,0.5470306,0.33576363,0.19240387,0.331991,0.362172,0.32444575,0.27917424,0.29426476,0.2263575,0.32067314,0.66020936,1.1431054,1.4826416,1.3355093,2.0108092,2.795515,3.5047686,4.478106,4.9232755,4.4215164,3.6254926,2.9086938,2.3654358,2.4484336,3.3312278,3.7499893,3.531177,3.6066296,3.127506,3.1463692,3.270866,3.1840954,2.637065,2.3993895,2.263575,2.4899325,3.0671442,3.712263,3.6443558,3.942393,4.0216184,3.9763467,4.5912848,4.447925,4.640329,5.028909,5.330719,5.0854983,5.0175915,5.1647234,5.010046,4.5950575,4.5422406,4.4818783,4.817642,4.7006907,4.3422914,5.0175915,5.3382645,6.0248823,6.700182,7.1378064,7.2887115,8.45068,9.1976595,9.857869,10.253995,9.718282,12.283667,14.735873,15.282904,14.147344,13.577678,13.6682205,12.755245,11.642321,10.748209,10.091772,10.842525,10.438853,9.986138,9.846551,9.65792,9.473062,11.234878,11.932813,12.098808,15.814844,15.999702,13.928532,11.989402,11.529142,12.849561,20.19109,34.659107,34.91942,20.489126,11.729091,13.630494,18.040693,19.032892,15.158407,9.457971,6.541732,5.745708,8.624221,12.645839,11.16697,9.835234,10.069136,10.0276375,9.650374,10.646348,12.736382,14.139798,15.596032,17.278622,18.7839,22.499935,23.322369,20.949387,16.592005,12.97783,11.5857315,11.740409,11.249968,10.080454,10.382264,10.114408,10.49167,11.193378,11.876224,12.193124,12.789199,13.573905,14.053028,13.656902,11.729091,11.759273,11.706455,11.102836,10.163452,9.748463,9.680555,9.914458,9.869187,9.242931,8.050782,7.5490227,7.4018903,7.726336,8.405409,9.073163,8.288457,8.850578,9.710737,10.246449,10.310584,10.823661,10.770844,10.393582,10.054046,10.216269,8.729855,8.22055,8.341274,8.412953,7.4282985,7.4999785,7.8508325,7.515069,6.6813188,6.700182,5.6325293,4.459243,3.8103511,3.8443048,4.2819295,5.040227,4.9044123,4.515832,4.327201,4.5950575,4.4818783,3.6141748,3.0143273,2.987919,3.138824,2.6068838,2.5201135,2.4484336,2.3013012,2.3314822,2.474842,3.1765501,3.7235808,3.8895764,3.9122121,3.8254418,4.2328854,4.6856003,5.13077,5.9305663,6.2851934,6.3531003,6.519096,6.907676,7.413208,7.1264887,6.228604,5.5457587,5.3194013,5.20245,4.647874,4.6290107,4.678055,4.534695,4.123479,3.4745877,2.6483827,2.0485353,1.81086,1.8297231,1.5958204,1.4562333,1.388326,1.2864652,0.98465514,0.7696155,0.6375736,0.4979865,0.3772625,0.4074435,0.392353,0.43007925,0.43007925,0.3961256,0.422534,0.422534,0.52439487,0.56212115,0.5055317,0.44894236,0.7054809,0.8111144,0.8111144,0.76584285,0.7582976,0.76584285,0.724344,0.70170826,0.7205714,0.76584285,0.95824677,1.2713746,1.4373702,1.4034165,1.3505998,1.5015048,1.6976813,1.8636768,1.9051756,1.7429527,1.7316349,1.6486372,1.5920477,1.6524098,1.9202662,1.690136,1.539231,1.7089992,2.0636258,2.1315331,1.8297231,1.9768555,2.625747,3.5575855,4.285702,4.9987283,5.5004873,5.5495315,5.270357,5.13077,5.666483,5.907931,6.1720147,6.511551,6.6850915,6.6058664,6.719045,6.6020937,6.1644692,5.6551647,1.9391292,1.8372684,1.9504471,2.2069857,2.535204,2.8822856,3.2142766,3.1840954,3.0445085,2.9011486,2.7125173,2.565385,2.3314822,2.1466236,2.0900342,2.1843498,2.3993895,2.4484336,2.7389257,3.308592,3.8443048,3.8103511,3.8593953,4.195159,4.715781,5.0062733,6.1833324,7.798016,9.95973,12.525115,15.116908,16.135517,17.335213,18.549997,19.651604,20.564579,23.62795,25.574625,30.358313,37.281082,41.01598,41.759186,47.335125,44.12085,30.422447,16.475054,14.275613,12.528888,9.97482,7.3000293,7.1566696,5.4174895,4.172523,3.4783602,3.1124156,2.584248,2.6031113,2.0145817,1.5241405,1.4147344,1.5241405,1.2902378,1.6524098,2.161714,2.372981,1.8485862,1.2223305,0.73566186,0.5319401,0.5696664,0.6187105,0.55457586,0.5772116,0.58098423,0.5281675,0.44894236,0.4376245,0.49044126,0.5319401,0.52439487,0.4678055,0.46026024,0.5055317,0.6526641,0.784706,0.6149379,0.95824677,1.0751982,0.784706,0.29049212,0.18485862,0.33576363,0.30935526,0.21503963,0.13204187,0.094315626,0.06790725,0.14713238,0.150905,0.0754525,0.071679875,0.07922512,0.08299775,0.071679875,0.05281675,0.05281675,0.0754525,0.056589376,0.033953626,0.05281675,0.13204187,0.24522063,0.32444575,0.4074435,0.4640329,0.392353,0.38480774,0.48666862,0.7582976,1.0638802,1.0940613,1.5543215,1.4373702,1.2223305,1.0940613,0.95447415,0.8639311,0.87147635,1.1204696,1.4750963,1.5128226,2.8747404,2.7087448,2.6672459,2.9916916,2.4786146,2.5691576,2.6295197,3.0105548,3.7348988,4.5196047,4.636556,5.8588867,6.6813188,6.9454026,7.8206515,8.507269,8.341274,8.6732645,10.095545,12.457208,10.26154,9.012801,8.926031,9.7296,10.650121,12.253486,13.494679,15.256495,17.248442,18.02183,18.127462,17.006994,14.641558,12.1101265,11.608367,9.416472,8.0206,7.605612,7.748972,7.435844,7.4169807,8.09228,8.6732645,9.009028,9.590013,9.529651,10.0276375,9.952185,9.26934,9.088254,9.133525,9.250477,9.442881,9.774872,10.370946,11.925267,13.030646,13.721037,14.139798,14.566105,14.596286,14.883006,14.483108,13.713491,14.158662,15.784663,16.418465,16.592005,16.961721,18.319866,20.23636,21.605824,21.028612,18.881989,17.320122,16.365646,15.924251,15.852571,15.580941,14.132254,13.985121,14.230342,14.667966,14.973549,14.7321005,14.671739,14.445381,14.358611,14.358611,14.030393,14.136025,14.7321005,16.203424,18.248188,19.908142,20.477808,19.455427,17.784155,16.625957,17.391802,19.99114,20.040184,19.1423,18.602814,19.47429,20.817345,22.586706,24.148573,24.95214,24.529608,21.496418,19.553514,18.346275,17.659658,17.425755,18.191597,18.848034,20.032639,22.050993,24.865372,25.736847,25.548216,25.340723,25.650078,26.525326,25.333178,24.250433,24.182526,24.92196,25.15209,21.353058,18.795218,17.769064,17.844517,17.912424,18.968758,19.798737,20.142044,20.289177,21.081429,21.74541,22.062311,23.488363,25.691576,26.521553,29.39252,31.4901,32.172947,31.599506,30.73935,30.346996,31.773048,36.658596,42.883427,44.56979,34.576107,25.876434,18.840488,13.5663595,9.891823,7.6320205,5.7909794,4.221567,2.9200118,2.003264,1.8146327,2.0598533,2.191895,2.3390274,3.3010468,6.9454026,14.037937,22.100037,29.811283,37.02077,32.976517,20.764528,10.702937,6.8473144,6.9982195,7.756517,5.455216,2.7841973,1.1544232,0.69793564,0.8601585,0.72811663,0.52439487,0.47535074,0.77338815,0.9393836,1.7429527,4.9345937,10.910432,18.704676,20.025093,17.225805,11.740409,6.379509,5.3156285,8.197914,12.027128,13.113645,11.691365,11.910177,13.355092,12.185578,9.608876,6.7152724,4.4705606,6.432326,6.587003,5.8400235,5.0779533,5.1647234,5.4174895,5.9003854,5.2364035,3.8971217,4.214022,4.9949555,4.8138695,4.195159,3.6028569,3.4179983,2.8181508,3.029418,3.7084904,4.3800178,4.45547,4.8138695,5.100589,5.934339,7.424526,9.175024,7.0246277,9.190115,9.510788,7.3453007,7.5603404,6.692637,7.488661,6.771862,4.8025517,5.27413,4.5988297,4.447925,3.6971724,2.8256962,3.8971217,4.45547,4.1197066,3.31991,2.8785129,3.9914372,3.4368613,1.6146835,0.3734899,0.15467763,0.0,0.0,0.0,0.13958712,0.3961256,0.5998474,0.3169005,0.32067314,0.27540162,0.124496624,0.07922512,0.3169005,0.38858038,0.58475685,0.8903395,0.9922004,0.6413463,0.6488915,0.6488915,0.482896,0.19994913,0.211267,0.24522063,0.2678564,0.26408374,0.26031113,0.2263575,0.362172,0.66020936,1.1091517,1.7278622,1.6335466,2.0485353,2.7691069,3.6669915,4.67051,4.9459114,4.45547,3.712263,3.0256453,2.4823873,2.565385,3.4255435,3.9386206,3.8254418,3.6330378,2.9766011,3.006782,3.308592,3.3727267,2.595566,2.4484336,2.0862615,2.1051247,2.71629,3.7462165,4.187614,4.327201,4.255521,4.244203,4.7346444,4.8440504,4.7572803,4.798779,4.8742313,4.4894238,4.927048,5.0741806,5.010046,4.7950063,4.4630156,4.5761943,4.7535076,4.504514,4.274384,5.4438977,5.1534057,5.3759904,5.764571,6.330465,7.424526,8.98262,9.352338,9.5183325,9.612649,8.907167,10.33322,13.038192,14.618922,14.4152,13.50977,12.408164,11.529142,11.016065,10.691619,10.069136,10.242677,10.163452,10.023865,9.8239155,9.344792,10.3634,11.615912,11.593277,11.076427,13.140053,14.324657,13.358865,11.117926,9.714509,12.47607,21.371922,31.384468,30.614851,19.708193,11.861133,14.996184,18.357594,17.448391,12.249713,7.2660756,4.708236,4.878004,7.624475,11.351829,13.011784,10.838752,10.329447,10.114408,9.857869,10.250222,11.170743,11.299012,11.431054,11.864905,12.404391,12.879742,13.671993,13.909668,13.445636,12.872196,12.540206,12.279895,11.6008215,10.846297,11.219787,10.638803,10.729345,11.072655,11.378237,11.476325,12.238396,12.770335,13.215506,13.20796,11.838497,11.710228,11.080199,10.49167,10.291721,10.597303,10.382264,10.93684,10.978339,10.140816,9.005256,8.99771,8.035691,7.5565677,8.152642,9.559832,9.378746,9.831461,10.11818,9.948412,9.544742,10.684074,11.189606,10.850069,10.272858,10.868933,9.650374,9.318384,9.627739,10.057818,9.831461,8.314865,8.329956,8.269594,7.696155,7.3151197,5.983383,4.8327327,4.1612053,4.093298,4.5724216,5.2364035,5.1798143,4.8440504,4.534695,4.429062,4.164978,3.2746384,2.6483827,2.6031113,2.8709676,2.3918443,2.2447119,2.2258487,2.2447119,2.3088465,2.4371157,2.969056,3.3123648,3.3274553,3.3463185,3.5349495,4.1612053,4.8025517,5.372218,6.092789,6.247467,6.2889657,6.379509,6.677546,7.3377557,6.858632,5.5570765,4.587512,4.3385186,4.406426,4.044254,4.0782075,4.044254,3.863168,3.8405323,3.4896781,2.7615614,2.1466236,1.8259505,1.6637276,1.3807807,1.3204187,1.2600567,1.1016065,0.8563859,0.77716076,0.62248313,0.5017591,0.44516975,0.41498876,0.4678055,0.46026024,0.44139713,0.4979865,0.7582976,0.7469798,0.69793564,0.6752999,0.7054809,0.784706,0.814887,0.8639311,0.84884065,0.79602385,0.83752275,0.7997965,0.7054809,0.67152727,0.73188925,0.83752275,1.0336993,1.2487389,1.418507,1.4864142,1.4109617,1.7278622,1.8863125,1.8900851,1.8259505,1.8561316,1.7844516,1.6825907,1.6712729,1.7919968,2.003264,1.81086,1.7769064,1.9051756,2.071171,2.033445,1.8900851,2.1579416,2.584248,3.0897799,3.7462165,4.779916,5.572167,5.7004366,5.342037,5.2892203,5.4438977,5.7079816,6.115425,6.673774,7.364164,7.149124,6.9567204,6.6322746,6.1644692,5.6778007,2.0183544,2.04099,2.2975287,2.71629,3.1539145,3.4255435,3.4029078,3.31991,3.2331395,3.108643,2.8521044,2.8596497,2.5917933,2.4408884,2.5125682,2.637065,2.7426984,2.7804246,2.9351022,3.2444575,3.6254926,3.6481283,3.8895764,4.29702,4.7836885,5.2175403,6.270103,7.6848373,9.963503,12.766563,14.909414,15.286676,16.173243,17.056038,17.87847,19.032892,22.609343,25.291677,30.313042,36.771774,39.623882,38.627907,47.16536,45.313,29.894281,14.50197,12.325166,11.46878,9.786189,7.364164,6.4964604,4.538468,3.5651307,3.1576872,3.0181,2.969056,2.806833,1.9768555,1.4411428,1.5279131,1.9051756,1.569412,1.7354075,1.9881734,1.961765,1.3317367,0.8299775,0.7582976,0.9205205,1.2713746,1.931584,1.2185578,0.9507015,0.8299775,0.7167987,0.62625575,0.58098423,0.5055317,0.45648763,0.4640329,0.5357128,0.52062225,0.51684964,0.5998474,0.7092535,0.63002837,1.0223814,1.0412445,0.7130261,0.2867195,0.21881226,0.34330887,0.32444575,0.23390275,0.13958712,0.1056335,0.071679875,0.08677038,0.08299775,0.06413463,0.11317875,0.1358145,0.17354076,0.13958712,0.049044125,0.033953626,0.056589376,0.06413463,0.08677038,0.13958712,0.22258487,0.543258,0.52439487,0.32821837,0.13958712,0.18485862,0.27917424,0.73188925,1.3128735,1.6524098,1.2525115,1.8485862,1.6033657,1.6712729,2.093807,1.780679,1.9127209,1.7769064,2.2258487,3.0558262,3.0218725,3.5575855,3.1652324,3.4142256,4.1498876,3.4972234,4.0178456,3.9159849,4.1008434,4.7308717,5.221313,5.4401255,6.3644185,6.790725,6.670001,7.0963078,7.454707,7.964011,9.027891,10.714255,12.762791,10.710483,9.461743,8.959985,9.242931,10.469034,12.37421,14.139798,17.101309,20.734346,22.628204,19.844007,17.365393,14.807553,12.479843,11.378237,9.208978,7.5075235,6.9680386,7.3000293,7.2472124,7.5716586,8.137552,8.82417,9.522105,10.140816,9.842778,10.457717,10.487898,9.865415,9.929549,10.265312,10.340765,10.099318,10.201178,12.042219,13.472044,14.434063,15.671484,16.980585,17.23335,17.165443,16.188334,14.754736,13.713491,14.339747,15.286676,16.177015,17.040947,18.03692,19.47429,21.326649,22.473528,22.07363,20.274086,18.202915,17.16167,17.067356,17.312576,17.1164,15.531898,14.8339615,14.698147,14.811326,15.203679,16.252468,16.878725,16.58446,16.063837,15.55076,14.830189,14.200161,14.298248,15.226315,16.984358,19.4592,21.1267,20.82489,19.67424,18.595268,18.301004,21.31533,21.436056,20.138271,19.047983,19.957186,21.4851,23.816582,26.023567,27.181763,26.34424,22.843245,20.583443,18.881989,17.546478,16.874952,17.629477,18.934805,20.858843,23.348776,26.22729,27.615616,28.339958,27.841972,26.921452,27.721249,27.19308,26.480055,26.374422,26.940315,27.532618,25.287905,22.341486,20.289177,19.61765,19.68933,20.621168,21.005976,20.945614,20.798481,21.1682,21.681276,21.83218,23.107328,25.370903,26.90636,31.210926,33.912125,34.330887,32.78411,30.577126,30.263998,30.905344,33.191555,36.104023,36.900043,30.645033,24.522062,18.723537,13.890805,11.121698,11.087745,8.171506,5.3194013,3.6783094,2.5691576,1.8599042,2.0636258,2.4069347,2.6597006,3.1199608,5.9682927,10.86516,16.275105,21.11161,24.722012,25.525581,18.629223,11.272603,7.567886,8.488406,10.985884,8.314865,4.485651,1.7882242,0.80734175,0.7469798,0.663982,0.5885295,0.63002837,0.9808825,1.3015556,1.3128735,2.6823363,5.832478,9.922004,8.941121,6.673774,4.9723196,4.768598,6.0739264,11.457462,16.923996,17.542706,13.664448,10.914205,10.484125,10.469034,9.774872,8.209232,6.458734,8.258276,7.9300575,6.6624556,5.696664,6.319147,5.5683947,4.6214657,3.9499383,3.7990334,4.172523,4.6554193,4.745962,4.172523,3.3123648,3.187868,2.5578396,2.425798,2.6785638,3.1539145,3.6481283,4.564876,5.7796617,7.1076255,8.36391,9.397609,9.416472,9.627739,8.677037,7.1076255,7.3453007,6.096562,9.386291,9.250477,5.1043615,3.742444,3.8971217,3.8858037,3.6858547,3.4368613,3.4330888,4.214022,4.738417,4.2706113,3.4670424,4.353609,3.4934506,1.7919968,0.5281675,0.10186087,0.0,0.0,0.06790725,0.17354076,0.32821837,0.6111652,0.32821837,0.33953625,0.3169005,0.1659955,0.02263575,0.120724,0.26031113,0.51684964,0.8639311,1.1619685,0.784706,0.7997965,0.7884786,0.573439,0.24899325,0.181086,0.1961765,0.23013012,0.241448,0.241448,0.24522063,0.36971724,0.6111652,1.0450171,1.8259505,1.7995421,2.003264,2.6936543,3.7613072,4.749735,4.7912335,4.45547,3.9310753,3.3048196,2.5767028,2.686109,3.4670424,3.9801195,3.9310753,3.6745367,2.9916916,3.0181,3.2972744,3.3576362,2.7087448,2.444661,2.04099,1.9806281,2.4861598,3.5085413,4.4403796,4.647874,4.6290107,4.6931453,4.979865,5.081726,4.8666863,4.6252384,4.3875628,3.9386206,4.534695,4.5196047,4.459243,4.5422406,4.561104,4.8327327,4.9044123,4.6290107,4.4139714,5.2175403,5.0213637,5.534441,5.617439,5.624984,7.413208,9.208978,8.9788475,8.873214,9.386291,9.367428,9.899368,11.091517,12.713746,13.966258,13.521088,11.487643,11.1782875,11.212241,11.019837,10.842525,10.31813,10.367173,10.152134,9.593785,9.367428,11.065109,11.502733,11.3971,11.438599,12.306303,12.615658,12.925014,10.906659,9.74469,18.150099,28.204145,27.310032,21.922724,16.180788,11.898859,15.441354,18.433046,17.482344,13.128735,9.854096,4.52715,3.8556228,5.7607985,8.733627,11.846043,11.936585,11.133017,10.257768,9.910686,10.484125,10.899114,10.699164,10.34831,10.065364,9.827688,10.963248,12.061082,12.638294,12.717519,12.785426,13.026875,12.551523,11.642321,10.933067,11.41219,11.114153,11.170743,11.234878,11.231105,11.351829,12.181807,12.166716,12.332711,12.709973,12.332711,11.506506,10.419991,9.937095,10.34831,11.355601,11.532914,12.151625,12.377983,11.7026825,9.955957,9.574923,8.654402,8.028146,8.235641,9.510788,10.174769,10.487898,10.31813,9.759781,9.110889,9.948412,10.461489,10.170997,9.718282,10.853842,10.902886,10.653893,10.842525,11.329193,11.09529,8.741172,8.43559,8.801534,9.035437,8.903395,6.488915,5.292993,4.7006907,4.5422406,5.1156793,5.4703064,5.270357,4.9459114,4.636556,4.183841,3.7047176,3.0256453,2.474842,2.2748928,2.5427492,2.263575,2.1202152,2.1390784,2.2711203,2.4182527,2.535204,2.867195,3.2557755,3.4896781,3.2935016,3.7198083,4.3649273,5.0741806,5.666483,5.926794,5.7796617,5.938112,6.149379,6.436098,7.115171,6.8435416,5.4288073,4.3196554,3.99521,3.953711,3.9876647,3.9650288,3.863168,3.7386713,3.7462165,3.6292653,3.1161883,2.444661,1.8259505,1.4260522,1.3430545,1.2261031,1.0487897,0.84884065,0.7092535,0.69039035,0.56212115,0.47157812,0.45648763,0.45648763,0.5055317,0.47535074,0.49044126,0.63002837,0.9016574,0.95824677,0.935611,0.98465514,1.1053791,1.1506506,0.87902164,0.91297525,0.9318384,0.86770374,0.8903395,0.80734175,0.7092535,0.7054809,0.8224323,1.0148361,1.1431054,1.2147852,1.2902378,1.4034165,1.5920477,2.022127,2.0108092,1.7542707,1.539231,1.7391801,1.7089992,1.7240896,1.81086,1.9164935,1.9429018,1.9957186,2.203213,2.3880715,2.4522061,2.3805263,2.3088465,2.5238862,2.7992878,3.1539145,3.874486,4.768598,5.587258,5.832478,5.5759397,5.455216,5.515578,5.7872066,6.2436943,6.9152217,7.8998766,7.6584287,7.175533,6.5643673,5.956975,5.511805,2.1315331,2.3390274,2.7011995,3.0331905,3.270866,3.4783602,3.2369123,3.1199608,3.0822346,2.9992368,2.686109,2.7351532,2.655928,2.704972,2.8634224,2.8445592,2.848332,3.1048703,3.1652324,3.0407357,3.187868,3.4255435,3.9197574,4.45547,5.0062733,5.7192993,6.4134626,7.647111,9.718282,12.2119875,13.966258,14.637785,15.00373,15.373446,16.192106,18.052011,21.771818,24.250433,27.92497,32.067314,32.791656,31.83341,42.574074,43.136196,29.294434,14.471789,11.570641,9.982366,8.213005,6.0626082,4.6252384,2.916239,2.463524,2.5691576,2.7804246,2.8898308,2.886058,2.2484846,2.071171,2.516341,2.8521044,3.1010978,2.6710186,2.1164427,1.6486372,1.1242423,1.1355602,1.3091009,1.629774,2.252257,3.500996,1.9579924,1.3619176,1.1355602,0.97333723,0.8526133,0.784706,0.56589377,0.452715,0.5357128,0.73566186,0.65643674,0.452715,0.3734899,0.44516975,0.48666862,0.845068,0.8941121,0.66020936,0.331991,0.26031113,0.30935526,0.33953625,0.29049212,0.181086,0.12826926,0.090543,0.056589376,0.03772625,0.049044125,0.10940613,0.16976812,0.23767537,0.19994913,0.10186087,0.1358145,0.16222288,0.21881226,0.29049212,0.362172,0.4376245,1.20724,1.1280149,0.66020936,0.27917424,0.452715,0.5017591,1.3958713,2.3126192,2.5729303,1.6410918,2.252257,2.1315331,2.8181508,3.9197574,3.1237335,3.7462165,3.048281,3.3312278,4.538468,4.236658,3.6368105,3.3727267,4.327201,5.5495315,4.255521,5.191132,5.142088,5.119452,5.2364035,4.727099,5.221313,5.3759904,5.455216,5.7607985,6.617184,7.5188417,8.605357,9.903141,11.046246,11.25374,10.314357,10.687846,10.70671,10.382264,11.378237,13.143826,15.071637,18.18028,21.809546,23.639269,19.376202,16.4411,14.422746,12.808062,10.993429,9.34102,7.8734684,7.3717093,7.6395655,7.4811153,8.228095,8.809079,9.7069645,10.570895,10.223814,10.329447,10.831206,10.93684,10.657665,10.808571,11.815862,11.740409,10.944386,10.808571,13.728582,15.07541,16.071383,17.723793,19.636513,20.025093,19.945868,17.769064,15.62244,14.724555,15.39231,15.871433,17.338985,19.130981,20.602304,21.138018,21.952906,22.137764,22.107582,21.420965,18.806536,17.953922,18.104828,18.817854,19.289433,18.350048,16.595778,15.7657995,15.169725,15.022593,16.452417,18.327412,18.85558,18.297232,17.105082,15.905387,14.713238,14.083209,14.283158,15.629986,18.451908,21.741638,21.979313,21.228561,20.606077,20.270313,22.069857,21.884998,20.892797,20.183544,20.75321,22.330168,25.02382,27.581661,28.702131,27.038403,23.190327,21.254969,19.727057,18.02183,16.490145,17.14658,18.919714,21.296469,23.775084,25.876434,27.770292,30.041412,30.131956,28.377686,28.004196,28.373913,28.362595,28.868126,29.76224,29.898052,30.241362,28.434275,25.789665,23.522316,22.745155,23.111101,23.114874,23.02433,23.031876,23.284641,23.190327,22.941332,23.58268,25.302996,27.438301,32.42194,36.620872,37.5678,35.21368,31.957907,29.747149,28.81531,29.24916,30.301723,30.35454,26.838455,22.281124,17.60684,13.800262,11.9064045,14.313339,10.601076,6.5341864,4.504514,3.5387223,2.2447119,2.4484336,2.897376,2.9954643,2.8030603,4.878004,7.7640624,10.933067,13.826671,15.860115,17.282394,14.4114275,9.812597,6.971811,10.299266,14.509516,11.41219,6.4436436,2.6898816,0.90920264,0.66775465,0.66020936,0.80734175,1.0940613,1.5731846,1.4524606,1.0223814,1.358145,2.6785638,4.3422914,3.5689032,2.7691069,3.0143273,4.3913355,6.006019,11.200924,17.36162,19.24416,16.546734,13.917213,10.306811,10.3634,10.665211,9.850324,8.627994,9.058073,8.288457,7.277394,6.8435416,7.699928,6.670001,4.5460134,3.99521,4.9987283,4.851596,4.3800178,4.4931965,4.168751,3.338773,2.9086938,2.969056,2.5389767,2.1315331,2.11267,2.674791,3.3274553,4.745962,7.303802,9.986138,10.359629,12.58925,9.993684,8.631766,9.348565,7.77538,5.523123,9.291975,10.536942,7.2962565,4.187614,3.6028569,2.886058,3.4179983,4.7535076,4.6252384,4.561104,5.160951,4.696918,3.470815,3.7990334,2.7615614,1.7693611,0.7696155,0.0,0.0,0.0,0.17354076,0.29426476,0.30181,0.3169005,0.24899325,0.32067314,0.38858038,0.331991,0.056589376,0.018863125,0.19994913,0.44139713,0.6828451,0.9393836,0.845068,0.9620194,0.9016574,0.5998474,0.32444575,0.20749438,0.20749438,0.21503963,0.20749438,0.21503963,0.26408374,0.32444575,0.59230214,1.0978339,1.690136,1.7014539,1.8033148,2.4559789,3.62172,4.7912335,4.429062,4.2706113,4.0103,3.451952,2.516341,2.6823363,3.470815,3.9348478,3.8405323,3.682082,3.1237335,3.0822346,3.150142,3.0822346,2.8030603,2.2447119,1.9542197,1.9730829,2.335255,3.078462,3.983892,4.504514,4.7836885,4.9647746,5.191132,4.8855495,4.715781,4.5120597,4.2027044,3.802806,4.123479,4.08198,4.06689,4.293247,4.798779,5.0854983,5.1873593,5.1156793,4.9534564,4.8629136,5.0251365,6.1644692,6.058836,5.292993,7.281166,8.624221,8.160188,8.20546,9.288202,10.155907,10.567122,9.944639,10.808571,12.921241,13.253232,11.083972,11.529142,11.725319,11.231105,12.00072,10.827434,10.601076,10.091772,9.208978,9.012801,11.117926,11.004747,11.193378,12.385528,13.479589,11.830952,13.592768,12.362892,12.774108,30.475266,37.647026,26.536644,14.928277,10.710483,11.876224,13.962485,17.172989,19.221525,18.878216,15.961976,8.375228,5.081726,5.7004366,7.9451485,7.6282477,11.563096,11.23865,10.095545,9.955957,11.042474,11.189606,11.197151,11.344283,11.457462,10.944386,11.970539,12.189351,12.012038,11.725319,11.510279,11.910177,11.793225,11.072655,10.284176,10.597303,10.846297,11.419736,11.559323,11.310329,11.551778,12.393073,12.419481,12.6345215,13.151371,13.177779,11.480098,10.748209,10.56335,10.834979,11.8045435,12.770335,13.238141,13.5663595,13.189097,10.650121,9.167479,8.843033,8.677037,8.518587,9.092027,10.246449,10.499215,10.31813,9.944639,9.374973,9.148616,9.171251,8.967529,8.952439,10.453944,11.732863,11.32542,11.223559,11.536687,10.49167,8.729855,8.473316,9.167479,10.182315,10.804798,7.2283497,5.855114,5.372218,5.191132,5.4212623,5.492942,5.0439997,4.7836885,4.659192,3.893349,3.2557755,2.897376,2.4823873,2.093807,2.2258487,2.1768045,2.1164427,2.1541688,2.335255,2.637065,2.8521044,3.1425967,3.651901,4.06689,3.6066296,4.146115,4.749735,5.458988,5.9418845,5.511805,4.961002,5.2552667,5.753253,6.2436943,6.9491754,6.8963585,5.5457587,4.5007415,4.1498876,3.6934,4.055572,4.006528,3.9084394,3.8405323,3.6330378,3.712263,3.4029078,2.6785638,1.7995421,1.2902378,1.388326,1.1732863,0.87147635,0.6413463,0.55080324,0.47912338,0.43007925,0.40367088,0.43007925,0.543258,0.58098423,0.6111652,0.70170826,0.84129536,0.9318384,1.2147852,1.50905,1.6939086,1.7089992,1.5430037,1.0525624,1.0110635,0.995973,0.8865669,0.8978847,0.814887,0.7884786,0.845068,0.9922004,1.2185578,1.267602,1.2751472,1.2110126,1.237421,1.7127718,2.1088974,2.0447628,1.6788181,1.3392819,1.5241405,1.6486372,1.841041,1.9844007,2.022127,1.9353566,2.2484846,2.6672459,2.9501927,3.0822346,3.2482302,3.2067313,3.2029586,3.3161373,3.6783094,4.496969,5.028909,5.674028,6.1305156,6.2021956,5.798525,5.9796104,6.119198,6.4511886,7.073672,7.9413757,7.726336,7.1868505,6.4511886,5.7570257,5.4665337,2.1202152,2.2673476,2.4672968,2.41448,2.2447119,2.565385,2.674791,2.674791,2.5276587,2.2711203,2.0145817,2.11267,2.1164427,2.1654868,2.2711203,2.3201644,2.1466236,2.5993385,3.0105548,3.127506,3.127506,3.9197574,4.349837,4.8629136,5.534441,6.0739264,6.670001,7.828197,9.303293,10.684074,11.3669195,12.868423,13.13628,13.830443,15.354584,16.82968,18.881989,20.877707,23.299732,25.246407,24.431519,28.422956,35.61735,35.40986,25.691576,12.849561,10.065364,8.088508,6.2021956,4.2706113,2.7313805,2.1466236,2.0258996,2.1164427,2.305074,2.6106565,3.610402,3.2935016,3.2935016,4.112161,5.111907,6.405917,5.6476197,4.4894238,3.3576362,1.4637785,2.6483827,2.3692086,1.9730829,1.841041,1.388326,0.65643674,0.7092535,0.965792,1.0223814,0.65643674,0.754525,0.68661773,0.68661773,0.8563859,1.1732863,1.1129243,0.66775465,0.34330887,0.3169005,0.42630664,0.7922512,1.0601076,0.91297525,0.45648763,0.19994913,0.29426476,0.41121614,0.4074435,0.2867195,0.21503963,0.1659955,0.1056335,0.08677038,0.09808825,0.060362,0.060362,0.1056335,0.19240387,0.3055826,0.42630664,0.47535074,0.55080324,0.6073926,0.5093044,0.0452715,0.76584285,0.83752275,0.7809334,1.026154,1.8938577,1.6976813,2.5540671,3.5236318,3.863168,3.0218725,4.1197066,5.300538,6.5341864,6.9944468,5.0666356,6.115425,4.4931965,3.6971724,4.0178456,2.5012503,4.6742826,4.7610526,4.779916,5.353355,5.7079816,3.9499383,4.2517486,4.961002,5.081726,4.2894745,5.300538,4.3083377,4.8025517,7.213259,8.91094,9.314611,9.405154,9.265567,8.948667,8.484633,9.435335,11.476325,12.272349,11.891314,12.815607,15.260268,16.418465,17.761518,18.829172,17.244669,14.532151,15.309312,15.494171,13.970031,12.604341,9.318384,8.390318,8.409182,8.375228,7.6886096,7.8961043,9.669238,10.9594755,10.944386,10.038955,10.759526,10.729345,11.457462,12.577931,11.872451,11.053791,10.555805,10.917976,12.079946,13.396591,15.897841,17.357847,17.799244,18.244415,20.723028,19.696875,17.727566,16.874952,17.014538,15.8676605,18.16519,18.663176,20.319359,22.88097,22.918697,22.760246,22.03213,21.651094,21.613369,21.02484,19.353567,19.15739,20.059048,21.145563,20.949387,17.897333,15.897841,15.309312,15.803526,16.403374,18.500954,19.794964,19.968504,19.017803,17.271078,15.124454,14.158662,14.781145,16.437326,17.60684,22.782883,23.088465,21.824636,21.11161,21.881226,21.27006,20.613623,20.802254,21.496418,21.119154,22.997923,25.774574,28.094738,28.78513,26.857317,21.375692,19.47429,18.666948,17.599297,16.03743,17.086218,18.757492,21.156881,23.741129,25.314314,25.363358,27.8382,29.268024,28.309778,25.75571,26.09902,27.064812,29.298206,31.923952,32.546436,34.21771,34.874146,33.048195,29.215208,25.770802,25.895298,25.97075,26.215971,26.642279,27.068584,25.578398,25.242634,25.763256,26.853544,28.245644,31.724003,38.14124,40.910347,38.32987,33.568817,27.600525,25.43881,25.744392,26.55928,25.314314,24.12971,21.043703,17.716248,15.629986,16.0827,13.81158,11.514051,8.601585,5.80607,5.172269,3.3915899,3.0897799,3.3840446,3.4632697,2.6106565,3.451952,5.3571277,6.9680386,7.888559,8.684583,9.74469,9.808825,8.514814,8.028146,13.045737,16.950403,13.819125,8.228095,3.4594972,1.4939595,0.77338815,0.56589377,0.8111144,1.3770081,2.0598533,1.267602,0.7092535,0.95447415,1.8636768,2.6106565,2.546522,1.7014539,1.0450171,1.20724,2.4408884,3.9574835,5.824933,8.518587,12.147853,16.478827,13.622949,13.788944,13.800262,12.193124,9.201432,7.0510364,7.888559,8.6581745,8.201687,7.2472124,6.1116524,4.8025517,4.191386,4.3649273,4.606375,3.5575855,3.772625,3.4859054,2.7389257,3.3727267,2.848332,2.3880715,2.093807,2.052308,2.335255,2.0183544,2.837014,3.7990334,5.0251365,7.7376537,8.7751255,7.356619,8.560086,11.487643,9.276885,6.0286546,7.707473,10.419991,10.801025,6.043745,3.4557245,3.4745877,4.8440504,6.858632,9.397609,6.3945994,3.2935016,1.5656394,1.2864652,1.1129243,0.6149379,0.1961765,0.0,0.0,0.0,0.0,0.17354076,0.28294688,0.2678564,0.24522063,0.14713238,0.08677038,0.03772625,0.00754525,0.030181,0.056589376,0.19994913,0.4074435,0.5998474,0.67152727,1.1242423,1.3166461,1.1091517,0.6413463,0.33576363,0.19994913,0.18485862,0.18485862,0.181086,0.23013012,0.26408374,0.30181,0.77338815,1.3958713,1.1883769,1.4939595,1.4449154,2.0296721,3.4481792,5.0968165,4.0706625,3.7235808,3.3953626,2.795515,2.0145817,2.4031622,3.2821836,3.8367596,3.8782585,3.8292143,3.3161373,2.9501927,2.8030603,2.776652,2.595566,1.6184561,1.539231,1.8184053,2.2258487,2.8219235,3.8254418,4.191386,4.3196554,4.459243,4.715781,4.06689,3.8782585,4.2328854,4.644101,4.0593443,4.5460134,4.9345937,5.0515447,5.0439997,5.3873086,5.3382645,5.342037,5.6476197,6.0324273,5.8136153,5.0213637,5.66271,5.7607985,5.6476197,7.964011,7.696155,7.7376537,8.397863,9.446653,10.133271,9.80128,9.846551,10.518079,11.570641,12.253486,10.691619,10.38981,10.306811,10.453944,11.917723,10.197406,9.446653,9.110889,8.586494,7.2170315,11.393328,11.155652,10.533169,11.344283,13.200415,10.868933,15.611122,16.0412,18.161417,45.392223,38.81654,23.959942,11.32542,6.9567204,12.434572,10.080454,16.15438,26.64605,33.048195,22.367893,20.036411,14.958458,12.67602,12.219532,6.1041074,10.291721,10.925522,10.065364,9.416472,10.344538,10.884023,10.853842,12.261031,14.826416,15.961976,14.70192,13.060828,12.189351,12.1101265,11.717773,11.476325,11.495189,11.227332,10.499215,9.522105,9.88805,11.664956,12.427027,11.574413,10.329447,11.465008,12.657157,13.498452,13.604086,12.604341,11.348056,12.057309,12.570387,12.3289385,12.3893,13.743673,13.762536,13.29473,12.577931,11.261286,9.661693,9.125979,8.601585,8.07719,8.590267,9.676784,10.570895,10.993429,10.816116,10.069136,8.850578,8.20546,7.9300575,8.231868,9.733373,10.163452,9.574923,9.556059,9.918231,8.695901,8.586494,8.586494,9.058073,9.9257765,10.695392,7.6584287,6.5040054,6.296511,6.156924,5.2628117,4.9723196,4.1197066,4.1498876,4.689373,3.5387223,2.9313297,2.595566,2.3126192,2.0787163,2.0900342,2.1503963,1.991946,2.003264,2.3428001,2.9313297,3.4670424,4.0970707,4.1574326,3.742444,3.6934,4.376245,5.2250857,5.907931,6.0248823,5.0968165,4.534695,4.9421387,5.7004366,6.458734,7.1566696,6.5455046,5.1760416,4.2894745,3.9989824,3.2670932,3.0822346,3.0746894,2.8596497,2.6332922,3.1576872,3.5990841,3.3425457,2.5125682,1.5958204,1.448688,1.3015556,1.1280149,0.94692886,0.7809334,0.67152727,0.4640329,0.4376245,0.48666862,0.56589377,0.70170826,0.94692886,1.1355602,1.2261031,1.2713746,1.418507,2.1164427,2.7653341,2.7389257,2.1805773,1.9844007,1.4222796,1.0789708,0.87147635,0.7884786,0.8865669,0.9695646,1.1016065,1.2110126,1.2789198,1.327964,1.3392819,1.3505998,1.3204187,1.3317367,1.6033657,1.7240896,2.003264,1.8787673,1.4411428,1.4034165,1.6863633,1.8561316,1.9957186,2.1315331,2.2296214,2.4823873,2.7691069,2.9200118,3.2105038,4.3347464,4.7120085,4.5120597,4.2706113,4.349837,4.957229,5.534441,6.217286,7.0510364,7.643338,7.141579,6.934085,6.571913,6.5228686,6.903904,7.4773426,7.232122,6.7680893,6.1644692,5.674028,5.723072,2.2899833,2.252257,2.3918443,2.4522061,2.4484336,2.6974268,2.9351022,2.9313297,2.7389257,2.493705,2.3918443,2.2183034,2.1768045,2.1768045,2.2296214,2.4672968,2.1956677,2.4031622,2.7992878,3.1350515,3.2142766,4.2328854,4.5912848,4.776143,5.1156793,5.7796617,6.983129,8.058327,9.050528,9.842778,10.148361,11.793225,11.774363,12.068627,13.132507,13.8870325,16.33924,19.572378,21.760502,23.499681,27.796701,36.926453,41.41588,35.96821,22.971514,12.479843,10.868933,8.820397,6.809588,5.251494,4.478106,3.0407357,2.3880715,2.2107582,2.2862108,2.463524,2.9954643,2.867195,2.9086938,3.180323,2.9992368,2.7992878,2.3428001,1.7580433,1.1846043,0.7582976,1.3241913,1.358145,1.2902378,1.3128735,1.388326,1.4750963,1.4713237,1.2562841,0.9507015,0.9242931,0.98465514,1.1695137,1.3996439,1.4298248,0.87147635,0.73188925,0.513077,0.41498876,0.452715,0.47535074,1.1921495,2.372981,2.2975287,0.97333723,0.16222288,0.32821837,0.4376245,0.4376245,0.331991,0.18863125,0.18863125,0.12826926,0.1056335,0.11317875,0.03772625,0.056589376,0.06413463,0.1659955,0.36971724,0.56212115,0.6488915,0.4640329,0.694163,1.2147852,1.0827434,1.1996948,1.1242423,1.1506506,1.5203679,2.4182527,5.3269467,6.7643166,6.3908267,5.3609,6.3153744,6.809588,5.96452,5.666483,6.1908774,6.224831,5.7419353,5.1571784,5.402399,6.1116524,5.6023483,7.2887115,7.220804,6.4474163,6.1003346,7.3905725,7.4094353,8.118689,8.639311,8.503497,7.6810646,7.0548086,6.934085,8.013056,9.540969,9.314611,8.907167,8.643084,8.854351,9.469289,10.020092,10.672756,10.917976,11.7894535,13.075918,13.328684,12.706201,14.452927,16.033657,16.41092,16.033657,16.03743,15.999702,15.965749,15.01882,11.310329,8.786444,8.084735,8.00551,7.9715567,8.0206,9.857869,10.808571,10.963248,10.499215,9.673011,10.657665,11.000975,11.7555,12.770335,12.687338,11.3820095,10.79348,11.849815,13.815352,14.264296,15.301767,17.082445,18.62545,19.263023,18.648085,17.904879,17.399347,17.369165,17.765291,18.23687,20.006231,19.934551,19.738375,20.085455,20.613623,23.511,23.892035,22.560297,20.26277,17.693611,20.043957,20.764528,20.719257,20.813572,21.97554,20.515535,19.047983,17.889788,17.320122,17.57666,18.002966,19.180025,20.300495,20.69662,19.859098,20.085455,19.727057,19.319613,19.180025,19.413929,24.110846,25.717985,26.15561,26.012249,24.556017,22.126446,20.519308,19.247932,18.670721,19.983595,21.707684,23.228052,24.846508,25.79721,24.269297,21.160654,18.840488,17.229578,16.392056,16.550507,17.512526,19.410156,21.383238,23.179008,25.144547,25.834936,26.231062,27.061039,27.80802,26.721502,25.548216,26.480055,29.068075,32.301216,34.572334,36.137974,36.74537,35.83994,33.346233,29.679241,28.207916,28.121147,28.287142,28.28337,28.400322,26.480055,26.110338,26.566826,27.604298,29.464201,32.818066,38.095966,42.287354,42.807976,37.499893,30.00746,26.148064,25.216225,25.544443,24.495655,23.254461,21.534143,18.832945,15.905387,14.766054,12.581704,10.782163,8.548768,6.19465,5.160951,4.0216184,3.7537618,3.7914882,3.7650797,3.4896781,3.3048196,4.961002,6.587003,7.1264887,6.326692,6.881268,6.971811,6.5756855,6.8850408,10.299266,12.623203,11.570641,8.52236,4.9534564,2.4220252,1.8184053,1.599593,1.6750455,1.931584,2.2069857,1.5203679,1.0374719,0.7432071,0.69793564,1.0223814,1.3732355,1.4750963,1.8485862,2.8106055,4.4931965,4.930821,4.7044635,5.553304,7.752744,10.095545,11.974312,16.026112,16.361876,12.740154,10.582213,9.9257765,8.880759,8.299775,8.273367,8.103599,7.164215,6.809588,6.809588,6.911449,6.85486,4.1536603,3.7499893,3.3840446,2.8332415,3.8971217,2.9916916,2.3993895,2.505023,2.897376,2.3578906,2.4899325,3.0331905,3.651901,4.3422914,5.4401255,5.100589,6.270103,7.7376537,8.514814,7.835742,6.688864,6.0814714,6.2889657,6.907676,6.8359966,5.4212623,4.2404304,4.191386,5.1043615,5.7381625,3.9273026,3.3915899,2.384299,0.8224323,0.26031113,0.12826926,0.0452715,0.00754525,0.0,0.0,0.0,0.06413463,0.1358145,0.23767537,0.48666862,0.43007925,0.32821837,0.21881226,0.13204187,0.06790725,0.16976812,0.633801,0.79602385,0.6073926,0.62248313,1.0336993,0.95824677,0.90543,0.9205205,0.55457586,0.27540162,0.19994913,0.17731337,0.16222288,0.23013012,0.34330887,0.392353,0.6187105,1.0110635,1.3015556,1.4298248,1.6109109,2.0598533,2.9615107,4.4743333,4.2291126,3.99521,3.5689032,3.0633714,2.916239,3.0143273,3.5387223,3.9914372,4.112161,3.8669407,3.6669915,3.2746384,2.7087448,2.191895,2.1541688,2.0258996,2.0145817,2.0749438,2.2899833,2.848332,3.4859054,3.7952607,3.9725742,4.1800685,4.5422406,4.5120597,4.2064767,4.3875628,4.821415,4.255521,4.587512,4.9723196,5.111907,5.028909,5.0553174,5.0854983,4.768598,4.9119577,5.6023483,6.1908774,5.6325293,5.9532022,6.168242,6.2097406,6.9265394,7.7640624,7.7301087,7.8508325,8.405409,8.922258,9.393836,9.25425,9.763554,10.985884,11.778135,11.993175,12.049765,11.114153,9.95973,10.978339,9.06939,8.179051,8.477088,9.06939,7.986647,10.884023,10.374719,10.593531,12.102581,11.917723,10.77839,13.513543,12.581704,13.656902,35.61735,32.086174,19.65915,11.234878,10.819888,13.547497,8.13378,10.525623,18.23687,23.654358,14.007756,17.448391,12.6345215,8.443134,8.058327,8.98262,9.910686,9.933322,9.397609,8.952439,9.590013,11.69891,11.246195,11.174516,12.393073,13.81158,13.0646,12.234623,12.095036,12.457208,12.181807,11.498961,11.219787,11.16697,11.212241,11.291467,10.193633,10.642575,11.578186,12.030901,11.136789,10.921749,11.299012,11.868678,12.151625,11.589504,10.891568,11.555551,12.1252165,12.004493,11.498961,11.9064045,12.67602,12.981603,12.536433,11.589504,10.020092,9.016574,8.601585,8.820397,9.714509,10.223814,9.854096,9.763554,10.012547,9.57115,9.246704,8.616675,8.333729,8.763808,9.989911,9.129752,8.356364,8.345046,8.778898,8.379,8.993938,9.291975,9.74469,10.099318,9.352338,7.194396,6.096562,5.5985756,5.5004873,5.885295,5.4778514,4.779916,4.2592936,3.9989824,3.712263,2.8256962,2.3428001,2.1202152,2.1277604,2.4333432,2.3956168,2.3654358,2.4031622,2.5804756,2.9916916,3.3236825,3.5990841,3.62172,3.5387223,3.85185,4.9044123,5.885295,6.1833324,5.832478,5.5004873,5.142088,5.1345425,5.304311,5.73439,6.752999,6.092789,4.7044635,3.8820312,3.7462165,3.229367,2.8407867,3.169005,3.410453,3.3915899,3.572676,3.308592,2.7615614,2.0372176,1.4600059,1.5580941,1.2751472,1.1053791,0.9393836,0.7469798,0.55080324,0.4678055,0.44516975,0.47535074,0.58475685,0.83752275,1.0299267,1.4071891,1.5618668,1.4750963,1.5052774,1.750498,2.3767538,2.6936543,2.3880715,1.5203679,1.2298758,0.9808825,0.814887,0.8299775,1.1544232,1.5920477,1.7354075,1.7882242,1.8033148,1.7052265,1.629774,1.599593,1.5845025,1.6184561,1.7957695,1.9278114,2.093807,1.9504471,1.5807298,1.4637785,1.4826416,1.5580941,1.9278114,2.4559789,2.6295197,2.6634734,3.5575855,4.2517486,4.3611546,4.187614,4.8402777,4.9949555,4.7610526,4.398881,4.323428,4.878004,6.1342883,7.273621,7.756517,7.322665,6.900131,6.960493,7.0774446,7.069899,6.9869013,6.519096,6.3644185,6.3229194,6.360646,6.6134114,2.7540162,2.595566,2.5238862,2.625747,2.8634224,3.0520537,2.9841464,3.0256453,2.9351022,2.7087448,2.595566,2.4107075,2.263575,2.1881225,2.161714,2.0900342,2.033445,2.2220762,2.6408374,3.0105548,2.7879698,3.8593953,4.1083884,4.1612053,4.478106,5.349582,6.3531003,7.0812173,7.7150183,8.326183,8.899622,9.842778,10.238904,10.895341,11.951676,12.868423,15.946886,18.218006,20.270313,24.065575,32.96897,39.72197,37.499893,28.68704,17.727566,11.117926,10.114408,8.314865,6.2436943,4.5460134,3.9876647,3.2482302,2.7615614,2.505023,2.535204,2.9652832,3.1048703,2.5578396,2.2220762,2.3201644,2.4069347,1.7618159,1.2298758,0.814887,0.5470306,0.47157812,0.62248313,0.69039035,0.77716076,0.90543,1.0299267,1.3543724,1.448688,1.4411428,1.4222796,1.4298248,1.3694628,1.3355093,1.3015556,1.1544232,0.663982,0.6451189,0.5093044,0.41498876,0.41876137,0.51684964,1.2336484,2.3578906,2.2975287,1.1053791,0.49044126,0.7469798,0.6451189,0.44139713,0.271629,0.15467763,0.13204187,0.116951376,0.1358145,0.16222288,0.120724,0.060362,0.026408374,0.116951376,0.32067314,0.5583485,0.52439487,0.35462674,0.5470306,0.995973,1.0035182,1.3468271,1.7580433,2.3578906,3.8292143,7.4018903,8.405409,8.07719,8.29223,9.276885,9.574923,8.446907,7.484888,8.039464,9.22784,7.9451485,7.141579,7.394345,7.7942433,7.745199,6.9567204,8.590267,7.4999785,6.058836,6.0324273,8.601585,9.567377,9.348565,9.1825695,9.107117,7.9715567,8.099826,9.5032425,10.578441,10.740664,10.412445,9.450426,8.688355,8.160188,8.156415,9.224068,10.201178,10.31813,11.18206,12.536433,12.242168,12.377983,14.34352,16.173243,17.225805,18.19537,16.91645,14.339747,12.864652,12.487389,10.785934,9.435335,8.586494,8.541223,9.178797,9.95973,11.834724,12.15917,11.348056,10.057818,9.208978,10.072908,10.993429,11.834724,12.672247,13.762536,12.943876,13.034419,13.585222,14.268067,14.909414,17.244669,18.976303,20.391039,20.873934,18.94235,17.852062,17.701157,18.45568,19.60256,20.16468,20.48158,19.779873,19.051756,18.836716,19.221525,21.594505,22.183035,21.794455,20.413673,17.21826,19.21398,21.798227,23.201643,23.231825,23.284641,22.598024,21.571869,20.341993,19.164934,18.43682,18.7839,19.572378,20.704166,21.839725,22.394302,24.35984,25.472763,25.876434,25.706667,25.084183,26.476282,27.498663,28.44182,28.924715,27.868382,25.235088,22.1189,19.425245,18.157644,19.406384,20.836208,21.715229,22.782883,23.80149,23.563816,21.768045,19.40261,17.77661,17.28994,17.437073,18.723537,20.775846,22.748928,24.442837,26.29897,27.917425,27.800474,28.475773,29.784874,28.913399,27.815563,28.434275,30.546946,33.583908,36.63596,38.050697,38.34496,37.97147,36.828365,34.26298,31.433512,30.599762,30.128183,29.524563,29.437794,28.192827,27.49489,27.581661,28.592726,30.584671,32.806747,36.76423,41.408333,44.154804,40.89903,33.64804,27.970242,25.231316,24.771055,23.918442,21.888771,21.149336,19.519562,16.788181,14.709465,12.1252165,9.978593,7.914967,6.0814714,5.1571784,4.3649273,4.0706625,3.9876647,3.874486,3.5424948,3.2784111,4.2781568,6.0286546,7.405663,6.6624556,6.3116016,5.4967146,5.2288585,6.3908267,9.752235,11.114153,10.246449,8.001738,5.3458095,3.3689542,3.1765501,2.7992878,2.6936543,2.7653341,2.3805263,1.5618668,0.98842776,0.69793564,0.66775465,0.7997965,0.98842776,1.3392819,1.6939086,2.2258487,3.4594972,5.100589,6.3908267,7.5188417,7.9413757,6.356873,11.457462,17.769064,19.715738,17.301258,16.124199,11.887542,10.623712,10.397354,10.208723,9.989911,8.748717,8.235641,8.311093,8.356364,7.2698483,4.6252384,3.9386206,3.308592,2.4408884,2.637065,2.4182527,2.463524,2.6597006,2.8521044,2.8407867,3.078462,2.9049213,2.8445592,3.1539145,3.85185,5.2326307,6.300284,6.3116016,5.824933,6.72659,6.4021444,6.006019,6.7114997,7.4018903,4.6629643,4.142342,4.3800178,4.6214657,4.1574326,2.3578906,1.9504471,1.8938577,1.3694628,0.43007925,0.026408374,0.003772625,0.003772625,0.00754525,0.00754525,0.0,0.0,0.10186087,0.24899325,0.33576363,0.21881226,0.19994913,0.34330887,0.33953625,0.20749438,0.2678564,0.2678564,0.52062225,0.7167987,0.7394345,0.6752999,0.87147635,0.8601585,0.80734175,0.7507524,0.5998474,0.36594462,0.25276586,0.19994913,0.18863125,0.24899325,0.32444575,0.4376245,0.5696664,0.754525,1.0789708,1.4298248,1.841041,2.4710693,3.3312278,4.2819295,4.29702,3.8707132,3.259548,2.9916916,3.8405323,3.9499383,4.2894745,4.5309224,4.466788,4.014073,3.8556228,3.5689032,2.9086938,2.1013522,1.8523588,1.9881734,2.0485353,2.1013522,2.293756,2.8445592,3.1954134,3.429316,3.7914882,4.285702,4.647874,4.3800178,4.2027044,4.13857,4.112161,3.953711,4.4743333,4.878004,5.100589,5.0666356,4.67051,4.7120085,4.6252384,4.8365054,5.3948536,5.983383,5.938112,6.115425,6.0286546,5.8173876,6.273875,7.2887115,7.3905725,7.5226145,8.00551,8.503497,9.789962,9.714509,9.808825,10.480352,11.034928,11.725319,12.113899,11.344283,10.061591,10.431308,9.371201,8.7751255,8.82417,9.009028,8.152642,10.227587,10.106862,10.801025,12.276122,11.442371,10.838752,12.457208,11.615912,13.619176,33.77631,27.087448,16.237377,9.846551,10.416218,14.302021,9.87296,12.668475,18.961214,22.232079,13.189097,11.581959,7.1868505,4.8100967,5.9117036,8.567632,9.944639,10.314357,9.955957,9.242931,8.639311,10.533169,11.45369,11.9064045,12.132762,12.076173,11.664956,11.623458,11.876224,12.249713,12.479843,12.464753,11.7894535,11.578186,11.947904,11.989402,11.2801485,11.193378,11.615912,12.102581,11.868678,11.52537,11.551778,12.030901,12.445889,11.695138,11.038701,11.3971,11.981857,12.121444,11.23865,10.751981,11.46878,12.2119875,12.419481,12.113899,10.827434,10.253995,9.971047,9.899368,10.295494,9.967276,9.21275,9.084481,9.563604,9.556059,9.208978,8.605357,8.307321,8.424272,8.60913,7.835742,8.069645,8.416726,8.541223,8.677037,9.469289,9.122208,9.171251,9.374973,7.707473,6.952948,6.009792,5.3382645,5.2326307,5.832478,5.342037,4.9044123,4.406426,3.9273026,3.7348988,2.8785129,2.3201644,2.0673985,2.1353056,2.5276587,2.7502437,2.8143783,2.8294687,2.938875,3.3350005,3.5424948,3.8405323,3.8405323,3.6858547,4.0480266,4.644101,5.2552667,5.50426,5.4363527,5.5080323,5.4438977,5.372218,5.5457587,6.1041074,7.0548086,6.149379,4.9044123,3.9612563,3.4594972,3.0445085,2.8332415,3.2255943,3.500996,3.4066803,3.1463692,2.516341,2.2371666,1.8825399,1.4411428,1.3317367,1.146878,0.91297525,0.754525,0.67152727,0.55457586,0.44139713,0.4640329,0.66775465,0.98842776,1.2638294,1.1317875,1.3317367,1.4034165,1.3241913,1.50905,1.6788181,2.1315331,2.4672968,2.372981,1.6033657,1.297783,1.116697,1.116697,1.2940104,1.6033657,1.9844007,2.1466236,2.2107582,2.214531,2.093807,2.1654868,2.04099,1.9806281,2.071171,2.2598023,2.2183034,2.263575,2.11267,1.841041,1.8749946,1.8485862,1.8146327,2.1466236,2.8030603,3.3274553,3.7575345,4.346064,4.927048,5.311856,5.2854476,5.6551647,5.643847,5.2137675,4.557331,4.1272516,4.4139714,5.5306683,6.72659,7.4018903,7.1038527,6.4021444,6.5040054,6.72659,6.5266414,5.511805,5.119452,5.194905,5.523123,5.9418845,6.3417826,2.867195,2.8445592,2.625747,2.655928,2.9464202,3.0445085,2.8747404,2.8785129,2.7917426,2.5993385,2.5427492,2.4182527,2.305074,2.252257,2.214531,2.0372176,2.305074,2.4823873,2.7351532,2.9313297,2.6597006,3.5236318,3.6707642,3.7613072,4.1989317,5.119452,5.5683947,6.0324273,6.620957,7.356619,8.152642,8.503497,9.042982,9.982366,11.389555,13.166461,16.682549,17.870924,20.858843,27.940062,39.56729,38.725994,30.599762,21.405874,14.34352,9.578695,8.13378,6.198423,4.1989317,2.6785638,2.293756,2.305074,2.1466236,2.022127,2.071171,2.3805263,2.6182017,2.263575,1.8787673,1.7957695,2.1164427,1.5807298,1.056335,0.7884786,0.77338815,0.7507524,0.8639311,0.8941121,0.8865669,0.8865669,0.90920264,1.1619685,1.2638294,1.3543724,1.4449154,1.4260522,1.2826926,1.0487897,0.8262049,0.6413463,0.452715,0.6828451,0.7130261,0.6828451,0.65643674,0.6488915,1.1619685,1.7655885,1.6637276,0.95447415,0.63002837,0.784706,0.5583485,0.3055826,0.18485862,0.14335975,0.17354076,0.14713238,0.1358145,0.13958712,0.12826926,0.041498873,0.02263575,0.11317875,0.30181,0.5357128,0.392353,0.35462674,0.7205714,1.2525115,1.1921495,1.2902378,1.6637276,2.3013012,3.742444,7.069899,7.2962565,7.4697976,8.590267,9.839006,8.59404,8.492179,8.469543,9.22784,10.091772,9.005256,8.024373,8.043237,8.126234,7.8961043,7.533932,7.956466,6.900131,6.224831,6.696409,8.013056,8.582722,8.6732645,8.703445,8.639311,7.9828744,9.205205,10.736891,11.083972,10.253995,9.767326,8.480861,7.8432875,7.7225633,8.235641,9.714509,9.982366,10.269085,11.057564,12.215759,13.004238,13.445636,14.5132885,15.758255,16.980585,18.233097,16.380737,12.570387,10.257768,10.401127,11.438599,10.902886,10.408672,10.378491,10.948157,12.00072,12.672247,12.351574,11.227332,9.774872,8.756263,9.2995205,10.174769,11.046246,11.853588,12.823153,12.672247,13.5663595,14.64533,15.7657995,17.497435,20.568352,21.888771,22.756474,23.077147,21.371922,19.881733,19.644058,20.613623,22.00195,22.296213,21.032385,20.330677,19.768555,19.293203,19.21398,20.941841,21.31533,21.4851,21.122927,18.421728,19.444109,21.911406,23.84299,24.639013,25.080412,24.340977,23.084692,21.55678,20.100546,19.161163,20.198635,20.673985,21.677504,23.337458,24.83519,27.208172,29.550972,31.026068,31.437284,31.218472,30.980797,30.45263,30.313042,30.592216,30.701622,29.456656,25.646305,21.70391,19.398838,19.851553,20.760756,21.23988,22.03213,23.145054,23.820354,22.8357,20.979568,19.61765,19.176252,19.164934,20.711712,22.49239,24.197617,26.117884,29.120892,30.920435,31.622143,32.240852,32.69357,31.773048,31.988087,32.45212,34.093212,36.930225,40.076595,42.004406,41.8535,41.33288,40.668896,38.593952,35.417404,33.81781,32.55021,31.40333,31.184519,30.580898,29.381203,29.079393,30.214954,32.39553,33.565044,36.485058,40.778305,43.99258,41.638462,34.338432,27.962696,24.050484,22.503708,21.609596,20.387266,20.775846,19.893051,17.169216,14.335975,11.574413,9.242931,7.33021,5.9494295,5.342037,5.0025005,4.617693,4.2819295,3.9725742,3.5424948,3.3274553,3.9612563,5.775889,7.809334,7.8395147,6.832224,5.572167,5.451443,7.1981683,10.872705,11.996947,10.661438,8.145098,5.6098933,4.0782075,3.92353,3.3764994,2.987919,2.7125173,1.9164935,1.1016065,0.60362,0.5281675,0.7432071,0.8903395,1.1053791,1.6637276,1.8485862,1.7957695,2.5012503,5.5457587,8.892077,11.2650585,11.031156,6.217286,10.0465,14.913187,18.685812,20.813572,22.337713,13.622949,11.800771,11.9064045,11.638548,11.348056,10.133271,9.544742,9.869187,10.061591,7.745199,5.2099953,4.0782075,3.0218725,1.8976303,1.7693611,2.0900342,2.565385,2.7087448,2.7087448,3.470815,3.7160356,3.078462,2.848332,3.2218218,3.2972744,5.1647234,6.6549106,6.779407,5.881522,5.6098933,6.0248823,6.6850915,8.480861,9.171251,3.4066803,3.4481792,4.466788,4.7535076,3.6141748,1.358145,0.95824677,0.7394345,0.6073926,0.42630664,0.00754525,0.0,0.0,0.00754525,0.018863125,0.0,0.0,0.13958712,0.26031113,0.29049212,0.24522063,0.23390275,0.3734899,0.392353,0.30181,0.422534,0.482896,0.56212115,0.7884786,1.0223814,0.845068,0.87147635,0.88279426,0.875249,0.8337501,0.754525,0.5281675,0.33576363,0.23013012,0.211267,0.23390275,0.29049212,0.4074435,0.5885295,0.7884786,0.91674787,1.358145,1.9693103,2.8709676,3.92353,4.727099,4.3007927,3.7235808,3.259548,3.3161373,4.432834,4.323428,4.6554193,4.8666863,4.7346444,4.3422914,4.0480266,3.7009451,2.9652832,2.052308,1.7354075,1.8297231,1.8636768,1.9768555,2.305074,2.9954643,3.3840446,3.6443558,4.036709,4.5007415,4.659192,4.172523,4.0216184,3.9159849,3.8178966,3.9348478,4.478106,4.738417,4.949684,4.9760923,4.3309736,4.6290107,4.7836885,4.9459114,5.191132,5.5004873,5.73439,6.1908774,6.175787,5.8400235,6.19465,6.937857,7.1302614,7.3981175,7.865923,8.160188,9.665465,9.80128,9.778644,10.11818,10.661438,11.204697,11.487643,11.102836,10.310584,10.0276375,9.465516,9.405154,9.265567,8.801534,8.126234,9.525878,9.906913,10.401127,10.95193,10.336992,10.782163,11.41219,12.030901,16.109108,30.811028,23.186554,14.800008,9.963503,10.79348,17.18808,17.21826,21.03993,24.284388,23.831673,17.814335,14.200161,8.590267,5.73439,6.7379084,9.050528,9.175024,10.076681,10.797253,10.672756,9.348565,10.005001,10.940613,11.92904,12.261031,10.744436,10.355856,10.944386,11.480098,11.732863,12.261031,12.762791,11.823407,11.442371,11.910177,11.819634,11.834724,11.887542,11.849815,11.830952,12.174261,11.853588,11.59705,11.796998,12.140307,11.59705,11.419736,11.408418,11.876224,12.438345,12.027128,11.212241,11.291467,11.559323,11.706455,11.800771,11.231105,11.197151,10.997202,10.616167,10.748209,10.005001,9.325929,9.239159,9.676784,10.012547,9.276885,8.473316,7.997965,7.911195,7.91874,7.647111,8.194141,8.484633,8.495952,9.26934,9.378746,8.311093,8.141325,8.533678,6.730363,6.802043,5.9607477,5.198677,5.089271,5.802297,5.2137675,4.8666863,4.4818783,4.014073,3.6669915,2.8747404,2.3088465,2.04099,2.0787163,2.3993895,2.8181508,2.8936033,2.938875,3.169005,3.7084904,4.0480266,4.4101987,4.4139714,4.274384,4.8138695,5.010046,4.8365054,4.8742313,5.191132,5.330719,5.5797124,5.915476,6.360646,6.8058157,6.9944468,6.1606965,5.292993,4.3121104,3.4255435,3.1312788,3.1614597,3.2746384,3.1916409,2.8709676,2.5125682,1.9542197,2.0070364,1.8334957,1.3015556,0.995973,0.9620194,0.7205714,0.59607476,0.6149379,0.5055317,0.42630664,0.5357128,0.7922512,1.1091517,1.3543724,1.3166461,1.4449154,1.4939595,1.4524606,1.5316857,1.8297231,2.1881225,2.4182527,2.335255,1.7655885,1.5543215,1.4335974,1.5920477,1.9881734,2.3428001,2.3163917,2.4484336,2.6483827,2.8030603,2.746471,2.9086938,2.9539654,3.187868,3.5839937,3.7650797,3.3236825,3.1425967,2.927557,2.7200627,2.897376,3.1463692,3.2444575,3.4179983,3.8141239,4.534695,5.3684454,5.5306683,5.6551647,5.983383,6.3342376,6.537959,6.3455553,5.8173876,5.194905,4.8968673,4.7535076,5.3609,6.3153744,7.009537,6.620957,5.956975,5.873977,6.0286546,5.855114,4.5233774,4.29702,4.504514,5.0439997,5.6551647,5.938112,2.6710186,2.8294687,2.6332922,2.546522,2.655928,2.6898816,2.7389257,2.6634734,2.5540671,2.4974778,2.595566,2.372981,2.354118,2.41448,2.463524,2.4182527,2.938875,3.0181,2.9426475,2.8785129,2.8822856,3.3350005,3.4368613,3.6745367,4.2328854,4.9723196,5.119452,5.4401255,6.138061,7.1076255,7.9526935,7.967784,8.514814,9.710737,11.846043,15.384765,19.28566,20.85507,26.525326,37.19431,48.2481,37.647026,26.302742,18.270823,13.547497,8.058327,5.692891,3.3576362,1.6222287,0.754525,0.70170826,0.87902164,0.8941121,0.9318384,0.9922004,0.8903395,1.4600059,1.8561316,1.7919968,1.4750963,1.6109109,1.2638294,0.98465514,1.0072908,1.2449663,1.2751472,1.5920477,1.6637276,1.4449154,1.1431054,1.1883769,1.2600567,1.237421,1.1393328,1.0186088,0.98465514,0.814887,0.58475685,0.41121614,0.331991,0.331991,0.90543,1.2185578,1.3732355,1.4034165,1.2525115,1.2789198,1.2336484,1.0336993,0.72811663,0.47535074,0.42630664,0.25276586,0.14713238,0.15467763,0.18863125,0.271629,0.1961765,0.1056335,0.060362,0.05281675,0.011317875,0.0452715,0.181086,0.3961256,0.6073926,0.4376245,0.5357128,1.1732863,1.9579924,1.8221779,1.20724,1.0072908,1.1053791,1.358145,1.599593,2.957738,5.2062225,6.477597,5.9984736,4.0970707,6.587003,7.665974,7.673519,7.4094353,8.126234,7.462252,6.8850408,6.990674,7.7376537,8.439363,7.01331,7.0170827,7.575431,7.779153,6.7152724,6.673774,8.103599,8.582722,7.9791017,8.443134,9.661693,9.982366,9.756008,9.152389,8.145098,6.537959,6.670001,8.235641,10.401127,11.8045435,10.823661,10.540714,10.967021,12.219532,14.520834,14.151116,13.966258,14.407655,15.331948,16.029884,15.131999,12.600568,11.02361,11.363147,12.958967,12.276122,12.219532,12.113899,12.1101265,13.196642,12.362892,11.363147,10.423763,9.578695,8.654402,8.544995,8.6732645,9.4127,10.38981,10.472807,10.963248,12.434572,14.928277,18.127462,21.334194,24.408884,25.306768,25.634987,25.842482,25.216225,23.537407,23.001694,23.277096,23.759993,23.575134,21.636003,21.511507,21.454918,21.05502,21.232334,22.7942,22.775337,22.258488,21.488873,19.87796,20.866388,21.519053,22.548979,24.307022,26.793182,25.763256,24.00144,22.137764,20.7268,20.258997,21.719002,22.07363,23.175236,25.310541,27.2044,28.8304,31.241108,33.02933,33.964943,35.017506,35.560764,33.8744,32.23708,31.807001,32.621887,33.089695,29.875418,25.385994,21.824636,21.1682,21.488873,21.617142,22.277351,23.492136,24.567333,24.352295,23.314823,22.235851,21.65864,21.888771,23.001694,24.148573,25.344494,27.355305,31.697596,33.361324,35.45136,36.179474,35.432495,34.760967,35.94557,36.59069,38.46191,41.729004,44.962143,47.79916,47.45962,46.5806,45.71667,43.336143,40.378407,37.775295,35.69658,34.225254,33.36887,32.919926,31.467464,31.048704,32.33894,34.65156,35.73053,37.748886,40.412357,41.849728,38.586407,30.897799,25.05023,21.164427,19.002712,17.984104,18.700903,19.911915,19.251705,16.41092,13.143826,10.63503,8.646856,6.983129,5.828706,5.7570257,5.956975,5.583485,4.9647746,4.3422914,3.8480775,3.470815,4.104616,5.753253,7.7225633,8.654402,7.466025,6.5455046,6.820906,8.729855,12.23085,13.543724,12.128989,9.250477,6.205968,4.353609,4.1083884,3.5538127,2.7728794,1.8599042,0.935611,0.3772625,0.17354076,0.30181,0.6073926,0.79602385,1.2449663,1.9994912,2.2409391,2.0862615,2.6295197,5.7419353,9.695646,13.717264,15.052773,8.986393,7.8395147,9.25425,14.053028,20.564579,24.620152,14.8339615,12.204442,11.898859,11.574413,11.378237,10.56335,10.291721,11.00852,11.400873,8.371455,5.66271,4.0404816,2.7992878,1.9164935,2.0485353,2.1805773,2.5427492,2.8181508,3.218049,4.436607,4.4215164,3.783943,3.7688525,4.183841,3.380272,3.9197574,6.6020937,8.194141,7.364164,4.7044635,5.541986,6.700182,8.552541,9.148616,4.217795,4.696918,4.9119577,4.7044635,3.8707132,2.1315331,0.875249,0.543258,0.6413463,0.6526641,0.0,0.0,0.0,0.011317875,0.018863125,0.0,0.060362,0.13204187,0.1358145,0.1961765,0.6451189,0.5772116,0.5017591,0.422534,0.38103512,0.48666862,0.69793564,0.9205205,1.1695137,1.3128735,1.0525624,1.1808317,0.97710985,0.9620194,1.1317875,0.95447415,0.7167987,0.43007925,0.2565385,0.21503963,0.20372175,0.29049212,0.3734899,0.6451189,0.97710985,0.9318384,1.2751472,1.9844007,3.0256453,4.293247,5.583485,4.425289,3.8178966,3.7386713,4.0895257,4.696918,4.063117,4.459243,4.8440504,4.8553686,4.7648253,4.3686996,3.731126,2.776652,1.8448136,1.7127718,1.6863633,1.6109109,1.7919968,2.3428001,3.2142766,3.8443048,4.2630663,4.561104,4.738417,4.6818275,4.2027044,3.8858037,3.893349,4.1498876,4.3686996,4.817642,4.745962,4.7610526,4.8327327,4.3347464,4.949684,5.0666356,4.927048,4.798779,4.983638,5.2892203,6.224831,6.651138,6.439871,6.48137,6.9189944,7.1906233,7.492433,7.748972,7.594294,8.695901,9.133525,9.435335,9.986138,11.046246,11.125471,10.917976,10.7218,10.438853,9.6051035,9.016574,9.276885,9.156161,8.477088,8.137552,8.812852,9.424017,9.4013815,8.899622,8.801534,10.306811,10.099318,12.445889,17.942604,23.492136,19.342249,14.720782,11.834724,13.057055,20.911661,24.20139,28.328642,28.834173,25.72553,23.48459,25.529354,16.437326,9.590013,9.450426,11.581959,8.858124,9.220296,10.95193,12.253486,11.197151,11.204697,10.340765,10.668983,11.646093,10.125726,9.533423,10.295494,10.955703,11.1782875,11.729091,12.366665,11.495189,11.09529,11.498961,11.393328,11.608367,12.042219,11.864905,11.336739,11.815862,11.310329,10.887795,10.812344,11.012292,11.0613365,11.751727,11.461235,11.668729,12.600568,13.226823,12.709973,12.079946,11.287694,10.653893,10.842525,11.034928,11.261286,11.129244,10.816116,11.09529,10.601076,10.023865,9.842778,10.148361,10.63503,9.654147,8.529905,7.8017883,7.7150183,8.262049,8.394091,8.235641,8.009283,8.20546,9.578695,8.601585,7.2283497,7.164215,7.865923,6.537959,6.771862,6.0286546,5.247721,5.1232247,6.0814714,5.485397,4.908185,4.432834,4.036709,3.5802212,2.7917426,2.2371666,1.9806281,1.9994912,2.1881225,2.565385,2.595566,2.7238352,3.150142,3.8556228,4.5761943,5.119452,5.300538,5.3344917,5.855114,5.855114,4.9232755,4.587512,5.05909,5.2099953,5.753253,6.620957,7.254758,7.2623034,6.4474163,5.9796104,5.4703064,4.557331,3.5538127,3.440634,3.5877664,3.3048196,2.7691069,2.252257,2.1051247,1.9391292,1.9768555,1.659955,1.0450171,0.76207024,0.79602385,0.6526641,0.6111652,0.6451189,0.41498876,0.45648763,0.62625575,0.7884786,0.935611,1.1959221,1.5279131,1.8334957,1.9730829,1.901403,1.6976813,2.142851,2.3993895,2.474842,2.3503454,1.9542197,1.901403,1.8485862,2.1579416,2.7691069,3.1539145,2.6898816,2.7992878,3.270866,3.772625,3.8254418,3.893349,4.2027044,4.8930945,5.66271,5.772116,5.028909,4.659192,4.3686996,4.134797,4.2102494,4.776143,5.13077,5.2062225,5.2250857,5.745708,6.6586833,6.6850915,6.4210076,6.319147,6.7077274,7.1038527,7.009537,6.5832305,6.1644692,6.2436943,5.8173876,5.7494807,6.0776987,6.368191,5.723072,5.617439,5.3910813,5.3458095,5.2779026,4.459243,4.4139714,4.67051,5.2250857,5.7607985,5.6551647,2.916239,2.6823363,2.6597006,2.5880208,2.4710693,2.595566,2.776652,2.795515,3.0030096,3.3915899,3.5839937,2.8030603,2.6106565,2.7540162,2.9049213,2.625747,3.1237335,3.048281,2.7917426,2.6408374,2.7615614,2.8219235,2.957738,3.3538637,3.9348478,4.349837,5.191132,5.247721,5.6476197,6.696409,7.8432875,7.1340337,8.790216,11.133017,14.517061,21.31533,26.27256,30.780848,41.20461,54.997326,60.697765,41.974224,29.052984,19.73083,12.415709,6.119198,4.006528,1.9579924,0.7130261,0.45648763,0.8224323,0.77338815,0.69793564,0.5696664,0.47535074,0.6111652,0.7696155,1.1921495,1.1619685,0.80734175,1.0978339,0.52439487,0.5998474,1.0148361,1.3845534,1.2525115,1.5580941,1.8523588,1.6260014,1.177059,1.6184561,1.4826416,1.358145,1.2487389,1.1431054,1.0223814,0.80356914,0.6187105,0.4979865,0.47912338,0.62625575,1.6373192,2.1466236,2.4408884,2.6898816,2.9615107,1.9353566,1.2562841,0.9205205,0.7432071,0.36594462,0.40367088,0.3470815,0.27917424,0.26408374,0.33576363,0.1659955,0.120724,0.09808825,0.06413463,0.0754525,0.0150905,0.08299775,0.30181,0.6187105,0.9016574,0.7432071,0.91297525,1.2713746,1.6524098,1.8448136,1.4071891,1.177059,1.1091517,1.1242423,1.0978339,0.965792,0.84129536,1.0148361,1.448688,1.7391801,2.5314314,3.9386206,4.6856003,4.466788,3.953711,5.8928404,6.6360474,8.318638,10.650121,10.895341,9.661693,9.737145,8.729855,7.1038527,8.179051,10.133271,10.929295,9.465516,7.164215,7.9791017,7.284939,7.2283497,8.492179,10.121953,9.537196,7.1679873,8.031919,10.56335,12.830698,12.513797,12.3893,10.080454,9.431562,10.819888,11.140562,11.823407,12.313848,13.7851715,15.90916,16.859861,15.347038,16.003475,16.852316,16.535416,14.32843,12.083718,10.842525,10.597303,11.363147,13.185325,12.049765,10.54826,9.473062,9.156161,9.461743,7.9338303,7.2698483,7.654656,8.850578,10.193633,11.668729,13.456953,15.686575,18.663176,22.873425,28.1966,29.36234,29.188799,29.135983,29.283115,27.585434,26.317833,24.83519,23.013012,21.254969,20.839981,21.066338,21.737865,23.148827,26.076384,25.699121,25.129456,23.22428,20.658894,19.927006,21.149336,21.802,22.801746,24.582424,27.083675,26.680004,25.544443,24.405111,23.492136,22.552752,22.918697,23.220507,24.601288,27.079903,29.569836,30.377176,30.980797,31.859818,33.074604,34.270527,34.991096,34.29316,33.53109,33.391502,33.90458,33.893265,32.09372,28.705904,24.854053,22.582933,22.631977,22.469755,22.7527,23.835445,25.785892,26.664913,26.080156,25.32186,25.087955,25.46522,24.63524,25.291677,26.457418,27.85329,29.890509,32.931244,35.734303,37.205627,37.360306,37.32258,36.371876,37.431984,40.782078,45.622353,50.062733,52.982746,53.36378,53.137424,52.66207,50.73426,46.92768,42.076088,39.027805,37.579117,34.455383,33.93099,33.176464,33.206646,34.312023,36.054977,38.71845,39.182484,37.831882,35.130684,31.61837,25.148317,20.02132,17.28994,16.520325,15.82239,16.373192,16.667458,16.075155,14.366156,11.7026825,9.556059,8.231868,6.6247296,5.270357,6.3342376,6.700182,6.779407,6.304056,5.3609,4.4101987,3.7877154,4.244203,5.342037,6.8133607,8.544995,7.4811153,6.9227667,7.484888,9.190115,11.476325,12.721292,12.479843,10.4049,7.0849895,4.0593443,4.7535076,4.5799665,3.3538637,1.5580941,0.33576363,0.13958712,0.23767537,0.4640329,0.6375736,0.56589377,0.7469798,1.0940613,1.4562333,1.8976303,2.71629,3.5689032,5.753253,11.861133,17.716248,12.344029,7.0472636,8.488406,12.559069,16.173243,17.25976,14.230342,12.740154,11.555551,10.423763,10.069136,9.276885,9.0957985,9.590013,9.737145,7.432071,5.270357,3.8065786,3.4142256,3.561358,2.7917426,2.0975795,2.052308,3.1727777,5.070408,6.439871,5.2779026,4.8629136,4.353609,3.5764484,2.9916916,3.5274043,5.5004873,6.156924,5.191132,4.776143,4.093298,4.002755,4.032936,4.304565,5.523123,6.7567716,5.983383,6.0814714,6.1229706,1.388326,1.0601076,0.6187105,0.4678055,0.47535074,0.0,0.0,0.0,0.0,0.0,0.0,0.29426476,0.14713238,0.1659955,0.48666862,0.7922512,0.5357128,0.6375736,0.55080324,0.32821837,0.59607476,0.5357128,1.2147852,1.539231,1.2864652,1.1129243,1.8448136,1.1883769,0.7469798,0.90543,0.80734175,0.784706,0.49421388,0.27917424,0.241448,0.23013012,0.31312788,0.5017591,0.7092535,0.88279426,0.9922004,1.4449154,2.033445,2.8822856,4.1762958,6.1795597,5.032682,4.29702,4.247976,4.696918,4.991183,3.9273026,4.221567,4.719554,4.9345937,5.0213637,4.8968673,3.904667,2.5691576,1.5279131,1.5430037,1.5052774,1.3845534,1.6675003,2.384299,3.127506,3.7499893,4.3649273,4.8327327,5.119452,5.2779026,4.5950575,4.06689,3.9461658,4.255521,4.8063245,5.6853456,5.2175403,4.8138695,4.957229,5.20245,5.485397,5.2628117,4.61392,4.06689,4.5912848,5.3382645,6.2663302,6.6850915,6.56814,6.530414,7.0057645,7.6395655,7.858378,7.5226145,6.911449,7.5226145,8.390318,9.190115,10.20495,12.3289385,11.548005,10.997202,10.733118,10.374719,9.0957985,8.971302,8.646856,8.107371,7.7112455,8.224322,8.07719,8.390318,8.597813,8.582722,8.66572,9.118435,9.020347,11.212241,14.656648,14.434063,14.094527,13.622949,13.166461,14.366156,20.387266,16.969267,21.470009,26.389511,27.430756,23.499681,34.251663,19.911915,9.175024,10.933067,14.268067,12.766563,9.752235,9.465516,11.6008215,11.306557,13.687083,11.427281,9.522105,9.782416,10.834979,10.174769,10.155907,10.438853,10.899114,11.657412,12.830698,12.51757,12.257258,12.321393,11.732863,11.393328,11.717773,11.536687,10.816116,10.680302,10.106862,10.11818,10.533169,10.985884,10.925522,11.84227,11.438599,11.359374,12.128989,13.151371,13.166461,12.555296,11.359374,10.269085,10.63503,10.710483,10.899114,10.963248,10.899114,10.985884,11.204697,10.26154,9.846551,10.340765,10.819888,10.208723,9.110889,8.360137,8.137552,7.9791017,8.345046,7.707473,7.2094865,7.515069,8.7751255,7.5527954,6.398372,6.4436436,7.17176,6.379509,7.073672,6.6624556,5.9607477,5.704209,6.5455046,6.2889657,5.1534057,4.3007927,3.983892,3.5538127,2.7879698,2.173032,1.9164935,1.991946,2.1503963,2.323937,2.3465726,2.493705,2.8936033,3.5387223,4.689373,5.9984736,6.8246784,6.828451,6.013564,5.485397,4.606375,4.22534,4.610148,5.4174895,6.2361493,6.952948,7.3000293,7.0963078,6.2399216,5.8513412,5.1043615,4.1310244,3.3576362,3.4783602,3.5274043,3.2557755,2.7804246,2.3126192,2.1654868,2.3616633,1.6976813,1.1053791,0.90920264,0.8224323,0.7507524,0.80734175,0.8903395,0.8526133,0.48666862,0.55080324,0.63002837,0.7997965,1.1091517,1.5882751,1.5882751,2.1541688,2.372981,2.1353056,2.1353056,2.5616124,2.2862108,2.1390784,2.354118,2.5616124,2.2107582,2.2748928,2.837014,3.519859,3.5085413,3.1312788,3.3953626,4.255521,5.2288585,5.3873086,5.191132,5.251494,5.772116,6.428553,6.3945994,6.149379,6.0512905,5.8437963,5.43258,4.881777,5.1647234,5.4363527,5.696664,5.855114,5.723072,6.3342376,6.5756855,6.466279,6.255012,6.439871,7.2094865,7.594294,7.3490734,6.8058157,6.8661776,6.8435416,5.96452,5.1534057,4.636556,3.953711,4.9421387,5.032682,4.8138695,4.6554193,4.715781,4.9232755,5.1835866,5.4703064,5.5457587,4.961002,3.1576872,2.8106055,2.5691576,2.4031622,2.3163917,2.3503454,2.505023,2.7502437,2.9992368,3.1652324,3.1350515,2.8785129,2.7125173,2.776652,2.9728284,2.9652832,3.0181,3.1350515,3.1161883,2.9803739,2.9954643,3.1237335,3.3312278,3.731126,4.274384,4.776143,5.832478,5.772116,5.7306175,6.3945994,8.001738,8.514814,10.955703,14.373701,20.23636,32.43703,37.5678,44.845192,57.03832,68.30715,64.20253,39.688015,24.423975,14.664193,8.179051,4.2630663,2.5502944,1.3958713,0.68661773,0.3961256,0.56589377,0.694163,0.6828451,0.543258,0.42630664,0.6451189,0.63002837,0.6149379,0.55457586,0.4678055,0.42630664,0.25276586,0.39989826,0.65643674,0.7884786,0.56589377,0.9318384,1.0601076,1.1657411,1.2826926,1.2638294,1.2562841,1.2789198,1.2713746,1.2487389,1.2902378,1.1280149,1.0412445,0.9695646,0.98465514,1.297783,2.142851,2.4069347,2.806833,3.4783602,3.9725742,2.7426984,1.6486372,0.84884065,0.41121614,0.3169005,0.2565385,0.30181,0.26031113,0.15845025,0.24899325,0.23390275,0.21881226,0.18485862,0.1358145,0.08677038,0.15467763,0.31312788,0.62625575,0.8601585,0.48666862,0.452715,0.7432071,1.1619685,1.5769572,1.9202662,2.0673985,1.5505489,1.1393328,1.1996948,1.720317,0.97333723,1.0374719,1.7014539,2.3201644,1.81086,2.1881225,2.6031113,2.7653341,3.0633714,4.561104,4.2781568,5.9984736,7.5263867,8.058327,8.186596,8.495952,10.121953,10.329447,9.261794,9.937095,8.499724,9.8239155,10.657665,10.084227,9.507015,8.322411,8.035691,9.756008,12.083718,11.087745,9.997457,11.393328,12.653384,12.902377,13.023102,13.419228,11.370691,9.756008,9.616421,10.137043,11.200924,13.057055,14.400109,14.852824,14.943368,14.875461,15.452672,15.878979,16.135517,17.014538,15.373446,14.117163,13.792717,14.441608,15.577168,12.97783,11.268831,10.182315,9.371201,8.43559,7.54525,7.7414265,8.560086,9.393836,9.495697,10.446399,11.532914,15.116908,20.541943,24.12971,27.675978,28.675722,29.513245,30.471493,29.709421,28.762493,27.042175,24.752193,22.684793,22.194353,22.57916,23.680767,25.431265,26.981813,26.698868,26.351786,25.661396,24.110846,21.934042,20.1345,21.96045,22.911152,23.182781,23.235598,23.812809,24.514517,24.767282,24.325886,23.4695,23.028103,24.186298,26.019794,28.023058,30.279089,33.451866,34.61006,34.225254,34.387478,35.349495,35.52681,33.75745,31.901318,31.214699,31.50142,31.135473,30.067822,30.188545,29.41893,27.460938,25.804754,24.107073,23.601542,24.186298,25.56708,27.27608,28.788902,31.022295,31.093975,29.128437,28.238098,27.574116,27.932516,28.747402,29.483065,29.64906,29.279343,31.052477,33.49714,35.209908,34.88169,33.421684,34.296932,36.66237,40.28409,45.5469,48.942265,51.635918,54.031536,55.114277,52.431942,48.436733,44.48302,41.423424,38.94858,35.590942,35.22877,33.93099,33.772537,35.364586,37.850746,40.98957,40.91412,38.00165,33.033104,27.174217,20.96825,17.467255,15.833707,15.207452,14.735873,13.920986,13.928532,13.223051,11.544232,9.895596,8.627994,8.27714,7.9791017,7.5490227,7.466025,7.9715567,8.345046,7.964011,6.7379084,5.093044,4.247976,3.8707132,4.3347464,5.6551647,7.5075235,8.360137,8.786444,9.205205,9.748463,10.253995,10.823661,9.556059,7.4509344,5.7419353,5.87775,5.0515447,3.8858037,2.4899325,1.1129243,0.17731337,0.116951376,0.16222288,0.18863125,0.17731337,0.211267,0.36594462,0.60362,0.8978847,1.3355093,2.1051247,4.032936,5.583485,7.8961043,10.001229,8.827943,8.043237,10.295494,12.185578,12.604341,12.755245,13.573905,12.81938,10.902886,9.020347,9.144843,9.103344,8.714764,7.9828744,7.696155,9.431562,7.281166,5.5570765,5.1458607,5.20245,3.1350515,2.1654868,1.7655885,2.0372176,2.837014,3.7537618,3.7273536,3.3274553,3.1576872,3.2142766,2.8936033,3.1765501,3.4745877,3.832987,4.6290107,6.6058664,5.59103,4.1310244,4.5422406,6.356873,6.3153744,8.967529,8.722309,8.967529,9.265567,5.379763,2.1805773,0.67152727,0.23390275,0.23013012,0.0,0.0,0.0,0.0,0.124496624,0.62248313,0.32067314,0.14335975,0.38858038,1.0072908,1.5731846,0.5357128,0.42630664,0.47535074,0.452715,0.694163,0.8563859,0.9922004,1.2185578,1.3241913,0.77338815,1.1619685,0.97333723,0.8903395,1.116697,1.3694628,1.0148361,0.55457586,0.271629,0.241448,0.32821837,0.35462674,0.5394854,0.7130261,0.87902164,1.2223305,1.4901869,2.0108092,2.7125173,3.7537618,5.5193505,4.6742826,4.1762958,3.7877154,3.640583,4.255521,3.9574835,4.376245,4.7950063,4.9647746,5.081726,5.221313,4.29702,2.7879698,1.4939595,1.5052774,1.5279131,1.327964,1.5618668,2.252257,2.7615614,3.6368105,4.4630156,4.640329,4.398881,4.7912335,4.3724723,4.123479,4.112161,4.4215164,5.1345425,5.828706,5.836251,5.5759397,5.1873593,4.5309224,4.98741,4.7233267,4.0404816,3.6179473,4.4818783,4.8666863,5.624984,6.0022464,6.092789,6.8359966,6.930312,7.2094865,7.756517,8.182823,7.6320205,7.432071,8.22055,8.6732645,8.956212,10.718028,10.902886,10.759526,10.495442,9.955957,8.654402,8.7751255,8.552541,7.937603,7.6093845,8.933576,7.8961043,7.6282477,7.61693,7.7187905,8.152642,8.537451,10.0276375,16.395828,21.94536,11.480098,7.7602897,5.772116,4.9987283,6.5455046,13.147598,13.196642,19.787418,23.978804,21.986858,15.184815,18.244415,12.709973,7.24344,5.704209,7.149124,11.800771,14.524607,13.528633,9.80128,7.0963078,11.763044,12.58925,10.940613,9.035437,9.967276,10.167224,10.510533,10.665211,10.589758,10.54826,11.45369,11.815862,12.336484,12.996693,13.0646,12.381755,11.566868,11.106608,11.038701,10.974566,10.850069,11.091517,11.129244,10.861387,10.646348,11.227332,11.495189,11.887542,12.344029,12.336484,12.31762,11.891314,11.310329,10.95193,11.306557,11.359374,11.246195,11.038701,10.872705,10.93684,11.363147,10.948157,10.352083,9.918231,9.669238,9.880505,9.457971,9.020347,8.718536,8.235641,8.152642,7.284939,6.6624556,6.700182,7.175533,5.8664317,5.323174,5.613666,6.296511,6.4511886,7.1566696,7.0548086,6.673774,6.3153744,6.0324273,5.7381625,4.9647746,4.349837,4.0103,3.5538127,3.380272,2.8936033,2.4672968,2.2409391,2.1277604,2.1692593,2.1503963,2.3880715,3.0256453,4.0178456,5.349582,6.4738245,7.281166,7.567886,7.0246277,5.3269467,4.8553686,4.708236,4.8025517,5.8928404,6.436098,6.952948,7.009537,6.628502,6.2889657,5.8513412,4.798779,3.802806,3.2482302,3.2331395,3.2444575,3.0860074,2.6936543,2.2371666,2.1315331,1.9429018,1.358145,1.0638802,1.0940613,0.8224323,0.83752275,0.84129536,0.69793564,0.46026024,0.3772625,0.8903395,1.2789198,1.7618159,2.3314822,2.757789,2.3692086,2.546522,2.505023,2.3503454,3.0520537,3.2255943,2.5993385,2.2183034,2.3692086,2.5880208,2.1843498,2.5917933,3.2067313,3.7198083,4.1083884,3.6028569,4.1498876,5.1156793,6.0739264,6.779407,7.3151197,7.484888,7.1000805,6.258785,5.342037,5.5683947,5.764571,6.1116524,6.609639,7.0548086,6.398372,5.492942,5.4665337,6.1908774,6.270103,6.6662283,6.7039547,6.7756343,7.194396,8.209232,9.507015,9.627739,8.4544525,6.8359966,6.587003,6.387054,6.2851934,6.1418333,5.8098426,5.1345425,5.2665844,5.3458095,5.379763,5.409944,5.5080323,5.726845,5.6891184,5.5382137,5.251494,4.666737,3.0105548,2.6672459,2.4672968,2.3918443,2.372981,2.2899833,2.2975287,2.4710693,2.5993385,2.6182017,2.5917933,2.5201135,2.5125682,2.625747,2.8332415,2.9954643,2.9124665,3.1425967,3.187868,2.9652832,2.8219235,3.218049,3.4972234,4.0593443,4.851596,5.3684454,6.458734,6.247467,6.187105,6.900131,8.197914,10.529396,14.2077055,19.210207,26.668686,38.880672,42.317535,49.402523,58.901993,63.663048,50.594673,28.762493,16.535416,9.25425,4.617693,2.674791,1.6260014,1.0487897,0.6526641,0.38103512,0.392353,0.58098423,0.6451189,0.62248313,0.55080324,0.4640329,0.38103512,0.35839936,0.4074435,0.51684964,0.67152727,0.4376245,0.43385187,0.51684964,0.6187105,0.754525,1.0525624,1.0412445,1.056335,1.1581959,1.1204696,1.0186088,1.086516,1.3317367,1.6146835,1.6675003,1.5505489,1.5769572,1.5807298,1.6486372,2.142851,2.384299,2.3126192,2.5502944,3.1765501,3.742444,2.897376,1.8863125,1.0035182,0.46026024,0.3772625,0.20372175,0.271629,0.34330887,0.32821837,0.26408374,0.32067314,0.28294688,0.26031113,0.2678564,0.21881226,0.43385187,0.76584285,1.0223814,1.1242423,1.086516,1.3996439,1.8485862,2.263575,2.6031113,2.9539654,3.108643,2.323937,1.4562333,1.0412445,1.2902378,0.7696155,0.8111144,1.3694628,2.1315331,2.546522,2.4408884,2.5427492,2.6219745,2.8256962,3.663219,3.4783602,4.3800178,5.6815734,6.722818,6.8850408,7.073672,8.782671,9.224068,8.303548,8.601585,8.654402,9.156161,10.11818,10.948157,10.472807,10.038955,9.405154,9.910686,11.155652,11.00852,11.54046,12.543978,13.407909,13.8870325,14.094527,14.117163,12.857106,11.966766,11.710228,10.9594755,11.649866,13.275867,13.973803,13.65313,14.000212,13.419228,12.883514,13.283413,14.509516,15.422491,14.5132885,14.313339,14.124708,13.815352,13.849306,12.736382,11.887542,11.136789,10.412445,9.725827,8.575176,8.382772,8.2507305,8.001738,8.186596,10.33322,12.940104,17.542706,23.443092,27.721249,28.377686,29.07562,29.637741,29.581152,28.121147,27.891016,27.011995,25.574625,24.51829,25.608578,24.66165,25.751938,27.227036,27.95515,27.332668,27.01954,25.634987,24.07312,22.877197,22.228306,23.767538,24.291933,24.084438,23.488363,22.911152,23.895807,24.884235,24.831417,23.990122,23.89958,25.201136,27.53639,29.898052,32.172947,35.12691,36.454876,36.08516,36.039886,36.828365,37.435757,36.654823,35.15332,33.334915,31.429739,29.479292,28.01174,28.445593,28.532362,27.615616,26.619642,24.997414,24.427748,25.238861,26.974268,28.373913,30.211182,33.576363,33.953625,31.271288,29.875418,29.603788,30.309269,30.62617,30.346996,30.429993,30.445084,30.026323,30.475266,31.610825,31.76173,30.294178,30.456402,31.505192,34.187527,40.75567,43.97749,47.829338,52.00186,54.672882,52.507393,48.225464,45.007416,42.14022,39.17871,35.938026,35.77203,34.444065,34.059258,35.5004,38.40155,41.008434,41.706367,38.79013,32.53512,25.174726,19.429018,16.195879,14.034165,12.698656,13.12119,11.638548,11.299012,10.367173,8.7751255,8.099826,8.337502,8.956212,9.092027,8.669493,8.382772,8.605357,9.352338,9.295748,8.009283,5.9418845,4.8855495,3.863168,4.093298,5.560849,7.001992,7.7301087,9.65792,10.638803,10.382264,10.442626,10.295494,7.835742,5.824933,5.1534057,4.821415,3.482133,2.5729303,1.6146835,0.6187105,0.08299775,0.10940613,0.13204187,0.1056335,0.06413463,0.1056335,0.23013012,0.543258,0.87147635,1.3392819,2.372981,5.2892203,8.182823,9.118435,8.190369,7.54525,7.4773426,9.442881,10.785934,11.212241,12.781653,15.184815,14.313339,11.5857315,9.020347,9.250477,8.801534,7.605612,6.643593,6.6624556,8.14887,6.247467,4.9421387,5.149633,5.8588867,4.115934,2.8898308,2.4295704,2.1805773,2.142851,2.8822856,3.1312788,3.2557755,3.350091,3.5160866,3.874486,2.7992878,2.2183034,2.4069347,3.5839937,5.9003854,5.492942,3.772625,4.063117,6.307829,7.073672,9.220296,9.846551,9.582467,8.284684,5.0515447,1.6976813,0.49044126,0.33576363,0.3961256,0.090543,0.25276586,0.3470815,0.362172,0.46026024,0.9808825,0.59230214,0.41498876,0.5772116,0.98465514,1.3128735,1.0525624,1.1846043,1.1129243,0.845068,0.9808825,1.086516,1.1619685,1.3732355,1.5807298,1.327964,1.2902378,1.086516,1.026154,1.116697,1.1091517,0.8224323,0.49044126,0.331991,0.36971724,0.4074435,0.42630664,0.5017591,0.5998474,0.754525,1.0978339,1.4298248,2.0296721,2.7351532,3.6254926,5.0251365,4.146115,3.953711,3.8971217,3.893349,4.349837,4.0782075,4.1083884,4.395108,4.8025517,5.0854983,4.8930945,4.13857,2.8521044,1.6825907,1.8976303,1.7731338,1.388326,1.5920477,2.41448,3.0558262,4.074435,4.478106,4.327201,4.093298,4.640329,4.323428,4.2781568,4.4894238,4.8742313,5.300538,5.3344917,5.194905,5.0779533,4.8855495,4.217795,4.6516466,4.187614,3.6707642,3.6443558,4.346064,4.6818275,5.27413,5.455216,5.455216,6.417235,7.062354,7.4471617,7.567886,7.5075235,7.454707,7.0510364,7.809334,8.5563135,9.159933,10.518079,10.834979,10.34831,9.669238,8.963757,7.960239,8.209232,7.699928,7.375482,7.745199,8.899622,7.1793056,7.232122,7.3113475,7.0963078,7.6886096,7.6207023,8.68081,13.607859,18.044466,10.540714,7.4018903,5.9532022,5.3609,7.5301595,17.086218,17.108854,18.549997,16.724047,11.668729,8.16396,12.359119,10.733118,7.6622014,5.745708,5.802297,7.809334,14.471789,17.003222,13.93985,11.159425,10.061591,12.113899,12.359119,10.253995,9.650374,10.050273,10.33322,10.450171,10.3634,10.03141,10.733118,11.706455,12.6345215,13.302276,13.607859,12.736382,11.563096,10.77839,10.665211,11.083972,11.129244,11.283921,11.027383,10.442626,10.216269,10.748209,11.087745,11.555551,11.932813,11.45369,11.193378,11.23865,11.4838705,11.7026825,11.529142,11.6008215,11.680047,11.3971,10.884023,10.770844,10.93684,10.484125,9.808825,9.193887,8.778898,9.612649,9.578695,9.058073,8.518587,8.529905,8.326183,7.3113475,6.439871,6.2135134,6.6549106,5.3609,5.089271,5.455216,6.089017,6.6247296,7.115171,7.232122,6.8133607,6.1116524,5.8136153,5.5457587,4.8968673,4.4101987,4.123479,3.5651307,3.3878171,2.938875,2.5729303,2.4559789,2.5502944,2.5427492,2.5389767,2.848332,3.5424948,4.5007415,5.66271,6.48137,6.990674,7.115171,6.6850915,5.485397,5.240176,5.1081343,4.983638,5.4891696,5.4891696,5.987156,6.2361493,6.1116524,6.1078796,5.907931,4.708236,3.6481283,3.259548,3.4745877,3.2859564,2.9049213,2.4974778,2.1579416,1.9202662,1.5203679,1.2261031,1.1053791,1.0714256,0.87147635,0.8186596,0.7054809,0.5998474,0.6149379,0.91674787,1.4109617,1.8938577,2.4295704,2.927557,3.1539145,2.7804246,2.9954643,3.0671442,2.9766011,3.4179983,3.2142766,2.7728794,2.565385,2.6672459,2.7389257,2.3918443,2.8936033,3.7009451,4.4516973,4.9534564,4.847823,5.5004873,6.2889657,6.85486,7.1000805,8.031919,8.269594,7.835742,6.9189944,5.87775,6.089017,6.273875,6.507778,6.8246784,7.213259,6.6020937,5.670255,5.5570765,6.198423,6.3531003,7.009537,7.24344,7.1868505,7.2283497,8.009283,9.220296,9.748463,8.944894,7.4018903,6.964266,7.115171,6.8737226,6.560595,6.319147,6.138061,5.847569,5.5570765,5.4891696,5.674028,5.945657,6.156924,6.0248823,5.7607985,5.5382137,5.4703064,2.8521044,2.686109,2.6295197,2.6823363,2.7125173,2.4597516,2.282438,2.2899833,2.3126192,2.282438,2.2258487,2.2598023,2.3956168,2.546522,2.6936543,2.886058,2.848332,3.0369632,3.0331905,2.8407867,2.8785129,3.2331395,3.4481792,4.036709,5.0251365,5.96452,6.9491754,6.507778,6.5643673,7.5112963,8.197914,11.415963,16.188334,22.552752,30.407358,39.533337,39.92569,45.51672,51.23979,49.98351,32.584164,16.912678,9.276885,5.2628117,2.7125173,1.7278622,1.1053791,0.8186596,0.6413463,0.49044126,0.44139713,0.5357128,0.63002837,0.69039035,0.6375736,0.35839936,0.33576363,0.32067314,0.40367088,0.63002837,1.026154,0.8337501,0.69039035,0.56589377,0.55080324,0.83752275,1.2789198,1.3505998,1.3128735,1.2826926,1.2223305,1.1242423,1.2298758,1.5958204,1.9994912,1.9240388,1.7316349,1.780679,1.8297231,1.9240388,2.4107075,2.6144292,2.5012503,2.3993895,2.493705,2.8332415,2.516341,1.8221779,1.086516,0.56589377,0.44516975,0.23013012,0.23013012,0.34330887,0.452715,0.44894236,0.4376245,0.33576363,0.271629,0.27917424,0.3169005,0.7092535,1.3241913,1.659955,1.6825907,1.81086,2.4371157,3.0331905,3.4481792,3.663219,3.8254418,3.7990334,3.169005,2.214531,1.3845534,1.297783,1.0412445,0.8601585,1.0450171,1.5731846,2.0862615,1.9202662,2.3201644,2.5389767,2.4823873,2.71629,3.3048196,3.1576872,3.7462165,5.081726,5.726845,5.6023483,6.749226,7.069899,6.485142,6.8963585,8.14887,8.024373,8.503497,9.673011,9.733373,11.348056,10.910432,10.435081,10.582213,10.691619,11.378237,11.747954,12.619431,13.694629,13.551269,13.539951,12.864652,12.826925,13.019329,11.348056,12.5326605,13.505998,13.498452,12.755245,12.540206,11.517824,10.287949,10.657665,12.245941,12.513797,12.506252,12.894833,13.158916,13.124963,12.992921,12.562841,12.2270775,11.608367,10.804798,10.355856,9.435335,9.020347,8.439363,7.964011,8.82417,11.487643,14.724555,18.765038,23.45441,28.245644,28.106056,28.622906,28.366367,27.03463,25.453901,25.548216,25.087955,24.869144,25.589716,27.841972,27.061039,27.804247,28.422956,28.230553,27.502436,27.215717,25.982069,24.85028,24.35984,24.556017,25.4954,25.419947,24.997414,24.529608,23.937305,23.84299,24.718239,25.174726,25.140774,25.857573,26.721502,28.607815,30.852528,33.187782,35.764484,37.541393,36.971725,36.353016,36.711414,37.809246,40.250137,41.125385,38.639225,33.595226,29.411385,27.030859,25.865116,25.5369,25.593489,25.480309,24.940825,24.85028,25.733074,27.343987,28.664404,30.580898,33.938534,34.20639,31.497646,30.588444,30.279089,31.112839,31.44483,31.078884,31.290152,31.497646,29.59247,28.238098,28.14001,28.057013,26.597006,25.61235,25.4954,27.611843,34.285618,37.94506,42.691025,48.27451,52.51494,51.3077,46.63342,43.80772,41.264973,38.303463,35.077866,35.538128,35.130684,34.613834,35.089184,38.016743,39.1523,40.521767,38.17142,31.708914,24.269297,19.440336,15.720529,12.600568,10.544487,10.982111,10.789707,9.122208,7.4697976,6.6322746,6.72659,7.673519,9.133525,9.4127,8.756263,9.329701,9.261794,9.982366,10.084227,8.963757,6.779407,5.515578,4.055572,4.104616,5.564622,6.507778,7.303802,9.6051035,10.646348,10.148361,10.303039,10.005001,6.9454026,4.8402777,4.38379,3.2218218,2.0108092,1.5920477,1.4411428,1.0940613,0.16222288,0.15845025,0.18863125,0.150905,0.0754525,0.10940613,0.24522063,0.5696664,0.8337501,1.1129243,1.7995421,4.6818275,7.2698483,8.00551,7.303802,7.5829763,6.8473144,7.752744,9.34102,11.385782,14.4114275,17.312576,15.8676605,12.826925,10.11818,8.827943,8.137552,7.043491,6.477597,6.7077274,7.352846,5.666483,4.7836885,5.270357,6.156924,4.9723196,3.7613072,3.199186,2.7125173,2.3880715,2.9652832,2.9237845,3.1765501,3.5575855,3.8556228,3.832987,2.4597516,1.6637276,1.4864142,2.0447628,3.5575855,4.2291126,3.338773,3.9688015,6.5266414,8.75249,9.7296,10.265312,8.3525915,4.715781,2.7992878,0.7997965,0.362172,0.47157812,0.5055317,0.23013012,0.3734899,0.47157812,0.4376245,0.46026024,0.98465514,0.7922512,0.68661773,0.8111144,1.056335,1.056335,1.1959221,1.3770081,1.3053282,1.0789708,1.177059,1.0374719,1.2864652,1.6448646,1.8976303,1.8900851,1.6146835,1.237421,1.026154,0.9997456,0.90543,0.633801,0.42630664,0.36594462,0.41121614,0.392353,0.44894236,0.47157812,0.5055317,0.6187105,0.91674787,1.3996439,2.2296214,3.2142766,4.0895257,4.5120597,3.9574835,4.044254,4.0706625,3.9725742,4.323428,4.0291634,3.953711,4.0782075,4.4101987,4.9949555,4.4818783,3.7235808,2.7426984,1.9391292,2.123988,2.093807,1.6486372,1.7995421,2.686109,3.591539,4.3422914,4.5233774,4.3309736,4.13857,4.52715,4.4139714,4.4215164,4.659192,5.070408,5.4212623,5.111907,4.7874613,4.617693,4.534695,4.2291126,4.5422406,3.8707132,3.5047686,3.7877154,4.1197066,4.5724216,4.817642,4.8025517,4.9760923,6.2889657,7.069899,7.3868,7.1264887,6.620957,6.6247296,6.466279,7.2660756,8.333729,9.314611,10.20495,10.702937,9.993684,8.922258,7.9828744,7.3075747,7.643338,7.149124,7.073672,7.7678347,8.661947,7.175533,7.5037513,7.432071,6.7454534,7.194396,7.0585814,7.360391,9.2844305,11.393328,9.612649,8.578949,8.201687,8.09228,11.302785,24.307022,22.258488,18.285913,12.513797,6.700182,4.214022,9.34102,9.805053,8.409182,6.903904,5.9984736,4.447925,10.435081,16.086473,17.320122,13.853079,9.333474,10.79348,12.170488,11.400873,10.393582,10.340765,10.480352,10.578441,10.484125,10.121953,10.646348,11.480098,12.091263,12.457208,13.041965,12.298758,11.423509,10.514306,9.967276,10.450171,10.744436,10.672756,10.397354,10.072908,9.846551,10.559577,10.876478,11.072655,11.151879,10.834979,10.408672,10.597303,11.231105,11.868678,11.793225,11.721546,12.042219,12.076173,11.61214,10.921749,10.574668,9.97482,9.224068,8.499724,8.073418,9.088254,9.491924,9.21275,8.692128,8.854351,8.431817,7.515069,6.5455046,5.9909286,6.33801,5.111907,4.8930945,5.300538,5.9607477,6.507778,6.771862,7.1302614,6.8359966,6.043745,5.824933,5.3948536,4.708236,4.191386,3.9008942,3.5085413,3.2255943,2.727608,2.4484336,2.5427492,2.867195,2.8106055,2.795515,3.199186,4.044254,5.0251365,5.938112,6.5002327,6.7341356,6.590776,5.945657,5.3986263,5.1798143,5.05909,4.949684,4.8855495,4.568649,4.859141,5.194905,5.4363527,5.8702044,5.7192993,4.557331,3.6179473,3.4066803,3.682082,3.429316,2.897376,2.4107075,2.0862615,1.81086,1.3128735,1.1732863,1.0676528,0.95824677,1.0601076,1.0186088,0.8865669,0.8299775,0.9393836,1.267602,1.7316349,2.3692086,2.8822856,3.180323,3.3651814,3.2105038,3.3840446,3.5764484,3.7160356,3.983892,3.8065786,3.4142256,3.1954134,3.1539145,2.897376,2.7653341,3.2444575,4.1272516,5.0741806,5.613666,5.775889,6.549277,7.277394,7.564113,7.2924843,7.854605,7.8508325,7.462252,6.9152217,6.458734,6.4511886,6.2851934,6.092789,5.96452,5.934339,5.798525,5.5080323,5.5759397,5.9607477,6.066381,6.673774,7.1302614,7.1604424,6.983129,7.3075747,8.371455,9.352338,9.1976595,8.00551,7.0246277,7.6207023,7.5188417,7.01331,6.5756855,6.881268,6.587003,6.2625575,6.145606,6.2399216,6.3116016,6.417235,6.273875,6.1795597,6.3455553,6.907676,2.686109,2.7728794,2.8558772,3.0331905,3.1312788,2.7238352,2.4031622,2.282438,2.2862108,2.3013012,2.1956677,2.3277097,2.4484336,2.5201135,2.565385,2.674791,2.7691069,2.8936033,2.9086938,2.9086938,3.229367,3.350091,3.4972234,3.9159849,4.7836885,6.2021956,6.9567204,6.3531003,6.5040054,7.6018395,7.914967,10.884023,15.894069,22.349031,29.037895,34.138485,31.542917,35.579628,38.952354,35.142002,18.448135,8.771353,4.859141,3.3425457,2.354118,1.50905,0.97333723,0.72811663,0.6828451,0.7167987,0.6790725,0.633801,0.6828451,0.6828451,0.5772116,0.3772625,0.44894236,0.3772625,0.3961256,0.6111652,1.0072908,1.0374719,0.90920264,0.7130261,0.573439,0.6488915,1.2110126,1.5279131,1.6410918,1.6033657,1.478869,1.5430037,1.7316349,2.0108092,2.203213,2.003264,1.7165444,1.7354075,1.8825399,2.1277604,2.595566,3.1425967,3.108643,2.6144292,2.003264,1.8599042,1.8259505,1.4034165,0.90543,0.5583485,0.4979865,0.27917424,0.19240387,0.24522063,0.41498876,0.6187105,0.5470306,0.3961256,0.26031113,0.21881226,0.34330887,0.80356914,1.7391801,2.323937,2.3314822,2.142851,2.8521044,3.591539,4.055572,4.1762958,4.142342,3.85185,3.5538127,2.8709676,2.071171,2.0749438,1.961765,1.5052774,1.2600567,1.1921495,0.694163,0.7884786,1.6335466,1.9655377,1.7391801,2.123988,2.897376,2.4672968,2.4333432,3.289729,4.432834,4.478106,5.172269,5.3910813,5.2288585,6.0324273,6.7567716,6.790725,7.0246277,7.635793,8.080963,11.514051,11.725319,11.472552,11.578186,10.940613,10.921749,10.93684,11.615912,12.445889,11.766817,12.185578,11.589504,11.480098,11.819634,11.038701,12.96274,13.521088,13.034419,12.012038,11.151879,10.20495,9.461743,9.725827,10.638803,10.695392,11.32542,11.631002,12.272349,13.230596,13.830443,13.004238,12.51757,11.827179,10.884023,10.103089,10.057818,9.891823,9.676784,9.839006,11.155652,13.162688,15.565851,18.055782,21.073883,25.800982,26.838455,27.230806,26.148064,24.09953,22.911152,23.303505,22.726294,23.303505,25.518036,28.1966,29.626425,30.184772,29.943325,28.985079,27.404348,26.962952,26.763002,26.653595,26.566826,26.498919,26.845999,26.219744,25.763256,25.785892,25.759483,24.193844,24.17121,24.959686,26.265015,28.256962,29.034122,30.056503,31.614597,33.70086,36.013477,38.62036,37.89979,36.65105,36.31906,37.00568,41.770504,45.45636,43.781315,37.216946,31.022295,26.872408,23.231825,21.851044,22.571615,23.31105,24.182526,24.92196,25.819845,26.97804,28.306005,30.011232,32.516254,32.61057,30.56958,30.143274,29.139755,29.822601,30.690304,31.063795,31.067568,30.101774,27.947605,26.182018,25.284132,24.623924,22.858335,20.504217,19.678013,21.549234,26.351786,31.071339,36.60201,43.426685,49.244076,48.99885,43.79263,40.699078,38.454365,36.13043,33.138737,35.055233,36.824593,36.503918,35.06655,36.398285,36.168156,37.19431,35.38345,30.02255,23.775084,19.806282,15.46399,11.714001,9.291975,8.695901,10.303039,7.333983,5.0477724,5.1232247,5.6325293,6.7756343,8.329956,8.526133,8.058327,10.069136,10.008774,10.461489,10.518079,9.616421,7.5301595,6.013564,4.38379,4.1989317,5.3609,6.1342883,7.6810646,8.922258,9.216523,8.846806,9.031664,9.314611,6.3945994,4.002755,3.150142,2.1088974,1.3015556,1.1431054,1.6071383,1.901403,0.45648763,0.47157812,0.42630664,0.271629,0.10940613,0.17354076,0.28294688,0.49044126,0.6149379,0.6073926,0.5394854,2.584248,3.1425967,4.093298,6.0776987,8.503497,7.4169807,6.6020937,7.9791017,11.498961,15.131999,17.757746,15.98084,13.422999,11.242422,8.130007,7.9526935,7.7187905,7.5301595,7.5075235,7.7942433,6.5832305,5.9532022,5.9532022,6.0814714,5.292993,4.5535583,3.85185,3.308592,3.0746894,3.3010468,2.837014,2.6823363,3.0897799,3.482133,2.4484336,2.2711203,1.690136,1.0487897,0.7394345,1.2223305,2.7540162,2.9916916,4.3875628,7.2623034,9.812597,10.227587,9.669238,5.9532022,0.9620194,0.62625575,0.20749438,0.30935526,0.43385187,0.42630664,0.4640329,0.35462674,0.3470815,0.2565385,0.23767537,0.76584285,0.76584285,0.8526133,1.1280149,1.3996439,1.1846043,1.0148361,0.995973,0.98842776,1.0110635,1.2261031,0.95447415,1.3053282,1.7882242,2.0787163,2.0108092,1.7354075,1.4637785,1.1657411,0.9318384,0.965792,0.62625575,0.422534,0.35085413,0.36594462,0.38103512,0.45648763,0.47157812,0.47535074,0.55080324,0.80734175,1.5241405,2.5540671,3.8556228,4.8063245,4.191386,4.425289,4.659192,4.285702,3.663219,4.123479,3.8858037,4.195159,4.221567,4.0706625,4.8138695,4.2291126,3.289729,2.5578396,2.233394,2.1805773,2.3654358,2.052308,2.214531,3.0671442,4.074435,4.3422914,4.689373,4.6629643,4.3385186,4.3196554,4.534695,4.466788,4.504514,4.8063245,5.292993,5.2326307,4.9685473,4.6252384,4.376245,4.4177437,4.504514,3.7235808,3.380272,3.6783094,3.6971724,4.3875628,4.2404304,4.1310244,4.7308717,6.4738245,6.6322746,6.63982,6.379509,5.8890676,5.372218,5.7192993,6.5643673,7.6923823,8.744945,9.208978,10.186088,9.639057,8.405409,7.2585306,6.9265394,7.1340337,7.1378064,7.2585306,7.665974,8.390318,7.865923,8.103599,7.809334,6.9491754,6.7643166,6.911449,6.911449,6.911449,7.1679873,8.069645,9.476834,9.22784,9.548513,14.418973,29.57738,26.219744,20.289177,14.241659,8.990166,3.9008942,6.8246784,8.254503,8.186596,7.1906233,6.4134626,4.142342,5.802297,11.725319,17.429527,13.63804,11.087745,9.876732,10.144588,11.200924,11.506506,10.751981,11.053791,11.242422,10.933067,10.49167,10.819888,11.00852,10.906659,10.868933,11.774363,11.329193,11.034928,10.310584,9.416472,9.454198,10.099318,9.793735,9.673011,9.891823,9.64283,10.676529,11.076427,10.868933,10.480352,10.714255,10.287949,10.231359,10.657665,11.404645,12.045992,11.861133,12.245941,12.725064,12.694883,11.431054,10.536942,10.005001,9.224068,8.254503,7.8206515,8.571404,9.382519,9.748463,9.556059,9.0957985,8.284684,7.5716586,6.7077274,5.907931,5.8513412,4.7233267,4.508287,4.9647746,5.674028,6.039973,6.19465,6.6850915,6.7379084,6.3116016,6.0814714,5.330719,4.504514,3.8443048,3.4632697,3.3274553,3.0218725,2.5276587,2.3277097,2.535204,2.916239,2.8030603,2.7917426,3.2972744,4.3611546,5.6363015,6.3229194,6.692637,6.779407,6.458734,5.451443,5.040227,4.666737,4.534695,4.5535583,4.3649273,4.123479,4.134797,4.3800178,4.878004,5.7079816,5.247721,4.214022,3.6066296,3.610402,3.5839937,3.4934506,3.0558262,2.4786146,1.9768555,1.7769064,1.3128735,1.1544232,1.0450171,1.0412445,1.5015048,1.4335974,1.3430545,1.2789198,1.267602,1.327964,1.9957186,2.7502437,3.1916409,3.3425457,3.6330378,3.7084904,3.783943,4.0216184,4.406426,4.7346444,4.8138695,4.247976,3.8367596,3.6745367,3.169005,3.3274553,3.7990334,4.5912848,5.5004873,6.1003346,6.296511,7.115171,7.854605,8.073418,7.605612,7.2358947,6.8963585,6.5266414,6.307829,6.673774,6.5040054,5.798525,5.168496,4.8138695,4.4894238,4.6856003,5.0553174,5.43258,5.692891,5.753253,5.9117036,6.4134626,6.760544,6.8774953,7.115171,8.118689,9.159933,9.265567,8.254503,6.7152724,7.6282477,8.103599,7.699928,6.937857,7.2924843,7.152897,7.1868505,7.254758,7.2057137,6.8737226,6.779407,6.651138,6.911449,7.643338,8.620448,2.1353056,2.3201644,2.5012503,2.8445592,3.127506,2.7615614,2.4182527,2.2899833,2.323937,2.4522061,2.546522,2.6219745,2.4295704,2.2748928,2.2598023,2.2598023,2.5389767,2.9011486,3.2935016,3.5462675,3.3878171,3.7914882,4.255521,4.5309224,4.7610526,5.492942,5.8966126,5.5495315,5.7192993,6.620957,7.4169807,10.148361,13.679539,17.580433,21.1267,23.284641,20.074137,23.337458,27.415667,25.978296,12.038446,5.9003854,3.8141239,3.0445085,2.3126192,1.7995421,1.3241913,0.9016574,0.8224323,0.9808825,0.8865669,0.90920264,0.80734175,0.5998474,0.3772625,0.3055826,0.3169005,0.38480774,0.40367088,0.38480774,0.45648763,0.45648763,0.59607476,0.814887,0.965792,0.80734175,0.68661773,1.0940613,1.4373702,1.5430037,1.6637276,1.8825399,2.2107582,2.2598023,2.052308,2.0145817,1.9542197,2.0560806,2.5691576,3.4594972,4.425289,4.327201,3.7462165,2.957738,2.1654868,1.478869,1.1732863,0.66775465,0.3772625,0.41121614,0.59607476,0.29049212,0.18485862,0.21503963,0.30181,0.35085413,0.52062225,0.4640329,0.36594462,0.331991,0.38103512,0.5281675,1.6260014,2.425798,2.4371157,1.9240388,2.3880715,3.308592,3.9197574,4.06689,4.22534,3.410453,2.7087448,2.173032,2.052308,2.806833,3.1614597,2.7011995,2.0372176,1.4147344,0.7167987,0.754525,1.3204187,1.5165952,1.2449663,1.2223305,0.73188925,1.20724,2.1805773,3.187868,3.7386713,4.3007927,5.3382645,5.564622,5.142088,5.692891,6.485142,7.115171,7.454707,7.677292,8.239413,10.167224,10.642575,11.838497,13.309821,11.978085,13.45318,13.72481,13.2607765,12.464753,11.657412,11.98563,11.091517,9.465516,8.756263,11.732863,11.781908,12.336484,11.714001,10.687846,12.479843,11.027383,11.974312,12.351574,11.661184,11.857361,11.917723,12.608112,12.6345215,12.193124,13.000465,13.890805,13.373956,12.989148,12.826925,11.521597,11.921495,11.649866,11.329193,11.41219,12.14408,13.6833105,15.769572,18.13878,21.187061,25.985842,26.729048,26.649822,25.05023,22.726294,21.956678,23.726038,23.978804,24.654104,26.47251,28.917171,32.07863,33.059513,32.331398,30.418674,27.894789,26.808273,27.14781,28.1966,29.026577,28.487091,28.279596,27.064812,26.58946,26.944088,26.566826,25.61235,24.220253,24.12971,25.936796,29.098257,31.965452,32.68225,33.021786,34.025307,36.024796,39.540882,40.476494,40.061504,39.09194,37.933743,39.09194,42.347717,43.336143,40.28409,34.010216,27.725021,23.12242,20.836208,20.65135,21.53037,23.593996,24.842735,25.982069,27.170444,28.000423,29.109575,29.928234,30.403585,30.033867,27.845745,25.721758,26.70264,27.989105,28.404093,28.381458,26.525326,24.525835,23.005466,22.428255,23.088465,20.500444,16.893814,15.931795,17.708702,18.7839,23.97126,29.56229,37.356533,44.920647,45.592175,39.635197,35.145775,32.9237,32.23708,30.807257,35.40986,40.778305,41.34797,36.91136,32.63698,33.138737,32.433258,30.924208,28.32487,23.650587,19.24416,14.754736,11.042474,8.488406,6.9869013,6.7680893,5.451443,4.187614,3.6669915,4.1197066,6.952948,6.7077274,6.1342883,6.9567204,9.88805,10.303039,11.065109,11.185833,10.216269,8.239413,6.3116016,4.8855495,4.5422406,5.304311,6.620957,8.356364,8.14887,7.466025,7.0170827,6.760544,8.088508,5.5759397,2.9954643,1.8146327,1.20724,0.7432071,0.6526641,0.6828451,0.7469798,0.9318384,1.4071891,0.98465514,0.4376245,0.18485862,0.32067314,0.18485862,0.27917424,0.41498876,0.51684964,0.62625575,2.3956168,2.674791,3.983892,6.964266,10.344538,10.235131,6.903904,5.983383,8.89585,12.864652,13.875714,13.023102,11.732863,10.570895,9.216523,10.193633,9.740918,9.009028,8.318638,7.17176,7.6093845,7.3717093,6.270103,4.9760923,5.036454,5.304311,4.7836885,4.2064767,3.802806,3.3274553,2.897376,2.4182527,1.9391292,1.5203679,1.1921495,2.3993895,2.1164427,1.4675511,1.1242423,1.297783,2.5540671,2.6597006,4.214022,6.651138,6.2097406,7.956466,6.5341864,3.3161373,0.30935526,0.1358145,0.150905,0.08677038,0.10186087,0.32821837,0.91674787,0.573439,0.5055317,0.52062225,0.5470306,0.65643674,0.5583485,0.97333723,1.4939595,1.7467253,1.4034165,1.478869,1.539231,1.1921495,0.76207024,1.3128735,1.5203679,1.5241405,1.6712729,1.8900851,1.6939086,1.4373702,2.161714,2.11267,1.1581959,0.7922512,0.7205714,0.4640329,0.3470815,0.45648763,0.62625575,0.6149379,0.482896,0.452715,0.5772116,0.7469798,1.8825399,2.7615614,3.8292143,4.798779,4.6554193,5.6778007,5.824933,5.0025005,4.014073,4.561104,4.063117,4.870459,5.036454,4.398881,4.606375,4.0103,3.0181,2.5314314,2.6446102,2.655928,2.5087957,2.3993895,2.837014,3.7198083,4.3196554,4.587512,5.0213637,4.9345937,4.3686996,4.0895257,4.52715,4.3913355,4.214022,4.2328854,4.3800178,4.9044123,4.9534564,4.6856003,4.3913355,4.5007415,4.172523,3.429316,2.9652832,2.927557,2.916239,4.036709,3.9159849,3.8669407,4.557331,5.9984736,5.4212623,5.4174895,5.379763,4.930821,3.904667,4.8100967,5.5306683,6.511551,7.575431,7.9036493,9.258021,8.948667,7.756517,6.696409,6.9869013,6.4134626,7.0963078,7.6923823,7.7904706,7.888559,7.960239,8.062099,8.337502,8.265821,6.6662283,6.6058664,6.6360474,6.971811,7.273621,6.651138,10.914205,8.424272,8.60913,16.014793,30.335678,30.592216,26.61587,19.768555,12.140307,6.560595,7.3679366,6.9265394,6.432326,6.7944975,8.635539,8.073418,6.541732,9.631512,15.946886,17.105082,17.591751,11.0613365,7.4471617,9.163706,11.091517,10.201178,11.389555,12.053536,11.408418,10.469034,10.552032,10.774617,10.518079,10.137043,10.955703,10.49167,10.450171,10.193633,9.673011,9.431562,10.212496,9.767326,9.57115,9.861642,9.64283,10.948157,11.431054,11.114153,10.627484,11.216014,10.884023,10.657665,10.612394,10.899114,11.7026825,12.0082655,12.257258,12.593022,12.725064,11.932813,10.736891,10.638803,10.076681,8.956212,8.650629,8.884532,9.608876,10.435081,10.608622,9.031664,7.960239,7.0849895,6.379509,5.802297,5.3269467,4.323428,4.266839,4.7421894,5.3080835,5.4778514,5.674028,5.8136153,6.0324273,6.349328,6.6662283,5.7419353,4.7308717,3.953711,3.4481792,2.9615107,2.6068838,2.4522061,2.4408884,2.5767028,2.9313297,2.795515,2.9992368,3.531177,4.5497856,6.3945994,6.7944975,6.8963585,6.8435416,6.511551,5.523123,4.889322,4.3007927,3.8669407,3.682082,3.8141239,3.8895764,4.115934,4.5497856,5.1345425,5.723072,4.719554,3.6934,3.4481792,3.7198083,3.1576872,3.3312278,3.2067313,2.565385,1.7165444,1.4939595,1.2864652,1.1996948,1.3656902,1.780679,2.3201644,1.7316349,1.478869,1.4939595,1.6561824,1.7542707,2.8407867,3.240685,3.429316,3.6330378,3.8292143,4.014073,4.432834,4.8440504,5.040227,4.881777,4.5912848,4.123479,3.9348478,4.0103,3.874486,4.1800685,4.8063245,5.5080323,6.187105,6.881268,7.333983,7.7376537,8.080963,8.152642,7.567886,6.5568223,6.530414,6.628502,6.6850915,7.2472124,7.1868505,6.1078796,5.292993,5.0741806,4.8666863,4.6252384,4.881777,5.3344917,5.753253,5.9984736,5.9117036,6.2663302,6.6813188,7.141579,7.9941926,8.75249,9.1976595,8.854351,7.8508325,6.911449,8.009283,8.586494,8.405409,7.7187905,7.277394,6.971811,7.1793056,7.6207023,7.9753294,7.888559,7.594294,7.496206,8.152642,9.4127,10.38981,2.3088465,2.354118,2.3993895,2.4484336,2.4371157,2.2371666,2.1088974,2.1277604,2.1579416,2.161714,2.1805773,2.372981,2.2899833,2.2786655,2.474842,2.806833,2.9992368,3.5085413,3.9574835,4.085753,3.742444,3.7650797,4.2064767,4.6290107,4.90064,5.2137675,6.1041074,5.8173876,5.983383,6.8397694,7.232122,9.039209,11.962994,15.98084,19.36111,18.670721,15.354584,21.107838,26.815819,25.910389,14.369928,9.352338,6.224831,4.112161,2.6031113,1.7391801,1.2449663,0.98465514,0.98465514,1.056335,0.8111144,0.814887,0.72811663,0.5998474,0.48666862,0.452715,0.452715,0.47535074,0.40367088,0.2867195,0.31312788,0.30181,0.49421388,0.7205714,0.7884786,0.5017591,0.6752999,1.3694628,1.7919968,1.9429018,2.6031113,2.3918443,2.704972,3.2218218,3.8405323,4.6629643,4.425289,4.214022,4.315883,4.9534564,6.2663302,5.8890676,5.05909,4.164978,3.2746384,2.1503963,1.2298758,0.63002837,0.47157812,0.5696664,0.41121614,0.26408374,0.38103512,0.41121614,0.27540162,0.1659955,0.3961256,0.38480774,0.32821837,0.32821837,0.35839936,0.3169005,0.6375736,1.0336993,1.4298248,1.9730829,2.5804756,3.3123648,3.5424948,3.1048703,2.2862108,1.6939086,1.327964,1.3807807,1.7278622,1.9164935,1.6260014,1.3996439,1.2864652,1.1846043,0.8526133,1.0035182,0.8903395,0.7394345,0.663982,0.66020936,0.66020936,1.1506506,1.9127209,2.806833,3.7877154,4.357382,4.9949555,5.1873593,4.9723196,4.9459114,6.1418333,7.273621,8.167733,8.99771,10.291721,10.499215,10.435081,11.016065,12.121444,12.577931,13.487134,14.456699,14.784918,14.490653,14.317112,13.807808,13.373956,12.494934,11.962994,13.905896,11.69891,11.400873,11.7894535,12.404391,13.543724,14.139798,12.774108,12.091263,12.249713,10.902886,12.498707,13.019329,13.641812,14.302021,13.671993,14.211478,14.373701,14.132254,13.63804,13.241914,13.000465,12.913695,13.068373,13.70972,15.271586,14.396337,16.094019,18.402864,20.440083,22.398075,23.84299,24.755966,24.891779,24.435291,23.959942,25.661396,26.698868,28.030603,29.856554,31.625916,33.195328,34.930737,35.047688,33.915897,34.044167,32.29367,31.51651,31.1732,30.961933,30.8563,30.520536,29.422703,28.192827,27.442074,27.73634,27.95515,26.280106,24.85028,25.072866,27.60807,28.377686,29.61888,30.335678,30.973251,33.425457,37.175446,36.930225,37.59798,40.13696,41.54792,40.978252,40.336906,40.01623,39.42016,36.95286,31.622143,27.66466,24.623924,22.711203,22.797974,24.190071,25.8123,26.800728,27.476028,29.332159,30.618624,29.73583,29.135983,28.754948,26.004704,22.816835,22.797974,23.80149,24.525835,24.499426,23.87317,22.598024,21.390783,20.587215,20.1345,17.87847,14.830189,13.65313,14.335975,14.219024,19.798737,28.472,34.75342,37.00568,37.462166,34.77983,31.799456,28.879444,26.917679,27.366621,34.213936,43.51346,46.886185,42.687252,36.03234,31.69005,28.189054,26.016022,24.56356,22.111355,18.742401,14.517061,11.091517,8.89585,7.17176,6.85486,4.779916,2.987919,2.546522,3.5349495,7.537705,6.7454534,5.983383,7.303802,9.948412,10.812344,12.347801,12.551523,11.02361,8.959985,6.85486,5.583485,5.3382645,5.881522,6.5228686,7.484888,6.8963585,6.2361493,5.9796104,5.5759397,6.828451,4.961002,2.5993385,1.1204696,0.65643674,0.44516975,0.67152727,0.8903395,0.9620194,1.0299267,1.5430037,1.5920477,1.3732355,1.0789708,0.91674787,0.66775465,0.52062225,0.5017591,0.58475685,0.68661773,1.3241913,1.9051756,2.9464202,4.3611546,5.4250345,7.99042,9.869187,10.080454,9.190115,9.2995205,11.91395,11.627231,11.32542,11.295239,9.22784,8.624221,8.948667,8.284684,6.741681,6.462507,6.7077274,6.304056,5.798525,5.5985756,5.96452,5.9682927,5.4212623,5.191132,5.0439997,3.6330378,2.795515,2.0485353,1.5920477,1.5165952,1.7995421,1.7316349,1.5958204,1.0751982,0.5583485,1.1506506,1.9768555,3.4972234,5.9532022,7.224577,2.8294687,2.9539654,2.5691576,1.5241405,0.38480774,0.41876137,0.10940613,0.19240387,0.1961765,0.21503963,0.9280658,1.1431054,0.8186596,0.5583485,0.5885295,0.76584285,0.9695646,1.0299267,1.2902378,1.5580941,1.0978339,1.2487389,1.7354075,1.7391801,1.3732355,1.6788181,1.3204187,1.2789198,1.2940104,1.3317367,1.5958204,1.6524098,1.8033148,1.7580433,1.5279131,1.4147344,0.73566186,0.452715,0.36594462,0.41498876,0.6752999,0.67152727,0.5281675,0.51684964,0.6526641,0.68661773,1.2147852,2.1353056,3.5047686,4.6290107,4.044254,5.353355,5.87775,5.3948536,4.4139714,4.172523,3.7877154,4.617693,5.13077,4.8365054,4.304565,3.470815,2.7917426,2.4899325,2.565385,2.8143783,2.704972,2.9049213,3.4594972,4.164978,4.587512,5.2175403,5.5268955,5.0213637,3.9612563,3.3576362,3.8367596,3.6330378,3.4972234,3.7084904,4.112161,5.221313,5.330719,4.9534564,4.5535583,4.52715,3.874486,3.4179983,3.0369632,2.7841973,2.8898308,3.8858037,3.7084904,3.451952,3.7047176,4.568649,4.5309224,4.45547,4.29702,4.08198,3.904667,4.564876,4.776143,5.4740787,6.5530496,6.8925858,8.394091,8.586494,7.7187905,6.72659,7.232122,7.175533,7.224577,6.911449,6.7567716,8.29223,8.167733,8.118689,8.224322,7.914967,5.983383,7.1340337,7.3490734,7.5301595,8.069645,8.8618965,11.080199,9.190115,12.4307995,22.096264,31.531599,25.027594,21.719002,14.434063,4.9647746,4.032936,7.0170827,8.243186,8.880759,9.408927,9.612649,7.0284004,5.1232247,6.009792,10.133271,16.263786,17.297485,17.727566,13.63804,7.8961043,10.1294985,10.0276375,10.585986,11.61214,12.2270775,10.846297,10.676529,11.348056,11.125471,10.246449,10.917976,10.834979,10.831206,10.740664,10.325675,9.273112,10.1294985,9.786189,9.627739,10.038955,10.374719,11.057564,11.234878,10.933067,10.63503,11.299012,11.695138,11.234878,11.151879,11.54046,11.348056,12.064855,11.706455,11.423509,11.3820095,10.785934,10.506761,10.740664,10.7218,10.340765,10.152134,9.857869,9.850324,9.748463,9.258021,8.190369,7.9753294,6.952948,6.115425,5.9305663,6.3153744,5.311856,4.749735,4.447925,4.3686996,4.5988297,4.9987283,5.2062225,5.6363015,6.1795597,6.205968,5.541986,4.7648253,4.093298,3.5839937,3.1539145,2.7238352,2.4559789,2.516341,2.8747404,3.2972744,3.3274553,3.6669915,3.9650288,4.5120597,6.258785,6.8850408,7.352846,7.6508837,7.356619,5.5985756,4.708236,3.8367596,3.4896781,3.5990841,3.5085413,4.2291126,4.45547,4.8402777,5.342037,5.2326307,4.496969,3.9876647,3.7914882,3.7688525,3.5500402,3.0445085,2.595566,2.093807,1.5769572,1.2034674,1.1883769,1.8033148,2.3880715,2.5502944,2.1466236,1.9353566,1.8636768,1.961765,2.2069857,2.546522,2.8747404,3.4029078,3.983892,4.376245,4.2706113,4.666737,4.6290107,4.776143,5.0025005,4.4931965,4.217795,3.6330378,3.2444575,3.3312278,3.9499383,4.293247,5.2665844,6.356873,7.152897,7.322665,8.103599,8.624221,8.650629,8.209232,7.54525,7.5075235,7.99042,8.243186,7.997965,7.454707,8.458225,8.27714,7.6886096,7.2396674,7.2472124,7.5112963,7.84706,7.756517,7.273621,6.960493,7.4207535,8.578949,9.65792,10.163452,9.876732,10.416218,10.3634,9.393836,7.9413757,7.1566696,8.5563135,9.673011,10.023865,9.424017,7.9489207,8.084735,8.6581745,9.22784,9.461743,9.122208,8.907167,8.66572,9.088254,10.167224,11.185833,2.4974778,2.6710186,2.6219745,2.4408884,2.2409391,2.1805773,2.1994405,2.1466236,2.1353056,2.1503963,2.0636258,2.11267,2.1768045,2.3013012,2.5125682,2.8181508,3.0407357,3.361409,3.591539,3.6481283,3.5651307,3.5953116,4.0593443,4.6856003,5.198677,5.3269467,5.6363015,5.8173876,6.2889657,7.0057645,7.4509344,9.891823,12.649611,15.384765,17.123945,16.252468,15.290449,22.043447,26.755457,24.17498,13.551269,8.763808,5.621211,3.5274043,2.161714,1.448688,1.3732355,1.3468271,1.2487389,1.0638802,0.8865669,0.90543,0.814887,0.66775465,0.5281675,0.452715,0.36971724,0.3169005,0.2678564,0.271629,0.422534,0.513077,0.65643674,0.73566186,0.69793564,0.55457586,0.8563859,1.3468271,1.6033657,1.7240896,2.323937,2.6672459,3.138824,3.4972234,3.7198083,3.9876647,3.663219,3.4330888,3.5462675,3.92353,4.183841,3.4029078,2.6597006,2.11267,1.720317,1.2562841,0.77716076,0.52062225,0.41121614,0.362172,0.26408374,0.24899325,0.3772625,0.42630664,0.32821837,0.15845025,0.27917424,0.27540162,0.25276586,0.2565385,0.2867195,0.47157812,0.7054809,1.0487897,1.4637785,1.81086,1.7391801,1.8900851,1.7882242,1.3619176,0.95824677,0.845068,0.754525,0.87902164,1.1581959,1.2713746,1.0827434,1.2298758,1.3091009,1.1619685,0.8563859,0.9808825,0.8262049,0.6790725,0.6413463,0.6111652,0.66020936,0.94692886,1.991946,3.4142256,3.9386206,2.9501927,3.7009451,4.779916,5.4174895,5.511805,6.960493,8.262049,10.080454,12.08749,12.96274,11.046246,11.16697,11.646093,11.947904,12.687338,12.381755,13.856852,14.268067,13.611631,14.728328,15.297995,16.218515,16.033657,14.864142,14.441608,14.373701,14.456699,14.720782,14.743419,13.65313,13.283413,13.422999,13.592768,13.411682,12.570387,13.223051,14.109617,14.924504,15.218769,14.396337,15.199906,15.614895,15.682802,15.30554,14.237886,13.287186,13.679539,14.78869,15.920478,16.290195,16.078928,17.825653,20.43631,22.40562,21.820864,22.53389,24.657877,25.880207,25.767029,25.759483,27.687294,28.377686,29.332159,30.91289,32.357803,32.59925,34.244118,35.549446,36.115337,36.900043,33.97626,32.440804,31.463692,30.91289,31.376923,31.478783,31.34674,30.56958,29.467974,29.109575,29.366114,28.739857,28.294687,28.351276,28.490864,27.740112,28.147554,28.653088,29.03035,29.875418,32.5238,34.45161,36.047432,37.52253,38.90708,40.272774,41.872364,41.238564,38.431732,36.05875,33.34246,31.324106,30.067822,29.215208,27.970242,27.343987,27.351532,27.826881,28.71345,30.048958,31.788137,31.226017,30.162136,28.954897,26.532871,24.152346,22.050993,20.772074,20.745665,22.266033,21.009748,19.696875,18.485863,17.41821,16.399601,15.071637,13.060828,12.079946,12.313848,12.427027,17.599297,25.253952,30.66767,32.274807,31.705141,28.871899,26.895044,25.031366,23.748674,24.737103,32.357803,43.38896,51.09643,50.711624,39.42393,29.80751,25.597261,23.450638,21.511507,19.429018,17.380484,14.962231,12.310076,9.756008,7.8131065,6.8246784,5.0439997,3.7688525,3.3764994,3.3123648,5.8400235,5.7683434,5.8211603,7.092535,9.039209,10.718028,12.936331,13.264549,11.472552,9.525878,7.537705,6.2021956,5.8437963,6.19465,6.40969,7.073672,6.439871,5.745708,5.3646727,4.7836885,5.885295,4.7346444,2.6672459,0.86770374,0.392353,0.21503963,0.3055826,0.452715,0.5998474,0.8337501,1.1317875,1.4109617,1.780679,2.1692593,2.3390274,1.569412,1.3204187,1.0638802,0.7167987,0.6451189,1.8523588,3.240685,4.9949555,6.5002327,6.375736,6.790725,9.035437,9.627739,8.194141,7.466025,8.480861,9.265567,10.295494,10.567122,7.6093845,7.6810646,7.7037,7.6131573,7.432071,7.273621,7.0548086,6.300284,5.926794,6.1833324,6.651138,6.0512905,5.6098933,5.1156793,4.2894745,2.8030603,2.2786655,2.0372176,2.2258487,2.7426984,3.2255943,1.9844007,1.2298758,0.65643674,0.452715,1.2789198,2.173032,2.8445592,5.168496,7.492433,4.6290107,2.2183034,1.4826416,1.2487389,1.0412445,1.0827434,0.44516975,0.6790725,0.7167987,0.4376245,0.694163,1.2449663,1.2147852,0.95824677,0.8186596,1.1317875,1.1431054,1.5920477,1.9202662,1.931584,1.7995421,1.6712729,1.5279131,1.6033657,1.8863125,2.1466236,1.418507,1.3807807,1.478869,1.4750963,1.4335974,1.6788181,1.9429018,2.052308,1.931584,1.5882751,0.935611,0.58475685,0.44139713,0.49421388,0.84129536,0.94315624,0.7432071,0.6073926,0.69793564,0.95447415,1.1808317,1.9466745,3.3840446,4.7006907,4.2027044,5.5080323,5.8173876,5.3948536,4.6214657,3.9914372,3.712263,4.6327834,5.349582,5.300538,4.7572803,3.8443048,3.3878171,3.1010978,2.9011486,2.9351022,3.1463692,3.4934506,3.8971217,4.304565,4.727099,5.1760416,5.349582,4.7535076,3.6066296,2.8256962,3.2859564,3.187868,3.0822346,3.2029586,3.4859054,5.191132,5.270357,4.5950575,3.9688015,4.1272516,3.7914882,3.561358,3.240685,2.9426475,3.0746894,4.063117,4.1197066,3.8443048,3.610402,3.5689032,3.5160866,3.4594972,3.3425457,3.4368613,4.3347464,4.2404304,4.195159,4.5837393,5.281675,5.666483,7.0510364,7.6131573,7.533932,7.1264887,6.85486,6.722818,6.56814,6.0286546,5.926794,8.265821,7.865923,7.567886,7.8734684,7.964011,5.6853456,7.3415284,7.224577,7.220804,8.001738,9.001483,9.789962,9.322156,11.3820095,17.652113,27.721249,29.36234,22.266033,12.494934,4.957229,3.4029078,6.9454026,9.14107,9.495697,8.786444,9.061845,7.964011,6.2323766,5.292993,6.326692,10.257768,13.539951,16.67123,14.750964,9.680555,10.125726,10.457717,10.438853,10.899114,11.781908,12.140307,10.925522,11.117926,10.744436,9.846551,10.487898,10.985884,10.884023,10.533169,10.03141,9.224068,10.20495,10.465261,10.589758,10.887795,11.393328,10.834979,10.944386,11.200924,11.332966,11.348056,10.79348,10.457717,10.842525,11.581959,11.442371,12.151625,11.759273,11.299012,11.046246,10.499215,10.163452,10.465261,10.702937,10.653893,10.574668,10.423763,9.948412,9.310839,8.605357,7.8696957,7.752744,7.1340337,6.537959,6.1531515,5.828706,5.3684454,4.8365054,4.478106,4.447925,4.798779,4.9949555,5.2099953,5.764571,6.304056,5.7872066,4.7044635,4.0706625,3.5575855,3.0897799,2.8294687,2.6936543,2.425798,2.4710693,2.8294687,3.059599,3.4745877,3.9084394,4.285702,4.9459114,6.647365,6.6360474,7.2924843,7.8696957,7.6886096,6.138061,5.1647234,4.2027044,3.8669407,4.063117,4.0103,4.6554193,4.738417,4.9949555,5.247721,4.3875628,4.032936,3.863168,3.7575345,3.682082,3.7009451,3.1614597,2.4786146,1.8863125,1.4600059,1.1204696,1.720317,2.625747,3.0331905,2.6597006,1.7391801,2.1503963,2.2296214,2.2786655,2.4974778,3.0030096,3.187868,3.3689542,3.7877154,4.376245,4.772371,5.093044,5.172269,5.2665844,5.2892203,4.8063245,4.236658,3.4632697,3.187868,3.663219,4.67051,4.8855495,5.674028,6.7831798,7.805561,8.16396,8.394091,8.635539,8.548768,8.013056,7.164215,7.069899,8.013056,8.654402,8.624221,8.495952,9.363655,9.480607,9.363655,9.156161,8.631766,8.729855,9.307066,9.359882,8.710991,7.9791017,8.050782,8.959985,10.061591,10.79348,10.665211,11.174516,10.967021,10.038955,8.9788475,8.975075,10.20495,10.774617,10.759526,10.103089,8.612903,8.986393,9.582467,10.016319,10.250222,10.56335,10.653893,10.33322,10.314357,10.872705,11.830952,2.4107075,2.6144292,2.5389767,2.3088465,2.1051247,2.1466236,2.282438,2.1541688,2.1654868,2.3126192,2.214531,2.1013522,2.214531,2.4597516,2.6710186,2.6219745,2.7087448,2.8747404,2.9992368,3.1312788,3.4896781,3.863168,4.327201,4.927048,5.492942,5.6476197,5.523123,6.175787,6.8473144,7.443389,8.526133,11.649866,14.011529,15.878979,16.840998,15.803526,16.867407,23.639269,26.44233,21.68505,11.849815,7.2924843,4.346064,2.5691576,1.6373192,1.3468271,1.5920477,1.5958204,1.3732355,1.0525624,0.90920264,0.995973,0.91297525,0.724344,0.52062225,0.41498876,0.27917424,0.19994913,0.2263575,0.35462674,0.543258,0.7130261,0.784706,0.70170826,0.573439,0.70170826,1.0827434,1.358145,1.5052774,1.6524098,2.082489,2.7351532,3.0935526,3.029418,2.6785638,2.425798,2.1277604,2.123988,2.4974778,2.8521044,2.2975287,1.3204187,0.7394345,0.5093044,0.52439487,0.63002837,0.5470306,0.5357128,0.4640329,0.32067314,0.21503963,0.24522063,0.2867195,0.31312788,0.29803738,0.2263575,0.23767537,0.24522063,0.23013012,0.22258487,0.31312788,0.58098423,0.754525,0.9808825,1.2298758,1.297783,0.995973,0.98465514,0.8563859,0.55080324,0.34330887,0.5319401,0.63002837,0.8111144,1.1280149,1.5165952,1.569412,1.6712729,1.5807298,1.2600567,0.9016574,0.98465514,0.9318384,0.8337501,0.754525,0.70170826,0.73566186,0.8601585,1.6675003,2.7841973,2.8936033,1.750498,2.6446102,3.9008942,4.67051,4.949684,6.228604,7.748972,10.080454,12.351574,12.257258,10.601076,10.759526,11.631002,12.510024,13.060828,13.087236,13.502225,13.773854,14.003984,14.954685,16.373192,17.663431,17.674747,16.535416,15.667711,17.342756,17.863379,17.772837,17.33144,16.486372,14.551015,16.014793,16.950403,16.13929,15.052773,14.079436,14.222796,14.588741,14.667966,14.354838,15.871433,16.237377,16.350557,16.173243,14.750964,14.460471,15.150862,16.350557,17.557796,18.248188,18.821627,20.300495,22.337713,23.978804,23.669449,23.914669,25.944342,27.159128,27.343987,28.683268,30.116865,29.969732,29.826374,30.403585,31.565554,30.950615,32.025814,33.697086,35.183502,36.024796,33.96117,32.557755,31.54669,30.99966,31.309015,31.807001,32.27858,32.274807,31.765503,31.161882,31.222244,31.972998,32.878426,33.45941,33.282097,31.37315,30.678986,30.230043,29.660378,29.20389,30.550716,32.761475,33.48582,32.901062,33.723495,37.979015,42.849476,43.811493,40.336906,35.9003,34.26298,33.78763,35.71167,38.77504,39.223984,35.09673,31.803228,30.584671,31.20338,31.901318,32.429485,32.195583,30.931753,28.977533,27.29494,25.453901,22.341486,19.806282,18.878216,19.798737,18.395319,17.41821,16.063837,14.339747,13.072145,12.408164,11.664956,11.287694,11.427281,11.940358,16.444872,22.315077,26.261242,27.113855,25.808527,23.458181,22.748928,22.548979,22.92247,25.12191,31.837183,41.487556,51.44729,55.612267,44.42266,31.15811,26.004704,23.4695,20.930523,18.644312,17.093763,15.663939,13.287186,10.054046,7.183078,6.3719635,5.1835866,4.293247,3.7952607,3.199186,4.134797,4.5724216,5.243949,6.405917,7.816879,10.370946,13.011784,13.570132,11.92904,10.03141,8.288457,6.8774953,6.3832817,6.6134114,6.590776,7.17176,6.7869525,6.013564,5.2250857,4.5950575,5.270357,4.9685473,3.218049,0.9242931,0.34330887,0.120724,0.10940613,0.35462674,0.7884786,1.2411937,1.3053282,1.6863633,2.3993895,3.2972744,4.06689,3.561358,3.3840446,2.6974268,1.8033148,2.161714,3.1237335,4.7421894,7.2396674,9.318384,8.122461,6.168242,6.039973,6.4511886,6.466279,5.492942,5.2288585,6.6813188,8.382772,8.801534,6.3153744,7.0548086,7.062354,7.405663,7.997965,7.594294,7.352846,6.5266414,6.2927384,6.7944975,7.145352,5.798525,5.3646727,4.7912335,3.7914882,2.8521044,2.6823363,2.6597006,2.7351532,2.8747404,3.048281,1.7844516,1.086516,0.8262049,1.0601076,1.9994912,2.3201644,1.9089483,3.3350005,5.764571,4.9459114,2.5502944,1.599593,1.2902378,1.2147852,1.3392819,0.84129536,1.0336993,1.0336993,0.7469798,0.8337501,1.056335,1.2034674,1.1619685,1.0450171,1.1921495,1.4373702,1.9655377,2.2598023,2.2069857,2.0862615,2.161714,1.9466745,1.9881734,2.3503454,2.6106565,1.9730829,1.8636768,1.9202662,1.9768555,2.0636258,2.4522061,2.746471,2.6597006,2.1843498,1.5845025,1.1053791,0.69793564,0.47535074,0.5319401,0.9205205,1.0638802,0.7922512,0.5696664,0.6526641,1.0827434,1.4298248,1.8900851,2.8521044,4.063117,4.5988297,5.802297,5.832478,5.5004873,5.0515447,4.187614,3.9612563,4.7610526,5.3873086,5.3986263,5.1345425,4.3121104,3.8820312,3.5160866,3.1539145,3.0105548,3.5500402,4.006528,4.244203,4.376245,4.745962,4.5837393,4.5761943,4.146115,3.2935016,2.5804756,2.9539654,3.0143273,2.938875,2.8936033,3.0030096,4.5460134,4.738417,4.1574326,3.561358,3.9197574,4.093298,3.8367596,3.3764994,2.9916916,3.0331905,3.874486,4.1762958,4.1008434,3.7462165,3.1425967,3.308592,3.2784111,3.3312278,3.6707642,4.432834,4.0593443,4.3007927,4.561104,4.659192,4.798779,5.775889,6.119198,6.5228686,6.8435416,6.1078796,5.692891,5.798525,5.485397,5.349582,7.4999785,7.2396674,6.7869525,7.273621,7.960239,6.228604,7.7301087,7.2283497,7.122716,8.0206,8.741172,9.186342,9.654147,9.646602,12.808062,26.913906,31.59196,22.801746,12.408164,6.221059,3.9876647,7.1000805,9.22784,9.454198,8.541223,8.933576,10.269085,8.401636,6.058836,4.957229,5.80607,7.7376537,11.544232,13.283413,12.223305,10.827434,10.70671,10.646348,10.585986,10.880251,12.306303,11.072655,10.978339,10.544487,9.797507,10.26154,10.582213,10.386037,10.099318,9.869187,9.57115,10.223814,10.887795,11.431054,11.785681,11.921495,10.661438,10.763299,11.272603,11.438599,10.702937,10.265312,10.265312,10.79348,11.431054,11.268831,11.774363,11.649866,11.415963,11.276376,11.114153,10.193633,10.1294985,10.287949,10.352083,10.310584,10.925522,10.216269,9.152389,8.243186,7.54525,7.2887115,6.983129,6.647365,6.2889657,5.9003854,5.5080323,4.9534564,4.640329,4.749735,5.240176,5.0968165,5.2779026,5.9192486,6.439871,5.564622,4.2404304,3.6745367,3.3010468,2.897376,2.565385,2.5993385,2.5125682,2.6182017,2.8936033,2.9728284,3.6971724,4.2404304,4.7648253,5.583485,7.1604424,6.809588,7.1981683,7.6584287,7.5075235,6.0701537,5.1835866,4.4630156,4.2819295,4.515832,4.515832,4.749735,4.938366,5.349582,5.5306683,4.315883,4.0404816,4.0782075,4.1197066,4.0895257,4.123479,3.5575855,2.727608,1.9655377,1.5279131,1.5882751,2.3428001,2.8445592,2.938875,2.637065,2.1051247,2.595566,2.6898816,2.7200627,2.886058,3.2520027,3.519859,3.7047176,4.074435,4.5724216,4.8138695,5.0854983,5.4740787,5.6513925,5.4778514,5.0025005,4.236658,3.3878171,3.2633207,4.0178456,5.160951,5.7909794,6.470052,7.284939,8.111144,8.616675,8.59404,8.560086,8.348819,7.8621507,7.0887623,6.85486,7.673519,8.431817,8.771353,9.0957985,9.608876,9.688101,9.703192,9.7069645,9.416472,9.367428,9.839006,10.080454,9.733373,8.854351,8.563859,8.956212,9.691874,10.438853,10.872705,11.370691,11.41219,10.963248,10.408672,10.518079,11.695138,11.740409,11.227332,10.533169,9.861642,10.265312,10.518079,10.827434,11.2650585,11.778135,11.898859,11.623458,11.359374,11.457462,12.253486,2.093807,2.1881225,2.2069857,2.1013522,1.9806281,2.1013522,2.3277097,2.1994405,2.233394,2.4559789,2.4031622,2.263575,2.3692086,2.6446102,2.8219235,2.4182527,2.3088465,2.4522061,2.6898816,3.048281,3.7499893,4.3913355,4.8742313,5.251494,5.6023483,6.0362,6.0626082,6.832224,7.5112963,8.284684,10.38981,13.196642,14.939595,17.1164,18.734856,16.324148,18.715992,25.993385,27.60807,21.11161,12.147853,7.605612,4.293247,2.3692086,1.6637276,1.6825907,1.9278114,1.7731338,1.418507,1.0601076,0.87147635,1.0601076,0.9695646,0.7205714,0.46026024,0.362172,0.32067314,0.3169005,0.39989826,0.5319401,0.58475685,0.7205714,0.754525,0.6187105,0.5093044,0.8978847,1.3317367,1.5052774,1.6486372,1.901403,2.2975287,2.7313805,2.727608,2.3880715,1.9806281,1.9240388,1.5845025,1.871222,2.584248,3.1199608,2.4597516,1.3430545,0.7696155,0.6375736,0.7469798,0.8186596,0.7507524,0.70170826,0.63002837,0.48666862,0.241448,0.24899325,0.211267,0.18863125,0.21881226,0.28294688,0.26031113,0.2867195,0.27540162,0.27540162,0.4640329,0.6187105,0.6187105,0.62248313,0.69039035,0.784706,0.8563859,1.1204696,1.1883769,0.90920264,0.3734899,0.72811663,0.95824677,1.2600567,1.7089992,2.2484846,2.335255,2.1013522,1.7467253,1.3996439,1.0827434,1.1846043,1.116697,0.94692886,0.77338815,0.7167987,0.79602385,0.88279426,1.026154,1.1959221,1.2487389,1.5128226,2.233394,2.7540162,3.0143273,3.5349495,4.447925,6.039973,7.9715567,9.318384,8.537451,9.024119,9.073163,10.502988,13.106099,14.649103,15.667711,14.166207,14.169979,15.83748,15.475307,16.769318,17.410664,17.112627,16.595778,17.603067,19.304522,19.734602,19.346022,19.002712,19.972277,17.738882,19.078165,20.345766,19.734602,17.28994,15.513034,13.947394,13.302276,13.532406,13.837989,15.769572,16.150608,16.18456,16.116653,15.23386,16.678776,17.282394,17.652113,18.58395,21.036158,21.666185,22.537663,23.307278,24.269297,26.34424,26.90259,28.01174,28.728539,29.464201,31.969225,32.17672,31.33165,30.25268,29.679241,30.290405,29.550972,30.143274,31.226017,32.26349,32.99915,33.255688,32.648296,32.1239,31.99186,31.89,32.58039,33.319824,33.949852,34.244118,33.912125,33.93099,35.545673,37.198082,38.47323,40.09923,37.718704,36.398285,34.783604,32.874653,32.040905,32.818066,32.89729,31.293924,29.000168,28.97376,34.715694,41.306473,45.82985,45.882664,39.582382,36.1342,35.315544,39.484295,47.47094,54.571022,50.51545,43.117332,37.254673,34.8666,34.91942,33.32737,32.776566,31.176973,28.754948,28.087193,25.661396,22.986605,20.858843,19.383747,17.976559,16.890041,16.165699,14.483108,12.027128,10.47658,9.982366,10.303039,10.7218,11.053791,11.631002,15.309312,19.836462,21.813318,20.843754,19.493153,19.353567,19.840235,21.624687,25.038912,30.060276,33.821583,38.941036,47.452076,54.959602,50.624855,35.99084,29.143528,25.631214,22.831926,19.957186,18.006739,16.003475,13.151371,9.476834,5.824933,5.541986,4.779916,3.863168,3.0897799,2.7238352,3.048281,3.5123138,4.3913355,5.6061206,6.749226,10.054046,12.96274,13.762536,12.415709,10.555805,9.009028,7.61693,7.0472636,7.17176,7.020855,7.5037513,7.598067,6.8058157,5.492942,4.8855495,4.9534564,5.7004366,4.2819295,1.237421,0.47912338,0.19994913,0.2565385,0.784706,1.5467763,1.9768555,1.8561316,2.2447119,2.9426475,3.953711,5.4740787,5.8890676,5.7192993,4.7346444,3.7952607,4.878004,4.3611546,5.281675,7.8923316,10.253995,8.258276,6.006019,3.4972234,3.1614597,4.353609,3.3840446,3.610402,4.9459114,6.25124,6.7680893,6.126743,6.6662283,7.032173,7.435844,7.6508837,7.0170827,7.2698483,6.930312,7.020855,7.5037513,7.2698483,5.379763,4.8063245,4.538468,4.187614,3.9612563,3.9197574,3.4481792,2.5917933,1.6750455,1.3355093,0.995973,1.0751982,1.5316857,2.2484846,3.0256453,2.3805263,1.4335974,1.6146835,2.686109,2.7653341,2.8143783,2.2560298,1.6335466,1.3317367,1.5882751,1.1431054,1.1129243,1.1053791,1.0789708,1.3656902,1.0525624,0.97710985,1.0525624,1.1091517,0.9242931,1.6637276,1.8976303,2.1390784,2.3465726,1.9202662,2.4597516,2.8294687,2.8445592,2.7540162,3.2029586,2.8898308,2.686109,2.584248,2.7691069,3.6330378,3.8669407,3.953711,3.5274043,2.6219745,1.6825907,1.237421,0.7432071,0.45648763,0.52062225,0.9318384,0.95447415,0.663982,0.45648763,0.5394854,0.91297525,1.6260014,1.9127209,2.2409391,3.1048703,4.9987283,6.19465,6.089017,5.855114,5.6815734,4.7648253,4.561104,4.9345937,5.2628117,5.2892203,5.1232247,4.534695,4.0291634,3.5387223,3.1425967,3.048281,3.821669,4.3422914,4.4931965,4.429062,4.6026025,3.9914372,3.7952607,3.5538127,3.1010978,2.5616124,2.7992878,2.9200118,2.886058,2.795515,2.897376,3.610402,4.0404816,3.9159849,3.5462675,3.8103511,4.3800178,4.014073,3.4066803,2.9803739,2.8936033,3.4972234,3.9763467,4.1272516,3.8669407,3.2482302,3.85185,3.8858037,4.1083884,4.459243,4.063117,3.99521,4.7572803,5.0741806,4.749735,4.6327834,5.028909,4.8100967,5.1458607,5.836251,5.3080835,4.8365054,5.4438977,5.5193505,5.20245,6.3644185,6.651138,6.2135134,6.590776,7.5792036,7.24344,8.114917,7.564113,7.5565677,8.394091,8.710991,9.646602,10.303039,9.1825695,11.227332,27.830654,26.397057,20.964478,14.252977,8.552541,5.7306175,7.756517,9.058073,9.344792,9.224068,10.212496,11.627231,10.016319,7.677292,6.0324273,5.670255,3.059599,6.224831,11.019837,13.890805,11.872451,10.529396,10.661438,10.446399,10.008774,11.400873,11.16697,11.295239,10.993429,10.329447,10.253995,9.922004,9.639057,9.680555,9.95973,10.005001,10.03141,10.914205,11.921495,12.404391,11.766817,10.574668,10.710483,11.080199,10.93684,9.88805,10.653893,10.880251,11.004747,11.034928,10.555805,11.050018,11.25374,11.419736,11.672502,12.034674,10.680302,10.110635,9.993684,10.023865,9.9257765,11.114153,10.412445,9.129752,7.986647,7.115171,6.930312,6.6624556,6.428553,6.417235,6.911449,5.9682927,5.2364035,4.870459,4.9534564,5.511805,5.1043615,5.304311,5.9682927,6.4511886,5.59103,4.4403796,3.8556228,3.5047686,3.1425967,2.6106565,2.6295197,2.7540162,2.9501927,3.1539145,3.2821836,4.183841,4.825187,5.4967146,6.398372,7.654656,7.3188925,7.2170315,7.3151197,7.062354,5.3759904,4.7233267,4.3649273,4.395108,4.6516466,4.7044635,4.659192,5.13077,5.7607985,5.9909286,5.0439997,4.6554193,4.7610526,4.821415,4.6931453,4.61392,3.9612563,3.1124156,2.2975287,1.9164935,2.5125682,2.7540162,2.5125682,2.4786146,2.8106055,3.1614597,3.1652324,3.127506,3.2142766,3.4255435,3.6028569,3.92353,4.4215164,4.8666863,4.979865,4.4177437,4.6818275,5.168496,5.3986263,5.2137675,4.745962,4.044254,3.380272,3.410453,4.217795,5.323174,6.6586833,7.443389,8.016829,8.52236,8.941121,9.144843,8.805306,8.22055,7.677292,7.466025,7.598067,7.8923316,8.371455,8.903395,9.201432,9.533423,9.510788,9.2995205,9.224068,9.763554,9.710737,9.703192,9.997457,10.291721,9.733373,9.374973,9.295748,9.522105,10.035183,10.774617,11.317875,11.815862,11.921495,11.631002,11.272603,12.785426,12.838243,12.15917,11.532914,11.819634,11.876224,11.570641,11.7894535,12.491161,12.706201,12.623203,12.449662,12.174261,12.042219,12.574159,1.9240388,2.0447628,2.3880715,2.4295704,2.2258487,2.3956168,2.6898816,2.5691576,2.3993895,2.293756,2.1202152,2.2183034,2.4522061,2.5201135,2.3805263,2.2598023,2.4031622,2.4861598,2.867195,3.5424948,4.164978,4.2404304,4.878004,5.20245,5.3269467,6.379509,6.7944975,7.0359454,7.7602897,9.461743,12.449662,13.355092,14.954685,18.316093,20.802254,16.06761,21.09652,31.803228,34.50443,26.883726,17.957695,11.891314,6.888813,3.9084394,2.8521044,2.546522,2.5616124,2.3163917,1.7429527,1.0940613,0.94692886,1.2525115,1.0072908,0.6149379,0.32821837,0.23013012,0.5470306,0.73566186,0.814887,0.7809334,0.6111652,0.55080324,0.6073926,0.65643674,0.7884786,1.3128735,1.7278622,1.6863633,1.6976813,2.003264,2.5804756,2.897376,2.7653341,2.757789,3.1539145,3.9348478,3.1199608,3.4632697,4.3724723,4.9987283,4.2404304,2.4220252,1.5203679,1.3619176,1.478869,1.0978339,1.0487897,0.8526133,0.633801,0.4376245,0.23013012,0.26408374,0.21881226,0.24522063,0.32067314,0.26031113,0.24899325,0.27917424,0.32444575,0.41498876,0.67152727,0.965792,1.0186088,1.0374719,1.0902886,1.1129243,1.1883769,1.4071891,1.4449154,1.20724,0.83752275,1.7165444,2.1013522,2.2560298,2.2598023,2.0296721,1.871222,1.7957695,1.6486372,1.4600059,1.448688,1.6071383,1.3996439,0.9997456,0.63002837,0.59607476,0.65643674,0.69793564,0.98465514,1.4071891,1.478869,2.0787163,2.0900342,2.1805773,2.8143783,4.2404304,5.353355,6.0626082,6.477597,6.647365,6.560595,7.232122,7.9225125,9.405154,12.608112,18.614132,17.308804,15.784663,15.116908,15.294222,15.181043,16.03743,16.818363,16.124199,15.196134,17.942604,20.104319,19.938324,18.949896,17.799244,16.31283,16.373192,17.595524,20.043957,21.790682,18.934805,18.41041,16.109108,14.302021,13.860624,14.252977,14.973549,16.048746,16.610868,16.516552,16.358103,18.602814,18.761265,18.663176,19.413929,21.375692,22.63575,23.243143,23.646814,24.608833,27.223263,28.211689,30.048958,31.441057,32.105038,32.776566,32.00695,31.210926,30.8148,30.690304,30.165909,30.335678,31.324106,31.769276,31.486328,31.448603,31.765503,31.614597,32.105038,33.319824,34.330887,35.285362,37.22449,38.303463,37.963924,36.926453,36.93777,38.2431,40.023777,41.845955,43.641727,42.332626,41.27629,39.518246,37.2509,35.81353,37.50744,37.23581,34.17998,29.607561,26.887499,30.694077,37.431984,46.66737,53.537323,48.74986,41.072567,36.737823,38.707134,48.83286,67.83934,77.68967,66.86978,50.677673,39.21644,37.398033,36.26247,35.447586,32.904835,29.822601,30.64126,26.951633,24.740875,22.963968,21.360603,20.432537,17.769064,15.135772,12.691111,10.4049,8.073418,7.6584287,8.22055,9.224068,10.18986,10.725573,13.057055,15.773345,16.716501,15.735619,14.709465,16.637276,16.837225,21.492645,31.097748,40.434994,38.68827,36.90759,40.67644,49.259163,55.61604,41.140476,33.101013,28.770039,25.51049,20.73812,18.417955,15.165953,11.570641,8.390318,6.5455046,4.738417,4.0480266,3.3312278,2.233394,1.2223305,1.5241405,2.5012503,3.9348478,5.372218,6.1041074,9.97482,13.36641,14.173752,12.593022,11.155652,9.578695,8.280911,7.6697464,7.5792036,7.2623034,7.4811153,8.186596,7.643338,5.983383,5.20245,4.847823,6.9567204,5.9003854,1.8599042,0.80734175,0.43007925,0.5470306,1.1431054,1.780679,1.5882751,1.2336484,1.5015048,2.11267,3.3010468,5.828706,6.379509,5.6363015,5.247721,5.7192993,6.439871,4.8402777,4.561104,6.224831,8.296002,7.0510364,6.5228686,4.991183,3.1312788,1.991946,3.006782,4.8742313,5.4703064,5.4703064,5.6023483,6.651138,6.651138,6.571913,6.832224,7.1981683,6.760544,7.443389,8.228095,8.710991,8.379,6.620957,4.889322,4.1612053,4.1762958,4.485651,4.485651,4.4743333,3.199186,1.8561316,1.0186088,0.6413463,0.7394345,0.965792,2.0636258,3.500996,3.4632697,3.1237335,1.7165444,0.8563859,1.2525115,2.71629,3.9386206,3.802806,3.4255435,3.31991,3.4179983,1.3430545,1.1619685,1.4562333,1.5845025,1.6939086,1.9881734,1.4298248,0.965792,0.8865669,0.83752275,1.0714256,1.5882751,2.3314822,2.9200118,2.6408374,2.6144292,2.8106055,2.8521044,3.029418,4.2894745,3.7990334,3.712263,3.712263,4.063117,5.5985756,4.7572803,4.8666863,4.8855495,4.112161,2.1805773,1.5241405,0.7922512,0.44894236,0.62625575,1.1129243,0.8337501,0.6451189,0.52062225,0.48666862,0.59607476,1.4260522,2.2447119,2.8256962,3.5575855,5.462761,6.952948,6.719045,6.2625575,6.058836,5.5683947,5.4363527,5.1345425,5.3382645,5.7079816,4.927048,4.659192,4.2706113,3.6141748,2.9766011,3.097325,4.025391,4.478106,4.5120597,4.3196554,4.2102494,4.38379,4.0970707,3.6669915,3.199186,2.5616124,2.674791,2.565385,2.5578396,2.776652,3.1425967,3.289729,3.802806,3.8895764,3.4330888,3.006782,3.7009451,3.6368105,3.4557245,3.4066803,3.3576362,3.9801195,4.6856003,4.678055,4.0291634,3.663219,4.1008434,4.349837,4.5309224,4.478106,3.7235808,3.772625,4.3686996,4.7233267,4.7912335,5.2779026,5.2062225,4.98741,4.98741,5.111907,4.8063245,5.0025005,5.885295,6.1644692,5.775889,5.873977,6.6322746,6.326692,6.156924,6.620957,7.5226145,7.6320205,7.6697464,8.096053,8.684583,8.514814,9.771099,10.661438,9.699419,10.11818,19.881733,15.158407,17.512526,19.719511,17.437073,9.186342,9.491924,10.106862,9.148616,8.322411,12.925014,8.016829,9.325929,10.314357,9.137298,8.635539,4.425289,4.8100967,9.035437,13.705947,12.800517,10.227587,9.684328,9.371201,9.363655,11.59705,11.548005,11.92904,11.849815,11.046246,9.88805,9.937095,9.454198,9.258021,9.491924,9.612649,9.5032425,11.1782875,12.619431,12.721292,11.291467,10.265312,10.631257,11.106608,11.083972,10.61994,10.985884,10.812344,10.378491,9.895596,9.507015,10.714255,11.080199,11.41219,11.876224,12.0082655,11.299012,10.838752,10.570895,10.38981,10.133271,10.182315,9.733373,8.903395,7.8734684,6.8963585,7.3717093,7.17176,6.85486,6.8737226,7.5829763,6.228604,5.541986,5.2175403,5.194905,5.6476197,5.1835866,5.6061206,6.168242,6.3342376,5.798525,4.881777,4.1612053,3.6028569,3.1840954,2.8521044,3.048281,3.078462,3.1539145,3.3651814,3.7084904,4.8553686,5.462761,6.3945994,7.6282477,8.239413,7.201941,7.145352,7.273621,6.828451,5.0968165,4.7535076,4.349837,4.214022,4.4101987,4.715781,5.081726,5.4665337,5.617439,5.5457587,5.5080323,5.409944,5.413717,4.9685473,4.2706113,4.2706113,3.942393,3.3123648,2.8106055,2.7540162,3.3425457,2.8898308,2.595566,2.7841973,3.3463185,3.7235808,3.440634,3.187868,3.3312278,3.8820312,4.515832,4.7610526,4.9685473,4.979865,4.708236,4.134797,4.146115,4.085753,4.0970707,4.183841,4.195159,3.7198083,3.610402,4.0178456,4.870459,5.8588867,6.983129,7.756517,8.801534,9.989911,10.469034,10.502988,9.405154,7.914967,7.0170827,7.91874,9.152389,9.4127,9.5183325,9.774872,9.993684,10.091772,10.208723,9.933322,9.457971,9.567377,9.21275,8.82417,9.367428,10.612394,11.121698,10.56335,9.880505,9.688101,10.03141,10.419991,11.32542,12.034674,12.23085,12.042219,12.053536,14.237886,14.747191,14.400109,13.95494,14.11339,13.185325,12.377983,12.321393,12.989148,13.671993,13.743673,13.505998,13.147598,12.913695,13.12119,2.2296214,2.173032,2.655928,2.9011486,2.6634734,2.1994405,1.9844007,2.0258996,2.1466236,2.2220762,2.1579416,2.4295704,2.4672968,2.4974778,2.584248,2.637065,2.6446102,2.7615614,3.187868,3.863168,4.447925,4.187614,4.466788,4.957229,5.624984,6.730363,6.307829,7.122716,8.884532,11.242422,13.792717,13.456953,14.7736,16.659912,17.225805,13.79649,23.514772,36.51901,38.035606,27.29117,17.520071,11.012292,6.8963585,4.323428,2.8143783,2.2560298,2.4522061,2.2183034,1.5618668,0.7997965,0.55457586,0.7130261,0.56589377,0.38480774,0.3055826,0.32821837,1.1695137,1.1242423,0.79602385,0.6187105,0.87902164,0.7582976,0.7432071,0.7432071,0.95824677,1.8749946,1.50905,1.2487389,1.3732355,1.6825907,1.5052774,1.9579924,2.2560298,2.9841464,4.0970707,4.938366,3.8254418,4.3385186,5.379763,5.7683434,4.2404304,2.5502944,1.6109109,1.2110126,1.0827434,0.9280658,0.97710985,0.70170826,0.38480774,0.19240387,0.181086,0.13958712,0.13204187,0.181086,0.2678564,0.331991,0.271629,0.2565385,0.331991,0.573439,1.0751982,1.8863125,2.41448,2.6823363,2.9464202,3.7009451,3.2784111,2.5502944,2.0070364,1.7316349,1.4147344,3.0633714,3.4859054,3.1237335,2.2975287,1.237421,0.9507015,0.9318384,0.9242931,0.9205205,1.1431054,1.3732355,1.327964,1.0035182,0.60362,0.5583485,0.5998474,0.6752999,0.83752275,1.0525624,1.1732863,1.4109617,1.8184053,2.1768045,2.4823873,2.9351022,4.5950575,5.6061206,6.149379,6.5002327,7.0510364,7.533932,8.001738,8.616675,9.563604,11.046246,11.763044,12.521342,12.857106,12.73261,12.54775,14.6302395,16.957949,18.146326,18.157644,18.297232,17.852062,16.509007,16.735365,17.829426,15.920478,18.255732,18.4255,18.938578,19.930779,19.1423,20.289177,18.938578,17.222033,16.048746,15.131999,15.441354,15.852571,16.018566,16.165699,17.08999,20.545715,20.372175,20.043957,20.485353,20.059048,22.93756,24.484337,25.506718,26.951633,29.905598,32.029587,33.448093,34.77606,35.274044,32.859562,30.969479,31.708914,31.810774,30.494127,29.471746,29.973505,30.25268,30.026323,29.37743,28.71345,29.188799,29.766012,31.176973,33.044422,33.881947,36.52278,38.680725,40.40481,41.86482,43.34746,43.155056,42.408077,41.51774,41.24988,42.71366,42.521255,42.728752,42.347717,41.41965,41.023525,40.004917,39.684242,37.907337,34.55347,31.535372,31.535372,33.391502,41.6196,54.880375,65.96435,53.93722,42.70989,37.484802,41.857273,57.807934,83.70323,91.84078,80.975624,59.3698,44.758423,41.796913,40.951843,38.793903,34.73833,31.05625,28.102283,26.480055,24.250433,21.507734,20.394812,17.440845,14.581196,12.479843,10.785934,8.122461,7.1981683,7.6282477,8.612903,9.58624,10.201178,10.140816,11.608367,13.230596,14.1058445,13.792717,15.663939,15.920478,23.111101,37.26599,49.89674,46.557964,38.75995,37.164127,44.513203,55.619812,45.799667,35.881435,30.309269,28.328642,23.993895,17.516298,13.690856,11.302785,9.352338,7.0585814,4.930821,3.7499893,2.6936543,1.5543215,0.7582976,1.0827434,1.6863633,3.1048703,4.9232755,5.7607985,8.431817,10.842525,12.200669,12.415709,12.106354,10.853842,9.201432,8.103599,7.673519,7.1906233,7.0774446,8.118689,7.858378,6.1229706,5.0213637,5.534441,6.696409,5.3948536,2.123988,0.965792,0.5885295,0.6828451,1.1732863,1.7278622,1.7580433,1.7165444,2.4371157,2.6219745,2.5238862,3.9386206,4.7006907,6.5455046,8.763808,9.733373,6.937857,5.6325293,5.0025005,5.7494807,6.688864,4.7308717,5.3269467,5.6513925,5.8513412,6.006019,6.1305156,6.0550632,5.05909,4.395108,4.67051,5.847569,6.4021444,7.111398,7.7942433,7.8395147,6.2097406,6.356873,6.360646,6.900131,7.496206,6.549277,7.032173,5.7381625,4.8327327,4.749735,4.191386,3.4670424,2.2484846,1.2223305,0.62248313,0.2263575,0.98842776,1.026154,1.9278114,3.5047686,3.8292143,2.5691576,3.308592,3.187868,2.505023,4.7308717,6.643593,8.959985,9.665465,8.201687,5.455216,2.9313297,2.1768045,1.9693103,1.7014539,1.3996439,1.0676528,0.6752999,0.814887,1.2751472,1.0714256,1.8599042,1.9202662,1.7316349,1.8259505,2.7879698,2.7502437,2.7841973,2.927557,3.2746384,3.9461658,4.2894745,4.61392,4.5912848,4.4101987,4.8063245,4.1197066,3.821669,4.0706625,4.1612053,2.535204,1.4675511,0.814887,0.55080324,0.69039035,1.2864652,1.2185578,0.7696155,0.47535074,0.5281675,0.76584285,0.9922004,2.5314314,3.6481283,4.436607,6.8171334,7.7602897,6.5945487,5.523123,5.409944,5.7419353,5.692891,5.3646727,5.583485,6.085244,5.5382137,5.191132,4.432834,3.5462675,2.916239,3.0369632,3.6330378,4.244203,4.538468,4.4441524,4.1498876,4.436607,3.874486,3.3236825,2.9916916,2.4182527,2.3918443,1.7278622,1.7014539,2.5276587,3.361409,3.0105548,3.2255943,3.3123648,3.0709167,2.7502437,3.1425967,3.1350515,3.0822346,3.169005,3.3953626,4.5724216,5.8136153,6.085244,5.2967653,4.285702,4.7346444,4.5497856,4.353609,4.217795,3.6858547,3.9801195,4.285702,4.285702,4.0593443,4.1083884,4.961002,5.670255,5.7381625,5.2099953,4.67051,4.908185,5.4703064,5.6061206,5.342037,5.458988,5.2779026,6.1908774,6.888813,6.820906,6.1908774,6.6624556,6.356873,6.609639,7.3377557,7.0510364,8.843033,10.623712,9.831461,8.0206,10.861387,13.306048,21.017294,20.413673,11.046246,5.5985756,5.511805,6.439871,6.089017,6.405917,13.59654,14.086982,9.337247,8.001738,11.012292,11.566868,6.8171334,7.3905725,10.925522,12.883514,6.5530496,8.284684,8.756263,8.616675,8.899622,11.034928,11.329193,12.00072,12.019584,11.197151,10.193633,10.299266,9.846551,9.680555,9.967276,10.186088,10.536942,11.92904,12.996693,13.000465,11.864905,10.8576145,10.506761,10.653893,10.899114,10.582213,10.589758,10.008774,9.416472,9.178797,9.480607,10.495442,10.593531,10.665211,10.970794,11.155652,11.423509,11.536687,11.536687,11.336739,10.718028,10.084227,9.7069645,8.835487,7.4811153,6.458734,7.6282477,7.4735703,6.9227667,6.560595,6.643593,5.560849,5.281675,5.3910813,5.643847,5.9494295,5.4288073,5.27413,5.292993,5.3873086,5.553304,4.708236,3.7877154,3.150142,2.9464202,3.1350515,3.1916409,3.0407357,3.0897799,3.5085413,4.221567,5.036454,6.0814714,7.115171,7.8131065,7.752744,6.930312,7.01331,7.073672,6.560595,5.304311,5.040227,4.564876,4.2064767,4.2064767,4.727099,5.6098933,5.7381625,5.6061206,5.6023483,5.9984736,6.0739264,5.081726,3.9876647,3.3727267,3.429316,3.772625,3.7650797,3.4859054,3.1727777,3.2331395,3.4066803,3.3236825,3.3236825,3.5236318,3.832987,3.5047686,3.2369123,3.2935016,3.8103511,4.798779,5.081726,5.1873593,5.010046,4.52715,3.8065786,3.5236318,3.7575345,4.1197066,4.323428,4.1612053,4.2781568,4.5535583,5.27413,6.3531003,7.3113475,7.654656,8.239413,9.073163,10.065364,11.027383,10.997202,9.963503,8.959985,8.484633,8.480861,8.952439,8.6581745,8.627994,9.125979,9.639057,10.450171,10.650121,10.378491,9.805053,9.103344,9.031664,8.816625,9.374973,10.431308,10.514306,10.751981,10.763299,10.265312,9.661693,10.03141,11.099063,11.793225,12.234623,12.808062,14.177525,16.31283,16.290195,15.490398,14.943368,15.347038,14.769827,13.513543,12.664702,12.838243,14.18507,15.411173,14.618922,13.419228,12.796744,13.109872,2.3956168,2.5314314,2.897376,2.8709676,2.4069347,2.04099,1.8334957,1.8221779,1.9391292,2.093807,2.203213,2.2409391,2.2975287,2.3465726,2.4371157,2.704972,2.9652832,3.2784111,3.7537618,4.349837,4.8742313,4.7950063,5.2062225,5.5004873,5.6551647,6.205968,6.326692,7.726336,9.239159,10.510533,12.015811,13.257004,15.807299,17.093763,16.784409,16.791954,26.58946,34.77606,32.63698,21.579414,13.117417,8.443134,6.089017,4.214022,2.4672968,1.9881734,2.2484846,1.7278622,1.0110635,0.47157812,0.27540162,0.38103512,0.39989826,0.35462674,0.29049212,0.29426476,0.8563859,0.9695646,1.0186088,1.20724,1.5958204,1.2864652,1.1808317,1.1016065,1.0751982,1.3166461,1.0148361,0.8526133,1.0827434,1.5241405,1.539231,2.2975287,2.7426984,3.9914372,5.5306683,5.243949,4.961002,5.553304,6.3832817,6.511551,4.719554,2.5804756,1.720317,1.4373702,1.267602,0.9507015,0.845068,0.49421388,0.23013012,0.150905,0.11317875,0.16976812,0.18485862,0.25276586,0.362172,0.38858038,0.43007925,0.4376245,0.58098423,0.95824677,1.6146835,2.3201644,2.9426475,3.4632697,4.036709,4.9534564,4.8138695,4.0593443,3.1124156,2.354118,2.1164427,3.5764484,4.2064767,3.8556228,2.746471,1.478869,1.3807807,1.2487389,0.95447415,0.6488915,0.7469798,0.845068,0.84884065,0.73566186,0.573439,0.5394854,0.6073926,0.7394345,0.87902164,0.9695646,0.9808825,0.9280658,1.1016065,1.3920987,1.7655885,2.2899833,3.7386713,4.3913355,5.093044,5.9230213,6.1908774,6.439871,7.092535,7.8734684,8.744945,9.895596,10.846297,11.970539,12.604341,12.823153,13.45318,14.886778,16.535416,18.082191,19.191343,19.523335,17.165443,15.452672,15.358356,16.463736,16.969267,19.391293,19.323385,18.780127,18.5085,18.014284,19.700647,20.26277,20.391039,19.957186,18.033148,17.667202,16.908905,16.897587,17.810562,18.836716,19.681786,21.013521,22.315077,22.956423,22.17549,23.428001,24.529608,25.838709,27.921198,31.539145,34.64779,36.1757,36.8095,36.409603,34.03662,32.9237,31.72023,30.211182,29.120892,30.120638,30.075367,29.426476,27.99665,25.959433,23.839218,25.170954,26.872408,28.67195,30.42622,32.12013,33.93099,36.71896,39.080624,41.10275,44.39248,46.10525,46.640965,46.11657,45.437496,46.290108,45.626125,44.833874,44.43398,44.14726,42.875885,41.729004,40.333134,38.925945,37.696068,36.756687,34.39125,33.644268,37.11886,46.614555,63.153744,63.659275,51.960365,40.706623,37.737568,46.05998,66.45479,85.88381,92.68962,83.22788,61.878593,50.764442,46.573055,43.543636,39.042896,33.565044,31.124157,28.841719,25.65385,22.07363,20.175999,17.097536,14.57365,12.894833,11.555551,9.239159,8.243186,8.627994,9.857869,11.050018,10.997202,9.9257765,10.091772,11.231105,12.774108,13.837989,15.297995,15.807299,22.1189,35.00996,49.259163,48.57632,40.64249,35.719215,39.129665,51.269974,48.91963,39.201347,31.467464,27.872154,23.363867,17.274849,13.4644985,10.989656,9.205205,7.7829256,4.957229,3.2482302,2.0900342,1.4071891,1.5920477,1.2940104,2.0598533,4.1083884,6.2436943,5.8588867,7.3792543,8.639311,10.061591,11.46878,12.08749,11.868678,10.729345,9.465516,8.465771,7.7225633,7.0284004,7.643338,7.61693,6.6360474,5.9984736,5.624984,5.2628117,3.904667,1.9127209,0.9997456,0.7809334,0.90543,1.20724,1.50905,1.6071383,1.6071383,2.2673476,2.8106055,3.078462,3.5085413,3.5802212,4.496969,6.039973,6.9793563,5.070408,6.356873,5.7909794,5.8702044,6.7944975,6.511551,6.387054,6.096562,6.0626082,6.013564,4.961002,5.353355,4.478106,3.6556737,3.5839937,4.3007927,5.832478,7.2358947,7.805561,7.3679366,6.300284,6.0362,6.1342883,6.3229194,6.462507,6.530414,6.9227667,5.9607477,5.624984,5.945657,4.979865,3.0746894,1.659955,0.80356914,0.39989826,0.1961765,1.3053282,1.056335,1.0978339,1.7316349,1.8976303,1.7354075,4.247976,4.5233774,2.4522061,2.7087448,5.330719,10.280403,13.158916,11.864905,6.617184,3.6481283,2.3465726,1.8825399,1.6675003,1.3468271,1.5316857,1.1280149,0.9016574,1.0789708,1.3505998,1.7354075,1.9881734,1.8636768,1.6863633,2.3465726,2.8822856,3.5160866,3.640583,3.3953626,3.640583,4.6742826,5.5004873,6.096562,6.462507,6.620957,5.674028,5.089271,4.851596,4.4743333,3.0256453,1.7467253,1.026154,0.6790725,0.67152727,1.116697,1.1996948,0.73566186,0.43385187,0.52439487,0.76207024,1.3128735,2.746471,4.123479,5.492942,7.914967,8.560086,7.0472636,5.613666,5.2099953,5.4891696,5.8890676,5.621211,5.6815734,6.047518,5.692891,5.4363527,4.425289,3.4368613,2.9426475,3.0860074,3.7084904,4.564876,4.9949555,4.8063245,4.2819295,4.3875628,3.9461658,3.4368613,2.9652832,2.2711203,2.2183034,1.6637276,1.6750455,2.4597516,3.3463185,3.1539145,3.006782,2.8822856,2.8294687,2.9615107,3.1010978,3.0520537,2.9803739,3.0369632,3.3651814,4.9421387,6.1531515,6.3719635,5.5985756,4.485651,5.451443,5.6061206,5.198677,4.4931965,3.8065786,3.7499893,4.315883,4.5007415,4.2291126,4.3347464,4.961002,5.5495315,5.617439,5.251494,5.1232247,5.0251365,5.2288585,5.100589,4.640329,4.478106,4.478106,5.6325293,6.3719635,6.092789,5.1534057,5.553304,5.481624,6.009792,7.0510364,7.333983,8.82417,10.193633,9.903141,9.122208,11.717773,18.372684,25.276588,21.896315,9.989911,3.6028569,3.85185,5.05909,5.5193505,6.4474163,11.970539,15.762027,8.986393,6.3945994,10.804798,13.087236,11.170743,11.849815,12.751472,11.751727,6.9680386,7.696155,8.27714,8.45068,8.718536,10.344538,11.257513,11.849815,11.608367,10.691619,9.929549,10.197406,10.106862,10.110635,10.295494,10.393582,10.77839,11.7026825,12.630749,13.0646,12.559069,11.646093,10.733118,10.435081,10.684074,10.710483,10.627484,10.231359,9.6201935,9.21275,9.767326,10.431308,10.408672,10.325675,10.401127,10.472807,10.744436,11.057564,11.133017,10.842525,10.186088,9.533423,9.122208,8.280911,7.1038527,6.4474163,7.462252,7.496206,7.2585306,6.983129,6.417235,5.564622,5.3948536,5.6853456,6.0814714,6.0626082,5.50426,5.2099953,4.8666863,4.564876,4.7874613,4.164978,3.7235808,3.350091,3.0935526,3.1765501,3.3350005,3.187868,3.1765501,3.561358,4.447925,5.036454,5.904158,6.439871,6.670001,7.273621,6.8473144,6.8774953,6.990674,6.730363,5.564622,4.063117,3.6028569,4.025391,4.9044123,5.534441,5.934339,5.9682927,5.9494295,5.8890676,5.485397,5.836251,5.1081343,4.0103,3.1010978,2.7804246,3.3953626,4.055572,3.9386206,3.3236825,3.5802212,3.9688015,3.8782585,3.572676,3.3350005,3.4594972,3.4745877,3.5047686,3.6254926,3.9989824,4.878004,5.292993,5.194905,4.82896,4.3083377,3.6028569,3.7688525,4.4705606,4.8968673,4.9232755,5.0666356,5.2552667,5.515578,6.2625575,7.201941,7.326438,7.7904706,8.235641,9.0957985,10.167224,10.638803,10.246449,9.688101,9.193887,8.83926,8.548768,8.98262,9.2844305,9.461743,9.87296,11.227332,11.529142,10.77839,10.012547,9.544742,8.986393,8.782671,8.793989,9.167479,9.7220545,9.940866,10.431308,10.616167,10.374719,10.050273,10.446399,10.963248,11.344283,11.631002,12.219532,13.875714,15.882751,16.048746,15.580941,15.211224,15.207452,14.543469,13.7851715,13.283413,13.328684,14.147344,15.07541,14.64533,13.826671,13.253232,13.245687,2.3767538,2.7351532,3.0935526,2.9841464,2.4597516,2.082489,2.04099,2.0145817,2.0183544,2.0862615,2.282438,2.1164427,2.2598023,2.3163917,2.3163917,2.7351532,3.2633207,3.7273536,4.2328854,4.7346444,5.032682,5.2288585,5.409944,5.4665337,5.5306683,5.975838,6.862405,8.514814,9.6051035,10.103089,11.299012,14.369928,18.221779,20.051502,19.94964,20.885252,27.947605,30.656351,25.348267,14.803781,8.216777,6.277648,5.142088,3.5839937,1.8297231,1.5618668,1.7693611,1.1280149,0.543258,0.3470815,0.32444575,0.331991,0.392353,0.422534,0.4074435,0.362172,0.58475685,0.8337501,1.1883769,1.6524098,2.1503963,2.3088465,2.4031622,2.1466236,1.690136,1.6184561,1.4600059,1.2487389,1.3430545,1.7127718,1.9466745,3.380272,3.8178966,4.485651,5.281675,4.798779,5.564622,6.0814714,6.458734,6.258785,4.4818783,2.6672459,2.093807,2.003264,1.8485862,1.2902378,0.95447415,0.55080324,0.27540162,0.181086,0.15467763,0.20749438,0.19240387,0.27540162,0.42630664,0.44139713,0.5583485,1.0072908,1.7316349,2.4371157,2.5616124,2.7691069,3.199186,3.682082,4.183841,4.7950063,4.908185,4.647874,4.244203,3.942393,3.9989824,5.111907,5.7570257,5.0854983,3.3048196,1.6712729,1.7391801,1.7429527,1.448688,0.98465514,0.83752275,0.86770374,0.7054809,0.59607476,0.5998474,0.5998474,0.84884065,0.9507015,0.9620194,0.90920264,0.77716076,0.58475685,0.5017591,0.62248313,0.9620194,1.4335974,2.4899325,2.757789,3.3048196,4.236658,4.6856003,4.561104,5.270357,6.356873,7.6320205,9.159933,10.93684,12.770335,14.011529,14.811326,16.120426,16.863634,17.4333,17.618158,17.603067,17.942604,15.645076,14.543469,14.173752,14.505743,15.946886,17.180534,16.825907,16.625957,17.101309,17.538933,18.863125,19.80251,20.628714,20.979568,19.859098,19.557287,17.991648,17.580433,18.500954,18.69713,19.055529,22.205671,24.66165,25.253952,25.140774,25.148317,25.672712,27.03463,29.460428,33.101013,35.530582,37.28485,37.48103,36.639732,36.654823,36.383194,34.025307,31.210926,29.641514,31.109066,30.199863,29.32084,27.600525,24.929506,21.937815,23.409138,24.257978,25.155863,26.770548,29.769783,30.94307,33.474503,35.722984,37.71493,41.140476,45.030052,48.16133,49.46666,49.628883,51.09266,50.95307,48.874355,47.387943,46.65228,44.45284,43.090923,40.842438,39.208893,38.71845,38.922173,36.726505,35.836166,36.1342,39.688015,50.726715,60.788307,56.619556,46.659824,38.563774,39.182484,49.49307,68.5486,86.404434,93.34983,79.926834,62.87834,53.427914,47.429443,41.600735,33.512226,31.641006,29.856554,26.793182,22.862108,20.228815,18.078419,15.592259,13.6833105,12.3289385,10.601076,9.899368,10.378491,11.442371,12.234623,11.631002,12.132762,11.072655,11.299012,13.324911,15.347038,16.309057,16.822134,20.489126,28.977533,42.00818,47.38417,43.3701,36.451103,33.67445,42.634434,48.082108,41.283836,32.316307,25.823618,20.994658,16.546734,12.570387,9.669238,7.914967,6.8171334,4.3309736,2.7313805,1.7278622,1.3732355,2.0636258,1.6750455,2.7238352,5.1345425,7.2396674,5.772116,6.6134114,7.122716,8.469543,10.525623,11.876224,12.698656,12.449662,11.087745,9.224068,8.099826,6.934085,6.9491754,7.0246277,6.820906,6.779407,5.6363015,4.3724723,2.9728284,1.6712729,0.9808825,1.1581959,1.177059,1.2110126,1.3015556,1.3656902,1.4600059,1.8448136,2.5201135,3.2670932,3.6179473,3.4783602,4.0970707,5.089271,5.6400743,4.478106,7.5490227,7.1604424,7.1264887,8.167733,7.8810134,6.8925858,6.25124,5.987156,5.715527,4.6327834,5.081726,4.6214657,4.2027044,4.285702,4.8666863,5.8626595,6.8925858,7.0774446,6.507778,6.258785,5.4967146,5.406172,5.3571277,5.194905,5.247721,5.0175915,5.0854983,5.3156285,5.2288585,4.002755,2.1692593,1.0525624,0.51684964,0.3470815,0.24522063,1.1657411,0.8186596,0.422534,0.3961256,0.3772625,0.77338815,3.2105038,4.538468,3.6971724,1.7354075,3.0030096,7.8998766,11.370691,10.740664,5.7306175,3.4330888,2.3880715,1.9994912,1.8033148,1.4675511,1.931584,1.3543724,0.88279426,1.0035182,1.5241405,1.3656902,1.7316349,2.082489,2.2862108,2.6219745,3.9801195,5.0062733,5.2779026,5.036454,5.20245,6.1003346,7.020855,7.8395147,8.288457,7.964011,7.1793056,6.809588,6.1606965,5.081726,3.9612563,2.282438,1.358145,0.8526133,0.6828451,1.0072908,1.2449663,0.8186596,0.482896,0.56589377,0.94692886,1.5731846,2.686109,4.002755,5.621211,8.031919,8.631766,7.2660756,5.783434,5.0666356,5.0439997,5.560849,5.6325293,5.7909794,6.017337,5.73439,5.3986263,4.214022,3.2859564,3.048281,3.2746384,3.9574835,4.7308717,5.1458607,4.9685473,4.191386,4.115934,3.9763467,3.5877664,2.8596497,1.7957695,1.9504471,1.7693611,1.81086,2.2296214,2.7653341,2.927557,2.757789,2.5729303,2.5804756,2.9237845,3.0709167,2.8936033,2.7125173,2.8030603,3.4029078,5.1760416,6.0211096,6.013564,5.481624,5.028909,5.9117036,6.356873,5.8664317,4.696918,3.8593953,3.5990841,4.1762958,4.564876,4.459243,4.2894745,4.7308717,4.9760923,4.9459114,4.8402777,5.111907,4.557331,4.7535076,4.7233267,4.2517486,3.8895764,4.5233774,5.194905,5.7004366,5.772116,5.0553174,5.1534057,5.251494,5.7909794,6.779407,7.7678347,8.816625,9.597558,9.665465,9.922004,12.596795,19.447882,25.623669,23.68454,13.717264,3.31991,3.9310753,5.1873593,6.3229194,7.5301595,9.989911,13.758763,9.771099,8.4544525,11.419736,11.449917,11.404645,10.993429,10.850069,10.378491,7.7225633,7.647111,7.8131065,8.039464,8.443134,9.446653,10.782163,11.287694,11.083972,10.423763,9.691874,10.072908,10.246449,10.38981,10.56335,10.710483,10.899114,11.389555,12.238396,13.091009,13.166461,12.351574,11.336739,10.748209,10.733118,10.955703,10.751981,10.514306,10.167224,9.854096,9.9257765,10.099318,9.95973,9.842778,9.827688,9.748463,10.0465,10.423763,10.650121,10.552032,10.005001,9.265567,8.835487,8.130007,7.250985,7.0170827,7.4735703,7.7414265,7.748972,7.4471617,6.8133607,6.319147,6.145606,6.205968,6.2625575,5.9418845,5.6513925,5.2665844,4.8968673,4.6554193,4.659192,3.8895764,3.7462165,3.5953116,3.3425457,3.451952,3.5236318,3.3538637,3.3161373,3.712263,4.772371,5.2364035,5.7079816,5.9418845,6.187105,7.1868505,6.6850915,6.6134114,6.790725,6.692637,5.4740787,3.361409,2.8936033,3.7198083,5.160951,6.2361493,5.772116,5.6589375,5.6891184,5.5382137,4.772371,4.9760923,4.8063245,4.1008434,3.1425967,2.6710186,3.218049,3.9650288,4.0782075,3.7575345,4.2404304,4.406426,4.08198,3.5575855,3.1463692,3.2142766,3.4594972,3.682082,4.044254,4.561104,5.1269975,5.2967653,4.9345937,4.3875628,3.8895764,3.5500402,4.349837,5.093044,5.383536,5.406172,5.945657,5.994701,6.560595,7.4999785,8.296002,8.028146,8.318638,8.431817,9.027891,9.944639,10.186088,9.876732,9.563604,9.333474,9.178797,9.012801,9.442881,10.054046,10.220041,10.401127,12.155397,12.00072,10.767072,10.012547,9.952185,9.450426,8.831716,9.009028,9.329701,9.514561,9.65792,10.26154,10.650121,10.665211,10.393582,10.152134,10.846297,11.114153,11.321648,12.012038,13.913441,15.418718,15.82239,15.618668,15.131999,14.543469,14.124708,13.920986,13.951167,14.203933,14.641558,14.943368,14.867915,14.652876,14.422746,14.177525,2.4371157,2.9464202,3.3312278,3.3463185,2.9615107,2.372981,2.4484336,2.5276587,2.5087957,2.4371157,2.4974778,2.335255,2.516341,2.546522,2.5238862,3.108643,3.5877664,3.9914372,4.5196047,5.0062733,4.9421387,5.270357,4.919503,4.9345937,5.6363015,6.617184,7.91874,9.559832,10.540714,11.133017,12.883514,17.150352,22.167944,25.476536,26.023567,24.156118,28.490864,28.479546,21.503962,10.684074,4.847823,4.949684,4.217795,2.727608,1.20724,1.0186088,1.0714256,0.6111652,0.30935526,0.38103512,0.56589377,0.4640329,0.44894236,0.5281675,0.62248313,0.55080324,0.7054809,0.935611,1.2751472,1.7429527,2.3126192,3.4179983,3.8254418,3.361409,2.6106565,2.897376,2.7011995,2.3163917,2.1579416,2.3277097,2.6106565,4.4177437,4.738417,4.2819295,3.832987,4.217795,5.349582,5.485397,5.342037,4.930821,3.5802212,2.8558772,2.686109,2.6823363,2.4710693,1.690136,1.177059,0.7696155,0.45648763,0.2678564,0.29426476,0.1961765,0.13204187,0.211267,0.3961256,0.5093044,0.7432071,1.81086,3.2935016,4.274384,3.3576362,3.3236825,3.5160866,3.5839937,3.5651307,3.8820312,4.134797,4.5460134,5.3873086,6.4511886,7.0774446,8.016829,8.360137,6.94163,4.1536603,1.9542197,1.8787673,2.1654868,2.2862108,2.0636258,1.6561824,1.539231,1.1129243,0.7469798,0.6111652,0.66775465,1.177059,1.1959221,1.0186088,0.7922512,0.52062225,0.34330887,0.211267,0.211267,0.3169005,0.392353,1.0714256,1.237421,1.4864142,2.1088974,3.0897799,2.8181508,3.451952,4.6818275,6.1041074,7.2283497,9.982366,12.740154,14.916959,16.739138,19.21398,19.719511,19.108345,17.421982,15.437581,14.694374,13.736128,13.59654,13.332457,12.936331,13.336229,13.0646,12.619431,13.377728,15.414946,17.486116,17.803017,17.972786,18.493408,19.281887,19.670467,19.806282,18.640541,18.274595,18.738628,17.969013,20.915434,25.231316,27.619389,27.78161,28.400322,28.796446,29.268024,30.388494,32.29367,34.655334,34.76474,36.496376,37.09245,37.062267,40.178455,40.174683,38.80145,36.156837,33.41791,32.848248,30.867619,30.245134,29.105803,26.898817,24.37493,24.412657,22.7527,21.964222,23.405365,27.23458,28.792673,30.46772,32.22199,34.14603,36.469967,41.04616,46.06375,49.49307,51.54915,54.691746,57.25713,55.397224,52.631893,50.31927,47.64448,45.524265,42.8872,40.423676,38.669407,37.990334,37.18299,37.416893,37.647026,37.779068,38.66186,47.161587,53.250603,51.586876,44.00767,39.52202,43.049423,53.718407,70.64618,87.20422,91.0108,74.69043,61.42588,51.89623,43.72095,31.456148,29.898052,29.471746,27.69484,24.235344,20.922977,20.345766,17.614386,14.849052,13.026875,11.970539,12.106354,12.5326605,12.796744,12.709973,12.3289385,15.071637,13.128735,12.804289,15.546988,17.935059,18.018057,18.059555,19.112118,23.035648,32.4823,43.788857,45.87889,39.09194,30.181,32.32008,43.08715,41.329105,33.11233,23.941078,18.734856,15.354584,11.151879,7.9338303,6.0626082,4.447925,3.240685,2.3163917,1.6109109,1.2902378,1.7542707,1.7919968,2.9916916,5.2628117,7.118943,5.6778007,6.126743,6.3342376,7.6131573,9.914458,11.827179,13.098554,13.747445,12.521342,9.906913,8.099826,6.6662283,6.2135134,6.217286,6.4021444,6.730363,5.5268955,4.2819295,2.897376,1.6222287,1.0336993,1.5430037,1.3732355,1.1959221,1.2185578,1.1883769,1.4109617,1.5430037,1.9164935,2.6068838,3.4368613,3.6481283,5.4703064,6.9793563,7.1906233,6.0626082,8.145098,7.8432875,8.280911,9.352338,7.6886096,6.356873,6.089017,6.0550632,5.885295,5.692891,5.6098933,5.2288585,5.534441,6.5002327,7.0963078,6.066381,6.058836,6.145606,6.0776987,6.300284,5.1571784,4.504514,4.3196554,4.236658,3.5424948,3.4142256,4.4403796,4.485651,3.1161883,1.5731846,0.84884065,0.422534,0.31312788,0.36594462,0.24522063,0.56589377,0.3772625,0.181086,0.14713238,0.09808825,0.2678564,1.086516,3.663219,6.066381,3.3463185,1.5769572,3.5538127,5.666483,5.798525,3.3425457,2.8521044,2.686109,2.4559789,2.0636258,1.6976813,1.7957695,1.1091517,0.84129536,1.237421,1.5731846,1.1846043,1.4109617,2.0900342,2.9615107,3.6481283,5.80607,7.115171,7.7602897,8.07719,8.5563135,8.714764,9.024119,9.246704,9.005256,7.7640624,7.5263867,7.5565677,7.092535,6.017337,4.82896,2.8709676,1.720317,1.0186088,0.7167987,1.0412445,1.3468271,0.97333723,0.6149379,0.69793564,1.4071891,1.6863633,2.41448,3.4368613,4.851596,6.9869013,7.854605,7.066127,5.824933,4.908185,4.644101,4.908185,5.2175403,5.6778007,6.0512905,5.7607985,5.168496,3.8443048,3.0331905,3.078462,3.410453,4.002755,4.447925,4.8138695,4.825187,3.8895764,3.7990334,3.8065786,3.5085413,2.6710186,1.237421,1.629774,1.7467253,1.81086,1.8749946,1.8297231,2.142851,2.3013012,2.335255,2.354118,2.5767028,2.9049213,2.5502944,2.233394,2.4484336,3.451952,5.3156285,5.7306175,5.4703064,5.27413,5.8437963,5.9532022,6.2851934,5.8664317,4.738417,3.9499383,3.6971724,3.85185,4.221567,4.402653,3.7877154,4.3649273,4.2706113,4.104616,4.191386,4.568649,3.7499893,4.3196554,4.749735,4.4630156,3.8405323,5.1043615,5.0251365,5.458988,6.3644185,5.832478,5.6287565,5.715527,5.9418845,6.477597,7.8131065,8.586494,9.21275,9.473062,9.612649,10.3634,15.399856,20.92675,23.284641,18.983849,4.6818275,4.7950063,5.6287565,7.201941,8.812852,9.031664,10.005001,10.8576145,12.513797,13.132507,8.122461,7.4094353,5.583485,6.5040054,9.005256,6.907676,7.575431,7.149124,7.2358947,8.096053,8.635539,9.857869,10.253995,10.465261,10.472807,9.6051035,10.042727,10.340765,10.521852,10.676529,10.985884,10.906659,11.133017,11.940358,13.015556,13.430545,12.770335,12.140307,11.555551,11.144334,11.140562,10.797253,10.506761,10.469034,10.453944,9.797507,9.525878,9.337247,9.265567,9.258021,9.186342,9.601331,9.940866,10.378491,10.725573,10.431308,9.42779,9.137298,8.654402,7.9413757,7.8432875,7.647111,7.960239,7.9753294,7.605612,7.4811153,7.356619,7.145352,6.820906,6.405917,5.96452,5.9796104,5.4740787,5.2892203,5.458988,5.2288585,4.1008434,3.832987,3.7084904,3.5764484,3.863168,3.651901,3.3350005,3.3274553,3.8971217,5.149633,5.572167,5.832478,6.115425,6.549277,7.2094865,6.349328,6.1342883,6.2625575,6.138061,4.8742313,3.270866,2.938875,3.651901,5.0741806,6.760544,5.413717,5.0741806,4.949684,4.6856003,4.353609,4.1498876,4.1536603,3.8254418,3.229367,3.0143273,3.2670932,3.7348988,4.1612053,4.4818783,4.8327327,4.5196047,3.9461658,3.4066803,3.1237335,3.2821836,3.4066803,3.5802212,4.168751,4.991183,5.300538,5.032682,4.4215164,3.7537618,3.3878171,3.7273536,4.851596,5.1873593,5.2665844,5.5382137,6.3342376,6.519096,7.6810646,8.812852,9.4127,9.473062,9.26934,9.058073,9.235386,9.740918,10.038955,10.170997,9.854096,9.665465,9.80128,10.072908,10.1294985,10.502988,10.487898,10.423763,11.710228,11.68382,10.816116,10.540714,10.850069,10.284176,9.378746,9.64283,10.069136,10.159679,9.918231,10.585986,11.2801485,11.385782,10.751981,9.703192,11.106608,11.589504,12.0082655,13.008011,15.015047,15.799753,16.244923,15.897841,14.883006,13.8870325,14.019074,14.007756,14.260523,14.822643,15.380992,15.482853,15.558306,15.663939,15.784663,15.826162,3.1576872,3.8895764,3.8254418,3.5047686,3.180323,2.837014,2.9124665,3.1576872,3.4142256,3.4632697,3.0369632,2.9992368,3.0633714,3.0822346,3.2935016,4.3196554,4.123479,4.1762958,4.7535076,5.4288073,5.0515447,5.330719,5.1081343,5.451443,6.628502,8.118689,9.495697,11.332966,12.377983,12.970284,15.045229,20.69662,27.76652,32.814293,33.161373,26.90259,32.38044,32.799202,24.744648,11.608367,3.6028569,3.199186,2.9615107,2.252257,1.1883769,0.6413463,0.47157812,0.27917424,0.1659955,0.21503963,0.52062225,0.482896,0.5357128,0.6451189,0.73566186,0.68661773,0.90543,1.1544232,1.5241405,1.9579924,2.2296214,3.6066296,3.7877154,3.3048196,2.886058,3.4481792,3.240685,3.0520537,3.0445085,3.3425457,4.014073,4.3686996,4.4101987,4.3121104,4.327201,4.7912335,4.6818275,3.9310753,3.4066803,3.3350005,3.3123648,3.1048703,3.1425967,3.0822346,2.6182017,1.4939595,0.9695646,0.63002837,0.5017591,0.49044126,0.38103512,0.17354076,0.150905,0.20372175,0.32821837,0.59607476,1.3166461,2.384299,3.591539,4.13857,2.625747,3.6745367,3.953711,3.3764994,2.7087448,3.6028569,4.515832,5.50426,7.043491,8.933576,10.299266,11.140562,10.985884,9.061845,5.9682927,3.663219,2.9049213,3.0181,3.5236318,3.8065786,3.097325,2.2183034,1.7618159,1.1016065,0.38858038,0.5357128,1.1317875,1.20724,1.026154,0.7054809,0.23013012,0.1659955,0.08677038,0.041498873,0.03772625,0.060362,0.24522063,0.56589377,1.0450171,1.5656394,1.8448136,2.4333432,3.3840446,4.8930945,6.458734,6.911449,7.4999785,8.899622,11.370691,15.430037,21.851044,21.692595,18.595268,17.112627,17.501207,15.731846,14.705692,14.468017,13.777626,12.898605,13.58145,12.51757,13.58145,13.788944,13.298503,15.411173,14.362384,15.901614,18.312323,19.840235,18.693357,17.923742,19.149845,21.088974,22.496162,22.156626,26.73282,31.116611,33.08215,32.916153,33.41791,34.72324,35.689034,36.10025,35.92671,35.338177,33.05574,34.236572,36.285107,38.725994,43.181465,43.44932,43.61909,42.551437,40.11055,37.171673,33.568817,32.350258,31.10152,29.39252,28.732311,25.499172,22.684793,21.183289,21.666185,24.597515,26.536644,28.61536,30.92798,33.25946,35.08164,37.15658,41.33665,46.42215,51.40956,55.510403,62.76139,64.22517,61.418335,56.676144,53.160057,51.500103,48.11983,43.939762,40.004917,37.492348,35.549446,35.67017,36.65105,37.318806,36.515236,35.892754,42.84193,49.689243,51.326565,45.21114,44.05294,49.621338,61.87105,77.14264,88.166245,79.572205,69.2918,59.58861,49.16485,33.187782,30.76953,29.543427,28.788902,27.125174,22.522572,22.473528,20.100546,16.678776,13.8719425,13.702174,15.607349,15.260268,14.2944765,13.93985,15.015047,15.63753,13.558814,13.924759,17.4333,20.33822,18.312323,17.395575,17.803017,20.240133,25.880207,36.756687,45.241318,42.99661,32.188038,25.499172,35.97198,39.514473,34.300705,24.069347,18.112373,14.879233,11.41219,7.9036493,4.8629136,3.127506,2.565385,2.0598533,1.5543215,1.2298758,1.50905,1.2525115,2.3805263,4.45547,6.4134626,6.5455046,6.092789,5.9909286,7.164215,9.507015,11.887542,12.498707,13.81158,13.532406,11.1631975,8.024373,6.379509,5.5985756,5.379763,5.5193505,5.934339,4.7044635,3.7801702,2.7502437,1.7165444,1.327964,1.4260522,1.2562841,1.1959221,1.2751472,1.1883769,1.1657411,1.2600567,1.4939595,1.8372684,2.2296214,2.1164427,4.2706113,5.832478,6.3945994,7.9791017,5.455216,5.089271,6.2851934,7.884786,8.179051,6.63982,5.6325293,4.889322,4.3385186,4.104616,5.3609,4.8629136,5.723072,7.707473,7.2170315,4.666737,4.7610526,5.8702044,6.971811,7.6282477,6.858632,6.221059,5.485397,4.749735,4.4101987,5.873977,6.4247804,5.5570765,3.4896781,1.1581959,0.41498876,0.1659955,0.18485862,0.2678564,0.24522063,0.049044125,0.08299775,0.1056335,0.049044125,0.0,1.2336484,0.97333723,3.108643,6.6058664,5.5080323,1.871222,0.5772116,1.3053282,2.5616124,1.6939086,3.097325,3.2746384,2.7200627,2.0372176,1.9542197,1.6222287,1.3505998,1.3053282,1.4600059,1.5731846,1.3996439,1.5769572,1.901403,2.5729303,4.195159,6.881268,9.540969,10.668983,10.642575,11.717773,11.668729,10.521852,9.544742,8.763808,6.9567204,6.749226,6.3342376,6.881268,7.3188925,4.304565,3.169005,1.9768555,1.0450171,0.6375736,0.9922004,1.0148361,0.8563859,0.7092535,0.91674787,1.9693103,2.2975287,2.252257,2.9803739,4.3875628,5.1571784,6.7077274,6.8925858,6.092789,4.98741,4.5460134,4.7912335,4.3121104,4.7346444,5.847569,5.613666,4.8968673,3.4066803,2.5767028,2.727608,3.0822346,3.399135,3.874486,4.398881,4.5988297,3.8292143,3.9159849,3.4594972,3.059599,2.6295197,1.4335974,1.5316857,1.6222287,1.7655885,1.7919968,1.267602,1.2298758,1.659955,2.0862615,2.3314822,2.5012503,2.8332415,2.3013012,1.8674494,2.1202152,3.2821836,5.330719,5.5797124,5.1835866,5.0854983,6.0286546,5.587258,5.50426,5.402399,5.070408,4.485651,3.863168,3.5877664,3.7952607,4.214022,4.164978,4.508287,3.742444,3.5274043,4.1272516,4.4101987,3.874486,4.8742313,5.6551647,5.2779026,3.6330378,5.3156285,4.9044123,5.715527,7.5527954,6.700182,6.466279,6.7643166,6.94163,7.0812173,7.9941926,8.544995,9.57115,10.27663,10.084227,8.605357,14.879233,13.585222,16.18456,19.844007,7.4169807,5.1081343,4.7346444,6.692637,9.5183325,9.87296,7.6131573,9.0807085,12.279895,13.588995,7.7678347,5.0439997,4.353609,5.9230213,8.028146,7.001992,7.175533,6.2927384,6.587003,8.073418,8.575176,8.967529,8.82417,9.314611,10.095545,9.337247,9.899368,10.552032,10.668983,10.352083,10.438853,10.144588,10.336992,11.257513,12.50248,13.015556,12.7477,12.770335,12.510024,11.812089,10.970794,10.763299,10.453944,10.144588,9.846551,9.507015,9.21275,9.314611,9.246704,9.065618,9.431562,9.159933,9.175024,9.6051035,10.235131,10.529396,9.612649,9.733373,9.510788,8.695901,8.14887,7.352846,7.1378064,7.2170315,7.4471617,7.8131065,7.677292,7.3151197,7.164215,7.194396,6.9265394,6.477597,6.0512905,5.8437963,5.7683434,5.462761,4.5950575,4.1612053,3.953711,3.8405323,3.7537618,3.4255435,2.867195,2.9313297,3.8292143,5.111907,5.5268955,6.217286,6.379509,6.1078796,6.379509,5.938112,5.3986263,5.2326307,5.1043615,3.8593953,2.9200118,3.2972744,4.5196047,6.1606965,7.858378,5.723072,5.2326307,4.9345937,4.436607,4.425289,4.398881,3.772625,3.259548,3.150142,3.2972744,3.187868,4.093298,4.8327327,4.957229,4.7610526,4.063117,3.663219,3.3689542,3.2067313,3.4029078,3.108643,3.108643,3.519859,4.1536603,4.5309224,4.508287,3.712263,3.097325,3.2255943,4.2894745,4.983638,4.983638,5.0025005,5.4174895,6.270103,7.5037513,8.809079,9.34102,9.239159,9.64283,9.752235,9.880505,10.26154,10.589758,10.038955,10.065364,10.106862,10.038955,10.170997,11.246195,10.453944,10.9594755,11.246195,10.989656,11.0613365,11.52537,11.174516,10.7557535,10.638803,10.834979,10.453944,10.789707,11.219787,11.332966,10.955703,11.408418,12.113899,12.370438,12.0724,11.717773,12.536433,13.328684,14.200161,15.113135,15.8676605,16.331694,16.776863,16.071383,14.437836,13.472044,13.585222,13.472044,13.645585,14.173752,14.709465,15.403628,15.98084,16.105335,16.180788,17.365393,3.4632697,4.0895257,3.9310753,3.5387223,3.2784111,3.338773,3.5575855,3.3576362,3.3651814,3.5802212,3.3764994,3.3236825,3.1237335,2.9728284,3.0633714,3.610402,3.6971724,4.195159,5.070408,6.0814714,6.7454534,6.7039547,6.2625575,6.7039547,7.9225125,8.43559,10.616167,12.989148,13.875714,14.177525,17.365393,23.348776,30.048958,33.942307,35.07032,37.02077,48.282055,46.23352,32.92747,15.471535,6.0286546,4.67051,3.6066296,2.565385,1.4864142,0.5055317,0.3961256,0.2867195,0.24899325,0.331991,0.56589377,0.452715,0.633801,0.8186596,1.0450171,1.7014539,2.3767538,2.6446102,3.0558262,3.772625,4.557331,4.727099,4.5535583,4.5497856,4.689373,4.398881,3.7160356,3.500996,3.7235808,4.1536603,4.3686996,4.644101,4.7044635,4.8968673,5.7306175,7.854605,6.270103,4.515832,3.0822346,2.1768045,1.7240896,2.6408374,3.8254418,3.8480775,2.6295197,1.4449154,0.8224323,0.49421388,0.38103512,0.3772625,0.34330887,0.18485862,0.20372175,0.33576363,0.6790725,1.4750963,2.0560806,3.0256453,4.29702,5.6287565,6.6020937,5.87775,4.659192,3.7009451,3.572676,4.640329,5.3382645,6.405917,7.8319697,9.152389,9.446653,9.495697,9.201432,8.213005,6.983129,6.7756343,4.8930945,3.5839937,2.8332415,2.7615614,3.6481283,3.832987,2.7841973,1.4562333,0.52439487,0.38858038,0.48666862,0.58475685,0.52439487,0.32067314,0.1659955,0.056589376,0.018863125,0.02263575,0.056589376,0.10940613,0.25276586,0.6375736,1.1883769,1.780679,2.2371666,2.8030603,3.8895764,4.957229,5.7607985,6.349328,7.141579,7.2094865,8.065872,10.699164,15.577168,17.429527,15.486626,14.241659,14.724555,14.48688,13.324911,12.958967,12.849561,12.857106,13.226823,13.12119,14.445381,15.264041,15.01882,14.543469,14.600059,14.7170105,15.935568,17.953922,19.119663,19.83269,20.251451,21.345512,23.499681,26.525326,29.882963,34.4667,37.952606,38.97876,37.175446,39.714424,38.235554,35.753166,34.342205,35.130684,32.418167,34.08944,36.63596,38.952354,42.35149,43.355007,43.622864,42.415623,40.106777,38.220463,35.55699,33.719723,32.357803,31.40333,31.075111,27.460938,24.959686,24.41643,25.404858,26.246153,30.188545,31.99186,33.41414,35.28159,37.458393,37.190536,40.25391,44.788605,49.421387,53.227966,61.15425,67.76012,69.55212,66.02848,59.69047,58.860497,54.4503,47.68598,40.434994,35.19482,32.327625,31.063795,31.788137,33.006695,31.350513,30.931753,33.27455,39.13344,46.16561,48.946037,47.248356,50.062733,59.305664,72.94748,85.016106,79.213806,71.23848,65.157005,58.72468,43.381416,35.24009,30.826118,28.736084,27.532618,25.733074,23.58268,22.49239,19.512016,15.316857,14.237886,16.086473,15.75071,14.498198,13.426772,13.4644985,15.143317,15.222542,15.803526,18.225552,23.073374,19.1423,17.527617,18.0671,20.032639,22.167944,30.807257,41.461147,44.418888,36.983044,23.446865,27.857063,32.82561,31.233562,23.620405,18.21046,13.743673,10.412445,6.934085,3.6556737,2.565385,2.123988,1.8334957,1.7618159,1.871222,2.0372176,1.8976303,2.2107582,3.4255435,5.040227,5.594803,5.934339,5.7570257,7.5188417,10.767072,12.14408,12.400619,13.63804,13.951167,12.294985,8.4544525,6.387054,5.4665337,5.5193505,5.9796104,5.885295,4.2328854,3.2067313,2.384299,1.7316349,1.5845025,1.388326,1.6373192,1.6448646,1.297783,1.056335,1.3053282,1.4901869,1.6335466,1.8070874,2.1164427,1.9693103,3.832987,5.3344917,5.9720654,7.1000805,6.379509,5.5306683,6.2436943,8.013056,8.130007,7.6282477,6.688864,5.832478,5.5797124,6.458734,5.3458095,4.719554,5.5759397,6.907676,5.715527,7.7640624,7.5075235,7.7602897,8.831716,8.533678,10.801025,9.027891,6.6134114,5.2288585,4.8365054,4.6327834,4.1272516,3.0633714,1.6373192,0.47535074,0.16222288,0.06413463,0.120724,0.19240387,0.060362,0.05281675,0.03772625,0.4640329,0.8978847,0.0,1.0186088,0.9318384,1.5920477,3.169005,4.142342,2.7691069,1.237421,0.7092535,1.0601076,0.875249,2.0070364,2.04099,1.8636768,1.7655885,1.4637785,1.9655377,1.991946,1.8184053,1.6524098,1.6448646,1.3770081,2.4823873,3.2142766,3.4594972,4.719554,7.3377557,9.084481,10.272858,10.970794,10.997202,11.125471,11.076427,10.710483,9.759781,7.835742,8.243186,8.156415,8.526133,8.503497,5.4363527,3.9612563,2.2899833,1.0978339,0.83752275,1.7467253,1.5769572,1.2298758,0.995973,1.056335,1.4939595,1.8523588,2.1353056,2.9501927,4.3385186,5.7796617,5.96452,6.3342376,5.824933,4.6742826,4.447925,4.564876,4.398881,4.640329,5.281675,5.613666,4.847823,3.169005,2.3578906,2.6219745,2.6068838,3.2369123,4.014073,4.6742826,4.957229,4.5988297,3.8141239,3.2369123,2.957738,2.7087448,1.8749946,1.8259505,1.7655885,1.961765,2.282438,2.2069857,1.5656394,1.5656394,1.8146327,2.0485353,2.11267,2.335255,2.2447119,2.1541688,2.546522,4.085753,4.7308717,4.708236,4.8553686,5.2665844,5.2590394,5.081726,4.8968673,4.7120085,4.323428,3.338773,3.3010468,3.2633207,3.3576362,3.5123138,3.4444065,4.0706625,3.5236318,3.2821836,3.802806,4.4818783,4.5724216,5.194905,5.5004873,5.323174,5.168496,5.2628117,4.3875628,4.7006907,6.0701537,6.0776987,5.9607477,6.3832817,6.9680386,7.5905213,8.397863,7.9526935,9.205205,9.771099,9.861642,12.291212,10.461489,10.823661,13.539951,14.566105,5.6476197,3.6028569,4.0103,5.847569,7.673519,7.6395655,6.960493,6.900131,7.779153,9.027891,9.171251,6.25124,5.040227,5.915476,7.5905213,7.1000805,5.904158,5.4212623,6.25124,7.7338815,7.9413757,8.29223,8.303548,8.948667,9.869187,9.374973,9.469289,9.857869,9.865415,9.49947,9.446653,9.0957985,9.763554,10.963248,12.076173,12.344029,12.728837,12.736382,12.608112,12.283667,11.363147,10.997202,10.834979,10.27663,9.548513,9.665465,9.839006,10.159679,10.137043,9.922004,10.295494,9.178797,8.627994,8.884532,9.65792,10.137043,9.631512,9.318384,9.133525,8.835487,8.013056,6.779407,6.3153744,6.3644185,6.809588,7.654656,7.665974,7.586749,7.647111,7.745199,7.4773426,7.201941,6.820906,6.40969,5.938112,5.292993,4.5233774,4.2517486,4.104616,3.893349,3.5839937,3.127506,3.0407357,3.3764994,4.0895257,5.0515447,5.621211,5.9682927,6.115425,6.156924,6.2814207,5.6853456,5.089271,4.432834,3.6292653,2.5804756,2.584248,3.470815,4.9421387,6.519096,7.5527954,6.119198,5.587258,5.1458607,4.659192,4.6554193,4.5724216,4.236658,3.7801702,3.482133,3.783943,3.7537618,4.376245,4.5422406,4.0895257,3.8443048,3.6179473,3.5651307,3.3651814,2.969056,2.6106565,2.71629,2.8332415,2.9086938,3.0445085,3.470815,2.987919,2.6295197,2.7200627,3.3048196,4.1536603,4.61392,4.7535076,4.8063245,5.3382645,7.2472124,8.695901,9.14107,9.0543,9.220296,10.70671,11.438599,11.219787,11.242422,11.472552,10.638803,11.121698,11.189606,10.917976,10.612394,10.804798,10.4049,10.208723,10.193633,10.367173,10.782163,10.876478,11.125471,11.208468,11.057564,10.884023,11.080199,11.457462,11.947904,12.253486,11.846043,11.898859,12.668475,12.996693,12.58925,12.012038,13.162688,13.743673,13.890805,13.849306,13.93985,15.0376835,15.437581,14.649103,13.336229,13.340002,13.389046,13.340002,13.543724,14.147344,15.07541,16.173243,16.637276,16.991903,17.621931,18.757492,3.832987,3.7499893,3.6481283,3.4179983,3.1652324,3.199186,3.2218218,3.059599,3.0407357,3.1048703,2.795515,2.837014,2.7200627,2.71629,2.9237845,3.2784111,3.591539,4.1083884,4.8629136,5.6815734,6.1833324,6.6020937,6.477597,6.779407,7.5829763,8.047009,10.133271,12.857106,14.588741,15.724301,18.648085,24.065575,28.249416,31.271288,35.160866,43.928444,55.38968,50.496586,35.300453,18.350048,10.691619,7.3717093,5.1232247,3.097325,1.2600567,0.4074435,0.422534,0.32821837,0.27540162,0.3169005,0.3961256,0.38103512,0.5055317,0.6526641,0.935611,1.7165444,2.2447119,2.5125682,2.969056,3.9386206,5.5985756,6.368191,6.722818,6.258785,5.142088,4.146115,3.651901,3.6292653,4.164978,4.9119577,5.05909,5.3382645,4.8025517,4.606375,5.247721,6.579458,6.217286,4.7874613,3.3048196,2.2786655,1.6939086,2.444661,4.2027044,4.8855495,3.9989824,2.6332922,2.2484846,1.8787673,1.6033657,1.418507,1.2147852,0.995973,0.8903395,0.8941121,1.0789708,1.5656394,2.0787163,2.776652,4.293247,6.507778,8.52236,7.7414265,5.194905,3.7801702,4.285702,5.409944,5.6551647,5.9796104,7.032173,8.314865,8.216777,7.5037513,6.7341356,6.1418333,6.1116524,7.1679873,5.5797124,4.930821,3.7537618,2.3390274,2.7125173,3.7801702,3.0218725,1.7391801,0.7997965,0.633801,0.33953625,0.23390275,0.211267,0.21503963,0.20749438,0.18863125,0.150905,0.14335975,0.16222288,0.15845025,0.16976812,0.3055826,0.62248313,1.0714256,1.5279131,2.2220762,3.3048196,4.353609,5.138315,5.613666,6.4511886,6.7831798,7.0284004,7.699928,9.4013815,10.834979,11.155652,10.982111,11.18206,12.875969,12.67602,12.0724,12.294985,13.381501,14.219024,13.898351,15.041456,15.950659,16.192106,16.59955,14.70192,15.275358,16.403374,17.625704,19.911915,19.923233,20.670212,21.892544,23.318596,24.688059,29.21898,35.60226,39.948326,41.04239,40.378407,40.29918,37.292397,34.32334,33.749905,37.32258,37.907337,38.680725,39.065533,39.56352,41.740322,43.40782,42.81552,41.928955,41.5781,41.438515,40.401043,38.507183,35.90407,33.08215,30.875162,28.24187,26.529099,26.800728,28.415411,29.011486,32.26726,34.379932,36.424694,38.480774,39.631424,39.60879,41.310246,44.07935,47.67089,52.216904,58.377598,64.88161,70.110466,72.245766,69.24276,63.327282,55.55945,46.844685,38.707134,33.28587,30.082912,27.936289,27.687294,28.449366,27.615616,27.313805,27.362848,30.546946,37.545162,46.90505,50.08537,53.054424,58.717136,68.322235,81.46229,80.19092,73.07952,67.28099,64.02899,58.62659,46.690006,36.398285,29.913143,27.245897,26.280106,23.533634,24.442837,23.08092,18.414183,14.317112,16.422237,16.912678,16.893814,16.271332,13.736128,14.490653,15.739391,17.165443,19.757236,25.816072,19.647831,17.184307,17.667202,19.564833,20.60985,26.917679,36.00216,41.06502,37.933743,25.065321,21.87368,23.284641,22.990377,19.323385,15.24895,12.095036,9.035437,6.0739264,3.640583,2.6182017,1.8749946,1.7127718,1.6637276,1.6675003,2.093807,2.848332,3.0822346,3.3236825,3.9310753,5.070408,5.6325293,5.5457587,7.0774446,10.559577,14.377474,14.758509,15.328176,15.015047,13.268322,10.069136,7.5112963,6.2436943,5.783434,5.836251,6.3153744,4.7308717,3.1614597,2.1051247,1.690136,1.6939086,1.4562333,1.6825907,1.7429527,1.478869,1.2525115,1.5920477,1.7391801,1.841041,1.9127209,1.8146327,1.9051756,4.6290107,5.9418845,5.111907,4.7044635,3.893349,3.9386206,4.666737,5.5004873,5.4363527,5.666483,5.4288073,5.6891184,6.7756343,8.405409,5.670255,5.0213637,5.3571277,5.8098426,5.7607985,7.443389,7.1906233,7.356619,7.888559,6.3417826,7.54525,6.1342883,4.6214657,4.266839,5.081726,3.7537618,2.2786655,1.1506506,0.5055317,0.13204187,0.049044125,0.033953626,0.06413463,0.08299775,0.00754525,0.02263575,0.011317875,0.23767537,0.47535074,0.0,1.0223814,1.2600567,1.056335,0.98842776,1.841041,2.9011486,1.9089483,0.9280658,0.7884786,1.0827434,1.5731846,2.0183544,2.4408884,2.6106565,2.0296721,2.1164427,3.2557755,3.270866,2.071171,1.6524098,1.3543724,1.9957186,3.0030096,4.3347464,6.507778,7.4471617,8.880759,10.585986,11.740409,10.93684,10.442626,10.616167,10.77839,10.510533,9.650374,9.465516,9.6051035,9.646602,9.012801,6.9869013,5.59103,3.3274553,1.5279131,0.9620194,1.8372684,1.9164935,1.7580433,1.5354583,1.4562333,1.7580433,1.8825399,2.1503963,2.704972,3.572676,4.67051,4.45547,4.8742313,4.8025517,4.134797,3.802806,4.406426,4.1800685,4.221567,4.7874613,5.2779026,4.6856003,3.1237335,2.2711203,2.4295704,2.5314314,3.138824,3.7877154,4.2894745,4.5799665,4.727099,3.9989824,3.3161373,3.1350515,3.1614597,2.3503454,2.2409391,2.1466236,2.0749438,2.0372176,2.0749438,1.8825399,1.8749946,1.9391292,1.9768555,1.8938577,2.033445,2.1805773,2.3616633,2.8785129,4.315883,4.606375,4.3800178,4.402653,4.738417,4.727099,4.4705606,4.093298,3.7348988,3.4179983,3.0331905,3.3350005,3.0860074,2.9351022,3.0860074,3.3312278,3.7386713,3.942393,3.8858037,3.8782585,4.6026025,4.8402777,5.4740787,5.7079816,5.4891696,5.5268955,4.9723196,4.930821,5.270357,5.6287565,5.4174895,6.0550632,6.4549613,7.009537,7.6508837,7.877241,7.7150183,8.643084,9.039209,9.827688,14.475562,10.808571,8.805306,9.193887,9.710737,5.1043615,5.13077,5.0439997,5.945657,7.3490734,7.1981683,6.017337,4.708236,4.7535076,6.7341356,10.344538,6.579458,5.194905,5.613666,6.5266414,5.8702044,5.2137675,5.5985756,6.2889657,6.9567204,7.654656,8.126234,8.20546,8.654402,9.382519,9.439108,9.420244,9.57115,9.514561,9.265567,9.246704,8.98262,9.49947,10.140816,10.657665,11.216014,11.932813,12.162943,12.366665,12.506252,12.034674,11.68382,11.563096,10.880251,9.963503,10.26154,10.63503,10.982111,10.902886,10.431308,10.008774,8.986393,8.578949,8.76758,9.288202,9.590013,9.65792,9.156161,8.729855,8.492179,8.016829,7.0246277,6.507778,6.470052,6.851087,7.5226145,7.835742,8.009283,7.91874,7.6131573,7.33021,7.0548086,6.63982,6.1305156,5.624984,5.292993,4.8742313,4.779916,4.61392,4.2064767,3.640583,3.048281,3.2218218,3.6783094,4.3083377,5.383536,5.926794,6.096562,5.926794,5.621211,5.560849,5.1458607,4.6252384,3.7462165,2.6182017,1.7165444,2.5540671,3.3764994,4.52715,5.753253,6.205968,5.0854983,4.7572803,4.825187,4.881777,4.5309224,4.266839,4.1197066,3.942393,3.9159849,4.557331,5.0779533,4.8742313,4.3347464,3.7613072,3.350091,2.9992368,3.0143273,3.0256453,2.7691069,2.071171,2.0673985,2.474842,2.7313805,2.6823363,2.6106565,2.3918443,2.655928,3.4217708,4.376245,4.8629136,5.0138187,5.0553174,4.859141,5.028909,6.8774953,8.650629,9.050528,9.0807085,9.714509,11.895086,11.672502,10.295494,9.805053,10.393582,10.419991,10.529396,10.427535,10.616167,10.9594755,10.687846,10.20495,9.820143,9.989911,10.601076,10.967021,10.47658,10.884023,11.415963,11.646093,11.480098,11.887542,12.381755,12.698656,12.611885,11.9064045,11.872451,12.649611,13.377728,13.332457,11.921495,11.959221,12.672247,13.215506,13.434318,13.841762,14.520834,14.747191,14.222796,13.536179,14.18507,14.1926155,14.049255,14.234114,14.871688,15.735619,16.45619,16.878725,17.7917,19.146072,20.066593,3.802806,3.3010468,3.2142766,3.138824,2.9728284,2.9237845,2.9652832,2.897376,2.806833,2.6597006,2.3126192,2.584248,2.5276587,2.584248,2.8898308,3.2972744,3.5953116,4.036709,4.6252384,5.2250857,5.564622,6.0550632,6.1644692,6.4436436,7.032173,7.673519,9.386291,11.615912,13.826671,16.275105,19.99114,24.827644,28.189054,30.735577,34.719467,43.988808,52.51494,45.77703,31.59196,17.912424,12.804289,8.27714,5.0666356,2.5993385,0.8563859,0.35462674,0.38103512,0.31312788,0.26408374,0.2867195,0.3734899,0.4376245,0.5885295,0.814887,1.1619685,1.7467253,2.071171,2.5276587,3.0671442,3.9386206,5.674028,6.4436436,7.1679873,6.587003,4.9949555,4.217795,4.4705606,4.8402777,5.2137675,5.4476705,5.372218,5.8626595,5.0138187,4.3875628,4.459243,4.606375,4.6742826,3.9084394,3.3538637,3.361409,3.6028569,3.5424948,4.678055,5.2250857,4.564876,3.2746384,2.686109,2.335255,1.9429018,1.4901869,1.2223305,1.1581959,1.086516,1.0525624,1.1544232,1.5580941,2.3692086,3.097325,4.5724216,6.7114997,8.529905,7.9300575,5.775889,4.798779,5.583485,6.5756855,6.4926877,6.673774,7.7376537,8.831716,7.594294,6.096562,5.6853456,6.270103,7.3490734,8.009283,7.062354,7.2887115,6.017337,3.4217708,2.5427492,4.085753,3.6028569,2.2786655,1.1204696,0.97710985,0.47912338,0.16222288,0.16222288,0.32444575,0.18863125,0.23390275,0.17731337,0.18863125,0.25276586,0.18863125,0.08299775,0.06413463,0.21881226,0.60362,1.2298758,1.9994912,2.9426475,4.0970707,5.2099953,5.7079816,5.794752,6.0776987,6.3342376,6.488915,6.620957,7.748972,9.684328,10.767072,11.076427,12.4307995,13.441863,12.808062,12.528888,13.415455,15.109364,14.871688,15.064092,15.667711,16.769318,18.534906,16.739138,18.357594,19.764782,20.266542,22.111355,22.152855,22.428255,23.039421,23.778856,24.114618,27.366621,33.72727,38.065784,39.540882,41.59319,40.89903,37.692295,34.77983,34.591198,39.186256,42.01195,41.917637,41.068794,40.94807,42.347717,43.400276,42.39676,41.944046,42.864567,44.21139,43.528545,41.502647,38.394005,34.76474,31.456148,29.683014,28.619133,29.041668,30.580898,31.708914,33.267006,34.87792,37.175446,39.631424,40.533085,41.366833,42.823067,44.905556,47.78407,51.760414,56.823277,62.365265,67.56771,71.37807,72.50985,64.82879,55.0841,45.369587,37.458393,32.765247,29.607561,27.01954,25.589716,25.1785,24.899324,24.838963,24.314568,25.32186,29.977278,40.529312,49.157303,54.808697,59.05667,64.64393,75.50154,79.1459,74.20376,67.948746,65.38714,69.235214,62.508625,50.907803,39.069305,30.25268,26.34424,23.903353,25.431265,25.306768,21.322876,14.698147,16.124199,16.867407,18.417955,19.247932,14.803781,14.2077055,16.233604,18.542452,21.368149,27.525072,21.31533,17.716248,17.670975,19.757236,20.179771,24.933279,30.55449,34.81001,34.572334,25.8123,18.448135,15.943113,15.362129,14.57365,12.2270775,10.035183,7.488661,5.3873086,4.0517993,3.2972744,2.757789,2.886058,2.3918443,1.4675511,1.7882242,3.0105548,3.3576362,3.048281,2.9237845,4.432834,6.017337,5.9682927,6.4738245,8.990166,14.25675,16.678776,17.067356,16.24115,14.641558,12.3289385,9.480607,7.635793,6.3719635,5.670255,5.9494295,5.0251365,3.429316,2.2673476,1.8749946,1.8297231,1.6184561,1.6863633,1.6712729,1.5354583,1.5731846,1.9278114,1.9957186,2.161714,2.5993385,3.2633207,2.5276587,5.1458607,6.432326,5.2326307,3.9273026,2.6672459,3.2670932,4.093298,4.3196554,3.9197574,4.8025517,4.568649,4.7836885,5.8966126,7.220804,5.7607985,5.481624,5.243949,5.032682,5.975838,6.1305156,6.1229706,6.398372,6.379509,4.447925,4.1083884,3.3953626,3.0105548,3.2520027,3.9763467,2.3126192,0.9205205,0.181086,0.049044125,0.056589376,0.06413463,0.041498873,0.03772625,0.0452715,0.0,0.0,0.0,0.0150905,0.030181,0.0,0.6375736,1.1506506,1.0110635,0.41876137,0.32067314,2.1315331,1.9164935,1.1732863,0.87147635,1.4449154,1.4864142,2.2786655,2.9992368,3.1199608,2.4333432,2.3428001,3.5085413,3.7235808,2.637065,1.7467253,1.5882751,1.8033148,2.9237845,4.919503,7.194396,7.745199,9.201432,10.884023,11.800771,10.680302,10.303039,10.691619,10.93684,10.823661,10.868933,10.616167,10.238904,9.846551,9.205205,7.7376537,6.5040054,4.4139714,2.4672968,1.4750963,2.052308,1.9542197,1.9278114,1.8184053,1.7089992,1.9278114,2.1277604,2.1881225,2.5880208,3.1652324,3.1463692,3.1048703,3.7160356,4.08198,3.893349,3.429316,4.0782075,3.9197574,4.032936,4.6327834,5.0741806,4.3347464,3.0407357,2.233394,2.1994405,2.4786146,2.9426475,3.451952,3.9273026,4.2592936,4.3196554,4.1612053,3.6669915,3.4896781,3.470815,2.6597006,2.6219745,2.565385,2.3088465,1.9806281,2.033445,2.0070364,2.0447628,2.093807,2.0598533,1.8334957,1.8938577,2.1843498,2.5804756,3.1010978,3.8895764,4.5196047,4.255521,3.9612563,3.983892,4.191386,3.893349,3.4142256,3.0633714,2.9652832,3.0520537,3.1954134,2.8822856,2.7426984,2.9841464,3.4029078,3.8065786,4.2630663,4.247976,4.063117,4.8100967,5.198677,5.692891,5.704209,5.2099953,4.768598,4.3121104,5.0062733,5.5004873,5.323174,4.8629136,5.885295,6.398372,6.881268,7.352846,7.356619,8.069645,8.3525915,8.047009,8.880759,14.441608,12.932558,11.374464,9.020347,6.587003,6.25124,6.971811,7.1906233,6.94163,6.7341356,7.5792036,6.013564,4.0216184,3.289729,4.496969,7.3188925,6.398372,5.6513925,5.7872066,6.2399216,5.168496,5.251494,6.066381,6.5266414,6.719045,7.911195,8.409182,8.303548,8.420499,8.850578,8.944894,8.937348,8.907167,8.805306,8.699674,8.763808,8.650629,8.899622,9.148616,9.386291,9.922004,10.616167,11.212241,11.857361,12.362892,12.189351,12.23085,12.147853,11.389555,10.382264,10.544487,10.997202,11.234878,11.129244,10.533169,9.314611,8.827943,8.744945,8.865668,9.103344,9.476834,9.805053,8.993938,8.152642,7.828197,7.9941926,7.432071,6.9755836,6.9152217,7.2358947,7.6131573,7.726336,7.9715567,7.7602897,7.175533,6.971811,6.851087,6.4021444,5.9494295,5.7117543,5.836251,5.2892203,5.0779533,4.817642,4.323428,3.5990841,2.9916916,3.4029078,3.8820312,4.2404304,5.0553174,5.5382137,5.7306175,5.6287565,5.406172,5.3948536,4.8327327,4.2328854,3.3274553,2.3201644,1.8900851,2.837014,3.3915899,4.134797,4.98741,5.198677,4.3611546,4.3309736,4.6252384,4.776143,4.3196554,4.063117,3.802806,3.8405323,4.2781568,5.0138187,5.3156285,4.779916,4.0404816,3.440634,3.0218725,2.6785638,2.6295197,2.6483827,2.4597516,1.7542707,1.8976303,2.5012503,2.806833,2.6408374,2.4182527,2.7087448,3.470815,4.4403796,5.27413,5.5382137,5.4665337,5.5683947,5.3948536,5.406172,6.983129,8.7751255,9.465516,9.782416,10.325675,11.589504,11.283921,9.933322,9.408927,9.9257765,10.054046,9.703192,9.680555,10.133271,10.638803,10.231359,9.880505,9.488152,9.869187,10.782163,10.906659,10.235131,10.79348,11.61214,12.042219,11.747954,12.264804,12.645839,12.762791,12.464753,11.5857315,11.442371,12.106354,13.102326,13.536179,12.1101265,11.189606,11.812089,12.608112,13.083464,13.611631,14.2944765,14.520834,14.181297,13.717264,14.136025,14.520834,14.618922,14.894323,15.418718,15.916705,16.429781,16.965494,17.987877,19.353567,20.315586,3.3312278,2.9916916,2.8558772,2.8294687,2.8256962,2.7917426,3.006782,2.9916916,2.8219235,2.584248,2.384299,2.7992878,2.6597006,2.584248,2.8219235,3.2859564,3.5047686,3.9348478,4.52715,5.1798143,5.726845,5.783434,5.8966126,6.2625575,6.8925858,7.6282477,8.907167,9.944639,11.951676,15.62244,21.149336,25.944342,29.93578,31.750412,32.75393,37.05095,41.717686,34.4667,22.97906,13.385274,10.284176,6.33801,3.2859564,1.4977322,0.80734175,0.51684964,0.44139713,0.392353,0.33953625,0.331991,0.5017591,0.60362,0.845068,1.1996948,1.6146835,2.0145817,2.3616633,3.1840954,3.8895764,4.436607,5.349582,5.3382645,5.783434,5.560849,4.7610526,4.696918,5.4891696,6.187105,6.149379,5.4967146,5.1043615,5.80607,5.1081343,4.425289,4.2328854,4.0480266,3.218049,2.8709676,3.4142256,4.7836885,6.428553,6.205968,6.0739264,5.511805,4.4818783,3.4557245,2.2183034,1.9202662,1.599593,1.0827434,1.0035182,1.2864652,1.1883769,1.0072908,1.0638802,1.6863633,3.048281,4.22534,5.3986263,6.530414,7.3679366,6.828451,6.198423,6.1003346,6.63982,7.424526,7.594294,8.375228,9.476834,9.782416,7.356619,5.6061206,6.307829,8.265821,9.895596,9.220296,8.605357,8.937348,8.0206,5.802297,4.346064,5.704209,4.9949555,3.3840446,1.9466745,1.6373192,0.8563859,0.43007925,0.44894236,0.6111652,0.23013012,0.18863125,0.1961765,0.241448,0.2678564,0.17354076,0.033953626,0.03772625,0.181086,0.5696664,1.4222796,2.4295704,3.4934506,5.05909,6.628502,6.760544,5.43258,5.304311,5.7683434,6.304056,6.477597,8.126234,10.785934,12.653384,13.20796,13.238141,14.694374,14.196388,13.215506,13.192869,15.554533,15.55076,14.520834,14.962231,17.365393,20.206179,20.194862,22.009495,23.356321,23.892035,25.227543,26.215971,25.235088,24.74842,25.58217,26.951633,26.536644,29.969732,33.297188,36.01725,41.080112,42.2534,40.148273,37.416893,36.60201,40.14073,42.81552,42.653297,42.42317,43.094696,43.837902,43.47573,43.026787,43.01547,43.868084,45.909073,44.705605,42.909836,40.495358,37.601753,34.53461,32.81052,31.916407,32.010723,33.02556,34.644016,34.949596,34.817554,36.036114,38.394005,39.66915,41.41965,43.958626,46.814503,49.54211,51.75664,56.498833,61.24102,63.806408,64.65525,66.88864,62.610485,54.005127,44.875374,37.72625,33.72727,30.99966,28.28337,25.948114,24.307022,23.609087,23.61286,23.273323,23.394047,25.687803,32.79543,44.226482,53.32228,58.947266,62.697254,68.90322,76.00707,74.42258,68.182655,63.851677,70.54431,74.85642,69.71056,55.70658,38.295918,27.762747,24.944597,25.087955,25.472763,23.307278,15.743164,15.47908,15.83748,18.135008,20.153362,16.135517,14.268067,16.358103,19.161163,22.133991,27.411894,23.182781,18.817854,18.368912,20.892797,20.443855,24.714466,27.611843,29.758467,29.95087,25.15209,17.546478,12.702429,10.846297,10.884023,10.427535,8.299775,6.3455553,5.062863,4.8138695,5.824933,5.372218,5.6400743,4.5988297,2.4974778,1.8599042,2.505023,2.7389257,2.323937,1.9881734,3.4368613,6.4738245,6.587003,6.092789,7.043491,11.219787,16.105335,17.184307,16.72782,15.803526,14.302021,11.589504,9.276885,7.3905725,5.975838,5.0553174,4.7308717,3.7047176,2.7653341,2.252257,2.0560806,1.8636768,1.7919968,1.6448646,1.5241405,1.841041,2.1692593,2.1692593,2.5502944,3.5990841,5.1571784,3.1425967,4.29702,5.4891696,5.409944,4.5460134,3.4745877,3.8443048,4.640329,5.0062733,4.2404304,5.560849,5.1345425,4.4177437,4.115934,4.164978,5.7117543,5.938112,5.3458095,4.870459,5.8702044,5.292993,5.406172,5.4438977,4.908185,3.5500402,2.9011486,2.7200627,2.7087448,2.535204,1.8146327,0.59607476,0.13204187,0.0150905,0.02263575,0.10940613,0.11317875,0.07922512,0.08299775,0.10186087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.52062225,0.94315624,0.875249,0.12826926,1.116697,1.4071891,1.1921495,0.97710985,1.599593,1.6373192,2.5276587,3.078462,2.867195,2.2673476,2.535204,2.7351532,3.0331905,3.1350515,2.2786655,1.8900851,2.0145817,3.108643,4.908185,6.436098,8.20546,9.971047,11.16697,11.378237,10.329447,10.718028,11.389555,11.295239,10.680302,11.076427,11.59705,10.344538,9.2844305,8.722309,7.303802,6.013564,4.8968673,3.6066296,2.5087957,2.6898816,1.8976303,1.720317,1.7089992,1.7014539,1.8334957,2.505023,2.384299,2.6936543,3.1916409,2.2107582,2.3692086,3.0520537,3.640583,3.7688525,3.3236825,3.6292653,3.731126,4.1008434,4.6818275,4.9044123,3.9801195,2.969056,2.2484846,2.0296721,2.3654358,2.674791,3.150142,3.742444,4.115934,3.6481283,4.055572,4.0480266,3.874486,3.5387223,2.806833,2.867195,2.8747404,2.6483827,2.3163917,2.3390274,1.991946,1.9693103,2.082489,2.123988,1.841041,1.841041,2.1654868,2.746471,3.2935016,3.2972744,4.085753,3.9574835,3.5764484,3.3878171,3.6028569,3.3727267,3.006782,2.8898308,3.0369632,3.1312788,2.9086938,2.8256962,2.8709676,3.0746894,3.4896781,3.92353,3.9876647,3.9310753,4.085753,4.870459,5.5080323,5.4174895,5.040227,4.5497856,3.8593953,3.5462675,4.353609,4.908185,4.8025517,4.617693,5.342037,5.8702044,6.432326,6.911449,6.828451,8.499724,8.45068,7.4207535,7.8508325,13.890805,14.290704,15.890297,11.951676,5.1534057,7.5716586,7.586749,9.088254,8.314865,6.1531515,8.103599,7.2396674,5.455216,4.0782075,3.4745877,3.0520537,6.1531515,5.9607477,6.043745,6.8058157,5.50426,5.794752,6.3644185,6.7077274,7.0812173,8.503497,8.771353,8.382772,8.137552,8.171506,7.9338303,7.8961043,7.7716074,7.665974,7.6508837,7.7716074,7.8131065,7.967784,8.280911,8.635539,8.771353,9.216523,10.084227,11.053791,11.778135,11.910177,12.370438,12.253486,11.480098,10.56335,10.593531,10.982111,10.963248,10.77839,10.284176,8.963757,8.914713,8.835487,8.831716,9.065618,9.7296,10.03141,8.865668,7.647111,7.2585306,8.028146,7.6697464,7.3717093,7.326438,7.4999785,7.6093845,7.3490734,7.54525,7.3717093,6.8435416,6.8435416,7.069899,6.587003,6.277648,6.3945994,6.587003,5.5457587,5.0062733,4.647874,4.195159,3.4142256,2.9766011,3.5500402,4.0216184,4.0782075,4.195159,4.5837393,4.870459,5.1458607,5.4476705,5.7683434,4.8365054,4.044254,3.2746384,2.7125173,2.8445592,3.2444575,3.5689032,4.112161,4.768598,5.0062733,4.432834,4.5497856,4.5837393,4.3083377,4.0782075,4.0216184,3.591539,3.7348988,4.485651,4.957229,4.3385186,4.0480266,3.610402,3.0105548,2.7125173,2.6483827,2.5314314,2.3578906,2.0975795,1.7089992,2.3767538,2.9426475,2.9841464,2.6672459,2.746471,3.482133,4.353609,4.9723196,5.300538,5.6853456,5.6400743,6.096562,6.25124,6.3455553,7.677292,9.114662,9.978593,10.412445,10.514306,10.329447,11.042474,10.925522,10.842525,10.804798,9.944639,9.431562,9.631512,9.967276,10.0465,9.646602,9.582467,9.322156,9.756008,10.646348,10.627484,10.238904,11.016065,11.838497,12.042219,11.400873,12.027128,12.264804,12.351574,12.2119875,11.449917,11.246195,11.574413,12.347801,12.996693,12.449662,11.216014,11.532914,12.238396,12.755245,13.098554,14.083209,14.385019,14.086982,13.502225,13.155144,14.064346,14.784918,15.343266,15.686575,15.675257,16.165699,16.72782,17.346529,18.18028,19.595015,2.806833,2.9049213,2.7540162,2.7125173,2.8294687,2.8521044,2.7087448,2.9539654,3.0520537,2.9086938,2.8822856,2.9086938,2.6597006,2.463524,2.444661,2.516341,3.1161883,3.6141748,4.432834,5.4703064,6.119198,6.1908774,6.3945994,6.6058664,6.9567204,7.8131065,8.446907,8.533678,10.382264,14.690601,20.53817,26.057522,27.819336,27.196854,25.989614,26.427238,28.28337,21.160654,12.053536,5.5382137,3.7537618,2.4710693,1.931584,1.8749946,1.8599042,1.237421,1.1016065,0.95824677,0.7432071,0.513077,0.42630664,0.66020936,0.76207024,0.94692886,1.3317367,1.9542197,2.5616124,3.6971724,4.7044635,5.2779026,5.4476705,5.885295,5.5193505,5.0553174,4.708236,4.195159,3.9650288,4.346064,4.67051,4.689373,4.5761943,4.919503,4.3385186,4.1536603,4.7308717,5.462761,4.8402777,4.4818783,4.5912848,5.515578,7.7376537,9.933322,9.631512,8.031919,6.217286,5.142088,3.5802212,3.218049,3.218049,3.2746384,3.6179473,4.055572,3.0935526,2.003264,1.4901869,1.7089992,3.3463185,5.1534057,6.307829,6.587003,6.379509,6.5228686,5.836251,5.168496,5.081726,5.873977,7.413208,8.439363,8.182823,6.94163,6.0739264,5.7683434,6.964266,8.0206,8.156415,7.462252,6.643593,6.1833324,6.858632,8.167733,8.299775,8.507269,7.001992,5.379763,4.274384,3.3727267,1.5543215,1.1242423,1.1506506,1.0714256,0.7167987,0.362172,0.7054809,0.68661773,0.19994913,0.0754525,0.0150905,0.0,0.030181,0.21503963,0.76207024,2.7653341,5.0213637,7.9526935,10.080454,8.039464,5.515578,6.4134626,6.828451,5.5759397,4.195159,6.0286546,9.789962,11.310329,11.016065,13.947394,13.909668,13.324911,13.264549,14.260523,16.31283,14.920732,13.747445,15.109364,19.251705,24.367384,21.964222,21.519053,21.805773,23.118647,27.268534,27.509981,26.502691,26.623415,28.309778,30.030094,28.539907,27.389257,28.622906,33.1576,40.78585,41.423424,41.242336,39.842693,38.820312,41.76296,44.00767,44.698063,45.207367,45.58463,44.56979,44.18121,44.815014,45.41486,46.044888,47.91234,48.048153,48.36505,46.87864,43.543636,40.23882,37.809246,36.568054,36.783092,38.111057,39.612564,40.35577,37.779068,36.50769,37.315033,37.09245,40.71794,44.73956,48.25942,50.89271,52.733753,55.053917,56.785553,58.113514,58.453053,56.487514,55.219913,50.64372,44.630154,38.963673,35.338177,33.666904,30.950615,28.430502,26.551735,24.963459,24.061802,23.303505,23.235598,24.578651,28.230553,38.22801,48.36128,56.68746,62.67839,67.23195,73.99249,73.96986,68.00911,61.20707,62.927383,70.66504,78.8705,72.076004,50.89271,31.995632,25.578398,23.201643,24.239115,24.740875,17.440845,15.524352,16.105335,17.225805,17.80679,17.686066,14.109617,14.275613,16.923996,20.85507,24.933279,21.809546,18.5085,19.247932,22.60557,21.53037,26.14429,30.501673,32.25217,30.656351,26.581915,18.68204,12.321393,8.643084,7.888559,9.416472,8.243186,6.549277,5.3910813,6.571913,12.649611,10.001229,9.367428,8.424272,6.330465,3.6934,2.6672459,2.2560298,1.6863633,1.2261031,2.1654868,4.949684,5.9305663,6.092789,6.5455046,8.499724,11.819634,14.188843,15.1395445,14.962231,14.694374,12.706201,10.725573,8.873214,7.1566696,5.4476705,4.2517486,3.5839937,3.0181,2.4974778,2.3503454,2.1654868,2.003264,1.8976303,1.8636768,1.8749946,2.0975795,2.0787163,2.8709676,3.9008942,2.9615107,1.7655885,1.4109617,1.6976813,2.3390274,2.9615107,3.169005,3.3651814,4.025391,4.666737,3.8593953,4.9459114,6.4926877,6.8737226,5.836251,4.4705606,6.300284,6.356873,5.715527,5.292993,5.8437963,5.455216,4.9534564,3.8782585,2.463524,1.6335466,1.7165444,2.0787163,2.071171,1.448688,0.35085413,0.120724,0.02263575,0.0,0.011317875,0.060362,0.02263575,0.16976812,0.27540162,0.21881226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.34330887,0.8111144,0.6413463,1.3355093,1.3656902,1.2600567,1.3430545,1.7089992,2.1353056,3.1048703,3.2369123,2.4522061,1.9391292,2.1956677,2.5238862,2.848332,3.218049,3.8292143,1.6335466,1.1657411,2.1164427,3.9574835,5.934339,8.243186,10.740664,12.162943,12.08749,10.940613,11.027383,11.321648,10.925522,10.231359,10.940613,11.989402,10.944386,8.695901,6.5341864,6.119198,4.3121104,4.134797,4.172523,3.8707132,3.5538127,2.2371666,1.6033657,1.4449154,1.6033657,1.9693103,3.127506,3.1161883,2.867195,2.746471,2.5616124,2.233394,2.0787163,2.384299,2.8596497,2.6408374,3.3840446,3.5538127,3.904667,4.3800178,4.074435,4.085753,3.2369123,2.3956168,2.071171,2.425798,2.5616124,2.897376,3.3425457,3.5990841,3.1576872,3.500996,3.9876647,4.093298,3.6745367,2.9916916,2.9539654,2.9803739,2.8332415,2.5314314,2.3503454,2.142851,1.9881734,1.9089483,1.8636768,1.7542707,1.7542707,1.8749946,2.6295197,3.6368105,3.6028569,3.0030096,3.0558262,3.2067313,3.2105038,3.1124156,2.795515,2.8332415,2.9954643,3.1425967,3.2670932,3.2784111,3.4255435,3.2746384,3.0520537,3.663219,3.0897799,2.8709676,3.1237335,3.712263,4.274384,4.9685473,3.8141239,3.3953626,4.2027044,4.6554193,3.3236825,3.9876647,4.432834,4.274384,4.957229,5.070408,4.776143,5.5382137,6.6662283,5.3269467,7.7301087,8.707218,8.412953,9.473062,16.969267,12.804289,13.219278,9.967276,4.0178456,5.5683947,6.6322746,8.654402,9.06939,8.028146,8.409182,9.031664,8.726082,8.409182,8.201687,7.4471617,6.349328,4.3875628,4.847823,6.983129,6.043745,6.224831,6.300284,6.4926877,7.175533,8.835487,8.552541,8.216777,7.5905213,6.9454026,7.0812173,6.8850408,6.771862,6.730363,6.760544,6.881268,7.0284004,7.356619,7.7225633,8.001738,8.088508,8.367682,9.031664,9.81637,10.751981,12.193124,12.14408,11.69891,11.091517,10.751981,11.336739,11.32542,10.789707,10.20495,9.831461,9.718282,9.439108,8.537451,8.382772,9.118435,9.64283,10.133271,9.092027,7.8696957,7.454707,8.469543,7.748972,7.7602897,7.5905213,7.0510364,6.6850915,7.17176,7.484888,7.364164,7.062354,7.352846,7.865923,7.273621,7.001992,7.1604424,6.5002327,5.5495315,4.9723196,4.5988297,4.172523,3.3425457,3.2557755,3.6028569,4.1008434,4.4177437,4.134797,4.221567,4.3800178,4.4818783,4.6931453,5.462761,4.8138695,4.085753,3.6292653,3.5047686,3.4783602,3.380272,3.6330378,4.3083377,5.0779533,5.1873593,4.515832,4.349837,4.115934,3.7462165,3.663219,3.6858547,3.7198083,4.0480266,4.52715,4.5761943,3.7348988,3.361409,3.0897799,2.7615614,2.3956168,2.4069347,2.3201644,2.1315331,1.9655377,2.0749438,3.1124156,3.399135,3.1237335,2.7087448,2.806833,3.7952607,4.1989317,4.1800685,4.2328854,5.172269,5.5759397,6.5568223,6.8850408,6.677546,7.3868,8.360137,8.8618965,9.129752,9.58624,10.819888,11.649866,12.019584,12.2270775,11.947904,10.238904,9.87296,9.763554,10.1294985,10.56335,10.023865,9.608876,9.854096,10.246449,10.56335,10.895341,10.759526,11.514051,11.947904,11.59705,10.740664,11.438599,12.196897,12.630749,12.585477,12.14408,12.449662,12.068627,11.887542,12.057309,12.0082655,10.484125,10.880251,12.015811,13.147598,13.977575,13.819125,13.7700815,13.679539,13.449409,13.045737,13.679539,14.992412,16.056292,16.36942,15.8676605,15.63753,15.55076,15.875206,16.920223,19.059301,2.674791,2.4484336,2.2107582,2.052308,2.0485353,2.2786655,2.0372176,2.11267,2.335255,2.5201135,2.4559789,2.4333432,2.263575,2.173032,2.1768045,2.1164427,2.6936543,3.180323,3.9386206,4.9534564,5.8136153,6.432326,6.9491754,7.2396674,7.33021,7.3868,7.677292,7.91874,9.21275,11.993175,16.033657,19.519562,20.526854,21.507734,25.238861,34.83642,32.935017,20.285404,8.495952,2.7691069,1.8749946,1.7354075,1.8674494,1.9353566,1.7957695,1.5052774,1.4562333,1.2940104,1.0450171,0.7922512,0.66020936,0.6752999,0.7205714,0.8865669,1.1657411,1.4147344,1.8599042,2.2975287,3.1350515,4.2064767,4.7874613,4.2894745,3.5500402,2.9954643,2.7917426,2.867195,3.180323,3.5387223,3.7009451,3.9008942,4.847823,4.7006907,5.8400235,8.065872,9.676784,7.4999785,5.832478,6.5266414,7.394345,8.047009,9.910686,9.488152,8.130007,6.4738245,5.0025005,4.055572,3.6368105,3.7047176,3.9499383,4.266839,4.7648253,5.4174895,4.8629136,3.9989824,3.3840446,3.2218218,3.821669,4.61392,5.1269975,5.198677,4.961002,5.6363015,5.111907,4.8742313,5.564622,6.971811,7.9262853,7.5603404,6.6586833,6.126743,6.9869013,7.454707,7.752744,8.001738,8.314865,8.790216,7.33021,5.9607477,5.613666,6.673774,8.99771,13.977575,16.867407,15.256495,10.106862,5.775889,2.335255,1.3732355,1.237421,1.3091009,2.0108092,0.7696155,0.38858038,0.25276586,0.116951376,0.10186087,0.17731337,0.12826926,0.090543,0.241448,0.7997965,2.3993895,5.028909,7.699928,9.454198,9.359882,7.1340337,6.2097406,5.1081343,3.8480775,3.953711,4.4177437,7.032173,8.171506,7.635793,8.661947,10.891568,12.50248,13.95494,14.84528,13.905896,15.297995,15.158407,16.331694,18.99894,20.692848,21.560553,22.760246,22.89606,22.88097,25.948114,23.714722,24.703148,27.189308,29.237844,28.724768,26.793182,31.576872,36.477512,38.94481,40.480267,42.14022,42.102493,41.295155,41.095203,43.324825,44.71315,45.422405,45.565765,45.93171,47.97647,49.01017,50.266457,51.258656,52.122585,53.601456,55.423634,56.302654,55.544357,52.9752,48.953583,45.79212,44.301937,44.656563,46.16184,47.25213,48.025517,44.76597,41.630917,40.42745,40.597218,41.695053,44.18121,47.338898,50.628628,53.673138,53.688225,54.58988,55.08787,54.32957,51.88491,48.15756,47.81425,46.044888,42.042133,39.012714,36.76423,34.213936,31.27506,28.264507,25.865116,25.276588,24.69183,24.80501,25.88398,27.76652,34.587425,43.211647,51.69251,59.309437,66.545334,74.120766,75.62604,69.6087,59.709335,54.665337,56.55542,64.30062,66.26616,56.974182,37.111313,29.071848,24.050484,22.620659,22.19058,17.003222,18.191597,17.814335,16.693865,16.290195,18.69713,15.433809,13.555041,15.147089,19.293203,22.100037,18.723537,17.199398,20.628714,26.07261,24.571106,28.128693,30.128183,30.358313,28.966215,26.47251,20.04773,12.781653,8.152642,7.2962565,9.001483,8.394091,6.579458,5.1873593,6.6360474,14.102073,7.7414265,7.3453007,9.623966,10.880251,7.01331,4.9723196,3.663219,2.5087957,1.6109109,1.750498,3.4896781,5.1534057,6.6058664,7.6320205,7.9262853,10.378491,12.264804,13.275867,13.762536,14.754736,14.075664,12.728837,11.446144,9.929549,6.862405,4.9534564,4.255521,3.9499383,3.4859054,2.6182017,2.3390274,2.022127,2.0560806,2.4371157,2.7804246,2.9313297,3.7160356,4.587512,4.738417,3.1048703,2.173032,1.9240388,1.6448646,1.3128735,1.5920477,1.4600059,2.2371666,3.2105038,3.9574835,4.3611546,4.979865,6.089017,6.828451,6.6624556,5.409944,6.579458,6.1229706,5.8437963,5.934339,4.991183,4.1008434,3.5424948,2.9086938,2.093807,1.3015556,1.8372684,1.7844516,1.3091009,0.6526641,0.120724,0.7469798,0.5093044,0.14713238,0.011317875,0.049044125,0.011317875,0.049044125,0.06790725,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46026024,1.1355602,1.0789708,0.90543,1.0035182,1.1129243,1.1506506,1.1959221,2.003264,2.8407867,3.029418,2.3918443,1.2525115,2.1353056,2.886058,3.1199608,3.1652324,4.036709,2.0258996,1.267602,1.7618159,3.5123138,6.5341864,7.707473,9.314611,10.484125,10.827434,10.453944,10.751981,10.642575,10.284176,10.016319,10.355856,11.657412,11.649866,9.390063,6.126743,5.300538,5.1345425,4.247976,3.682082,3.6368105,3.4444065,2.4295704,1.7429527,1.6109109,2.0447628,2.8219235,3.6594462,3.874486,3.6556737,3.229367,2.867195,2.4710693,2.6483827,2.8709676,2.8709676,2.6521554,3.6292653,3.5575855,3.682082,4.0593443,3.5500402,3.5990841,3.1576872,2.474842,1.961765,2.1692593,2.7917426,3.0369632,3.1237335,3.1576872,3.1576872,3.4217708,3.7952607,3.832987,3.519859,3.2972744,3.0746894,2.987919,2.7728794,2.5012503,2.5804756,2.6068838,2.5427492,2.3314822,2.1315331,2.3163917,2.686109,2.655928,2.6898816,2.9124665,3.1010978,2.8558772,2.7087448,2.8030603,2.9615107,2.6974268,2.8407867,3.059599,3.350091,3.5538127,3.361409,2.6634734,2.795515,2.8558772,2.8558772,3.712263,3.1463692,2.897376,3.3161373,4.0216184,3.8707132,4.0178456,3.1840954,2.8294687,3.138824,2.9954643,2.9124665,3.7160356,4.0970707,4.0103,4.666737,5.05909,4.9044123,5.7192993,6.832224,5.3609,7.5037513,8.201687,7.7942433,8.141325,12.596795,9.510788,12.1101265,9.808825,3.4142256,5.13077,5.2062225,6.4549613,7.2962565,7.413208,7.7602897,8.7751255,10.555805,11.555551,10.884023,8.299775,9.556059,5.847569,4.112161,5.4288073,5.0062733,5.666483,6.1305156,6.5455046,7.1566696,8.296002,8.13378,7.5565677,6.719045,6.1418333,6.7152724,6.692637,6.5756855,6.515323,6.5341864,6.4926877,6.598321,7.073672,7.5565677,7.8244243,7.7829256,7.9262853,8.601585,9.2995205,10.035183,11.348056,11.653639,11.348056,10.884023,10.623712,10.850069,11.257513,11.370691,11.257513,11.050018,10.940613,10.299266,9.310839,8.8769865,9.137298,9.495697,9.944639,9.578695,8.858124,8.43559,9.125979,8.533678,8.20546,7.7716074,7.405663,7.8319697,7.752744,7.4584794,7.2283497,7.224577,7.488661,7.6886096,7.537705,7.462252,7.2924843,6.2436943,5.5080323,5.0439997,4.5196047,3.92353,3.561358,3.6896272,3.99521,4.3347464,4.4931965,4.172523,3.8556228,3.651901,3.85185,4.4101987,4.927048,4.2592936,3.7160356,3.6481283,3.893349,3.7613072,3.7990334,4.3309736,4.859141,5.040227,4.7120085,4.274384,4.1008434,4.08198,4.093298,3.9688015,3.9122121,4.191386,4.666737,5.0477724,4.870459,3.7273536,3.3123648,3.0143273,2.6144292,2.2975287,2.173032,2.052308,1.901403,1.8674494,2.2711203,3.2218218,3.3161373,3.0331905,2.8181508,3.1010978,3.6292653,3.904667,4.187614,4.6629643,5.4174895,6.25124,6.858632,7.575431,8.246958,8.2507305,8.29223,8.548768,8.89585,9.691874,11.793225,12.887287,13.298503,12.925014,11.883769,10.506761,10.061591,10.144588,10.419991,10.34831,9.193887,8.605357,8.914713,9.748463,10.850069,12.064855,12.2270775,12.245941,11.981857,11.5857315,11.510279,12.344029,13.377728,13.943622,13.792717,13.098554,12.728837,12.061082,11.834724,12.027128,11.849815,11.495189,11.857361,12.204442,12.385528,12.804289,12.804289,12.932558,12.992921,12.853333,12.46098,13.27964,14.618922,15.897841,16.712729,16.795727,16.505234,16.625957,16.931541,17.57666,19.108345,3.4179983,3.2218218,2.7389257,2.252257,1.9579924,1.9429018,1.9693103,2.1579416,2.372981,2.4823873,2.3578906,2.4672968,2.354118,2.2560298,2.2899833,2.425798,2.7502437,3.187868,3.7047176,4.349837,5.243949,5.9796104,6.3455553,6.620957,6.934085,7.2698483,8.09228,8.420499,8.793989,10.314357,14.641558,16.535416,17.99542,22.548979,31.595734,44.403797,36.613327,20.764528,8.401636,3.3576362,1.7316349,1.2147852,1.116697,1.0827434,1.0299267,1.1506506,1.3166461,1.3468271,1.237421,1.0336993,0.83752275,0.66020936,0.60362,0.69039035,0.88279426,1.0714256,1.3770081,1.6260014,2.3654358,3.361409,3.5990841,2.8596497,2.335255,1.9994912,1.9051756,2.2107582,2.071171,2.093807,2.2711203,2.6106565,3.1463692,2.9011486,4.146115,6.187105,7.5188417,5.8513412,4.4931965,5.492942,7.2887115,8.865668,9.756008,9.559832,8.68081,7.786698,7.201941,6.888813,7.1868505,6.8058157,6.3417826,6.089017,6.039973,5.9494295,5.20245,4.353609,3.772625,3.6556737,3.7650797,3.6669915,3.4330888,3.108643,2.7389257,3.8103511,4.164978,5.0854983,6.820906,8.601585,8.235641,6.9567204,6.0022464,6.4210076,9.039209,9.733373,9.235386,8.458225,7.9413757,7.8621507,7.454707,6.5832305,6.326692,7.2283497,9.307066,14.517061,17.682293,15.682802,10.103089,7.220804,3.8141239,2.082489,1.841041,2.1843498,1.5015048,0.5583485,0.2263575,0.211267,0.45648763,1.1431054,1.2940104,1.5203679,2.0183544,2.5917933,2.6483827,2.957738,4.123479,5.0515447,5.3986263,5.5985756,4.8930945,4.168751,3.4632697,3.0897799,3.663219,3.7198083,5.0515447,6.2021956,7.0246277,8.703445,10.929295,12.438345,13.358865,13.65313,13.094781,15.577168,16.788181,17.278622,17.48989,17.753973,20.270313,23.175236,23.839218,22.745155,23.4695,23.05074,25.593489,28.351276,29.811283,29.698105,30.637487,35.02505,38.016743,38.492092,39.024033,39.891735,40.246365,39.944553,40.001144,42.562756,45.69026,48.18774,49.2818,50.18723,54.13717,56.27625,57.872066,58.818996,59.47166,60.652493,58.792587,56.834595,54.231483,51.0738,48.082108,47.829338,47.546394,47.727478,48.485775,49.538338,52.201813,51.281292,48.40278,45.780804,46.188248,45.452587,46.20334,47.829338,50.062733,53.012928,53.378872,53.31851,53.08838,52.190495,49.361027,44.373615,44.12085,44.660336,44.030308,42.238308,39.442795,36.239838,32.72752,29.550972,27.894789,26.321604,25.92925,26.219744,26.819592,27.476028,32.003178,38.990078,46.788094,54.869057,63.813953,73.94722,79.43639,74.10944,60.686447,50.756897,46.33538,48.251873,52.31499,52.405533,40.487812,30.501673,23.601542,21.579414,22.024584,18.327412,20.960705,20.040184,17.248442,15.354584,18.184053,15.230087,12.593022,13.641812,17.587978,19.462973,16.55428,15.886524,20.640032,27.596752,27.144037,25.642532,24.02785,22.598024,21.783136,22.149082,18.131235,12.434572,8.326183,7.1378064,8.246958,7.5565677,5.5268955,4.293247,5.6778007,11.159425,5.983383,6.0550632,9.548513,12.789199,10.269085,7.073672,6.2135134,5.342037,3.9084394,3.1576872,4.2027044,5.5193505,6.9869013,8.175279,8.341274,10.178542,11.216014,11.981857,12.887287,14.222796,14.04171,13.645585,12.97783,11.619685,8.790216,6.485142,5.247721,4.6516466,4.2781568,3.712263,2.8785129,2.2786655,2.214531,2.776652,3.8556228,3.187868,3.8556228,4.274384,3.92353,3.3538637,2.5767028,1.9202662,1.388326,1.2902378,2.2296214,1.2336484,1.4109617,2.093807,2.957738,4.002755,4.8025517,5.3684454,5.847569,6.1795597,6.1305156,8.009283,7.152897,5.5985756,4.29702,3.108643,2.886058,2.4333432,1.7618159,1.1996948,1.3845534,1.9730829,1.4335974,0.6790725,0.5583485,1.8372684,0.935611,0.35839936,0.094315626,0.09808825,0.26408374,0.331991,0.14713238,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14713238,0.52439487,0.7507524,0.814887,1.0638802,1.3317367,1.3015556,1.4373702,1.961765,2.8709676,3.0860074,3.6028569,3.361409,2.2748928,1.237421,2.3578906,3.4142256,3.6443558,3.1954134,3.1199608,1.5769572,1.1732863,1.8938577,3.9574835,7.816879,8.827943,9.073163,9.1825695,9.559832,10.355856,11.25374,10.38981,9.34102,9.163706,10.382264,11.076427,10.801025,9.58624,7.7037,5.66271,5.9532022,4.98741,3.6481283,2.6672459,2.6031113,2.2258487,1.8787673,1.9391292,2.5578396,3.6783094,3.4217708,3.6896272,3.9688015,3.9914372,3.7047176,3.0558262,2.9728284,3.2784111,3.7575345,4.183841,4.5120597,4.1498876,3.832987,3.731126,3.4632697,3.591539,3.3161373,2.6634734,1.9844007,1.9579924,2.8445592,3.1652324,3.187868,3.1576872,3.3048196,3.2935016,3.4632697,3.4255435,3.2105038,3.2520027,3.0445085,2.5729303,2.3578906,2.5389767,2.8596497,2.7313805,2.5917933,2.4522061,2.3428001,2.3201644,2.5276587,2.5427492,2.6597006,2.8256962,2.637065,2.8521044,2.9351022,3.0445085,3.1614597,3.097325,3.4859054,3.2067313,3.218049,3.5274043,3.1765501,2.6408374,3.0935526,3.2972744,2.9841464,2.8445592,2.8898308,3.0143273,3.4444065,3.8405323,3.2821836,3.3048196,2.9426475,2.7540162,2.776652,2.5427492,3.4632697,3.9650288,3.9084394,3.7801702,4.7120085,5.0062733,4.6629643,5.2175403,6.330465,5.772116,6.9982195,7.7112455,6.9793563,6.066381,8.439363,6.356873,10.212496,8.963757,3.3727267,6.017337,4.7912335,9.001483,11.106608,9.446653,8.22055,8.892077,7.3151197,7.164215,8.571404,8.14887,9.480607,5.8702044,4.1762958,5.515578,5.2590394,5.9003854,6.3153744,6.5455046,6.7567716,7.2585306,6.7869525,6.119198,5.5193505,5.3986263,6.300284,6.4436436,6.156924,5.9984736,6.0550632,5.96452,6.1041074,6.511551,6.960493,7.3377557,7.624475,7.9828744,8.684583,9.295748,9.861642,10.899114,11.204697,10.93684,10.570895,10.480352,10.929295,11.676274,11.959221,11.978085,11.846043,11.574413,11.457462,10.895341,10.223814,9.654147,9.276885,9.363655,9.442881,9.529651,9.612649,9.65792,8.695901,8.145098,7.9451485,7.9225125,7.805561,7.383027,7.496206,7.77538,7.956466,7.888559,7.3868,7.326438,7.092535,6.4738245,5.6476197,5.251494,4.8968673,4.436607,3.9612563,3.7914882,4.0103,4.247976,4.504514,4.5950575,4.134797,3.7575345,3.7386713,4.104616,4.534695,4.3800178,3.9574835,3.5764484,3.5651307,3.821669,3.7914882,3.742444,4.2819295,5.036454,5.481624,4.930821,4.7572803,5.0175915,4.9459114,4.402653,3.8405323,3.9801195,4.2592936,4.5761943,4.738417,4.4403796,3.591539,3.2255943,2.867195,2.4031622,2.052308,1.7429527,1.7957695,1.8938577,2.0636258,2.6936543,3.8292143,3.731126,3.3764994,3.3048196,3.6028569,3.783943,4.142342,4.7535076,5.523123,6.2097406,7.039718,7.8131065,8.533678,8.99771,8.790216,8.98262,8.677037,8.66572,9.7296,12.679792,15.339493,14.7736,13.12119,11.634775,10.657665,10.582213,10.914205,10.9594755,10.3634,9.125979,8.269594,8.503497,9.020347,9.718282,11.189606,11.846043,12.095036,12.0082655,11.8045435,11.857361,12.566614,13.558814,14.015302,13.671993,12.815607,12.057309,11.808316,11.68382,11.581959,11.68382,11.642321,11.962994,12.272349,12.521342,12.97783,13.124963,12.985375,12.849561,12.7477,12.449662,13.12119,14.200161,15.101818,15.607349,15.882751,16.712729,17.769064,18.346275,18.459454,18.836716,4.4931965,4.146115,3.4745877,2.7691069,2.2748928,2.1881225,2.3201644,2.4484336,2.655928,2.7841973,2.4371157,2.5087957,2.505023,2.5427492,2.6634734,2.8219235,2.8634224,3.240685,3.5689032,3.8971217,4.7120085,5.5457587,5.6476197,5.836251,6.439871,7.273621,8.390318,8.793989,8.786444,9.789962,14.362384,15.78089,18.429274,25.601034,35.855026,43.007923,30.286634,16.535416,7.5188417,4.0593443,2.052308,0.97333723,0.5583485,0.422534,0.422534,0.6375736,0.7922512,0.8978847,0.9318384,0.88279426,0.73188925,0.56589377,0.66020936,0.80356914,0.91297525,1.0148361,1.3392819,1.7995421,2.3654358,2.806833,2.6898816,2.4371157,2.3654358,2.282438,2.1541688,2.1202152,2.003264,1.8372684,1.8372684,1.9127209,1.6675003,1.4147344,2.0749438,3.1237335,3.8254418,3.2633207,3.6028569,5.3571277,7.884786,10.253995,11.249968,12.287439,12.438345,12.555296,12.789199,12.58925,12.049765,10.269085,8.103599,6.217286,5.070408,4.557331,4.0178456,3.5160866,3.1727777,3.150142,3.1010978,2.6785638,2.1692593,1.7467253,1.4713237,2.3503454,3.4632697,5.4778514,7.8432875,8.793989,7.6508837,6.8850408,6.907676,8.14887,11.053791,11.00852,9.367428,7.5490227,6.2097406,5.2326307,6.960493,7.9036493,8.492179,9.099571,10.0465,14.132254,16.569368,15.116908,10.887795,8.367682,5.3344917,3.500996,2.7125173,2.4295704,1.7278622,0.72811663,0.35462674,0.4376245,0.90920264,1.8259505,2.5012503,3.048281,3.9273026,4.9685473,5.3646727,5.036454,4.255521,3.3236825,2.5540671,2.2748928,2.323937,2.3465726,2.4823873,2.8256962,3.410453,3.6858547,4.6026025,6.617184,9.235386,11.004747,12.257258,13.106099,14.286931,15.324403,14.558559,16.520325,17.297485,17.452164,17.30503,16.939087,20.836208,22.764019,22.888515,21.949133,21.277605,23.616632,26.763002,29.056757,30.184772,31.180746,35.504173,37.631935,38.51473,38.548683,37.55648,38.069557,37.990334,37.386715,37.43953,40.438766,45.21114,49.444023,52.262173,54.782288,60.120552,63.142426,64.681656,63.82904,61.637146,61.116524,55.89521,51.526512,48.229237,46.11657,45.192276,46.65605,47.195538,47.6143,48.742313,51.413334,55.55945,57.249584,56.20834,53.718407,52.620575,50.711624,50.53054,50.945526,51.662327,53.250603,54.620064,54.518204,54.216393,53.514687,50.722942,45.57331,43.92467,44.39248,45.290363,44.6377,41.513966,37.786613,33.851765,30.475266,28.754948,26.87618,26.581915,26.740366,26.879953,27.211945,30.105547,35.82862,43.253147,51.75287,61.22593,71.061165,81.87728,81.009575,66.92259,49.19503,39.386204,34.96846,36.541645,41.053707,41.80446,30.92798,22.518799,19.651604,20.7268,19.481836,22.167944,21.68505,19.346022,16.77309,15.8676605,13.166461,11.857361,13.264549,16.116653,16.550507,14.939595,14.139798,18.293459,25.28036,26.713957,20.247679,17.078674,16.086473,16.25624,16.663685,14.5132885,10.789707,7.9262853,6.85486,7.01331,6.541732,4.7308717,3.6745367,4.5007415,7.3717093,5.4891696,5.583485,8.424272,12.181807,12.442118,8.963757,9.224068,9.258021,7.6810646,5.6853456,6.5530496,7.677292,8.903395,9.835234,9.81637,11.317875,12.034674,12.396846,12.872196,13.93985,13.426772,13.573905,13.860624,13.434318,11.136789,8.511042,6.673774,5.3948536,4.568649,4.217795,3.3915899,2.7728794,2.757789,3.2670932,3.7763977,3.0030096,3.3312278,3.7009451,3.8593953,4.3724723,2.8030603,1.9391292,1.6260014,1.8033148,2.516341,1.6146835,1.2487389,1.5052774,2.282438,3.2859564,4.5422406,4.979865,5.142088,5.4740787,6.368191,7.8432875,6.3417826,3.99521,2.323937,2.2598023,2.5578396,1.9089483,1.0374719,0.6149379,1.2751472,1.4335974,0.8262049,0.24522063,0.3772625,1.8146327,0.573439,0.1358145,0.13958712,0.2678564,0.24899325,0.32821837,0.13958712,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14713238,0.52439487,0.5583485,0.42630664,1.0751982,1.5958204,1.6184561,2.0145817,2.8634224,3.440634,3.4444065,3.640583,3.3463185,2.6031113,2.1541688,2.9464202,4.0216184,4.395108,3.6594462,2.0145817,2.425798,2.535204,2.625747,3.8971217,8.477088,9.695646,9.310839,8.560086,8.397863,9.495697,10.510533,9.891823,8.926031,8.820397,10.687846,10.933067,9.97482,9.378746,8.956212,6.7756343,6.3945994,5.2288585,3.482133,1.9089483,1.81086,1.7165444,1.7240896,2.142851,2.9916916,3.9876647,3.0445085,3.380272,4.0103,4.323428,4.1083884,3.8405323,3.4745877,3.8895764,4.8138695,4.8440504,4.9647746,4.7950063,4.3196554,3.7650797,3.5839937,3.6783094,3.259548,2.6144292,2.0598533,1.9353566,2.7125173,3.1576872,3.289729,3.2520027,3.3048196,2.886058,2.8709676,2.916239,2.927557,3.0445085,2.637065,1.9240388,1.7618159,2.3013012,3.006782,2.8143783,2.6182017,2.5087957,2.474842,2.3993895,2.293756,2.3880715,2.6597006,2.8558772,2.4710693,2.6219745,2.8785129,3.029418,3.006782,2.8822856,3.4972234,3.0860074,2.9313297,3.2369123,3.138824,2.7087448,3.3161373,3.62172,3.1954134,2.5201135,3.029418,3.180323,3.3689542,3.4330888,2.6295197,3.0105548,3.0520537,2.9237845,2.704972,2.3956168,3.7763977,4.115934,3.7688525,3.4594972,4.2781568,4.7120085,4.4215164,4.878004,5.994701,6.145606,6.198423,6.7341356,6.145606,4.9044123,5.5457587,5.2779026,7.914967,7.0284004,3.572676,5.907931,5.3646727,10.4049,11.925267,8.654402,7.1340337,7.5565677,4.1762958,2.6974268,4.244203,5.3269467,7.356619,6.6020937,5.6023483,5.4174895,5.6287565,5.9682927,6.2021956,6.300284,6.2889657,6.2361493,5.7607985,5.240176,4.930821,5.0854983,5.9418845,6.156924,5.7607985,5.455216,5.4288073,5.372218,5.7419353,6.092789,6.515323,7.032173,7.586749,8.065872,8.616675,9.114662,9.616421,10.33322,10.676529,10.54826,10.453944,10.676529,11.276376,12.1101265,12.272349,12.204442,12.113899,11.959221,12.31762,12.223305,11.476325,10.336992,9.559832,9.567377,9.80128,10.050273,10.084227,9.665465,8.575176,7.997965,7.7301087,7.537705,7.141579,6.8397694,7.2924843,7.809334,7.99042,7.7225633,6.9793563,6.94163,6.5040054,5.6023483,5.2288585,5.0062733,4.6856003,4.3385186,4.063117,3.9914372,3.8895764,3.8141239,3.953711,4.2102494,4.2064767,4.0103,4.2781568,4.6629643,4.7648253,4.1612053,3.8593953,3.6254926,3.6669915,3.8820312,3.8556228,3.7235808,4.3724723,5.3910813,6.224831,6.187105,5.726845,5.7306175,5.342037,4.5988297,4.4403796,4.6026025,4.5422406,4.478106,4.3385186,3.7688525,3.3312278,2.8407867,2.3993895,2.0787163,1.9127209,1.659955,1.8561316,2.252257,2.7351532,3.361409,4.315883,4.247976,3.8782585,3.6858547,3.9084394,3.9273026,4.3800178,5.1156793,5.983383,6.8133607,7.865923,8.907167,9.49947,9.484379,9.016574,9.22784,8.688355,8.288457,9.024119,12.004493,14.947141,14.385019,12.808062,11.570641,10.917976,11.276376,11.438599,11.046246,10.242677,9.631512,9.0543,9.144843,9.374973,9.752235,10.819888,11.631002,12.219532,12.362892,12.091263,11.717773,12.408164,13.45318,13.924759,13.521088,12.570387,11.514051,11.012292,10.751981,10.770844,11.431054,11.306557,11.729091,12.47607,13.249459,13.694629,13.7700815,13.283413,12.73261,12.400619,12.340257,12.823153,13.513543,14.154889,14.667966,15.131999,16.867407,18.478317,19.18757,19.01403,18.780127,4.7346444,4.402653,3.8820312,3.2821836,2.8219235,2.8521044,2.8143783,2.6936543,2.8332415,3.0218725,2.4710693,2.3805263,2.5201135,2.7502437,2.927557,2.8936033,2.7879698,3.097325,3.3538637,3.572676,4.244203,5.1835866,5.168496,5.3269467,6.058836,7.0359454,8.065872,8.699674,9.012801,10.167224,14.407655,16.31283,20.598532,28.339958,35.236317,31.60328,16.65614,8.409182,4.719554,3.3425457,1.931584,0.9242931,0.58098423,0.47535074,0.3961256,0.35839936,0.33953625,0.35462674,0.422534,0.5093044,0.513077,0.49044126,0.88279426,1.237421,1.3996439,1.5165952,1.8863125,2.5125682,2.7313805,2.5087957,2.41448,2.9351022,3.3312278,3.4934506,3.308592,2.6823363,2.9539654,2.7615614,2.3616633,1.8938577,1.3958713,1.0223814,1.1317875,1.5543215,2.0749438,2.41448,5.243949,8.526133,12.053536,15.373446,17.780382,20.002459,21.051247,21.590733,21.277605,18.75372,15.30554,11.472552,7.598067,4.3121104,2.5314314,2.3126192,2.4031622,2.4710693,2.4031622,2.3163917,2.2711203,2.2183034,2.071171,1.8485862,1.6524098,1.9429018,3.289729,5.621211,7.696155,7.1340337,6.405917,7.284939,8.922258,10.695392,12.2119875,11.208468,8.382772,5.6589375,3.8443048,2.6446102,6.379509,9.076936,10.574668,11.1631975,11.59705,14.815099,16.573141,16.207197,13.58145,9.092027,6.2323766,4.9987283,3.4783602,1.9353566,2.795515,1.2525115,0.6828451,0.76584285,1.1996948,1.6976813,2.8898308,3.4934506,4.2592936,5.4250345,6.6850915,7.2358947,5.50426,3.5349495,2.2258487,1.3355093,1.0827434,1.50905,2.0862615,2.625747,3.2859564,3.9461658,5.089271,8.14887,12.038446,13.13628,14.245432,15.030138,16.856089,18.76881,17.497435,17.523844,16.935314,17.689838,19.31584,18.919714,22.416937,21.78691,21.14179,21.594505,21.262514,24.084438,27.072357,29.317068,30.803484,32.387985,38.34496,38.974987,39.246616,39.76724,36.80573,37.737568,36.851,35.647533,35.504173,37.669662,43.51723,48.930946,53.412827,57.600437,63.300877,66.87733,68.22415,64.836334,58.268192,54.118305,48.372597,44.260437,42.766476,43.57759,45.064007,46.50515,47.229492,48.368824,50.771988,54.967148,58.615276,61.882366,63.39519,62.56144,59.554657,56.593147,56.18193,56.212112,55.842396,55.502857,57.07227,58.015427,58.385143,57.668346,54.804924,50.277775,47.131405,45.739307,45.622353,45.42995,42.660843,39.00517,35.100502,31.44483,28.407866,26.936543,26.66114,26.502691,26.40083,27.336441,29.309525,34.11585,41.551693,50.598446,59.422615,65.87758,80.164505,87.18536,78.44797,52.050907,36.179474,26.895044,24.435291,28.788902,39.699333,29.815056,21.179516,17.040947,17.369165,18.87067,20.477808,20.813572,20.504217,18.734856,13.253232,10.70671,11.087745,13.068373,14.694374,13.396591,13.664448,12.268577,14.434063,19.87419,22.801746,14.320885,12.00072,13.249459,14.743419,12.438345,10.770844,8.303548,6.760544,6.300284,5.50426,5.6815734,4.7836885,3.8971217,3.7688525,4.817642,7.001992,6.5341864,7.515069,10.650121,13.268322,10.876478,12.042219,12.864652,11.61214,8.741172,9.439108,10.797253,11.978085,12.396846,11.736636,12.936331,13.913441,14.034165,13.611631,13.894578,13.026875,13.196642,14.286931,15.124454,13.490907,10.868933,8.548768,6.33801,4.568649,4.1008434,3.742444,3.3538637,3.4783602,3.7763977,3.0181,2.8143783,2.9992368,3.6934,4.6554193,5.2892203,3.240685,2.5917933,2.6710186,2.8106055,2.3163917,2.022127,1.5316857,1.5279131,2.0749438,2.6144292,4.315883,5.032682,4.957229,4.7950063,5.772116,5.59103,3.6443558,1.7769064,1.2449663,2.7238352,2.837014,1.7693611,0.8601585,0.65643674,0.9280658,0.46026024,0.15845025,0.02263575,0.0,0.0,0.0452715,0.090543,0.24522063,0.35085413,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026408374,0.150905,0.49421388,1.2034674,1.5731846,1.780679,2.3616633,3.0030096,2.5616124,2.8445592,2.8898308,2.8785129,2.9313297,3.0897799,3.289729,4.217795,4.8968673,4.395108,1.8033148,4.2630663,4.749735,3.8405323,3.572676,7.4207535,8.60913,8.986393,8.563859,7.9262853,8.216777,8.5563135,8.9788475,8.98262,9.046755,10.623712,10.484125,9.424017,8.944894,8.922258,7.6131573,6.1305156,4.640329,3.029418,1.690136,1.50905,1.2147852,1.3317367,2.0447628,3.0897799,3.7462165,2.8785129,3.1840954,3.7273536,3.9688015,3.7952607,4.2517486,3.9310753,4.4516973,5.462761,4.644101,4.9685473,5.2364035,4.930821,4.2064767,3.8820312,3.8103511,3.0633714,2.4107075,2.1503963,2.1013522,2.5502944,3.097325,3.4217708,3.4142256,3.1954134,2.3692086,2.2371666,2.463524,2.7238352,2.686109,1.8863125,1.2449663,1.1732863,1.7731338,2.8445592,2.867195,2.7238352,2.5993385,2.5917933,2.7502437,2.4107075,2.4672968,2.625747,2.6785638,2.5314314,2.1843498,2.4333432,2.5993385,2.4295704,2.082489,2.7653341,2.806833,2.7351532,2.8294687,3.1350515,2.837014,3.2029586,3.4934506,3.3878171,2.987919,3.4179983,3.289729,3.1576872,3.0030096,2.2296214,3.1576872,3.2821836,3.0860074,2.8256962,2.546522,3.5575855,3.7650797,3.3463185,2.8445592,3.169005,4.032936,4.3083377,4.9760923,5.956975,6.1078796,5.3382645,5.485397,5.3986263,4.772371,4.164978,5.5985756,5.455216,4.4818783,3.7613072,4.7044635,6.488915,8.858124,8.356364,5.485397,4.7006907,4.8138695,2.9464202,1.4071891,1.1393328,1.7240896,4.5497856,7.303802,7.0963078,4.9232755,5.692891,5.670255,5.7004366,5.772116,5.764571,5.4401255,5.3873086,5.20245,5.0854983,5.1873593,5.621211,5.783434,5.4363527,5.062863,4.90064,4.927048,5.511805,5.8966126,6.3531003,6.9491754,7.537705,7.9489207,8.311093,8.729855,9.205205,9.623966,10.099318,10.265312,10.616167,11.231105,11.7555,12.283667,12.181807,11.974312,11.981857,12.306303,12.604341,12.555296,11.766817,10.552032,9.940866,10.3634,10.687846,10.510533,9.88805,9.325929,8.526133,7.9225125,7.1868505,6.511551,6.590776,6.590776,6.930312,7.194396,7.213259,7.0472636,6.6058664,6.5568223,6.017337,5.142088,5.119452,4.8025517,4.4516973,4.1612053,3.99521,3.9763467,3.4330888,3.0030096,3.0030096,3.4896781,4.22534,4.3422914,4.8327327,5.0741806,4.8440504,4.2781568,3.8556228,3.7499893,3.92353,4.1574326,4.032936,4.0291634,4.8100967,5.80607,6.7379084,7.5829763,6.651138,5.798525,4.9723196,4.515832,5.1873593,5.2137675,4.7950063,4.395108,4.025391,3.2369123,2.938875,2.2862108,1.8259505,1.7580433,1.9240388,1.9051756,2.1541688,2.848332,3.7047176,4.0103,4.266839,4.45547,4.187614,3.6858547,3.772625,3.8858037,4.496969,5.304311,6.1795597,7.183078,8.601585,9.714509,10.212496,10.008774,9.26934,9.0957985,8.744945,8.228095,8.265821,10.27663,11.6008215,11.989402,11.925267,11.740409,11.593277,12.102581,11.774363,10.914205,10.103089,10.193633,10.235131,10.359629,10.729345,11.223559,11.457462,11.887542,12.494934,12.608112,12.045992,11.140562,11.944131,13.20796,13.875714,13.562587,12.559069,11.306557,10.054046,9.544742,10.008774,11.144334,10.925522,11.480098,12.6345215,13.849306,14.211478,14.283158,13.634267,12.736382,12.106354,12.310076,12.702429,13.057055,13.728582,14.664193,15.388537,17.237123,18.761265,19.470518,19.43279,19.24416,2.3805263,3.440634,3.7613072,3.7084904,3.5085413,3.2670932,3.0822346,2.9539654,2.7351532,2.4220252,2.1654868,2.252257,2.4107075,2.4899325,2.4672968,2.4408884,2.4522061,2.6672459,2.8822856,3.108643,3.5839937,4.2706113,4.485651,4.8629136,5.5080323,5.9984736,7.4018903,8.703445,9.484379,10.804798,15.211224,17.557796,23.835445,30.8563,33.399048,24.231571,10.182315,4.085753,2.022127,1.3807807,0.87147635,0.8224323,1.1204696,1.1883769,0.90920264,0.6413463,0.72811663,0.7469798,0.6790725,0.6111652,0.73188925,0.67152727,1.0412445,1.5882751,2.2258487,3.006782,3.1048703,3.0369632,2.674791,2.3163917,2.6710186,3.3161373,4.1197066,4.7044635,4.7950063,4.195159,3.500996,3.0256453,2.3088465,1.6524098,2.0900342,1.4071891,1.50905,2.2371666,3.62172,5.904158,10.785934,15.826162,21.934042,28.256962,32.15031,35.236317,36.65105,35.938026,31.705141,21.620914,13.272095,7.4207535,3.8443048,2.2296214,2.1654868,2.4371157,2.6483827,2.7087448,2.5729303,2.2447119,2.2183034,3.0558262,3.640583,3.4481792,2.5314314,2.655928,3.7575345,4.9534564,5.5004873,4.7912335,5.692891,7.7678347,10.438853,12.479843,12.053536,11.823407,8.816625,5.3684454,3.1237335,3.0369632,6.809588,8.5563135,10.008774,11.891314,13.917213,16.52787,16.641048,15.811071,13.777626,8.469543,5.8437963,5.0854983,3.640583,1.7316349,2.3805263,1.0638802,0.87147635,0.9922004,1.0751982,1.2223305,1.5128226,1.5430037,1.7995421,2.3880715,3.0218725,6.1342883,6.089017,4.3913355,2.3578906,1.1129243,0.9318384,1.1431054,1.50905,2.1164427,3.3727267,3.983892,4.557331,7.0472636,10.95193,13.321139,17.399347,19.266796,18.51227,17.142809,19.606333,16.62973,17.550251,20.168453,22.669704,23.620405,20.594759,20.734346,22.53389,24.620152,25.74062,23.692085,26.638506,30.211182,32.387985,33.523544,37.62439,38.31101,37.488575,36.685005,37.062267,37.61307,37.541393,37.190536,36.451103,34.730785,42.81175,49.70056,54.620064,57.9777,61.36929,64.851425,66.51515,63.214104,55.140686,45.852486,41.740322,41.215927,43.026787,46.139202,49.72697,53.122334,54.721924,56.47997,58.58132,59.449024,59.71688,63.647957,67.29231,68.62405,67.54885,62.606712,61.4787,61.456062,60.94676,59.494297,59.581066,61.92764,63.274467,61.874825,57.479713,53.831585,49.183712,45.795895,44.24912,43.441776,42.42694,39.446568,36.27379,33.206646,29.068075,26.834682,26.597006,26.502691,26.581915,28.717222,30.8148,34.481792,41.344196,50.289093,57.479713,61.64092,72.242,86.894875,92.55381,65.50409,38.2846,24.67674,20.647577,23.477045,31.754185,25.054003,19.65915,15.588487,13.607859,15.245177,14.890551,14.64533,15.294222,15.852571,13.59654,11.106608,9.2844305,10.325675,12.577931,10.529396,12.642066,11.317875,11.747954,14.784918,16.969267,11.034928,9.359882,11.812089,14.807553,11.291467,8.473316,6.3644185,5.6891184,5.7079816,4.255521,4.8063245,5.511805,5.1269975,4.014073,4.134797,11.23865,10.050273,9.14107,11.242422,13.245687,13.29473,14.075664,14.324657,13.513543,11.84227,11.193378,12.551523,13.758763,13.800262,12.785426,13.226823,14.260523,14.766054,14.320885,13.200415,13.649357,13.792717,14.252977,14.969776,15.150862,13.5663595,10.77839,7.537705,4.991183,4.7006907,4.0782075,3.7009451,3.5990841,3.7009451,3.8593953,3.3350005,3.7273536,4.142342,4.1272516,3.6783094,4.825187,4.561104,4.478106,4.659192,3.7084904,2.1956677,1.448688,1.4977322,2.003264,2.2748928,4.2404304,5.0854983,4.587512,3.561358,3.8895764,3.048281,2.0787163,1.4260522,1.5656394,3.006782,2.444661,1.3694628,0.91674787,1.1091517,0.8526133,0.23013012,0.030181,0.0,0.0,0.0,0.21881226,0.15467763,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12826926,0.76207024,1.4939595,1.1280149,2.0070364,2.071171,1.6939086,1.5958204,2.8521044,2.7540162,2.969056,2.625747,1.8938577,1.9542197,2.0749438,3.0935526,4.255521,4.745962,3.7084904,4.3422914,4.9421387,5.191132,4.8553686,3.7688525,4.0517993,6.6850915,8.801534,9.205205,8.360137,7.4811153,7.986647,8.567632,8.816625,9.231613,7.5603404,8.058327,8.537451,7.9941926,6.5756855,4.8666863,3.682082,2.595566,1.7429527,1.8146327,1.267602,1.1280149,1.5731846,2.4861598,3.4632697,2.987919,2.7389257,2.8332415,3.1124156,3.1727777,3.2972744,3.4745877,4.1762958,5.2665844,6.013564,5.534441,5.5004873,5.2665844,4.772371,4.515832,4.247976,3.31991,2.5578396,2.2862108,2.335255,2.6634734,3.2859564,3.8292143,3.953711,3.3425457,2.2899833,2.1390784,2.3767538,2.5012503,2.0145817,1.086516,0.7432071,0.7997965,1.2336484,2.1956677,2.5993385,2.625747,2.6521554,2.8332415,3.127506,2.7011995,2.5012503,2.3088465,2.1654868,2.4107075,1.9353566,2.2447119,2.3503454,2.093807,2.1654868,2.3126192,2.7691069,2.795515,2.425798,2.4861598,3.500996,3.2331395,3.187868,3.572676,3.2821836,3.048281,3.1840954,3.0860074,2.7200627,2.6106565,3.572676,3.218049,2.9954643,3.3764994,3.8895764,3.4142256,2.7540162,2.0787163,1.6448646,1.8146327,2.9011486,4.1989317,5.2175403,5.643847,5.3269467,4.8968673,4.919503,4.749735,4.2404304,3.7386713,4.06689,2.916239,2.6898816,3.7763977,4.5309224,7.3151197,6.6360474,6.205968,6.3342376,3.9688015,2.5767028,2.1013522,2.3126192,2.7615614,2.7615614,2.5314314,4.3686996,5.5193505,5.4363527,5.753253,5.5570765,5.3156285,5.0854983,4.889322,4.7308717,5.05909,5.243949,5.3156285,5.304311,5.2175403,5.194905,5.040227,4.889322,4.8440504,4.991183,5.221313,5.66271,6.1720147,6.6850915,7.232122,7.635793,8.258276,8.763808,9.050528,9.246704,9.661693,10.148361,10.914205,11.815862,12.3893,12.098808,11.732863,11.559323,11.819634,12.709973,12.393073,11.472552,10.329447,9.378746,9.046755,10.182315,11.053791,10.933067,10.008774,9.397609,8.922258,7.835742,6.820906,6.4436436,7.141579,6.7869525,6.900131,6.862405,6.643593,6.790725,6.5341864,6.2323766,5.6891184,5.1081343,5.0968165,4.485651,4.1498876,3.821669,3.4896781,3.4029078,3.1840954,2.9615107,2.9766011,3.259548,3.663219,4.112161,4.8666863,5.0138187,4.561104,4.425289,3.7763977,3.7537618,3.9914372,4.214022,4.22534,4.7044635,5.0968165,5.523123,6.1078796,6.971811,6.7039547,5.704209,4.617693,3.893349,3.783943,3.9688015,3.904667,3.682082,3.3953626,3.127506,2.4182527,2.052308,1.8259505,1.7316349,1.9391292,1.8900851,2.233394,3.2972744,4.447925,4.1197066,3.4481792,3.9122121,3.893349,3.2105038,3.1124156,3.6254926,4.8063245,6.1305156,7.24344,7.964011,9.088254,9.880505,10.4049,10.585986,10.208723,9.9257765,9.748463,9.563604,9.5183325,9.993684,9.152389,9.325929,10.382264,11.872451,13.045737,13.106099,12.664702,11.706455,10.570895,9.948412,9.910686,10.661438,11.604594,12.106354,11.521597,11.216014,11.52537,11.548005,11.019837,10.299266,10.997202,12.377983,13.196642,12.947649,11.887542,10.751981,9.982366,9.737145,10.084227,10.985884,11.012292,11.317875,12.117672,13.185325,13.8719425,14.762281,14.324657,13.5663595,13.151371,13.396591,13.739901,14.045483,14.652876,15.546988,16.32792,17.769064,19.108345,20.14959,20.647577,20.29295,2.806833,2.9803739,3.2784111,3.4557245,3.3538637,2.886058,2.5880208,2.5993385,2.5201135,2.2598023,2.033445,1.8938577,1.931584,2.052308,2.1881225,2.282438,2.2447119,2.2786655,2.444661,2.7841973,3.3161373,3.874486,4.4177437,4.991183,5.492942,5.6778007,7.484888,8.771353,9.491924,10.597303,14.030393,15.856343,20.043957,24.544699,25.736847,18.433046,7.5263867,3.531177,2.173032,1.2789198,0.73566186,0.87147635,0.7696155,0.6752999,0.6790725,0.70170826,0.845068,0.9922004,0.95824677,0.76207024,0.6111652,0.5998474,0.76584285,1.1393328,1.6637276,2.1994405,2.161714,2.11267,2.252257,2.625747,3.0860074,3.7613072,4.0895257,4.304565,4.5535583,4.8930945,4.878004,4.5950575,4.9723196,6.1003346,7.254758,7.115171,7.1378064,7.405663,9.348565,15.731846,22.4773,29.06053,34.97978,39.07685,39.533337,37.10754,33.57259,28.8304,22.341486,13.140053,6.5568223,3.4972234,2.2409391,1.8334957,2.093807,2.4408884,2.7917426,3.0331905,3.0407357,2.6710186,2.704972,3.0558262,3.5877664,4.063117,4.1310244,4.2819295,4.9685473,5.451443,5.6061206,5.915476,7.413208,9.14107,11.310329,13.102326,12.664702,12.970284,11.54046,8.27714,5.1345425,6.1116524,10.03141,10.914205,10.70671,11.027383,13.170234,15.871433,12.996693,10.974566,10.816116,8.103599,5.9192486,4.4215164,3.361409,2.5238862,1.7467253,0.66020936,0.59230214,0.62248313,0.55080324,0.8903395,0.9507015,1.7165444,2.3880715,2.6144292,2.5087957,4.7308717,5.1835866,4.2517486,2.5502944,0.8941121,1.0902886,1.6109109,2.3805263,3.1954134,3.6896272,4.8855495,5.723072,7.375482,9.876732,12.136535,15.343266,17.172989,18.025602,18.949896,21.65864,19.655376,19.263023,19.923233,21.156881,22.560297,18.055782,18.150099,20.19109,22.39053,23.824127,25.650078,26.302742,25.966978,26.04243,29.128437,32.342712,33.91967,35.209908,36.91136,39.065533,38.197826,39.1108,39.310753,37.42821,33.229282,38.439278,44.99987,49.78733,52.548893,55.902756,57.91734,59.320755,57.177906,51.349197,44.460384,41.068794,40.548172,42.276035,46.195793,52.839386,57.69853,60.784534,63.866768,66.288795,64.97592,61.79937,62.180405,63.417828,64.51943,66.20957,65.45504,65.05138,65.26264,65.39845,63.84036,59.75461,59.93192,60.671356,59.554657,55.453815,49.900513,45.463905,42.921154,41.95159,41.14802,40.08414,38.635452,36.685005,33.968716,30.105547,28.25319,27.792929,27.24967,27.260988,30.607307,33.410366,35.538128,40.740578,48.904537,56.06498,59.796104,65.98321,80.07397,92.94616,80.873764,48.165104,28.68704,20.043957,20.160908,27.287397,19.255478,15.671484,13.70972,12.996693,15.596032,15.271586,13.981348,13.924759,15.026365,14.924504,11.615912,8.959985,9.0807085,10.736891,9.318384,13.422999,14.9358225,15.135772,14.864142,14.539697,9.808825,8.088508,9.65792,12.336484,11.487643,7.7112455,4.919503,4.5196047,5.4363527,4.112161,4.1612053,4.447925,4.285702,3.8367596,4.134797,7.032173,8.507269,9.201432,10.016319,12.132762,13.472044,13.792717,13.109872,12.257258,12.879742,11.627231,11.732863,12.189351,12.393073,12.140307,13.721037,14.901869,14.988639,14.11339,13.234368,13.792717,14.622695,15.543215,16.365646,16.859861,16.32792,12.898605,9.963503,8.224322,5.6778007,4.8968673,4.2328854,4.1310244,4.398881,4.214022,4.0216184,4.3347464,4.376245,4.115934,4.2517486,3.5349495,3.1425967,2.8181508,2.3956168,1.8146327,1.4637785,0.9808825,0.87902164,1.2336484,1.6863633,8.809079,9.122208,6.511551,4.0970707,4.221567,3.3576362,2.6974268,2.3126192,2.2220762,2.384299,1.539231,0.724344,0.42630664,0.51684964,0.23013012,0.06790725,0.011317875,0.0,0.0,0.0,0.16976812,0.10940613,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19240387,0.7394345,1.2864652,0.9695646,1.448688,1.5882751,1.9994912,2.5201135,2.1956677,1.961765,1.9051756,1.4939595,0.87147635,0.8563859,0.6073926,1.5316857,3.3689542,5.1081343,4.991183,4.8440504,4.425289,3.8782585,3.3010468,2.7426984,4.3121104,6.187105,8.039464,9.220296,8.741172,6.79827,6.096562,6.0701537,6.379509,6.911449,5.2967653,5.458988,5.5797124,5.0439997,4.429062,4.6931453,4.014073,2.969056,2.0070364,1.4373702,1.3845534,1.3807807,1.9806281,3.0520537,3.7575345,3.3764994,3.059599,2.8181508,2.8822856,3.6745367,3.591539,3.1954134,3.4557245,4.5912848,6.096562,6.0814714,5.3910813,5.0779533,5.198677,4.798779,3.874486,3.4632697,3.0633714,2.6106565,2.493705,3.029418,3.4594972,3.7198083,3.6745367,3.1237335,2.1692593,1.8787673,1.9957186,2.1013522,1.6222287,0.9205205,0.6413463,0.7130261,1.0676528,1.6712729,1.9768555,1.9655377,2.0598533,2.4408884,3.0671442,2.7087448,2.2183034,1.8938577,1.8825399,2.203213,2.1881225,1.9957186,2.04099,2.3277097,2.4597516,2.565385,2.7502437,2.8332415,2.8445592,3.0256453,3.531177,3.4066803,3.2859564,3.2482302,2.8294687,3.0181,3.3727267,3.5877664,3.6481283,3.8405323,3.6934,2.9351022,2.8030603,3.2859564,3.1350515,2.5201135,1.9806281,1.6788181,1.6637276,1.8523588,2.3428001,3.0445085,3.8820312,4.5460134,4.4705606,4.093298,4.1612053,4.085753,3.6254926,2.9086938,2.1353056,1.2902378,1.5769572,2.9464202,4.093298,5.753253,4.8440504,4.564876,5.1458607,3.8820312,3.2821836,3.0671442,3.2142766,3.3953626,2.9954643,2.9464202,3.0746894,3.572676,4.266839,4.5912848,4.3083377,4.406426,4.5988297,4.7233267,4.7308717,5.4401255,5.798525,5.594803,5.093044,5.0477724,4.927048,4.798779,4.749735,4.7950063,4.9044123,5.372218,5.9682927,6.3153744,6.428553,6.696409,7.333983,8.028146,8.367682,8.341274,8.329956,9.009028,9.989911,11.148107,11.996947,11.68382,11.174516,10.914205,10.876478,10.985884,11.125471,11.197151,11.02361,10.514306,9.967276,10.099318,10.910432,11.261286,11.012292,10.465261,10.352083,9.280658,8.160188,7.4282985,7.0812173,6.6662283,6.8397694,6.8850408,6.8435416,6.7077274,6.4247804,6.3719635,6.0211096,5.6815734,5.3986263,4.938366,4.4139714,4.123479,3.7273536,3.2821836,3.2444575,3.308592,3.3915899,3.3123648,3.2557755,3.7952607,4.353609,4.7346444,4.568649,4.036709,3.863168,3.440634,3.6254926,4.13857,4.7233267,5.1647234,5.7607985,5.715527,5.6476197,5.9230213,6.643593,6.1003346,5.0025005,3.9197574,3.3048196,3.4670424,3.5538127,3.6896272,3.4972234,2.9728284,2.516341,1.8976303,1.8070874,1.81086,1.7580433,1.7919968,1.9768555,2.674791,3.821669,4.7950063,4.376245,3.6858547,3.8669407,3.9122121,3.6254926,3.6254926,4.304565,5.4174895,6.560595,7.533932,8.345046,8.782671,9.325929,9.918231,10.314357,10.061591,9.831461,9.846551,9.827688,9.771099,9.933322,10.193633,10.072908,10.378491,11.480098,13.328684,13.43809,12.596795,11.61214,10.982111,10.887795,11.223559,11.664956,12.204442,12.366665,11.216014,10.344538,10.502988,10.819888,10.853842,10.593531,11.170743,11.989402,12.694883,12.89106,12.14408,10.782163,9.876732,9.669238,10.167224,11.155652,11.532914,11.491416,11.638548,12.279895,13.392818,14.441608,14.286931,13.973803,13.9888935,14.252977,14.584969,14.762281,14.901869,15.32063,16.520325,17.572887,18.368912,19.357338,20.402355,20.772074,3.783943,4.123479,4.006528,3.7348988,3.4142256,2.938875,2.505023,2.4220252,2.4786146,2.5276587,2.474842,2.2560298,2.1164427,2.142851,2.2598023,2.1956677,2.2786655,2.4220252,2.6446102,2.9539654,3.350091,3.8178966,4.5120597,5.194905,5.6551647,5.692891,6.7454534,7.745199,8.639311,9.827688,12.15917,13.094781,15.380992,17.870924,18.534906,14.464244,6.5002327,3.3953626,2.3314822,1.6335466,0.7469798,0.7167987,0.5017591,0.38858038,0.47157812,0.6451189,0.7432071,0.8563859,0.84129536,0.70170826,0.6073926,0.84884065,1.2525115,1.5279131,1.5731846,1.478869,1.2147852,1.3958713,1.7127718,2.0862615,2.6483827,2.7917426,2.8181508,3.0256453,3.5802212,4.52715,5.534441,5.5382137,6.1116524,7.6697464,9.469289,12.14408,13.147598,13.4644985,14.905642,20.111864,24.797464,27.151583,28.007969,27.728794,26.212198,23.145054,19.60256,15.920478,12.053536,7.575431,4.123479,2.546522,2.033445,1.9806281,1.991946,2.3088465,2.625747,2.6295197,2.384299,2.3277097,2.4220252,2.8445592,3.7386713,4.8402777,5.492942,6.119198,6.4926877,5.9532022,4.983638,5.2137675,6.2625575,7.462252,9.42779,11.736636,12.909923,13.355092,11.785681,9.186342,7.0510364,7.3679366,9.522105,9.623966,8.827943,8.311093,9.258021,9.733373,8.75249,7.8131065,7.3905725,6.94163,6.470052,5.7306175,4.708236,3.7084904,3.3727267,0.91297525,0.5583485,0.7507524,0.83752275,1.1204696,0.84129536,1.4449154,2.0787163,2.41448,2.6182017,4.006528,4.266839,3.8669407,2.9841464,1.4977322,1.5052774,1.9240388,2.7389257,3.7650797,4.6554193,6.971811,7.7904706,8.156415,8.959985,10.944386,12.842015,15.16218,16.659912,18.082191,22.171717,19.76101,19.466745,21.398329,23.58645,22.01704,16.965494,16.263786,17.425755,18.7839,19.500698,21.609596,22.428255,22.613113,23.273323,25.978296,27.272306,29.366114,31.927725,34.817554,38.08465,37.2509,38.058243,38.08465,36.658596,34.847736,36.270016,40.114323,44.373615,47.723705,49.545883,50.3155,51.27752,51.024754,48.6895,43.939762,42.81552,42.249626,43.260693,46.418377,51.79814,55.668854,58.47946,62.142677,65.83608,66.002075,62.80666,60.543087,58.762405,57.856976,59.090626,62.508625,64.83256,65.37959,64.59111,64.03654,60.14319,58.841633,58.03429,56.200794,52.394215,47.957607,43.932217,41.827095,41.038616,38.84295,37.643253,36.986816,35.768257,33.583908,30.73935,28.754948,27.966469,27.385485,28.079647,33.187782,36.00593,36.71896,39.33339,45.01496,52.092407,58.098427,61.474926,69.78224,81.58679,86.46479,56.63842,32.83693,19.4592,17.53139,24.695602,15.599804,12.657157,11.634775,11.393328,13.856852,14.70192,13.35132,12.585477,12.777881,11.9064045,10.054046,8.639311,9.144843,10.461489,8.880759,12.619431,15.105591,14.400109,11.404645,9.903141,7.062354,7.4207535,9.148616,11.050018,12.551523,8.695901,5.081726,3.983892,4.666737,3.3764994,3.108643,3.0030096,3.3312278,4.0291634,4.7308717,8.918486,9.861642,9.64283,9.880505,11.774363,12.717519,13.679539,13.894578,13.830443,15.226315,13.109872,12.608112,12.777881,12.951422,12.736382,14.539697,15.905387,15.954432,14.894323,14.030393,14.837734,16.146835,17.625704,18.791445,19.036665,17.712475,13.947394,10.740664,8.722309,6.1305156,5.7381625,5.1760416,4.979865,5.081726,4.8063245,4.8855495,4.9647746,4.7874613,4.425289,4.266839,3.440634,3.218049,2.9426475,2.4559789,2.082489,1.5467763,0.87147635,0.55080324,2.1353056,8.262049,7.2585306,6.643593,6.1531515,5.704209,5.372218,3.8858037,2.5238862,1.8749946,1.901403,1.9730829,1.0714256,0.41876137,0.15467763,0.15845025,0.041498873,0.011317875,0.003772625,0.0,0.0,0.0,0.08677038,0.049044125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13958712,0.5583485,1.146878,1.5430037,1.599593,1.4524606,1.7127718,2.1466236,1.6825907,1.6976813,1.3958713,0.90543,0.4376245,0.27917424,0.13204187,0.79602385,2.6332922,4.851596,5.4665337,5.1156793,4.3649273,3.742444,3.3651814,2.9539654,4.5837393,5.191132,5.798525,6.6058664,7.01331,6.6624556,6.375736,5.987156,5.6061206,5.6287565,4.3121104,4.3196554,4.4101987,4.2291126,4.274384,5.0251365,4.164978,3.0030096,2.161714,1.5543215,1.3920987,1.3845534,1.901403,2.806833,3.4179983,3.4142256,3.519859,3.1350515,2.565385,3.029418,3.2482302,3.1350515,3.3123648,4.06689,5.330719,5.8626595,5.3571277,5.2137675,5.560849,5.2628117,3.8367596,3.4783602,3.2784111,2.9615107,2.8898308,3.3010468,3.4255435,3.519859,3.5462675,3.1765501,2.1541688,1.871222,1.9164935,1.8334957,1.1242423,0.63002837,0.5772116,0.9922004,1.6184561,1.8976303,1.8485862,1.7957695,1.8900851,2.1503963,2.4559789,2.0862615,1.8636768,1.7844516,1.8448136,2.033445,2.3880715,2.1051247,2.191895,2.7540162,2.9728284,2.5729303,2.5729303,2.7917426,3.0407357,3.1237335,2.9652832,3.138824,3.259548,3.1463692,2.8332415,3.0256453,3.5538127,3.8669407,4.0404816,4.798779,4.5837393,3.9348478,3.5123138,3.3350005,2.7615614,2.3277097,1.7882242,1.5203679,1.6184561,1.8787673,2.11267,2.4672968,3.108643,3.8292143,4.036709,3.6858547,3.6292653,3.4783602,3.0369632,2.2899833,1.5316857,1.0638802,1.3656902,2.4672968,3.9461658,4.557331,4.45547,4.5535583,4.8666863,4.5007415,4.1197066,3.832987,3.5500402,3.2444575,2.9426475,2.8596497,2.7691069,3.029418,3.5500402,3.7990334,3.942393,4.429062,4.7572803,4.8365054,4.9949555,5.6098933,5.8626595,5.5495315,4.9157305,4.640329,4.557331,4.5837393,4.6214657,4.689373,4.919503,5.613666,6.168242,6.398372,6.387054,6.488915,7.0284004,7.6508837,7.877241,7.756517,7.865923,8.858124,10.065364,11.227332,11.883769,11.378237,10.970794,10.895341,10.921749,10.887795,10.710483,10.740664,10.529396,10.359629,10.518079,11.268831,11.627231,11.6875925,11.408418,11.00852,10.948157,10.310584,9.35611,8.424272,7.598067,6.7114997,7.001992,6.881268,6.4549613,5.9532022,5.7004366,5.8098426,5.7419353,5.7419353,5.6023483,4.6327834,4.191386,3.9122121,3.6028569,3.2821836,3.2218218,3.2972744,3.4444065,3.5160866,3.7047176,4.5422406,4.851596,4.696918,4.3347464,3.9574835,3.6971724,3.5349495,4.0178456,4.847823,5.6853456,6.1342883,6.3116016,6.013564,5.881522,6.039973,6.1229706,4.9345937,3.7763977,3.2444575,3.2972744,3.259548,3.519859,3.4330888,2.9803739,2.3616633,2.0070364,1.6524098,1.7580433,1.9202662,1.9806281,2.0108092,2.7011995,3.3727267,4.002755,4.398881,4.191386,3.651901,3.7047176,3.7688525,3.7575345,4.1197066,4.7610526,5.534441,6.4511886,7.413208,8.190369,8.729855,9.2844305,10.023865,10.578441,10.016319,10.0465,10.110635,10.016319,9.767326,9.590013,10.593531,11.148107,11.212241,11.185833,11.9064045,12.012038,11.830952,11.374464,10.797253,10.401127,10.56335,11.140562,11.827179,12.253486,12.00072,11.608367,11.793225,11.966766,11.857361,11.498961,11.747954,12.37421,13.041965,13.257004,12.336484,10.846297,9.982366,9.876732,10.450171,11.41219,11.77059,11.736636,11.974312,12.67602,13.558814,13.970031,13.849306,14.0983,14.837734,15.399856,15.47908,15.546988,15.599804,15.954432,17.240896,17.655886,17.765291,18.263277,19.281887,20.394812,4.9421387,5.553304,4.8742313,4.2102494,3.9461658,3.561358,3.0407357,2.795515,2.7615614,2.897376,3.187868,3.1312788,2.9313297,2.7011995,2.5012503,2.3390274,2.4786146,2.6823363,2.9916916,3.3689542,3.6934,4.0178456,4.5422406,5.119452,5.6589375,6.149379,6.692637,7.2585306,8.043237,9.276885,11.200924,11.498961,12.619431,13.532406,13.475817,11.940358,6.149379,3.3350005,2.3993895,2.082489,0.9620194,0.56212115,0.38480774,0.4074435,0.55457586,0.7167987,0.6187105,0.68661773,0.7469798,0.7432071,0.7432071,1.0940613,1.6146835,1.7580433,1.5128226,1.3920987,1.2600567,1.8221779,2.1843498,2.173032,2.323937,2.384299,2.8521044,3.1652324,3.4066803,4.3196554,7.17176,6.9152217,6.63982,7.4471617,8.458225,10.808571,11.819634,12.487389,13.547497,15.467763,17.60684,17.689838,16.45619,14.664193,13.083464,10.970794,9.016574,7.454707,6.187105,4.798779,3.3425457,2.5314314,2.263575,2.2598023,2.071171,2.5389767,2.5993385,2.2484846,1.8221779,2.003264,2.4559789,3.380272,4.610148,5.8098426,6.48137,7.17176,7.2660756,6.360646,5.036454,4.8440504,6.039973,7.4169807,9.046755,11.031156,13.475817,14.622695,11.378237,8.68081,8.182823,8.288457,8.469543,7.5792036,6.349328,5.674028,6.620957,6.296511,6.2361493,6.175787,6.126743,6.4021444,6.198423,5.621211,4.6931453,3.8669407,4.032936,1.056335,0.5885295,0.8903395,1.0789708,1.1204696,0.724344,1.327964,2.142851,2.7691069,3.187868,2.9615107,2.546522,2.5578396,2.6898816,1.7316349,1.5958204,2.082489,2.7728794,3.62172,4.9421387,7.3981175,7.960239,7.7678347,7.6923823,8.318638,9.940866,12.1252165,14.517061,17.040947,19.889278,16.252468,17.4333,20.662666,22.631977,19.478064,15.871433,14.969776,14.943368,14.916959,14.954685,17.21826,19.534653,20.873934,21.432283,22.647068,22.624432,24.435291,27.317577,30.761984,34.511974,34.123394,34.719467,35.191048,35.02505,34.300705,34.459156,36.530327,40.269,44.17744,45.54313,44.39625,43.524776,43.528545,43.6455,41.744095,42.830612,42.615574,43.377644,45.758167,48.746086,50.97948,53.774998,57.67589,61.689964,63.28956,61.13916,57.10245,52.60171,49.61002,50.666355,55.3595,58.283283,59.55843,59.980965,61.029755,58.58132,56.85723,54.537067,51.247337,47.576572,45.561993,43.249374,41.340424,39.454113,36.137974,34.730785,34.447838,33.44432,31.456148,29.830147,28.079647,27.468483,27.298714,28.562544,33.94608,35.52681,35.621124,37.017,41.13293,48.00288,56.415833,58.943493,62.799114,71.25734,83.65796,60.5959,35.662624,19.312067,15.199906,20.183544,13.283413,11.046246,10.110635,9.846551,12.321393,12.510024,11.691365,10.729345,9.763554,8.201687,8.541223,10.518079,11.438599,10.540714,8.98262,12.166716,14.158662,12.147853,7.4735703,5.624984,5.455216,8.314865,9.767326,9.684328,12.264804,9.7296,5.907931,3.9310753,3.8141239,2.474842,2.1881225,1.961765,2.5880208,3.85185,4.5422406,9.537196,10.944386,10.446399,10.012547,11.895086,11.846043,13.192869,14.6151495,15.671484,16.788181,15.309312,15.30554,15.39231,15.045229,14.600059,16.758,17.410664,16.863634,15.731846,14.958458,16.776863,18.387774,19.666695,20.534397,20.960705,18.248188,14.11339,10.521852,8.122461,6.2399216,5.9909286,6.0701537,6.1342883,5.87775,5.0439997,5.1043615,5.0439997,4.9987283,4.817642,4.0517993,3.7499893,3.5575855,3.3689542,3.108643,2.7200627,1.7618159,1.0223814,0.62248313,2.727608,11.563096,5.885295,6.6247296,7.232122,5.8588867,5.342037,3.3010468,2.0183544,1.7316349,2.1390784,2.3692086,0.9318384,0.271629,0.0452715,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.05281675,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.116951376,0.1659955,0.32821837,0.7582976,1.5618668,1.5543215,1.4675511,1.539231,1.6410918,1.3015556,1.4034165,1.0110635,0.5357128,0.20372175,0.05281675,0.049044125,0.7507524,2.2560298,4.1762958,5.6287565,4.847823,4.255521,4.123479,4.0517993,2.9615107,4.164978,3.85185,3.4255435,3.6669915,4.7233267,6.0286546,6.0739264,5.753253,5.462761,5.0968165,4.1008434,3.983892,4.255521,4.561104,4.67051,4.9345937,3.7537618,2.637065,2.123988,1.8033148,1.569412,1.4335974,1.780679,2.4559789,2.7389257,2.7313805,3.4632697,3.6292653,3.1463692,3.127506,3.150142,3.361409,3.6934,4.142342,4.749735,5.0439997,5.0741806,5.0779533,5.149633,5.247721,3.9914372,3.4859054,3.2746384,3.1727777,3.2746384,3.4632697,3.3048196,3.3048196,3.4330888,3.1350515,2.0485353,1.7618159,1.7316349,1.5203679,0.7809334,0.5281675,0.6488915,1.1883769,1.8749946,2.1164427,1.7580433,1.7693611,1.8599042,1.8599042,1.750498,1.50905,1.5618668,1.7957695,2.0485353,2.1013522,2.335255,2.3201644,2.516341,2.927557,3.0822346,2.6710186,2.7426984,2.938875,3.0746894,3.097325,2.595566,2.8634224,3.1312788,3.0746894,2.8106055,3.1048703,3.7160356,4.1762958,4.5196047,5.3080835,5.0025005,4.4516973,3.7763977,3.0822346,2.444661,2.3616633,1.9202662,1.6448646,1.7052265,1.9391292,2.1956677,2.3654358,2.6898816,3.150142,3.4444065,3.410453,3.259548,3.029418,2.6710186,2.022127,1.6260014,1.3392819,1.4750963,2.2447119,3.7688525,4.3686996,5.2288585,5.0025005,4.093298,4.636556,5.1534057,5.142088,4.478106,3.5424948,3.229367,3.1425967,3.31991,3.4255435,3.451952,3.712263,4.08198,4.768598,5.1760416,5.194905,5.198677,5.4740787,5.6513925,5.43258,4.8327327,4.187614,4.1310244,4.4403796,4.6290107,4.6629643,4.961002,5.772116,6.33801,6.519096,6.4436436,6.519096,6.888813,7.194396,7.273621,7.201941,7.2924843,8.424272,9.748463,10.944386,11.661184,11.506506,11.332966,11.3669195,11.204697,10.77839,10.355856,9.971047,9.891823,10.253995,11.016065,11.921495,11.763044,11.747954,11.46878,11.083972,11.295239,11.11038,10.155907,8.967529,7.8432875,6.8737226,6.9454026,6.5266414,5.8136153,5.20245,5.292993,5.2099953,5.383536,5.6363015,5.534441,4.3875628,4.025391,3.8103511,3.6481283,3.500996,3.3878171,3.4142256,3.5274043,3.7235808,4.1197066,4.9459114,5.0968165,4.666737,4.221567,3.9763467,3.7763977,4.0480266,4.8063245,5.7683434,6.5455046,6.6586833,6.092789,6.1644692,6.432326,6.3116016,5.0968165,4.3611546,3.5424948,3.2255943,3.3840446,3.3878171,3.4859054,3.029418,2.3993895,1.8825399,1.6788181,1.5769572,1.6335466,1.7919968,2.0673985,2.5804756,3.3123648,3.6292653,3.6556737,3.5877664,3.6858547,3.350091,3.3651814,3.6179473,4.0517993,4.6554193,5.0666356,5.798525,6.5643673,7.2283497,7.7942433,8.416726,9.005256,9.793735,10.502988,10.314357,10.359629,10.506761,10.416218,10.080454,9.812597,10.585986,11.099063,11.038701,10.687846,10.940613,11.32542,11.59705,11.461235,10.93684,10.344538,10.3634,10.744436,11.442371,12.245941,12.800517,13.174006,13.234368,13.177779,12.989148,12.438345,12.272349,12.932558,13.622949,13.739901,12.883514,11.465008,10.502988,10.34831,10.955703,11.898859,12.2270775,12.457208,12.838243,13.328684,13.600313,13.6682205,13.9888935,14.671739,15.528125,16.090246,15.950659,15.814844,15.878979,16.380737,17.640795,17.542706,17.312576,17.527617,18.376457,19.644058,5.349582,5.832478,4.957229,4.395108,4.5007415,4.293247,3.8103511,3.500996,3.2633207,3.2105038,3.6707642,3.7990334,3.7198083,3.3048196,2.7804246,2.7011995,2.8181508,2.957738,3.270866,3.6971724,3.9725742,4.195159,4.4931965,4.889322,5.5306683,6.670001,7.224577,7.6131573,8.103599,9.050528,10.884023,11.498961,12.083718,11.68382,10.616167,10.469034,6.6813188,3.772625,2.4484336,2.1805773,1.1921495,0.5055317,0.4640329,0.77716076,1.056335,0.84129536,0.59607476,0.6828451,0.8601585,0.9620194,0.9016574,1.1204696,1.4449154,1.4260522,1.2223305,1.6184561,1.8863125,2.6219745,2.9237845,2.6936543,2.637065,2.795515,3.7575345,4.172523,4.025391,4.6327834,8.571404,7.865923,6.7680893,6.7114997,6.330465,5.8890676,6.1720147,7.356619,8.620448,8.114917,8.258276,8.710991,8.8618965,8.537451,7.986647,6.730363,6.149379,5.704209,5.0138187,3.8858037,2.8898308,2.4710693,2.3993895,2.4371157,2.3126192,2.9124665,2.6974268,2.2258487,2.0145817,2.5314314,3.5123138,4.9345937,6.224831,7.0849895,7.4773426,7.914967,7.9451485,7.4584794,6.696409,6.25124,7.907422,9.495697,10.299266,10.895341,13.162688,14.762281,10.33322,7.3000293,7.7640624,8.507269,7.3113475,5.7796617,4.4101987,4.0593443,5.9682927,6.6322746,5.451443,5.20245,6.138061,6.0022464,5.0666356,4.0404816,3.4066803,3.2029586,3.0445085,1.1053791,0.784706,1.0525624,1.2298758,0.9808825,0.8224323,1.7769064,2.9766011,3.9008942,4.3686996,2.3692086,1.0940613,1.3128735,2.8294687,4.4894238,2.5427492,2.4107075,2.704972,3.097325,4.315883,5.775889,5.975838,6.1003346,6.255012,5.485397,7.865923,9.476834,12.276122,15.271586,14.50197,11.283921,14.181297,17.157898,17.508753,15.863888,14.864142,14.3095665,13.415455,12.408164,12.555296,15.007503,17.942604,19.327158,19.036665,18.821627,18.787672,19.945868,22.450891,25.993385,29.799965,29.143528,29.830147,31.459919,32.72752,31.425966,31.882454,33.30096,36.194565,39.846466,42.276035,39.872875,37.115086,35.870117,36.35679,37.145267,39.1108,39.77101,41.295155,43.879402,45.743076,46.942772,50.251366,54.02399,57.132633,58.947266,57.411808,52.164085,45.950573,41.86482,43.309734,46.06375,47.546394,49.809967,53.250603,56.61201,55.53681,53.341145,49.806194,45.595947,42.26849,42.219448,41.925182,39.948326,36.371876,32.791656,31.097748,30.761984,29.652832,27.76652,27.19308,26.423466,26.638506,27.072357,28.29846,32.22576,32.218216,32.618114,34.428974,38.250645,44.283073,53.95608,57.423126,60.743034,66.68869,74.74702,58.70582,36.383194,20.036411,14.011529,14.694374,11.823407,10.729345,9.627739,8.933576,11.249968,9.307066,9.137298,8.741172,7.515069,6.258785,8.160188,13.736128,14.954685,11.283921,9.684328,13.660675,15.041456,11.676274,5.7079816,3.5387223,5.4212623,9.344792,9.952185,7.986647,10.321902,9.6201935,6.4964604,4.104616,3.1010978,1.6561824,1.7127718,1.5882751,2.1277604,3.1539145,3.4632697,7.937603,10.902886,11.287694,10.423763,12.061082,11.449917,12.136535,13.845533,15.739391,16.42601,17.056038,17.795471,17.84829,17.210714,16.686321,19.372429,19.278114,17.942604,16.614641,16.25624,19.123436,21.05502,21.473782,21.149336,22.209444,18.565088,14.030393,10.212496,7.884786,6.971811,6.043745,6.730363,7.33021,6.8963585,5.243949,5.311856,4.9723196,4.98741,5.1043615,4.055572,4.085753,3.8669407,3.6934,3.500996,2.8332415,1.7542707,1.750498,2.5238862,4.4743333,8.703445,5.7494807,8.926031,8.6581745,4.2064767,3.682082,1.7919968,1.6222287,2.1541688,2.6597006,2.704972,0.8111144,0.1659955,0.030181,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.0,0.060362,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2867195,0.2867195,0.20749438,0.30935526,0.90543,1.1204696,1.4373702,1.6184561,1.50905,1.0299267,0.90543,0.58475685,0.24522063,0.02263575,0.0150905,0.026408374,0.8903395,1.9164935,3.1425967,5.353355,4.164978,4.044254,4.315883,4.1083884,2.372981,3.1916409,2.6974268,1.9693103,1.8485862,2.9652832,4.7610526,4.6742826,4.768598,5.379763,5.1345425,3.8971217,3.6783094,4.1574326,4.719554,4.4516973,4.1197066,2.897376,2.0673985,1.9994912,2.1579416,1.9579924,1.7391801,1.9353566,2.3616633,2.2069857,1.9806281,3.0671442,3.9612563,4.1310244,3.9914372,3.338773,3.5764484,4.0480266,4.4177437,4.659192,4.3800178,4.870459,4.8327327,4.3385186,4.8327327,4.093298,3.4670424,3.2105038,3.3350005,3.5839937,3.6254926,3.3236825,3.2670932,3.3915899,2.9992368,1.9655377,1.569412,1.3996439,1.1506506,0.6413463,0.6073926,0.83752275,1.2336484,1.6637276,1.9542197,1.6712729,1.8297231,1.871222,1.629774,1.3317367,1.327964,1.4373702,1.8221779,2.3088465,2.384299,2.293756,2.625747,2.886058,2.9124665,2.8747404,2.8936033,3.0709167,3.059599,2.8747404,2.916239,2.595566,2.7011995,2.8936033,2.9426475,2.7426984,3.2821836,3.9801195,4.7044635,5.2892203,5.564622,4.851596,4.236658,3.4557245,2.625747,2.233394,2.372981,2.071171,1.7995421,1.7769064,1.9504471,2.2975287,2.4107075,2.4107075,2.4333432,2.625747,2.9916916,2.8596497,2.6483827,2.4408884,1.9881734,1.841041,1.6146835,1.7844516,2.5314314,3.7462165,4.7836885,5.9230213,5.119452,3.3048196,4.398881,5.572167,5.9192486,5.300538,4.2064767,3.7499893,3.802806,4.187614,4.2102494,3.9725742,4.3875628,4.5837393,5.2099953,5.6513925,5.6815734,5.451443,5.3910813,5.541986,5.4703064,4.961002,4.0480266,3.874486,4.4177437,4.8327327,4.9345937,5.191132,5.987156,6.677546,6.862405,6.6586833,6.696409,6.937857,6.828451,6.700182,6.6813188,6.692637,7.756517,9.152389,10.450171,11.404645,11.944131,12.136535,12.083718,11.457462,10.480352,9.9257765,9.242931,9.627739,10.536942,11.495189,12.083718,11.589504,11.642321,11.434827,11.0613365,11.510279,11.231105,10.186088,9.020347,7.967784,6.8774953,6.4964604,5.8702044,5.2552667,4.9459114,5.247721,4.878004,5.100589,5.353355,5.1873593,4.2706113,3.9650288,3.8292143,3.7990334,3.8065786,3.7688525,3.7650797,3.8895764,4.1498876,4.504514,4.8402777,4.9119577,4.4403796,4.0291634,3.9273026,4.044254,4.779916,5.7079816,6.519096,6.900131,6.5228686,5.541986,6.2021956,6.8359966,6.3116016,4.025391,4.376245,4.146115,3.7499893,3.5085413,3.6669915,3.2067313,2.5125682,1.9579924,1.6712729,1.5430037,1.7089992,1.5354583,1.569412,2.1315331,3.3161373,3.572676,3.4142256,3.0445085,2.7879698,3.1048703,3.0407357,3.138824,3.712263,4.610148,5.240176,5.3194013,6.19465,6.881268,7.145352,7.5075235,8.088508,8.726082,9.488152,10.344538,11.155652,10.789707,10.95193,10.978339,10.714255,10.499215,10.423763,10.159679,9.978593,10.125726,10.79348,11.52537,11.7894535,11.819634,11.672502,11.223559,11.151879,11.065109,11.529142,12.494934,13.283413,13.966258,13.656902,13.422999,13.502225,13.306048,12.887287,13.607859,14.241659,14.222796,13.641812,12.3289385,11.038701,10.601076,11.170743,12.242168,12.913695,13.58145,13.958713,13.958713,13.679539,13.977575,15.098045,15.965749,16.252468,16.395828,16.109108,15.645076,15.648849,16.305285,17.380484,17.20317,17.08999,17.45971,18.301004,19.161163,3.4934506,3.410453,3.470815,3.6481283,3.8782585,4.074435,3.8556228,3.7348988,3.6179473,3.451952,3.218049,3.0369632,3.1916409,3.1727777,2.9803739,3.127506,3.3236825,3.4444065,3.519859,3.5349495,3.4481792,3.874486,4.5309224,5.13077,5.6589375,6.379509,6.647365,7.786698,8.492179,8.601585,9.065618,11.714001,11.668729,9.929549,8.360137,9.688101,9.446653,5.8702044,2.7200627,1.4147344,1.0223814,0.5583485,0.77338815,1.5241405,1.9768555,0.6111652,0.7432071,0.90543,1.1091517,1.1959221,0.8526133,0.8186596,0.80734175,0.7054809,0.63002837,0.94692886,1.2638294,1.3166461,1.3091009,1.7957695,3.663219,2.5502944,2.1164427,2.6597006,3.9008942,4.9760923,5.583485,5.59103,5.9984736,6.9265394,7.598067,8.612903,9.955957,11.766817,13.570132,14.268067,11.619685,8.722309,6.8661776,6.1908774,5.692891,5.070408,5.379763,4.9760923,3.7499893,3.127506,2.7389257,2.4107075,2.3390274,2.4597516,2.4710693,2.4974778,2.4295704,2.4899325,3.0822346,4.7912335,5.938112,7.0774446,8.084735,8.869441,9.367428,10.284176,10.925522,10.906659,10.416218,10.208723,10.378491,9.989911,9.1976595,8.52236,8.865668,8.122461,6.828451,5.5495315,4.957229,5.798525,3.712263,3.308592,3.3161373,3.4179983,4.274384,4.7120085,4.0517993,3.3161373,3.048281,3.3425457,4.2706113,4.2819295,4.036709,3.5689032,2.2899833,1.8259505,1.5354583,1.7316349,2.0900342,1.6637276,2.04099,3.006782,4.104616,5.2326307,6.6360474,4.745962,2.8256962,2.8030603,6.722818,16.769318,7.284939,3.5764484,2.776652,3.059599,3.6330378,4.2064767,4.13857,4.52715,5.523123,6.3153744,9.039209,11.16697,11.204697,9.178797,6.6549106,9.850324,12.498707,13.6833105,13.996439,15.531898,15.569623,14.498198,13.479589,13.396591,14.86037,14.373701,13.777626,14.441608,15.792209,15.30554,16.316603,17.742655,19.794964,22.647068,26.44233,23.58645,24.491882,26.86109,29.279343,31.218472,28.181509,27.045948,27.706158,29.90937,33.278324,33.80649,33.002922,31.61837,30.62617,31.248653,31.788137,33.651814,36.983044,41.151794,44.75465,46.21843,49.09317,51.945274,54.261665,56.457333,54.431435,47.957607,41.566784,37.81679,37.292397,37.13395,39.457886,42.430714,46.30897,53.43546,54.073032,48.802677,43.943535,41.60828,39.703106,39.42393,38.29969,35.790894,32.206898,28.702131,26.638506,25.446356,24.378702,23.48459,23.605314,24.44661,25.8123,26.4876,26.928997,29.237844,29.626425,30.860073,32.92747,35.81353,39.472977,49.262936,54.752106,60.0451,64.54207,62.942474,51.443516,34.88169,22.062311,15.999702,13.902123,11.068882,11.076427,10.427535,8.7600355,8.820397,6.964266,7.032173,7.9300575,8.4544525,7.3075747,8.956212,14.366156,16.746683,14.517061,11.306557,18.361366,21.307787,16.950403,8.333729,4.745962,5.1835866,6.7039547,7.115171,6.719045,8.329956,7.707473,5.987156,4.1310244,2.535204,1.0223814,1.7429527,1.629774,1.7882242,2.3880715,2.6710186,9.556059,11.219787,11.52537,11.962994,11.657412,11.876224,10.668983,10.759526,12.521342,13.962485,16.376965,15.894069,15.905387,16.991903,16.905132,19.300749,21.088974,20.432537,18.417955,19.029121,20.907888,23.58268,23.503454,21.473782,22.658386,19.38752,14.769827,10.993429,9.314611,10.069136,7.2887115,7.24344,8.065872,8.246958,6.620957,7.598067,6.1418333,5.0968165,5.1534057,4.8365054,4.496969,4.776143,4.5799665,3.6292653,2.4559789,1.4939595,3.8065786,9.016574,12.291212,4.3347464,2.6974268,4.285702,4.504514,2.5691576,1.4939595,1.0299267,1.7769064,2.0447628,1.3996439,0.6413463,0.19994913,0.0452715,0.00754525,0.0,0.0,0.0,0.026408374,0.056589376,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2678564,0.32821837,0.36971724,0.47912338,0.62625575,0.80734175,1.146878,1.5241405,1.6033657,0.8224323,0.44516975,0.21503963,0.071679875,0.003772625,0.0150905,0.0150905,0.34330887,0.77716076,1.6524098,3.874486,3.6443558,4.146115,3.5387223,2.0296721,1.8448136,2.6295197,2.6672459,2.161714,1.720317,2.3805263,3.6368105,3.8782585,4.3686996,5.2665844,5.643847,2.6785638,2.505023,2.9766011,3.0369632,2.7313805,2.927557,2.1881225,1.750498,2.082489,2.916239,2.354118,2.4333432,2.565385,2.535204,2.4861598,2.8294687,3.3463185,3.5764484,3.5538127,3.783943,3.0030096,3.1010978,3.338773,3.6481283,4.6252384,5.2326307,5.73439,5.3910813,4.587512,4.8063245,3.8065786,3.2444575,3.3161373,3.7763977,3.9386206,3.9989824,3.8103511,3.7198083,3.6594462,3.1576872,2.3277097,1.7014539,1.237421,0.87147635,0.52062225,0.55457586,0.97710985,1.4449154,1.6712729,1.4034165,2.003264,2.1956677,2.033445,1.6976813,1.5241405,1.5618668,1.6071383,1.8448136,2.2598023,2.6408374,2.9803739,3.2142766,3.3161373,3.289729,3.1425967,2.9351022,2.7011995,2.4371157,2.2183034,2.1805773,2.535204,2.4597516,2.4899325,2.7804246,3.097325,3.5990841,4.6026025,5.572167,6.149379,6.149379,5.172269,4.5422406,3.6292653,2.625747,2.5616124,2.3314822,1.871222,1.4750963,1.3656902,1.6939086,1.8146327,2.0560806,2.0560806,1.8825399,2.0296721,2.1390784,2.11267,2.0560806,1.9881734,1.8297231,1.6712729,1.7882242,2.637065,3.9197574,4.5761943,4.3347464,4.2819295,4.4894238,4.8742313,5.20245,3.7009451,3.2369123,3.4594972,3.8480775,3.6783094,3.99521,4.432834,4.7233267,4.961002,5.583485,5.534441,5.96452,6.1720147,6.096562,6.3153744,6.156924,6.043745,5.873977,5.5004873,4.7308717,4.217795,4.564876,5.2250857,5.7909794,5.9984736,6.7039547,7.515069,7.707473,7.281166,6.9265394,7.062354,6.828451,6.458734,6.2889657,6.790725,7.7187905,9.122208,10.246449,11.091517,12.419481,13.275867,12.883514,11.657412,10.38981,10.253995,10.314357,10.868933,11.517824,12.049765,12.449662,12.219532,12.351574,12.438345,12.242168,11.717773,10.718028,9.982366,9.34102,8.401636,6.5455046,5.6287565,5.3382645,5.349582,5.342037,4.991183,5.0515447,5.2137675,5.1345425,4.7346444,4.2102494,3.893349,3.6971724,3.7009451,3.9386206,4.3800178,4.3196554,4.6327834,5.1081343,5.3646727,4.851596,4.425289,3.712263,3.4632697,3.8593953,4.5309224,5.3382645,6.2436943,6.7077274,6.511551,5.7683434,5.7796617,6.0286546,5.956975,5.3080835,4.134797,3.7914882,3.7273536,3.9348478,4.08198,3.4934506,2.565385,2.04099,1.8033148,1.7014539,1.5580941,2.2296214,1.9202662,1.9202662,2.6936543,3.8895764,3.7462165,3.3764994,2.8709676,2.516341,2.8219235,3.2369123,3.6971724,4.38379,5.20245,5.8136153,5.6287565,6.043745,6.590776,7.115171,7.752744,8.75249,9.669238,10.555805,11.506506,12.679792,11.593277,11.34051,11.302785,11.09529,10.559577,10.38981,10.246449,10.152134,10.099318,10.023865,10.416218,10.989656,11.876224,12.615658,12.178034,11.566868,11.623458,12.068627,12.796744,13.8719425,13.675766,12.864652,12.445889,12.951422,14.464244,14.332202,14.864142,15.128226,14.739646,13.8870325,12.298758,10.582213,9.688101,10.03141,11.521597,13.3626375,14.566105,15.067864,15.0376835,14.875461,15.486626,16.984358,17.799244,17.580433,17.225805,16.667458,15.784663,15.611122,16.195879,16.588232,17.074902,17.252214,18.002966,19.210207,19.76101,3.0897799,3.5538127,3.3123648,3.048281,2.957738,2.7313805,2.8634224,2.957738,3.2369123,3.62172,3.7198083,3.2935016,3.1463692,3.0256453,2.8709676,2.8106055,3.1237335,3.470815,3.7273536,3.821669,3.7650797,3.9386206,4.4441524,5.0025005,5.6325293,6.647365,6.7869525,7.564113,8.179051,8.348819,8.296002,10.86516,10.091772,9.650374,11.0613365,13.679539,12.713746,8.239413,4.4441524,2.897376,2.535204,2.372981,1.8863125,1.4034165,0.97333723,0.36594462,0.46026024,0.68661773,0.8299775,0.77716076,0.513077,0.5357128,0.6149379,0.87902164,1.3958713,2.142851,3.1614597,3.874486,4.8553686,5.9682927,6.360646,5.9532022,6.017337,6.560595,7.533932,8.831716,9.186342,8.941121,9.148616,10.072908,11.174516,13.615403,14.1058445,14.132254,13.656902,11.129244,7.9262853,5.7607985,4.8327327,4.7610526,4.5912848,4.293247,4.4705606,4.561104,4.5007415,4.738417,5.372218,4.9232755,4.3309736,3.9725742,3.6330378,4.2404304,4.8629136,5.5457587,6.432326,7.7829256,8.439363,9.046755,9.6201935,10.227587,10.978339,11.378237,11.846043,11.872451,11.332966,10.487898,9.144843,8.114917,7.0284004,6.013564,5.692891,5.6325293,5.13077,4.5422406,4.2706113,4.7610526,3.610402,2.6936543,2.3578906,2.7426984,3.783943,3.4142256,3.0143273,2.6898816,2.4220252,2.0598533,2.1768045,2.3616633,2.7691069,3.2067313,3.1048703,1.7731338,1.4411428,1.841041,2.3616633,2.04099,3.5047686,5.062863,6.0362,6.983129,9.665465,4.851596,3.4859054,4.0593443,6.3455553,11.363147,7.745199,5.7117543,4.255521,3.3425457,3.874486,4.6931453,5.142088,5.3269467,5.6325293,6.7077274,8.179051,8.499724,7.5905213,6.485142,7.3377557,8.601585,11.140562,13.079691,13.966258,14.750964,13.422999,12.332711,11.344283,10.967021,12.336484,12.860879,13.381501,14.735873,16.293968,15.950659,16.524097,17.452164,18.263277,19.078165,20.60985,20.330677,21.1267,22.432028,23.650587,24.17498,22.22076,22.454664,24.163664,26.649822,29.237844,30.143274,30.316814,29.882963,29.694332,31.324106,32.444576,35.572083,38.767494,40.910347,41.69128,45.743076,48.878128,50.232502,50.341908,51.12284,49.115807,44.93951,40.118095,36.33038,35.375904,34.327114,35.191048,37.46594,41.706367,49.530792,53.944763,50.10046,44.388706,39.83892,36.126656,32.350258,30.954388,29.177483,26.355558,23.918442,22.997923,22.22076,21.65864,21.402102,21.553007,23.209188,24.899324,26.121656,27.23458,29.441565,29.188799,29.886736,30.36963,31.041159,33.88572,43.498367,50.266457,56.385654,60.754353,58.988766,51.59819,38.484547,27.113855,20.006231,14.694374,11.646093,11.642321,10.650121,8.201687,7.4018903,6.1041074,6.0776987,7.2924843,8.624221,7.84706,8.243186,13.158916,15.441354,13.758763,12.58925,20.806026,23.609087,19.440336,11.072655,5.5985756,6.205968,6.881268,6.741681,6.089017,6.3908267,6.0022464,4.851596,3.6556737,2.6332922,1.50905,1.4298248,1.358145,1.5958204,2.1390784,2.6823363,11.510279,15.214996,17.063583,17.071129,12.012038,12.015811,9.963503,8.926031,10.408672,14.32843,15.086727,14.988639,15.920478,17.961468,19.410156,19.927006,21.032385,20.643805,18.987621,18.599041,19.04421,21.420965,21.719002,20.145817,21.145563,20.051502,16.939087,13.302276,10.672756,10.61994,8.880759,8.20546,8.062099,7.911195,7.194396,6.8359966,5.613666,5.032682,5.3080835,5.3609,4.930821,4.9119577,4.7610526,4.115934,2.7879698,1.7240896,5.798525,7.3415284,4.825187,2.8822856,1.9391292,2.123988,2.0108092,1.2826926,0.72811663,0.573439,0.68661773,0.7205714,0.5281675,0.150905,0.0452715,0.030181,0.02263575,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23013012,0.3055826,0.2263575,0.2678564,0.9922004,0.754525,0.965792,1.3241913,1.4637785,0.94692886,0.28294688,0.1358145,0.09808825,0.018863125,0.003772625,0.003772625,0.26031113,0.543258,1.1129243,2.7389257,2.7728794,2.746471,2.161714,1.2940104,1.1996948,2.7992878,3.4029078,3.3878171,3.0181,2.4786146,2.8747404,2.6182017,3.199186,4.346064,4.0103,1.8523588,1.5316857,1.6410918,1.5241405,1.267602,1.6675003,1.4939595,1.6825907,2.4371157,3.2067313,3.308592,3.3350005,3.2746384,3.059599,2.5729303,3.218049,3.8141239,4.5007415,5.1081343,5.1760416,3.9273026,3.8480775,3.772625,3.5349495,3.9650288,5.7570257,6.1418333,5.4891696,4.617693,4.8063245,4.0782075,3.440634,3.4896781,4.104616,4.436607,4.1083884,3.8669407,3.7650797,3.6896272,3.3538637,2.463524,1.7693611,1.1846043,0.72811663,0.52062225,0.7696155,1.237421,1.5015048,1.4637785,1.3430545,1.8636768,1.8033148,1.4864142,1.2411937,1.4034165,1.5279131,1.5882751,1.871222,2.4408884,3.1539145,3.1425967,3.0822346,2.8256962,2.5276587,2.655928,2.848332,2.5389767,2.2899833,2.2786655,2.2786655,2.6521554,2.6182017,2.5427492,2.6898816,3.2331395,4.036709,4.9459114,5.6778007,6.066381,6.0776987,4.776143,4.191386,3.7763977,3.3727267,3.2331395,2.4371157,1.9429018,1.6561824,1.5316857,1.5958204,1.599593,1.5769572,1.5241405,1.5241405,1.750498,1.8787673,1.8863125,1.9730829,2.1843498,2.4182527,2.5804756,2.9011486,3.338773,3.85185,4.38379,4.7346444,4.67051,4.979865,5.413717,4.689373,4.0782075,3.9122121,3.8556228,3.8103511,3.9348478,4.738417,5.0553174,5.4212623,5.8890676,6.0248823,5.926794,5.915476,6.0512905,6.2625575,6.3644185,6.432326,6.579458,6.3832817,5.87775,5.5495315,5.3382645,5.643847,6.2361493,6.7831798,6.862405,7.356619,7.707473,7.816879,7.6848373,7.4282985,7.201941,6.7379084,6.3719635,6.307829,6.643593,7.141579,8.224322,9.367428,10.499215,12.004493,12.294985,11.717773,11.019837,10.582213,10.450171,11.329193,12.053536,12.600568,13.04951,13.600313,13.132507,12.887287,12.706201,12.419481,11.815862,10.884023,10.27663,9.49947,8.152642,5.934339,5.353355,5.0175915,4.9534564,5.028909,4.9760923,5.1458607,5.0062733,4.7535076,4.3649273,3.5764484,3.4745877,3.5651307,3.7160356,3.9763467,4.561104,4.881777,5.2552667,5.534441,5.492942,4.8025517,3.9650288,3.561358,3.8065786,4.5007415,5.0553174,6.0286546,6.7341356,6.6360474,5.832478,5.05909,4.927048,5.081726,5.119452,4.772371,3.904667,3.4557245,3.9008942,4.2592936,3.9989824,3.0445085,2.1541688,1.720317,1.6184561,1.6825907,1.7014539,1.9164935,2.233394,2.5917933,3.1916409,4.4630156,3.9876647,3.4632697,2.9916916,2.746471,2.9803739,3.6896272,4.22534,4.4931965,4.8629136,6.156924,6.3342376,6.515323,6.7077274,7.0963078,8.031919,8.612903,9.344792,10.514306,11.623458,11.3971,11.053791,11.11038,11.080199,10.748209,10.182315,10.38981,10.751981,11.042474,10.993429,10.291721,10.155907,11.02361,12.049765,12.574159,12.113899,11.242422,10.514306,10.653893,11.593277,12.50248,12.687338,12.928786,13.430545,14.094527,14.5132885,13.822898,13.822898,14.075664,13.8870325,12.298758,10.684074,10.197406,10.676529,11.7894535,13.034419,15.211224,16.0412,15.905387,15.343266,15.049001,15.735619,17.255987,17.836971,17.176762,16.433554,16.086473,16.026112,16.524097,17.41821,18.112373,18.542452,18.961214,19.21398,19.18757,18.806536,3.2029586,3.6896272,3.3878171,2.9992368,2.7804246,2.5691576,2.6710186,2.8709676,3.2369123,3.5877664,3.5160866,3.380272,3.2784111,3.2105038,3.150142,3.0256453,3.2859564,3.6443558,3.863168,3.9348478,4.08198,4.3913355,4.8629136,5.4438977,6.1116524,6.8699503,7.1264887,7.6848373,8.239413,8.526133,8.311093,9.420244,9.137298,9.805053,11.691365,12.985375,11.170743,8.273367,5.613666,3.904667,3.2444575,3.1237335,1.9579924,0.94315624,0.5319401,0.43385187,0.47535074,0.73188925,0.784706,0.5696664,0.39989826,0.38480774,0.49421388,0.7469798,1.1544232,1.7467253,2.3767538,3.0143273,3.9197574,4.776143,4.6818275,5.342037,5.9192486,6.7567716,7.858378,8.888305,10.668983,10.665211,10.416218,10.582213,10.933067,11.306557,10.646348,9.442881,7.786698,5.3910813,3.62172,2.71629,2.7426984,3.5047686,4.538468,4.2027044,4.1083884,4.255521,4.715781,5.6287565,6.8925858,7.2283497,7.2170315,7.122716,6.888813,7.9828744,9.058073,10.163452,11.427281,13.041965,13.690856,13.79649,13.162688,11.944131,10.631257,10.499215,10.601076,10.650121,10.423763,9.782416,8.243186,7.152897,6.507778,6.609639,8.09228,6.4964604,5.828706,4.534695,3.169005,4.3913355,3.0218725,2.425798,2.1692593,2.0862615,2.2711203,2.0636258,1.9957186,2.003264,1.9391292,1.5845025,2.071171,2.5767028,3.0822346,3.3048196,2.6898816,1.9806281,2.2598023,2.5389767,2.4408884,2.2371666,3.7273536,6.3644185,7.1793056,6.983129,10.340765,4.708236,3.5689032,3.7160356,4.323428,6.934085,6.485142,9.703192,9.1976595,4.9987283,4.5422406,5.6400743,5.96452,6.1644692,6.749226,8.088508,8.031919,8.013056,7.1000805,5.975838,6.9491754,7.4735703,10.008774,12.310076,12.958967,11.351829,9.884277,9.891823,9.865415,9.876732,11.548005,13.045737,13.355092,13.6682205,14.143571,13.898351,15.648849,17.006994,18.206688,19.164934,19.470518,21.50019,21.383238,21.296469,21.28515,19.266796,18.606586,19.383747,21.24365,23.416683,24.740875,26.438557,27.438301,28.245644,29.645287,32.697342,35.043915,37.914883,39.91437,40.631172,40.668896,43.528545,46.04866,47.237038,47.029545,46.29388,44.158577,42.09872,39.352253,36.307743,34.474247,33.021786,32.79543,34.315796,37.89979,43.65682,49.821285,48.8819,44.52075,39.30698,34.71192,30.00746,26.393284,23.94485,22.537663,21.851044,20.330677,20.266542,20.647577,20.787165,20.345766,21.922724,23.89958,25.895298,27.819336,29.87919,28.796446,28.02683,27.5213,27.800474,29.932007,36.54919,42.027042,47.719933,52.609257,53.32228,52.231995,44.89801,34.383705,23.793945,16.25624,12.268577,10.653893,9.171251,7.303802,6.2625575,5.6891184,5.613666,6.4436436,7.605612,7.5490227,7.9715567,11.117926,12.3289385,11.3971,12.562841,20.036411,23.552498,20.557034,12.875969,6.7114997,6.858632,7.91874,7.5603404,5.8173876,5.081726,4.957229,4.0291634,3.1576872,2.5012503,1.5052774,1.1959221,1.3845534,1.81086,2.293756,2.757789,6.820906,11.031156,14.305794,15.460217,13.215506,12.815607,10.114408,8.469543,9.74469,14.302021,14.679284,15.147089,16.991903,19.579924,20.36463,20.647577,22.183035,22.756474,21.869907,20.745665,18.708447,23.035648,23.593996,19.821371,20.756983,20.360857,18.104828,14.924504,12.245941,11.98563,10.831206,9.6051035,8.763808,8.273367,7.6320205,6.7831798,6.0248823,5.3458095,4.9534564,5.281675,4.678055,4.432834,4.2819295,3.9084394,2.9501927,1.9730829,3.5047686,3.6141748,1.9429018,1.6939086,1.1732863,0.91674787,1.3091009,1.7014539,0.43385187,1.2525115,4.315883,4.055572,0.6526641,0.011317875,0.003772625,0.0754525,0.11317875,0.0754525,0.018863125,0.018863125,0.030181,0.02263575,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.20372175,0.21503963,0.24899325,0.69039035,0.95447415,1.0186088,0.90543,0.69039035,0.52062225,0.23390275,0.1056335,0.0452715,0.011317875,0.0,0.0,0.16222288,0.3169005,0.76584285,2.2748928,4.032936,3.410453,2.5540671,2.1013522,1.1921495,3.270866,4.878004,4.564876,2.938875,2.674791,2.6974268,2.305074,3.0860074,4.647874,4.617693,2.2899833,1.1355602,0.7054809,0.663982,0.77338815,1.1883769,1.6109109,2.3390274,3.399135,4.5535583,4.515832,3.7575345,3.4632697,3.5953116,2.897376,3.5651307,4.06689,4.715781,5.515578,6.145606,5.7079816,4.881777,4.036709,3.5651307,3.8820312,5.6023483,6.2361493,6.0286546,5.4288073,5.100589,4.285702,3.7650797,3.8782585,4.4101987,4.5988297,3.9159849,3.7914882,3.863168,3.7688525,3.1539145,2.5314314,1.8297231,1.2185578,0.7809334,0.5017591,0.90920264,1.418507,1.5845025,1.4034165,1.3091009,1.539231,1.4524606,1.2336484,1.1204696,1.4109617,1.4901869,1.5769572,1.8334957,2.323937,3.006782,2.7615614,2.5125682,2.252257,2.0560806,2.11267,2.3390274,2.0975795,1.9164935,1.9655377,2.0560806,2.5616124,2.6144292,2.5767028,2.7011995,3.138824,3.8858037,4.938366,5.938112,6.470052,6.058836,5.1534057,4.5950575,3.9725742,3.3425457,3.229367,2.6785638,2.2296214,1.9466745,1.8146327,1.7542707,1.6410918,1.4600059,1.3053282,1.2789198,1.4939595,1.8334957,2.0787163,2.2183034,2.4031622,2.938875,2.757789,3.3538637,3.8707132,4.002755,4.002755,4.534695,4.5120597,5.198677,6.149379,5.2137675,4.991183,5.081726,5.0477724,4.9345937,5.2628117,5.836251,5.828706,5.8626595,6.0550632,5.9796104,6.0211096,6.217286,6.3945994,6.519096,6.670001,6.507778,6.6662283,6.7077274,6.549277,6.477597,6.4511886,6.809588,7.3000293,7.673519,7.647111,7.7414265,7.854605,7.9036493,7.8734684,7.809334,7.111398,6.515323,6.1720147,6.1531515,6.4247804,6.7039547,7.4773426,8.703445,10.148361,11.3971,11.763044,11.291467,10.838752,10.763299,10.899114,11.732863,12.845788,13.698401,14.173752,14.588741,13.947394,13.494679,12.966512,12.23085,11.291467,10.638803,10.201178,9.265567,7.6131573,5.5193505,5.2288585,4.881777,4.5724216,4.5309224,5.119452,5.168496,4.9534564,4.7535076,4.459243,3.591539,3.3463185,3.6669915,4.0706625,4.3686996,4.6554193,5.149633,5.4967146,5.5382137,5.1873593,4.425289,3.8593953,4.0103,4.610148,5.4212623,6.2323766,7.0170827,7.1604424,6.485142,5.481624,5.323174,5.100589,4.8629136,4.534695,4.2328854,4.266839,4.142342,4.4101987,4.376245,3.7650797,2.7389257,1.8938577,1.4373702,1.3920987,1.5845025,1.6373192,1.8033148,2.4408884,3.0218725,3.500996,4.3422914,3.5462675,3.059599,2.8709676,2.938875,3.1954134,3.5802212,4.085753,4.398881,4.8553686,6.4134626,6.6020937,6.964266,7.3868,8.047009,9.420244,9.529651,9.752235,10.453944,11.18206,10.676529,10.661438,10.510533,10.484125,10.533169,10.295494,10.023865,10.340765,10.970794,11.434827,11.057564,10.823661,11.604594,12.623203,13.162688,12.566614,11.25374,10.253995,10.661438,12.147853,12.985375,13.573905,14.068119,14.464244,14.6151495,14.234114,13.909668,13.675766,13.6682205,13.59654,12.725064,11.849815,12.091263,13.019329,14.27184,15.535669,17.282394,17.399347,16.644821,15.735619,15.347038,15.841252,17.176762,17.723793,17.120173,16.263786,16.048746,16.437326,17.150352,17.931286,18.53868,19.021576,19.191343,19.274342,19.429018,19.73083,3.7763977,4.06689,3.7688525,3.3312278,3.0143273,2.867195,3.1916409,3.350091,3.5500402,3.7160356,3.4896781,3.2520027,3.1765501,3.2067313,3.2520027,3.2029586,3.2972744,3.5424948,3.663219,3.7348988,4.191386,4.779916,5.349582,5.8928404,6.3945994,6.8397694,7.33021,8.348819,9.533423,10.378491,10.223814,10.159679,10.989656,11.830952,12.064855,11.336739,12.619431,11.947904,9.352338,5.783434,3.108643,2.6521554,1.388326,0.513077,0.40367088,0.6451189,0.7130261,0.73566186,0.66020936,0.513077,0.4074435,0.41876137,0.51684964,0.6526641,0.8224323,1.0374719,1.2713746,1.7542707,2.3692086,2.8332415,2.6898816,3.6669915,4.719554,5.8588867,6.907676,7.5301595,9.88805,9.654147,8.873214,8.412953,7.9753294,6.8699503,5.904158,4.8100967,3.7914882,3.500996,2.4559789,2.9313297,4.274384,5.832478,6.94163,6.670001,6.7567716,7.0359454,7.6282477,8.971302,11.314102,12.657157,13.185325,12.940104,11.830952,12.498707,14.0983,16.188334,18.23687,19.63274,19.621422,18.595268,16.769318,14.50197,12.30253,10.9594755,10.125726,10.038955,10.272858,9.74469,8.703445,8.669493,8.401636,7.8395147,8.080963,6.0512905,4.847823,3.4217708,2.3201644,3.6896272,2.686109,2.323937,2.0636258,1.720317,1.4449154,1.3355093,1.2826926,1.3468271,1.418507,1.2298758,1.9579924,2.4069347,3.108643,3.8141239,3.500996,2.474842,2.4786146,2.7502437,2.8747404,2.7615614,4.3007927,6.8661776,7.911195,8.145098,11.498961,5.1760416,3.2142766,2.8256962,3.1048703,5.036454,6.296511,11.348056,11.966766,7.7338815,6.0362,6.1305156,5.926794,6.2663302,7.4207535,9.107117,8.552541,7.809334,6.587003,5.5306683,6.221059,8.13378,10.823661,12.306303,11.581959,8.661947,8.280911,8.356364,8.843033,9.533423,10.0276375,11.231105,11.548005,11.902632,12.657157,13.641812,14.683057,16.244923,18.297232,20.29295,21.179516,22.854563,22.01704,20.75321,19.63274,17.72002,17.41821,18.23687,19.798737,21.432283,22.19058,24.133482,25.687803,27.34776,29.788647,33.855537,36.545418,38.59018,39.98228,40.72926,40.88771,40.521767,41.200836,42.389214,43.38519,43.321053,41.679962,40.540627,39.042896,36.900043,34.410114,32.55398,31.682505,32.85202,35.855026,39.23153,43.637955,44.886692,43.351234,39.49561,33.881947,29.41893,24.476791,21.477554,20.741892,20.470263,18.987621,19.28566,20.006231,20.360857,20.145817,21.545462,23.726038,26.09902,28.192827,29.652832,28.464457,26.461191,25.208681,25.257725,26.1292,30.086685,33.98758,39.024033,44.388706,47.289856,52.605484,49.74206,40.06905,27.683523,19.406384,13.155144,10.510533,8.929804,7.277394,5.828706,6.017337,5.9230213,6.149379,6.7152724,7.066127,7.7678347,8.899622,8.933576,8.495952,10.359629,16.373192,21.409647,20.987112,15.056546,7.997965,6.439871,7.654656,7.635793,5.715527,4.5761943,4.0216184,3.270866,3.0218725,2.9803739,1.8749946,1.2525115,1.4034165,1.8900851,2.4333432,2.886058,3.7009451,6.8246784,9.922004,11.774363,12.264804,13.392818,10.967021,9.137298,10.186088,14.558559,14.958458,15.894069,18.12369,20.745665,21.202152,20.979568,24.616379,25.416174,22.843245,22.511253,18.976303,22.767792,23.307278,19.591242,20.194862,19.57615,17.629477,15.192361,13.396591,13.679539,12.657157,11.219787,9.767326,8.567632,7.7225633,6.858632,6.85486,6.043745,4.5535583,4.2894745,3.742444,3.7801702,3.85185,3.6292653,2.9992368,2.2371666,1.6637276,1.2336484,0.9393836,0.80734175,0.5583485,0.35462674,0.814887,1.3656902,0.24522063,1.7127718,4.7912335,4.221567,0.5281675,0.0,0.003772625,0.211267,0.573439,0.76584285,0.18485862,0.07922512,0.0452715,0.02263575,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18485862,0.33576363,0.3961256,0.47157812,0.87902164,1.116697,0.8941121,0.41498876,0.35839936,0.36594462,0.17731337,0.030181,0.0,0.0,0.0,0.10186087,0.1961765,0.633801,2.2107582,3.772625,4.115934,4.376245,4.247976,1.9693103,4.1008434,6.436098,5.8702044,3.1199608,2.7389257,2.674791,2.1013522,2.546522,4.0178456,4.9949555,2.8558772,1.327964,0.5281675,0.41498876,0.76584285,1.0789708,1.8938577,3.0633714,4.2706113,5.036454,4.644101,3.8480775,3.6858547,4.0706625,3.7688525,4.398881,4.508287,4.738417,5.323174,6.0739264,7.3905725,6.2135134,4.696918,3.9499383,4.0480266,5.304311,6.205968,6.326692,5.832478,5.4703064,4.447925,4.2592936,4.515832,4.745962,4.38379,3.6971724,3.682082,3.8292143,3.6934,2.886058,2.5389767,1.8976303,1.2864652,0.84884065,0.543258,1.0676528,1.448688,1.4901869,1.3015556,1.3204187,1.3694628,1.3468271,1.2336484,1.1581959,1.3958713,1.4109617,1.6109109,1.9353566,2.3503454,2.8596497,2.3956168,2.1164427,1.9994912,1.9730829,1.9089483,2.0447628,1.9240388,1.81086,1.871222,2.1843498,2.546522,2.5540671,2.5616124,2.8181508,3.440634,4.0970707,5.251494,6.466279,7.118943,6.3945994,5.80607,5.353355,4.5120597,3.5538127,3.5387223,3.169005,2.7841973,2.4823873,2.2711203,2.082489,1.9240388,1.7089992,1.5015048,1.4071891,1.569412,1.8976303,2.354118,2.6446102,2.8181508,3.2746384,3.1463692,3.6783094,4.1800685,4.3800178,4.432834,4.6742826,5.0666356,5.670255,6.326692,6.651138,6.6247296,6.5945487,6.5228686,6.515323,6.8171334,6.9152217,6.5455046,6.1795597,6.058836,6.168242,6.519096,6.881268,7.0170827,6.9189944,6.8246784,6.5756855,6.696409,6.8963585,7.009537,7.001992,7.118943,7.4811153,7.7829256,7.854605,7.6584287,7.647111,7.7829256,7.8508325,7.798016,7.7225633,6.790725,6.304056,6.1003346,6.089017,6.25124,6.48137,7.032173,8.345046,10.016319,10.804798,11.129244,10.846297,10.714255,11.065109,11.796998,12.344029,13.370183,14.252977,14.735873,14.939595,14.57365,13.815352,12.951422,12.0724,11.042474,10.612394,10.155907,9.122208,7.496206,5.7909794,5.304311,4.8968673,4.5988297,4.5837393,5.1647234,4.9044123,4.745962,4.6742826,4.496969,3.8103511,3.500996,3.874486,4.3121104,4.5120597,4.52715,4.9157305,5.198677,5.062863,4.5535583,4.0706625,4.085753,4.6554193,5.4363527,6.2323766,7.001992,7.4697976,7.0963078,6.2625575,5.594803,5.9796104,5.485397,4.889322,4.429062,4.3649273,4.979865,5.0477724,4.8440504,4.1197066,3.0709167,2.335255,1.7127718,1.358145,1.3619176,1.5731846,1.5845025,1.8976303,2.7087448,3.5990841,4.187614,4.1536603,3.0218725,2.6219745,2.7011995,2.9992368,3.218049,3.3312278,3.651901,4.1310244,4.9157305,6.349328,6.7077274,7.2283497,7.8319697,8.612903,9.876732,9.865415,10.03141,10.608622,11.227332,10.917976,11.200924,10.978339,10.914205,11.068882,10.884023,9.906913,9.812597,10.378491,11.11038,11.23865,11.272603,11.876224,12.638294,12.97783,12.121444,11.461235,11.053791,11.763044,13.215506,13.792717,14.358611,14.637785,14.656648,14.392565,13.762536,13.913441,13.815352,13.864397,14.022847,13.837989,13.373956,13.732355,14.747191,16.060064,17.105082,18.029375,17.923742,17.05981,15.961976,15.377219,16.048746,17.248442,17.67852,17.139036,16.561823,16.150608,16.452417,17.16167,17.946377,18.459454,18.7839,18.976303,19.500698,20.349539,21.043703,4.2706113,4.29702,4.0216184,3.7235808,3.4934506,3.229367,3.8065786,3.7650797,3.7198083,3.8141239,3.7160356,3.0520537,2.8407867,2.8898308,3.0181,3.059599,3.0030096,3.2067313,3.410453,3.6669915,4.3385186,4.9760923,5.59103,6.0022464,6.2399216,6.571913,7.424526,9.352338,11.631002,13.358865,13.445636,13.20796,14.909414,15.203679,13.611631,12.54775,19.711966,19.779873,14.784918,7.673519,2.3126192,1.4977322,0.7884786,0.38858038,0.38103512,0.7130261,0.8111144,0.5470306,0.41876137,0.49421388,0.43007925,0.51684964,0.5885295,0.6790725,0.7582976,0.72811663,0.8601585,1.2864652,1.7429527,2.0636258,2.1843498,2.8747404,4.244203,5.5268955,6.3908267,6.937857,8.329956,7.673519,6.8397694,6.428553,5.7570257,4.644101,3.9499383,3.5575855,3.8178966,5.5683947,4.7346444,6.379509,8.786444,10.612394,10.880251,11.378237,11.838497,11.940358,12.1252165,13.592768,16.244923,17.723793,18.225552,17.652113,15.62244,15.46399,17.40689,20.243906,22.582933,22.828154,21.688822,19.606333,17.425755,15.697892,14.68683,12.245941,10.631257,10.33322,10.763299,10.269085,10.155907,11.778135,11.532914,8.60913,4.991183,3.9688015,2.5125682,1.9542197,2.4182527,2.8332415,2.757789,2.282438,1.8448136,1.629774,1.5430037,1.3091009,1.1242423,1.2223305,1.4449154,1.2223305,1.6448646,1.7014539,2.625747,4.266839,5.1043615,3.5160866,2.3201644,2.335255,3.2029586,3.3689542,5.247721,7.0170827,8.726082,10.612394,13.128735,5.9418845,2.727608,2.4069347,3.7575345,5.3986263,7.069899,9.507015,10.593531,9.80128,8.175279,6.7454534,5.523123,5.5004873,6.749226,8.446907,8.273367,6.8661776,5.7607985,5.704209,6.670001,10.736891,13.468271,13.645585,11.785681,10.144588,10.159679,8.843033,9.016574,10.174769,8.45068,8.246958,9.027891,10.487898,12.50248,15.154634,14.520834,15.535669,17.746428,20.428764,22.586706,22.126446,21.326649,19.651604,17.991648,18.678267,17.874697,18.557543,19.73083,20.85507,21.854816,23.624178,25.39354,27.460938,30.245134,34.315796,35.91539,37.45462,39.242844,40.982025,41.732777,38.665634,37.15281,38.111057,40.917892,43.441776,43.08715,41.857273,40.246365,38.2431,35.349495,32.859562,31.580645,32.527573,35.134457,37.27731,37.877155,39.344707,40.37086,39.310753,34.198845,29.852781,24.888006,21.700138,20.587215,19.753464,19.097027,19.383747,19.87796,20.402355,21.345512,22.643295,24.552244,26.491373,27.974014,28.607815,27.67975,24.95214,23.431774,23.522316,23.046967,25.940569,29.430248,34.33466,39.661606,42.589165,51.72646,51.066254,42.72498,31.139246,23.065828,14.154889,11.189606,9.748463,7.9036493,6.228604,6.722818,6.6549106,6.477597,6.4021444,6.4021444,7.0284004,6.832224,6.258785,5.983383,6.9227667,11.046246,17.23335,19.76101,16.42601,8.563859,5.2590394,6.039973,6.541732,5.406172,4.2592936,3.0105548,2.5880208,3.5236318,4.647874,3.1048703,1.7693611,1.5279131,1.9579924,2.6597006,3.2482302,4.22534,5.4740787,7.066127,8.782671,10.121953,12.966512,11.830952,10.38981,10.95193,14.471789,15.905387,16.98813,18.851807,21.107838,21.854816,21.066338,25.751938,25.4954,20.526854,21.752956,18.38023,19.002712,19.229069,18.146326,18.297232,17.320122,15.686575,14.264296,13.815352,14.977322,13.6833105,12.344029,10.608622,8.75249,7.696155,6.8774953,7.3377557,6.4511886,4.134797,2.837014,2.5993385,3.2142766,3.663219,3.531177,3.0105548,2.546522,1.8636768,1.1242423,0.52062225,0.29049212,0.24899325,0.25276586,0.25276586,0.23390275,0.2263575,1.3770081,1.3543724,0.754525,0.32821837,0.95824677,0.26408374,0.40367088,1.0299267,1.3996439,0.38858038,0.13958712,0.041498873,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20372175,0.42630664,0.56212115,0.60362,0.55457586,0.98465514,1.0336993,0.6488915,0.5772116,0.56212115,0.27917424,0.056589376,0.0,0.0,0.0,0.071679875,0.14713238,0.5319401,1.931584,1.9164935,4.1762958,6.5945487,7.122716,3.7877154,4.8553686,8.235641,8.307321,4.7874613,2.7426984,2.5880208,1.8334957,1.5279131,2.282438,4.2517486,2.9049213,1.7693611,0.90920264,0.49044126,0.7432071,0.94315624,1.8787673,3.2746384,4.485651,4.485651,4.183841,4.055572,4.1989317,4.5460134,4.8327327,5.251494,4.9459114,4.7535076,4.949684,5.2288585,7.8998766,7.164215,5.6815734,4.825187,4.7006907,5.2364035,5.9418845,5.975838,5.455216,5.455216,4.5535583,4.779916,5.13077,4.961002,3.9612563,3.572676,3.561358,3.6066296,3.410453,2.704972,2.4182527,1.8448136,1.267602,0.8601585,0.663982,1.2713746,1.4109617,1.2902378,1.1619685,1.3241913,1.4034165,1.4109617,1.3241913,1.2411937,1.388326,1.3770081,1.7316349,2.1881225,2.584248,2.8785129,2.2862108,2.022127,1.9806281,2.0183544,1.9429018,2.0787163,2.1051247,2.0749438,2.1692593,2.6974268,2.6182017,2.4295704,2.4597516,2.9124665,3.874486,4.768598,5.8437963,6.94163,7.5829763,6.9567204,6.0324273,5.6287565,4.991183,4.236658,4.323428,3.6896272,3.3236825,3.0218725,2.704972,2.3993895,2.3013012,2.161714,2.0183544,1.9768555,2.203213,2.323937,2.8143783,3.2670932,3.5085413,3.6028569,3.8782585,4.0895257,4.5120597,5.1647234,5.772116,5.485397,6.3531003,6.530414,6.349328,8.345046,8.254503,7.854605,7.6584287,7.748972,7.805561,7.6923823,7.183078,6.617184,6.326692,6.628502,7.2698483,7.6093845,7.6584287,7.432071,6.937857,6.8850408,7.0472636,7.24344,7.3453007,7.2698483,7.284939,7.3792543,7.383027,7.24344,7.043491,7.2472124,7.537705,7.6622014,7.541477,7.2585306,6.33801,6.0701537,6.1078796,6.25124,6.4511886,6.6322746,6.9869013,8.254503,9.963503,10.469034,10.378491,10.231359,10.484125,11.34051,12.766563,13.313594,13.856852,14.320885,14.6151495,14.622695,14.864142,13.875714,12.883514,12.208215,11.291467,10.804798,10.144588,9.167479,7.9225125,6.6662283,5.80607,5.3080835,5.2062225,5.270357,5.0062733,4.5007415,4.38379,4.3875628,4.3007927,3.9688015,3.8367596,4.085753,4.2630663,4.236658,4.172523,4.327201,4.5120597,4.3686996,4.014073,4.074435,4.5233774,5.2099953,5.9532022,6.579458,6.952948,7.152897,6.63982,6.149379,6.1003346,6.560595,5.5985756,4.8365054,4.659192,5.0477724,5.594803,5.6098933,4.8855495,3.5085413,2.1051247,1.871222,1.5882751,1.4524606,1.5052774,1.6825907,1.7919968,2.3314822,3.270866,4.3385186,4.889322,3.904667,2.5880208,2.3616633,2.6521554,3.0256453,3.199186,3.3651814,3.5538127,4.1083884,5.093044,6.270103,6.9567204,7.4471617,7.997965,8.6732645,9.34102,9.416472,9.922004,10.797253,11.627231,11.619685,12.079946,12.113899,12.045992,11.898859,11.359374,10.054046,9.507015,9.64283,10.201178,10.740664,10.948157,11.393328,11.846043,11.910177,11.031156,11.932813,12.449662,13.102326,13.86817,14.173752,14.290704,14.143571,13.849306,13.498452,13.13628,13.490907,13.822898,14.252977,14.634012,14.547242,14.053028,14.211478,15.290449,16.807045,17.50498,17.686066,17.757746,17.172989,16.116653,15.509261,16.644821,17.738882,17.859608,17.154125,16.82968,16.177015,16.286423,17.048492,18.070873,18.663176,18.49718,18.980076,20.14959,21.4851,21.892544,3.6481283,3.3425457,3.2105038,3.682082,4.266839,3.5689032,3.3764994,2.987919,2.8898308,3.1539145,3.4481792,3.0935526,2.686109,2.565385,2.6823363,2.6106565,2.6219745,3.1199608,3.9197574,4.7421894,5.2175403,5.168496,5.3948536,5.6400743,5.873977,6.300284,7.7904706,10.057818,12.785426,15.131999,15.716756,16.033657,17.240896,17.429527,17.369165,20.50799,29.954643,26.823364,17.033401,6.5228686,1.2525115,0.8865669,0.9318384,0.7469798,0.31312788,0.21503963,0.1056335,0.18485862,0.29426476,0.35839936,0.38103512,0.38103512,0.482896,0.6149379,0.76584285,0.9620194,0.8262049,0.97710985,1.237421,1.6976813,2.686109,3.942393,5.2628117,6.4964604,7.6923823,9.110889,9.0957985,9.34102,9.884277,10.386037,10.114408,8.103599,6.628502,5.2175403,4.3347464,5.3873086,7.3151197,9.673011,11.310329,12.1252165,13.075918,15.811071,15.716756,14.079436,12.713746,13.947394,12.849561,12.1252165,12.136535,12.679792,12.985375,13.422999,14.724555,15.75071,15.697892,14.0983,12.842015,11.849815,11.057564,10.672756,11.185833,10.012547,9.601331,9.303293,9.073163,9.476834,10.819888,13.140053,12.736382,9.216523,5.492942,4.2706113,3.5387223,3.7198083,4.1762958,3.1727777,2.806833,2.2484846,1.7844516,1.5052774,1.297783,1.4562333,1.7316349,2.546522,3.361409,2.7011995,2.7125173,2.6898816,3.0746894,3.7763977,4.164978,5.594803,3.7462165,2.0485353,1.9768555,3.0520537,5.028909,7.77538,10.223814,11.785681,12.359119,5.534441,2.546522,3.4142256,5.983383,5.934339,5.7909794,6.1116524,6.7944975,8.00551,10.178542,9.578695,6.417235,4.3611546,4.395108,4.821415,4.285702,5.028909,7.1906233,9.759781,10.589758,13.932304,15.977067,16.565596,16.87118,19.425245,15.297995,12.408164,12.064855,12.857106,10.63503,9.461743,10.084227,10.884023,11.714001,13.8870325,15.99593,15.784663,16.316603,18.131235,19.240387,18.983849,19.1423,18.402864,17.493662,19.164934,18.323639,19.017803,19.97605,20.783392,21.881226,24.224026,25.891525,28.479546,31.946589,34.60629,34.11962,36.311516,38.69959,40.52554,42.77025,40.91412,38.9599,39.80874,43.611546,47.776524,49.081852,48.134922,45.320545,41.468693,37.8432,34.459156,32.50871,32.38044,33.91967,36.42092,35.56831,34.97978,35.534355,37.06604,38.36005,32.855793,27.166672,23.065828,21.31533,21.681276,20.545715,21.051247,21.854816,22.733839,24.567333,25.397312,25.842482,26.306515,26.872408,27.313805,25.408628,21.839725,21.35683,23.646814,23.314823,26.121656,30.980797,36.756687,41.2612,41.2612,48.36505,49.372345,43.268234,32.7577,24.261751,14.766054,10.201178,8.29223,7.54525,7.277394,6.779407,6.828451,6.790725,6.2323766,4.9119577,4.927048,4.919503,4.779916,4.6629643,5.0062733,6.1908774,10.853842,14.234114,13.287186,6.6850915,4.67051,5.1269975,5.3458095,4.3196554,2.746471,2.11267,2.2560298,4.847823,7.8017883,5.2628117,2.8332415,2.2899833,2.7879698,3.6179473,4.22534,4.323428,4.568649,5.342037,7.375482,11.732863,10.868933,11.457462,11.400873,10.834979,12.113899,17.682293,18.395319,19.236614,21.09652,20.768301,21.65864,20.341993,18.0671,16.380737,17.150352,14.894323,14.181297,13.924759,13.758763,14.037937,13.585222,13.226823,13.106099,13.513543,14.894323,13.000465,11.812089,10.751981,9.540969,8.209232,7.0510364,6.485142,5.2099953,3.2859564,2.1503963,2.1994405,2.8332415,3.3840446,3.4896781,3.097325,2.9615107,2.516341,1.7165444,0.7922512,0.23013012,0.422534,0.573439,0.6413463,0.69039035,0.8865669,0.44516975,0.34330887,0.55080324,1.6410918,4.7912335,1.2751472,0.5696664,0.44894236,0.13204187,0.29049212,0.071679875,0.071679875,0.06413463,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.150905,0.482896,0.8865669,0.59230214,0.27917424,0.15845025,0.28294688,0.56589377,0.49044126,0.21503963,0.026408374,0.0,0.0,0.0,0.0,0.0,0.08677038,0.44139713,1.9693103,4.2630663,7.4735703,9.7069645,7.032173,4.617693,11.2650585,13.739901,8.786444,3.097325,2.425798,1.991946,1.3996439,1.237421,3.0671442,2.2975287,1.7580433,1.086516,0.3772625,0.18485862,0.40367088,1.2826926,2.4786146,3.6556737,4.485651,5.4250345,5.119452,4.9685473,5.2364035,5.0666356,4.6629643,4.5988297,4.6252384,4.6554193,4.776143,6.0701537,6.349328,6.25124,6.25124,6.651138,5.6287565,5.040227,4.847823,4.768598,4.3196554,4.561104,5.0062733,5.1534057,4.7308717,3.6934,3.5085413,3.3727267,3.2557755,3.059599,2.595566,1.9957186,1.3807807,0.995973,0.87147635,0.80734175,1.4562333,1.5165952,1.3317367,1.1657411,1.1883769,1.3958713,1.3128735,1.237421,1.327964,1.5731846,1.6071383,1.9844007,2.4031622,2.6823363,2.7313805,2.3654358,1.9089483,1.6335466,1.5882751,1.6033657,2.0296721,2.282438,2.4220252,2.5880208,2.9916916,2.5012503,2.1503963,2.2258487,2.7011995,3.2520027,5.142088,5.9532022,6.6134114,7.2472124,7.1868505,4.9157305,4.13857,4.3347464,4.847823,4.8968673,3.6783094,3.2067313,2.9501927,2.6672459,2.4107075,2.5087957,2.505023,2.5729303,2.8747404,3.5689032,3.7273536,3.9989824,4.285702,4.4705606,4.4101987,4.274384,4.4630156,5.3910813,6.700182,7.2472124,6.700182,7.164215,7.5263867,7.7829256,9.061845,8.231868,7.8244243,7.7338815,7.7338815,7.4773426,7.9791017,7.8923316,7.537705,7.115171,6.7152724,7.273621,7.7716074,7.997965,7.914967,7.6584287,7.7338815,8.080963,8.280911,8.22055,8.088508,7.281166,6.511551,6.1342883,6.2625575,6.7756343,7.1038527,7.3981175,7.496206,7.333983,6.94163,5.9532022,5.587258,5.8702044,6.6360474,7.537705,7.4169807,7.4018903,8.258276,9.752235,10.665211,10.069136,9.910686,10.238904,11.16697,12.864652,14.094527,14.634012,14.588741,14.252977,14.083209,14.607604,14.124708,13.449409,12.755245,11.59705,10.582213,9.763554,9.092027,8.409182,7.4471617,7.152897,6.6586833,6.3719635,6.0286546,4.7006907,4.466788,4.2102494,4.085753,4.0782075,3.9688015,4.1498876,4.2064767,4.0480266,3.7801702,3.7084904,3.8895764,3.9084394,4.014073,4.304565,4.745962,4.9421387,5.485397,5.9192486,6.1229706,6.3153744,6.439871,6.398372,6.5002327,6.719045,6.6850915,5.2779026,4.52715,4.689373,5.3609,5.4476705,5.5193505,4.3309736,2.7313805,1.5656394,1.6637276,1.5769572,1.50905,1.5354583,1.8033148,2.546522,3.3538637,4.425289,4.870459,4.3347464,2.9916916,2.0145817,2.2560298,2.8521044,3.3463185,3.663219,4.1008434,4.6516466,5.138315,5.7570257,7.066127,7.7112455,8.039464,8.601585,9.367428,9.718282,9.416472,9.752235,10.419991,11.083972,11.351829,11.351829,11.672502,11.812089,11.480098,10.589758,9.869187,9.295748,9.06939,9.386291,10.438853,9.899368,10.133271,10.680302,11.155652,11.216014,12.936331,13.321139,13.290957,13.4644985,14.158662,13.830443,13.264549,12.623203,12.174261,12.283667,12.626976,13.460726,14.079436,14.2077055,14.022847,13.902123,14.237886,15.486626,17.237123,18.187824,18.263277,17.904879,17.225805,16.644821,16.874952,17.976559,18.663176,18.361366,17.244669,16.218515,16.124199,16.912678,18.119919,19.323385,20.142044,19.21398,19.512016,20.458946,21.488873,22.062311,2.9766011,2.7879698,2.6483827,2.7804246,3.0445085,2.9351022,2.9652832,2.7087448,2.5767028,2.6068838,2.4597516,2.505023,2.2711203,2.203213,2.354118,2.3767538,2.4861598,2.7728794,3.6066296,4.772371,5.462761,4.9949555,4.983638,5.2552667,5.726845,6.398372,6.7152724,8.265821,10.212496,11.996947,13.336229,14.562332,15.746937,16.920223,18.71222,22.326395,24.012758,18.79899,11.000975,4.2064767,1.2864652,1.0978339,1.0487897,0.90543,0.6149379,0.31312788,0.58098423,0.7884786,0.7130261,0.5093044,0.7092535,1.1016065,1.2864652,1.3845534,1.3996439,1.1921495,1.0412445,1.0223814,1.2298758,1.7769064,2.795515,4.217795,5.485397,6.5040054,7.1604424,7.3151197,6.94163,7.220804,7.6395655,7.7716074,7.2472124,5.8588867,5.9117036,6.5756855,7.383027,8.216777,8.329956,8.311093,7.8696957,7.352846,7.7187905,8.654402,9.650374,9.582467,8.643084,8.329956,7.8961043,8.503497,9.25425,9.556059,9.14107,9.14107,9.2995205,9.424017,9.635284,10.340765,12.061082,11.306557,9.884277,9.009028,9.318384,8.563859,7.605612,7.2623034,7.9262853,9.548513,10.208723,10.661438,10.585986,9.337247,5.956975,4.063117,3.6254926,3.4972234,3.4859054,4.3686996,3.338773,2.425798,2.0636258,2.1353056,1.9579924,1.5769572,1.2525115,1.297783,1.6825907,2.0296721,2.704972,2.987919,2.7200627,2.2786655,2.5427492,3.1010978,2.7125173,2.8785129,4.1272516,5.994701,7.6886096,8.137552,9.507015,11.231105,10.0276375,5.451443,3.3010468,3.8367596,5.523123,5.0439997,5.062863,6.692637,7.699928,7.779153,8.567632,7.020855,5.2175403,3.85185,3.3010468,3.6481283,4.1008434,4.606375,6.326692,9.092027,11.393328,12.261031,13.917213,15.954432,16.965494,14.566105,12.774108,11.551778,11.59705,12.151625,11.012292,11.608367,11.54046,11.864905,12.81938,13.800262,16.01102,16.588232,17.818108,19.70442,19.987368,18.87067,18.006739,17.614386,17.4333,16.712729,16.739138,19.006485,20.1345,19.33093,18.391546,21.952906,25.355812,29.109575,32.82561,35.191048,35.09673,37.590435,40.97448,44.098213,46.384426,43.74736,41.955364,42.374123,44.607517,46.49383,51.843414,53.473186,51.59819,47.074814,41.41965,36.424694,33.62918,32.935017,33.897038,35.726757,34.73456,33.738586,34.236572,35.707897,35.624897,31.448603,28.290915,25.012505,22.167944,21.986858,21.183289,20.730574,22.035902,24.842735,27.238352,27.355305,27.491117,27.702385,28.32487,29.973505,27.649569,24.148573,23.522316,25.03514,23.182781,24.503199,31.37315,37.95638,39.75215,33.568817,39.589928,45.109276,42.792885,32.70866,22.307531,14.2944765,9.480607,6.771862,5.572167,5.802297,5.613666,6.2814207,7.2170315,7.4811153,5.7909794,5.2288585,5.481624,5.451443,5.511805,7.496206,6.94163,10.084227,13.257004,13.381501,7.9753294,5.904158,6.0701537,6.25124,5.3873086,3.5764484,2.3163917,2.0183544,3.2859564,5.191132,5.2892203,4.217795,3.640583,4.0178456,4.930821,5.093044,5.2099953,4.991183,6.3455553,9.684328,13.905896,11.046246,10.77839,11.321648,11.879996,12.653384,16.22606,17.565342,19.647831,22.401848,22.70743,22.926243,21.888771,19.708193,17.320122,16.467508,14.335975,14.211478,13.5663595,12.223305,12.377983,12.249713,12.868423,13.211733,13.091009,13.170234,12.208215,11.514051,10.759526,9.695646,8.160188,7.0887623,6.0022464,4.6554193,3.259548,2.505023,2.2711203,2.535204,2.8822856,3.0709167,3.0105548,2.8181508,2.4672968,1.8221779,0.9922004,0.362172,0.38103512,0.39989826,0.41498876,0.6526641,1.5807298,2.4484336,2.6106565,2.6408374,2.686109,2.4371157,1.2147852,1.6675003,1.4750963,0.3470815,0.056589376,0.0150905,0.07922512,0.094315626,0.030181,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.1659955,0.5319401,0.422534,0.7884786,0.80356914,0.422534,0.38103512,0.55080324,0.38103512,0.150905,0.011317875,0.0,0.0,0.0,0.0,0.08299775,0.4074435,1.3958713,4.508287,9.016574,11.52537,5.9607477,4.4894238,10.970794,14.332202,10.725573,3.5123138,3.0671442,2.2862108,1.5165952,1.1996948,1.8599042,2.1051247,2.2447119,1.8561316,0.9997456,0.21881226,0.2263575,0.6451189,1.5203679,2.6446102,3.5839937,4.8930945,4.719554,4.447925,4.6629643,5.1269975,5.20245,4.3800178,4.3385186,5.0968165,4.983638,5.798525,5.9117036,6.2323766,6.6586833,6.115425,4.9723196,4.7006907,4.7120085,4.7044635,4.67051,4.7610526,5.160951,5.349582,4.9044123,3.4972234,3.169005,3.127506,2.9766011,2.6823363,2.5691576,2.0108092,1.5430037,1.1732863,0.9620194,1.0299267,1.2751472,1.3619176,1.2789198,1.1695137,1.3015556,1.478869,1.4222796,1.3091009,1.3015556,1.5467763,1.5354583,1.7089992,2.0296721,2.4371157,2.8181508,2.8407867,2.4522061,1.9579924,1.6033657,1.5656394,1.991946,1.9089483,1.961765,2.3277097,2.7238352,2.3013012,2.0787163,2.2107582,2.6219745,3.006782,5.1534057,5.8211603,6.149379,6.519096,6.5643673,5.59103,5.1458607,5.149633,5.2552667,4.8365054,3.802806,3.3576362,3.218049,3.229367,3.361409,3.3538637,3.1312788,2.9200118,2.886058,3.1425967,3.9461658,4.191386,4.402653,4.738417,5.0213637,5.402399,5.8513412,6.79827,7.745199,7.2472124,7.5188417,8.541223,8.967529,8.669493,8.771353,8.967529,8.907167,8.469543,7.6810646,6.730363,7.575431,8.035691,8.031919,7.6622014,7.201941,7.3453007,7.54525,7.888559,8.439363,9.258021,9.967276,9.654147,9.118435,8.75249,8.537451,7.4207535,6.7869525,6.8661776,7.3679366,7.4697976,7.4773426,7.5716586,7.586749,7.4811153,7.333983,6.4021444,6.3719635,6.94163,7.707473,8.160188,7.7150183,7.7187905,8.333729,9.246704,9.654147,9.318384,9.714509,10.612394,11.966766,13.936077,14.758509,14.558559,13.815352,13.249459,13.792717,14.483108,14.743419,14.3095665,13.200415,11.717773,11.019837,10.801025,10.408672,9.7296,9.216523,9.050528,8.492179,7.8206515,6.971811,5.553304,4.425289,4.1612053,4.266839,4.425289,4.4931965,4.587512,4.5309224,4.304565,3.9688015,3.6707642,3.5990841,3.7160356,3.9159849,4.187614,4.5988297,4.727099,5.070408,5.413717,5.7192993,6.1078796,6.485142,6.3832817,6.096562,5.798525,5.534441,5.4778514,5.406172,5.2854476,4.930821,4.0178456,3.5764484,3.0822346,2.4295704,1.8561316,1.9429018,1.4373702,1.4071891,1.7655885,2.4069347,3.169005,3.9650288,4.6554193,4.3724723,3.199186,2.161714,1.9768555,2.6332922,3.2331395,3.4142256,3.3689542,4.3649273,5.0553174,5.4363527,5.8588867,7.0284004,8.201687,8.514814,8.677037,9.031664,9.559832,9.469289,9.076936,9.548513,10.804798,11.521597,11.348056,11.815862,12.570387,13.143826,12.958967,11.193378,9.880505,8.918486,8.492179,9.0957985,10.140816,10.876478,11.502733,12.030901,12.276122,12.698656,12.804289,12.808062,12.811834,12.792972,12.434572,12.306303,11.996947,11.619685,11.808316,12.15917,12.955194,13.671993,14.015302,13.902123,14.2944765,15.531898,16.995676,18.206688,18.787672,18.52736,18.085964,17.674747,17.63325,18.451908,18.504726,17.795471,16.708956,15.735619,15.46399,16.195879,17.25976,18.58395,19.806282,20.251451,19.94964,20.689075,21.915178,22.790428,22.224533,2.5804756,2.4182527,2.3126192,2.5087957,2.9464202,3.2633207,3.6858547,3.2670932,2.71629,2.3390274,2.0485353,2.1277604,2.0749438,2.0673985,2.142851,2.191895,2.5087957,2.837014,3.5990841,4.6290107,5.1835866,4.9685473,5.0439997,5.1835866,5.4250345,6.085244,6.1078796,7.798016,9.42779,10.536942,11.917723,14.366156,16.0412,18.304777,21.217243,23.522316,18.372684,11.951676,6.439871,2.8822856,1.1883769,0.754525,0.79602385,0.8978847,0.8337501,0.573439,0.98465514,1.0412445,0.935611,0.9318384,1.3430545,2.2183034,2.6483827,2.757789,2.546522,1.8825399,1.4977322,1.3920987,1.9089483,3.1237335,4.881777,5.9230213,6.168242,6.571913,7.375482,8.137552,8.420499,8.088508,7.9036493,7.8131065,6.94163,7.073672,7.835742,8.050782,7.5037513,6.930312,6.8246784,6.217286,5.66271,5.4401255,5.534441,5.9796104,6.900131,7.352846,7.3981175,8.118689,8.971302,10.287949,10.816116,10.310584,9.540969,8.9788475,8.280911,7.594294,7.2623034,7.835742,9.420244,9.042982,8.544995,8.684583,9.125979,9.107117,8.59404,8.469543,9.352338,11.581959,11.45369,11.25374,10.642575,9.333474,7.062354,4.4630156,3.7688525,3.3274553,2.8634224,3.4330888,3.0558262,2.505023,2.1315331,1.9655377,1.7014539,1.237421,1.1657411,1.2638294,1.3732355,1.3958713,2.1353056,2.4220252,2.082489,1.4901869,1.5580941,1.8297231,2.7087448,4.2894745,6.1418333,7.322665,8.390318,8.065872,8.612903,9.35611,6.688864,4.327201,3.1048703,3.2557755,3.9122121,3.138824,4.164978,5.7796617,6.828451,7.220804,7.960239,7.277394,5.828706,4.123479,2.7992878,2.6144292,2.7313805,3.2520027,4.7912335,7.2887115,9.97482,9.81637,10.212496,11.819634,13.373956,11.714001,11.223559,10.646348,10.767072,11.359374,11.18206,12.879742,13.192869,13.604086,14.634012,15.875206,17.040947,17.463482,18.319866,19.553514,19.870417,19.308294,18.221779,17.297485,16.761772,16.373192,16.939087,18.334957,18.519815,17.870924,19.202662,21.564325,24.431519,28.456911,32.919926,35.753166,36.541645,40.01623,44.59997,48.97622,52.08486,47.85952,44.464157,42.174175,41.457375,42.951336,46.829594,52.05468,54.706837,52.722435,45.89021,39.001396,35.821075,33.75745,32.47098,33.866856,35.334404,34.11585,33.176464,33.512226,34.14603,32.38044,30.116865,26.725275,23.22428,22.29244,21.881226,21.666185,23.216734,26.208426,28.404093,29.094484,30.429993,31.146791,32.29367,37.22072,34.515747,29.094484,25.989614,25.374676,22.560297,23.571362,29.705648,33.938534,32.603024,25.374676,32.46721,37.616844,37.541393,31.5731,21.700138,14.464244,9.582467,6.436098,4.927048,5.485397,5.172269,6.3832817,7.8696957,8.4544525,7.0359454,6.255012,6.1531515,5.9796104,5.8890676,6.964266,6.519096,9.718282,12.593022,12.543978,8.356364,6.255012,6.270103,6.3644185,5.6287565,4.29702,3.2746384,2.2975287,2.3654358,3.4444065,4.432834,4.5799665,4.1800685,4.0782075,4.3913355,4.504514,4.6856003,4.708236,6.477597,9.635284,11.574413,10.099318,9.869187,11.031156,13.29473,15.916705,18.304777,20.477808,23.537407,26.408375,25.838709,25.982069,23.98635,21.949133,20.240133,17.50498,15.143317,14.04171,12.811834,11.529142,11.725319,11.604594,12.581704,13.347548,13.479589,13.445636,12.427027,12.042219,11.18206,9.559832,7.707473,6.6813188,5.983383,4.825187,3.3953626,2.8596497,2.5314314,2.4220252,2.5540671,3.2255943,5.0213637,3.1954134,2.3767538,1.7919968,1.177059,0.76207024,0.63002837,0.47535074,0.32444575,0.3169005,0.70170826,1.1959221,1.3128735,1.3128735,1.2223305,0.8111144,0.633801,1.0336993,3.0181,4.4403796,0.00754525,0.06790725,0.0754525,0.05281675,0.0150905,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21503963,0.4376245,0.5885295,0.7092535,0.5093044,0.7922512,0.80356914,0.47912338,0.44516975,0.56589377,0.44139713,0.26408374,0.120724,0.0,0.0,0.0,0.0150905,0.060362,0.15845025,0.6526641,4.398881,8.986393,10.79348,4.961002,4.0178456,9.680555,12.200669,8.8769865,4.0480266,3.3689542,2.5238862,1.7919968,1.418507,1.629774,1.8070874,2.0787163,2.4559789,2.3314822,0.45648763,0.21881226,0.41498876,1.0072908,1.8599042,2.7087448,4.617693,4.8025517,4.3913355,4.1574326,4.538468,4.821415,4.4818783,4.7308717,5.492942,5.409944,5.6363015,5.934339,6.375736,6.692637,6.2851934,4.659192,4.5950575,4.8327327,4.8100967,4.6327834,5.3910813,5.7796617,5.624984,4.7648253,3.0633714,2.6898816,2.9011486,2.9124665,2.5729303,2.3805263,1.9542197,1.6222287,1.2826926,0.9922004,0.965792,1.1619685,1.1619685,1.0601076,1.0148361,1.2449663,1.2562841,1.1996948,1.1581959,1.1921495,1.3505998,1.5354583,1.7052265,1.9164935,2.214531,2.625747,2.3013012,2.0372176,1.8599042,1.7995421,1.9051756,2.0108092,1.7316349,1.720317,2.0787163,2.3805263,2.071171,2.0145817,2.233394,2.6408374,3.0181,4.538468,5.3080835,5.723072,5.945657,5.9230213,5.7306175,5.832478,5.8098426,5.5080323,5.0138187,3.863168,3.4594972,3.4444065,3.5462675,3.610402,3.5424948,3.4670424,3.3048196,3.1350515,3.1539145,3.9574835,4.353609,4.8666863,5.485397,5.6287565,6.085244,6.7077274,7.3000293,7.413208,6.379509,7.1679873,8.756263,9.759781,9.797507,9.484379,9.7296,10.061591,9.6201935,8.311093,6.7831798,6.9567204,7.7716074,8.356364,8.382772,8.084735,8.318638,8.541223,8.884532,9.446653,10.299266,10.902886,10.469034,9.756008,9.216523,9.001483,8.118689,7.575431,7.6584287,8.107371,8.084735,8.122461,8.239413,8.16396,7.9300575,7.8810134,7.4018903,7.413208,7.8017883,8.258276,8.269594,8.024373,8.171506,8.465771,8.865668,9.5183325,9.725827,10.284176,11.216014,12.50248,14.079436,14.7170105,14.27184,13.404137,12.940104,13.8719425,14.569878,15.098045,14.769827,13.528633,11.951676,11.102836,10.797253,10.801025,10.801025,10.419991,9.473062,9.020347,8.394091,7.2057137,5.3458095,4.093298,3.9310753,4.134797,4.3875628,4.768598,4.7044635,4.515832,4.236658,3.8858037,3.440634,3.380272,3.5802212,3.8254418,4.08198,4.4630156,4.534695,4.7535076,5.0666356,5.5004873,6.156924,6.1229706,5.9003854,5.73439,5.6098933,5.240176,5.50426,5.670255,5.3344917,4.4177437,3.187868,3.1539145,2.916239,2.5616124,2.2183034,2.0673985,1.6033657,1.7316349,2.3088465,3.0671442,3.610402,4.617693,4.6554193,3.7801702,2.5201135,1.9089483,2.0296721,2.704972,3.2670932,3.4896781,3.5990841,4.353609,4.9534564,5.1156793,5.2099953,6.258785,7.413208,8.307321,8.461998,8.209232,8.68081,9.148616,8.922258,9.7296,11.348056,11.631002,11.570641,12.845788,14.268067,14.928277,14.188843,11.144334,9.661693,8.827943,8.469543,9.133525,10.559577,11.555551,12.513797,13.249459,12.992921,12.774108,12.6345215,12.6345215,12.608112,12.193124,11.212241,11.068882,11.344283,11.785681,12.30253,12.487389,13.196642,13.781399,14.030393,14.181297,14.815099,16.614641,18.5085,19.813826,20.243906,18.738628,18.304777,18.546225,18.995167,19.1008,17.957695,16.542961,15.414946,14.973549,15.475307,16.592005,18.002966,19.051756,19.58747,19.97605,19.462973,20.108091,21.432283,22.60557,22.454664,2.1956677,2.2220762,2.1994405,2.4559789,2.987919,3.4934506,4.3422914,3.904667,3.1199608,2.4786146,2.022127,1.931584,1.9579924,1.9957186,2.0372176,2.1805773,2.6898816,2.938875,3.4934506,4.274384,4.5497856,4.6290107,4.7874613,4.817642,4.8968673,5.5985756,5.9494295,8.096053,10.016319,11.23865,12.830698,16.233604,17.603067,19.225298,21.300241,21.937815,14.04171,7.6886096,3.7952607,2.082489,1.0714256,0.56212115,0.7130261,0.8865669,0.83752275,0.694163,1.0223814,1.0412445,1.1204696,1.4109617,1.8485862,3.0030096,3.682082,3.7801702,3.3840446,2.7426984,2.3616633,2.5125682,3.308592,4.851596,7.224577,8.016829,8.443134,8.990166,9.759781,10.469034,11.223559,9.986138,9.073163,9.088254,8.952439,10.416218,10.231359,8.869441,7.1679873,6.319147,5.9305663,5.2854476,4.825187,4.98741,6.2021956,6.888813,7.462252,8.152642,9.261794,11.144334,11.853588,12.193124,11.861133,10.899114,9.684328,8.069645,7.0359454,6.4134626,6.066381,5.9003854,6.628502,6.628502,6.7756343,7.3981175,8.296002,9.001483,9.310839,9.710737,10.61994,12.404391,11.721546,10.665211,9.107117,7.586749,7.3415284,5.168496,3.8556228,2.9954643,2.41448,2.1994405,2.214531,2.0787163,1.8561316,1.5920477,1.3204187,1.3920987,1.6825907,1.7995421,1.6561824,1.4864142,1.8448136,1.9806281,1.7052265,1.2600567,1.3166461,1.7354075,3.3048196,5.5382137,7.586749,8.239413,8.941121,8.307321,7.7716074,7.0284004,4.0593443,3.169005,2.7615614,2.8181508,3.0369632,2.806833,4.244203,5.783434,6.749226,7.250985,8.175279,8.473316,7.092535,5.2062225,3.572676,2.5238862,2.5087957,2.848332,3.8254418,5.406172,7.2283497,7.213259,7.5075235,9.050528,10.884023,10.148361,11.623458,12.932558,13.532406,13.50977,13.58145,15.939341,16.652367,16.45619,16.033657,16.0412,16.580687,16.882498,17.882242,19.421474,20.258997,19.719511,18.365139,17.18808,16.852316,17.716248,17.972786,18.161417,17.874697,17.874697,20.066593,21.326649,24.193844,28.166418,32.42194,35.817303,38.41287,42.898518,47.45962,51.002117,53.14497,48.440506,44.347206,41.242336,39.778557,40.910347,42.70989,47.678436,52.333855,53.83913,49.9986,43.59268,39.804966,35.217453,30.509218,30.448856,33.62541,33.45941,32.47098,32.188038,33.165146,33.293415,31.74664,28.702131,25.159636,22.92247,23.41291,23.424229,24.540926,26.793182,28.634224,30.154593,33.051968,34.821327,36.70764,43.736042,38.914627,32.07863,27.03463,24.601288,22.598024,25.22377,28.709677,28.422956,23.85808,18.632996,29.411385,33.059513,32.946335,30.05273,22.975286,15.697892,10.56335,7.0774446,5.2552667,5.6098933,5.4250345,7.1302614,8.68081,9.06939,8.311093,7.805561,7.5112963,7.8961043,8.643084,8.677037,7.0812173,9.2995205,11.355601,11.1631975,8.544995,6.398372,6.255012,6.356873,5.8702044,4.8968673,4.432834,2.9313297,2.1315331,2.584248,3.6481283,4.3800178,4.168751,3.7348988,3.4972234,3.5651307,3.7650797,4.187614,6.205968,8.7751255,8.443134,9.118435,9.371201,10.789707,13.777626,17.565342,20.75321,24.242887,27.85329,30.362085,29.494383,28.619133,25.706667,23.409138,21.77559,18.26705,15.905387,13.864397,12.079946,10.978339,11.476325,11.925267,12.513797,12.785426,12.792972,13.106099,12.574159,12.449662,11.6008215,9.80128,7.7150183,6.560595,6.8774953,5.8966126,3.6783094,3.108643,2.7011995,2.425798,2.4559789,3.150142,5.0854983,3.3350005,2.5201135,2.093807,1.7731338,1.539231,1.1393328,0.7432071,0.72811663,0.83752275,0.15845025,0.15467763,0.14713238,0.15845025,0.1659955,0.09808825,0.15845025,0.39989826,2.6182017,4.5837393,0.033953626,0.41121614,0.52439487,0.32067314,0.003772625,0.011317875,0.003772625,0.060362,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21503963,0.4376245,0.55457586,0.5319401,0.5998474,0.7205714,0.80734175,0.80356914,0.67152727,0.5093044,0.40367088,0.28294688,0.13204187,0.00754525,0.0,0.0,0.0150905,0.060362,0.15845025,0.73188925,3.5349495,6.881268,8.201687,4.063117,3.6292653,7.586749,8.5563135,5.6325293,4.395108,3.4066803,2.727608,2.1654868,1.7919968,1.9391292,1.8523588,1.9278114,2.6031113,2.9011486,0.43385187,0.18485862,0.35085413,0.8262049,1.5052774,2.2786655,4.0782075,4.515832,4.1310244,3.5877664,3.6971724,3.9348478,4.1536603,4.5535583,5.13077,5.666483,5.674028,5.73439,6.1003346,6.6134114,6.700182,5.1458607,4.8327327,4.908185,4.8855495,4.6214657,6.0248823,6.428553,5.9192486,4.640329,2.795515,2.5767028,2.848332,2.8521044,2.474842,2.2447119,1.8863125,1.6825907,1.3732355,0.9997456,0.8903395,1.0751982,0.9620194,0.845068,0.8941121,1.1431054,1.0827434,1.0223814,1.0902886,1.2449663,1.2638294,1.4222796,1.659955,1.8372684,1.9240388,2.0372176,1.7089992,1.5807298,1.7089992,1.9957186,2.203213,2.022127,1.6260014,1.5618668,1.8749946,2.123988,2.0258996,2.0636258,2.2220762,2.5427492,3.1463692,4.13857,4.817642,5.2665844,5.5268955,5.594803,5.6287565,5.7607985,5.8136153,5.6891184,5.3684454,4.3121104,3.9574835,3.8443048,3.7952607,3.9197574,3.8858037,3.640583,3.31991,3.1048703,3.2331395,3.8141239,4.4101987,5.1043615,5.7607985,6.039973,6.417235,7.1906233,7.5037513,7.2094865,6.8963585,7.8244243,9.26934,10.291721,10.480352,9.967276,9.831461,10.121953,9.876732,8.918486,7.877241,7.586749,8.16396,8.850578,9.22784,9.250477,9.590013,9.869187,10.186088,10.540714,10.801025,11.027383,10.589758,9.971047,9.548513,9.590013,9.092027,8.59404,8.514814,8.7751255,8.797762,8.820397,8.975075,8.98262,8.771353,8.477088,8.213005,8.14887,8.360137,8.643084,8.537451,8.43559,8.771353,9.024119,9.2844305,10.257768,10.7218,11.197151,12.0082655,13.041965,13.754991,13.973803,13.547497,13.068373,13.041965,13.898351,14.388792,14.679284,14.219024,13.0646,11.853588,10.982111,10.453944,10.393582,10.536942,10.223814,9.242931,8.790216,7.9828744,6.5455046,4.8138695,3.9574835,3.832987,3.9763467,4.191386,4.5309224,4.4894238,4.3196554,4.0782075,3.772625,3.350091,3.4255435,3.6254926,3.8669407,4.134797,4.466788,4.6327834,4.9421387,5.2779026,5.643847,6.1531515,5.783434,5.43258,5.372218,5.4967146,5.311856,5.4778514,5.50426,4.957229,3.9273026,3.0218725,3.0030096,2.8445592,2.6408374,2.4522061,2.293756,2.142851,2.3692086,2.9237845,3.6443558,4.244203,4.5422406,3.9989824,2.9728284,1.9994912,1.8221779,2.2069857,2.474842,2.897376,3.4444065,3.7763977,4.1498876,4.504514,4.5497856,4.5988297,5.5570765,6.63982,8.00551,8.492179,8.254503,8.7600355,9.473062,9.454198,10.216269,11.45369,11.050018,11.725319,13.671993,15.286676,15.531898,13.947394,10.7557535,9.333474,8.643084,8.420499,9.208978,10.272858,11.714001,13.200415,14.045483,13.185325,12.513797,12.276122,12.355347,12.400619,11.853588,10.567122,10.035183,10.352083,11.404645,12.826925,13.3626375,14.007756,14.234114,14.166207,14.558559,15.667711,17.437073,19.364883,20.836208,21.107838,19.685556,19.440336,19.681786,19.678013,18.644312,17.112627,15.520579,14.5132885,14.509516,15.70921,17.255987,18.780127,19.478064,19.48938,19.859098,19.006485,19.296976,20.489126,21.949133,22.654613,1.8787673,2.2069857,2.3805263,2.5993385,2.9237845,3.2859564,4.2592936,3.9914372,3.361409,2.8219235,2.372981,2.0673985,2.052308,2.161714,2.3201644,2.5276587,2.9766011,3.0105548,3.2935016,3.821669,3.942393,4.115934,4.2291126,4.2404304,4.395108,5.2137675,6.017337,8.296002,10.646348,12.562841,14.449154,17.852062,17.972786,17.448391,17.21826,16.524097,10.26154,5.5306683,2.795515,1.7165444,1.1280149,0.8865669,1.1695137,1.20724,0.87902164,0.724344,0.80734175,0.90920264,1.2789198,1.9240388,2.6295197,4.323428,5.1647234,5.040227,4.285702,3.6896272,3.6368105,4.5120597,5.802297,7.356619,9.390063,10.106862,11.672502,12.872196,12.996693,11.830952,12.057309,10.18986,8.8618965,9.103344,10.344538,12.1101265,10.70671,8.635539,7.3905725,7.4811153,6.40969,5.7306175,5.111907,5.240176,7.8244243,8.756263,9.205205,9.7069645,10.834979,13.204187,12.359119,10.985884,10.125726,9.661693,8.326183,6.017337,5.3684454,5.7004366,6.1078796,5.485397,5.670255,5.9230213,5.881522,5.8437963,6.7567716,7.6886096,8.612903,9.491924,10.212496,10.604849,9.7069645,7.9413757,5.87775,4.587512,5.6476197,5.032682,3.6896272,2.7087448,2.2560298,1.5882751,1.3317367,1.4071891,1.4298248,1.2864652,1.1242423,1.841041,2.4710693,2.3993895,1.8900851,2.0560806,1.9844007,2.0560806,1.9391292,1.7278622,1.9504471,2.6446102,4.4177437,6.439871,8.065872,8.83926,9.922004,8.956212,7.118943,5.081726,3.0105548,2.6483827,2.969056,3.199186,3.4745877,4.8629136,5.2250857,6.7643166,7.5716586,7.586749,8.60913,8.929804,8.122461,6.8435416,5.3684454,3.5802212,3.7462165,3.7537618,3.942393,4.4101987,5.0213637,5.553304,6.6850915,8.503497,10.140816,9.80128,12.789199,16.90136,18.938578,18.376457,17.354074,18.531134,19.451654,19.11589,17.38803,14.996184,15.961976,16.056292,16.859861,18.693357,20.606077,19.57615,17.693611,16.667458,17.23335,19.119663,18.780127,18.063328,18.191597,19.383747,20.836208,22.341486,25.887753,29.117119,31.750412,35.587173,40.321815,45.478996,49.002625,50.191,49.72697,46.391968,43.498367,42.019497,41.887455,42.042133,42.381668,43.479504,46.6221,50.771988,52.59794,49.504387,44.656563,37.315033,29.754694,27.257215,29.630198,31.010977,31.354286,31.327879,32.316307,33.32737,33.195328,31.350513,28.117374,24.699375,25.68403,25.555761,26.080156,27.687294,29.479292,31.131702,34.75342,37.488575,39.763466,45.320545,39.39375,33.451866,27.947605,24.141027,24.103302,28.434275,27.989105,22.782883,15.875206,13.355092,27.800474,31.686277,31.339195,29.467974,25.167181,18.09351,12.223305,8.213005,6.187105,5.7079816,6.0286546,8.107371,9.205205,8.873214,8.98262,8.518587,8.590267,10.269085,12.570387,12.46098,9.476834,9.65792,10.253995,10.042727,9.363655,7.0887623,6.651138,6.670001,6.349328,5.458988,5.560849,3.7952607,2.4710693,2.516341,3.482133,4.3422914,4.1008434,3.482133,2.9916916,2.9049213,3.138824,3.9763467,5.8437963,7.6093845,6.5568223,9.148616,9.899368,10.831206,13.045737,16.697638,21.643549,26.521553,30.445084,32.618114,32.346485,30.203636,27.008223,24.008986,21.296469,17.833199,15.490398,13.29473,11.351829,10.295494,11.299012,12.438345,12.245941,11.378237,10.718028,11.363147,12.147853,12.4307995,12.132762,11.00852,8.677037,7.2094865,7.8998766,6.8737226,4.172523,3.742444,2.867195,2.493705,2.474842,2.686109,3.0331905,3.0445085,2.7917426,2.584248,2.4484336,2.1654868,1.5882751,1.7844516,2.0485353,1.7995421,0.5583485,0.5319401,0.392353,0.3169005,0.29049212,0.10186087,0.033953626,0.33576363,0.8186596,1.0940613,0.56589377,0.79602385,1.0450171,0.7054809,0.003772625,0.02263575,0.003772625,0.124496624,0.14713238,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06413463,0.06413463,0.0,0.0,0.67152727,0.784706,0.935611,1.1431054,0.84884065,0.56589377,0.5281675,0.35085413,0.060362,0.0754525,0.018863125,0.003772625,0.003772625,0.071679875,0.34330887,1.2562841,2.2107582,3.7763977,4.927048,3.0445085,3.9273026,5.8437963,5.560849,3.5764484,4.146115,3.2444575,2.9464202,2.5691576,2.1013522,2.1956677,2.003264,1.9542197,2.2258487,2.1390784,0.13958712,0.08677038,0.3055826,0.8224323,1.5580941,2.3163917,3.3350005,3.7386713,3.5047686,2.9954643,2.957738,3.2670932,3.6368105,3.9612563,4.4215164,5.481624,5.745708,5.409944,5.4476705,6.0512905,6.6322746,5.873977,5.2062225,4.949684,5.028909,4.961002,6.258785,6.696409,6.1305156,4.689373,2.8030603,2.7615614,2.886058,2.7238352,2.335255,2.323937,1.9202662,1.7731338,1.4826416,1.0601076,0.9016574,0.9808825,0.7997965,0.7394345,0.8941121,1.0789708,1.0714256,0.995973,1.1355602,1.3996439,1.3392819,1.2411937,1.5430037,1.7278622,1.6184561,1.388326,1.4071891,1.3770081,1.599593,2.0258996,2.2409391,1.9429018,1.4977322,1.3920987,1.6675003,1.9278114,2.003264,2.052308,2.093807,2.323937,3.1312788,3.8895764,4.398881,4.8100967,5.191132,5.5495315,5.511805,5.1345425,5.0515447,5.323174,5.4665337,4.859141,4.534695,4.22534,4.0178456,4.3611546,4.3309736,3.6745367,3.0256453,2.806833,3.2142766,3.6179473,4.353609,4.9723196,5.4401255,6.1229706,6.5266414,7.4999785,7.7716074,7.5792036,8.66572,9.265567,9.922004,10.329447,10.284176,9.688101,9.382519,9.367428,9.280658,9.125979,9.261794,9.280658,9.476834,9.857869,10.31813,10.642575,10.899114,10.955703,11.09529,11.231105,10.910432,10.70671,10.257768,9.88805,9.81637,10.174769,9.922004,9.465516,9.26934,9.405154,9.556059,9.461743,9.574923,9.793735,9.827688,9.175024,8.684583,8.477088,8.597813,8.8618965,8.892077,8.816625,9.363655,9.891823,10.340765,11.234878,11.714001,12.140307,12.872196,13.634267,13.521088,13.098554,12.781653,12.853333,13.27964,13.721037,13.966258,13.79649,13.102326,12.095036,11.314102,10.808571,10.242677,9.786189,9.439108,9.042982,8.82417,8.058327,6.7756343,5.323174,4.357382,4.002755,3.8103511,3.7952607,3.8707132,3.8669407,4.0895257,4.1272516,3.9688015,3.682082,3.4029078,3.5500402,3.663219,3.9197574,4.304565,4.61392,4.859141,5.3609,5.7570257,5.8966126,5.847569,5.4476705,5.0666356,4.949684,5.13077,5.406172,5.4288073,5.100589,4.432834,3.6556737,3.2331395,2.7011995,2.584248,2.535204,2.4974778,2.704972,2.8294687,3.0633714,3.410453,3.8858037,4.5309224,3.6368105,2.8256962,2.0862615,1.6146835,1.8033148,2.263575,2.2107582,2.5276587,3.2670932,3.640583,3.9499383,4.266839,4.432834,4.617693,5.311856,6.3945994,7.8621507,8.778898,9.144843,9.88805,10.427535,10.397354,10.687846,11.091517,10.306811,11.653639,13.604086,14.762281,14.43029,12.623203,10.4049,9.216523,8.431817,8.050782,8.722309,9.473062,11.45369,13.332457,13.992666,12.521342,11.5857315,11.517824,11.796998,11.917723,11.3820095,10.382264,9.491924,9.371201,10.457717,12.970284,14.139798,14.622695,14.437836,14.094527,14.592513,16.486372,18.063328,19.768555,21.266287,21.409647,21.624687,21.300241,20.526854,19.266796,17.372938,16.31283,14.916959,14.04171,14.268067,15.890297,17.818108,19.225298,19.80251,19.734602,19.70442,18.85558,19.08571,20.130728,21.522825,22.598024,2.0145817,2.4295704,2.9992368,3.3123648,3.2482302,3.006782,3.2746384,3.059599,2.8256962,2.8634224,3.2670932,2.8521044,2.727608,3.0633714,3.5651307,3.4783602,3.2331395,3.3010468,3.4179983,3.5651307,3.9688015,4.1989317,4.191386,4.2064767,4.4818783,5.2628117,5.9117036,7.2358947,9.065618,10.948157,12.132762,13.815352,12.736382,10.842525,9.076936,7.356619,4.5233774,3.1010978,2.4484336,2.0673985,1.6184561,1.7769064,2.3918443,2.354118,1.5882751,1.0525624,0.845068,0.7922512,1.2864652,2.6068838,4.9119577,8.635539,9.548513,8.6581745,6.8397694,4.8365054,5.1647234,7.2358947,10.069136,12.306303,12.223305,12.442118,13.449409,14.124708,13.026875,8.379,6.670001,5.198677,4.3007927,4.3007927,5.5080323,5.9003854,6.6662283,7.356619,7.7376537,7.8131065,6.651138,6.089017,5.9003854,6.1041074,6.9567204,7.2283497,7.888559,6.7039547,5.0741806,8.028146,6.304056,5.4740787,6.0286546,7.3113475,7.5075235,6.8963585,7.541477,8.944894,10.035183,9.171251,8.83926,9.042982,8.737399,7.7338815,6.6850915,6.696409,7.4584794,8.039464,7.8206515,6.515323,5.6363015,5.3986263,4.5761943,2.9124665,1.1280149,2.071171,2.9464202,3.108643,2.4899325,1.5882751,1.1846043,1.4222796,1.3920987,0.9922004,0.9318384,1.237421,2.6483827,2.71629,1.569412,1.9240388,1.9957186,2.4371157,2.9237845,3.3161373,3.6481283,4.2328854,6.3116016,7.3377557,7.1793056,8.13378,10.70671,9.446653,6.7077274,4.315883,3.5689032,3.1425967,4.353609,4.561104,4.508287,8.314865,5.7909794,6.428553,6.9227667,6.7643166,8.254503,7.1793056,8.296002,8.488406,6.9982195,5.3873086,4.749735,4.7950063,4.927048,5.1835866,6.19465,6.4511886,6.8737226,6.964266,7.643338,11.231105,11.378237,16.293968,21.138018,22.49239,18.357594,13.449409,15.052773,18.621677,20.560806,18.218006,20.368402,18.915941,15.901614,14.381247,18.433046,18.406637,16.131744,14.777372,15.565851,17.77661,18.18028,16.03743,16.682549,21.009748,25.450129,28.528591,30.94307,31.414648,31.558008,35.90407,41.555466,46.91259,50.21741,50.74935,48.85927,48.346188,47.85952,47.38417,46.803185,45.897755,42.9702,41.917637,44.16235,48.813995,52.6583,53.94099,47.806705,39.688015,32.82561,28.260735,27.125174,27.902334,28.200373,28.400322,31.648552,33.134964,35.394768,34.960915,31.731548,28.962442,27.717476,27.596752,28.853037,31.12793,33.448093,33.68954,35.93048,38.51473,39.9521,38.925945,40.1445,38.5185,33.044422,26.921452,27.555252,29.252934,24.00144,16.03743,9.337247,7.6282477,19.945868,27.841972,31.93527,31.773048,25.800982,21.394556,14.094527,9.092027,7.3453007,5.5985756,6.307829,8.507269,8.616675,7.0284004,8.103599,5.881522,6.900131,9.703192,12.400619,12.679792,13.241914,12.932558,11.6008215,10.38981,11.717773,9.129752,8.190369,7.537705,6.7152724,6.1795597,6.790725,4.7912335,3.1199608,3.029418,4.104616,5.485397,4.749735,3.5651307,2.8332415,2.686109,3.1614597,4.727099,5.583485,5.59103,6.2851934,11.193378,12.015811,11.363147,11.8045435,15.8676605,20.274086,25.533127,30.064049,32.63698,32.39553,31.686277,28.736084,24.955914,20.922977,16.358103,13.026875,11.34051,10.167224,9.639057,11.140562,11.321648,10.808571,9.574923,8.484633,9.276885,11.242422,12.321393,13.407909,13.705947,10.725573,8.869441,7.0246277,5.5797124,4.9987283,5.828706,3.5085413,2.5917933,2.323937,2.323937,2.595566,2.6898816,2.7351532,2.5389767,2.0787163,1.478869,1.3468271,4.82896,4.7912335,1.2185578,1.20724,1.267602,0.91674787,0.49421388,0.23390275,0.26031113,0.124496624,0.2565385,1.177059,2.4333432,2.595566,0.56589377,0.4376245,0.41121614,0.0,0.0,0.0,0.0,0.1056335,0.20749438,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32821837,0.32821837,0.0,0.0,0.91674787,0.98842776,0.7884786,0.6413463,0.6413463,1.1431054,1.3128735,0.84884065,0.150905,0.32067314,0.0754525,0.02263575,0.02263575,0.041498873,0.1358145,0.5017591,1.3920987,2.3314822,2.6446102,1.4335974,5.692891,6.56814,6.3417826,5.511805,2.776652,2.9728284,3.2670932,2.897376,1.9994912,1.6335466,1.3505998,1.8297231,1.4901869,0.3470815,0.030181,0.056589376,0.18863125,0.7997965,1.7542707,2.425798,3.0256453,3.0746894,2.8332415,2.5917933,2.6408374,3.8480775,4.187614,4.515832,4.919503,4.7006907,5.43258,5.8437963,5.081726,3.983892,5.081726,5.251494,5.1760416,5.2854476,5.6325293,5.8890676,5.7306175,6.2323766,6.096562,4.8666863,2.916239,2.595566,2.6898816,2.5804756,2.335255,2.7011995,2.2598023,1.9391292,1.6184561,1.2525115,0.9016574,0.8639311,0.73566186,0.77338815,0.9808825,1.1280149,1.0789708,0.965792,1.0525624,1.3015556,1.388326,1.2789198,1.6071383,1.7014539,1.4864142,1.50905,1.1204696,1.0940613,1.358145,1.7391801,1.9844007,1.6675003,1.3128735,1.1732863,1.3053282,1.5882751,1.4637785,1.5165952,1.7731338,2.1805773,2.595566,2.8143783,3.7462165,4.45547,4.7950063,5.4174895,5.515578,4.8063245,3.8178966,3.3538637,4.5007415,4.5007415,4.146115,3.983892,4.142342,4.2894745,3.983892,3.4481792,2.9464202,2.7502437,3.127506,3.5424948,4.2064767,4.768598,5.2062225,5.828706,6.587003,7.8734684,8.201687,7.907422,9.14107,8.884532,8.918486,9.024119,9.027891,8.820397,9.295748,9.507015,9.250477,8.858124,9.201432,10.227587,11.1782875,11.732863,11.947904,12.253486,12.313848,11.521597,10.974566,10.948157,10.910432,10.178542,9.876732,9.955957,10.223814,10.344538,10.065364,9.710737,9.582467,9.748463,10.054046,10.03141,10.042727,10.340765,10.653893,10.178542,9.273112,8.744945,8.5563135,8.563859,8.514814,8.820397,9.639057,10.469034,11.016065,11.200924,12.064855,12.879742,13.611631,14.094527,14.007756,13.215506,12.996693,13.132507,13.377728,13.487134,13.841762,13.585222,12.887287,11.861133,10.544487,10.714255,10.419991,10.057818,9.590013,8.529905,8.311093,6.752999,5.2326307,4.3686996,4.0291634,3.7235808,3.4557245,3.31991,3.2935016,3.218049,3.7952607,4.13857,3.9688015,3.4632697,3.2821836,3.1954134,3.1840954,3.6028569,4.3347464,4.7610526,4.61392,5.062863,5.5080323,5.564622,5.0666356,4.640329,4.504514,4.4139714,4.504514,5.311856,5.323174,4.6742826,4.187614,3.9197574,3.1727777,2.6597006,2.5691576,2.4408884,2.4107075,3.2029586,3.1425967,3.4481792,3.6179473,3.4444065,3.006782,2.4333432,1.841041,1.5165952,1.5958204,2.0598533,1.6825907,2.4182527,3.006782,3.0897799,3.2520027,4.055572,5.2099953,5.802297,5.692891,5.5080323,6.375736,7.7716074,8.816625,9.473062,10.559577,10.963248,11.042474,11.249968,11.476325,11.0613365,11.355601,12.362892,12.577931,11.84227,11.351829,9.839006,9.224068,8.484633,7.6584287,7.8432875,9.442881,11.45369,12.966512,12.996693,10.484125,9.95973,10.469034,11.034928,11.102836,10.529396,10.016319,9.540969,9.397609,10.197406,12.849561,13.762536,13.698401,13.3626375,13.264549,13.702174,16.33924,18.693357,20.77962,22.315077,22.703657,24.254206,22.620659,20.1345,17.961468,16.06761,15.456445,14.479335,14.034165,14.558559,16.03743,17.56157,18.99894,19.930779,19.938324,18.568861,18.327412,19.591242,20.960705,21.73032,21.926497,2.795515,2.7502437,3.1350515,4.304565,5.6023483,5.3382645,3.8480775,3.259548,3.0181,2.886058,2.9351022,3.1954134,3.270866,3.2255943,3.0030096,2.4295704,2.3692086,2.535204,2.6936543,2.9011486,3.4783602,4.063117,4.327201,4.561104,4.9949555,5.8136153,6.3832817,7.7225633,8.635539,8.7751255,8.650629,8.971302,8.601585,7.748972,6.6360474,5.5004873,3.5839937,2.5540671,2.1654868,2.0975795,1.9466745,2.4974778,2.5804756,2.323937,1.8674494,1.3694628,1.3392819,1.7467253,2.7841973,4.357382,6.096562,7.6622014,8.284684,6.9227667,4.61392,4.459243,5.089271,6.488915,7.8508325,8.503497,7.888559,7.835742,7.273621,6.6850915,6.047518,4.8138695,5.583485,6.198423,7.5716586,9.06939,8.511042,7.3188925,6.9793563,6.3531003,5.292993,4.6629643,4.7421894,4.7233267,5.2628117,6.1606965,6.3719635,6.4549613,6.4210076,5.4703064,4.29702,5.0854983,4.878004,4.7950063,5.4967146,6.6360474,6.858632,7.001992,7.092535,7.01331,6.8737226,7.020855,6.3908267,5.6589375,5.081726,4.6554193,4.1310244,4.6931453,5.1156793,5.194905,5.149633,5.613666,5.1043615,4.146115,3.1840954,2.493705,2.1654868,2.8634224,2.9652832,2.535204,1.8297231,1.3053282,1.3241913,2.1277604,2.0372176,1.3166461,2.1654868,1.7769064,2.2258487,2.2220762,1.6486372,1.5430037,2.191895,3.3538637,5.0553174,6.7341356,7.2585306,7.564113,8.311093,8.416726,8.182823,9.280658,9.922004,7.805561,4.6742826,2.1881225,1.9089483,1.599593,1.8221779,2.584248,4.315883,7.888559,4.5912848,5.1571784,7.111398,8.778898,9.280658,9.574923,9.088254,7.5792036,5.8136153,5.5683947,5.6853456,5.836251,5.7607985,5.515578,5.4740787,5.4288073,4.9685473,4.878004,5.594803,7.1906233,7.5905213,12.400619,16.097792,16.0412,12.510024,8.793989,9.880505,13.70972,17.123945,15.863888,14.388792,13.35132,13.528633,14.5283785,14.781145,15.852571,17.142809,17.80679,18.429274,21.058792,21.100292,20.187317,22.077402,26.838455,30.822346,35.636215,36.87741,37.53762,39.416386,43.117332,45.037598,50.65881,54.869057,57.05341,61.0788,63.229195,60.305412,55.18596,49.6402,44.31325,39.5937,38.86558,45.305454,58.13615,72.615486,68.29206,57.664574,45.837395,35.953117,29.211435,25.585943,25.963205,27.287397,28.558771,30.829891,36.526554,41.344196,43.12865,40.808483,34.40634,31.361832,31.10152,32.282352,33.957397,35.5834,34.33466,37.03586,39.197575,38.47323,34.666653,39.389977,39.88042,34.315796,27.898561,32.818066,32.893517,22.213217,11.827179,8.07719,12.608112,15.943113,23.861853,30.818573,33.206646,29.354795,23.141281,15.433809,10.785934,9.58624,8.065872,8.069645,8.650629,8.22055,7.4735703,9.397609,5.4174895,4.5460134,5.2062225,6.6247296,8.846806,11.351829,11.714001,10.03141,8.329956,10.559577,10.148361,8.956212,7.624475,6.7831798,7.0472636,6.330465,4.5761943,3.2105038,2.987919,3.983892,4.610148,3.9574835,3.0218725,2.4371157,2.4672968,3.1576872,4.425289,6.9152217,8.884532,6.2021956,10.005001,12.004493,11.98563,11.638548,14.551015,17.855835,21.77559,26.348013,31.071339,34.9081,33.847992,31.256199,27.230806,22.945105,20.66644,16.81459,14.890551,13.472044,12.196897,11.774363,11.3820095,10.687846,9.895596,9.450426,10.057818,9.952185,11.378237,13.083464,13.781399,12.128989,10.099318,8.137552,6.3719635,5.070408,4.6214657,4.1272516,4.82896,5.323174,5.5193505,6.6586833,3.7877154,2.9803739,2.7540162,2.323937,1.5882751,1.2902378,1.7769064,1.6335466,0.7997965,0.58475685,0.4979865,0.5696664,0.55457586,0.392353,0.22258487,0.87902164,1.4713237,2.0183544,2.3013012,1.8749946,1.1657411,0.5017591,0.1056335,0.00754525,0.03772625,0.124496624,0.124496624,0.08677038,0.0452715,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.56212115,0.8337501,0.6488915,0.56212115,0.7432071,0.7092535,0.86770374,1.1883769,1.177059,1.6109109,1.478869,1.1355602,0.87147635,0.8941121,0.4640329,0.211267,0.17731337,0.25276586,0.17354076,0.58098423,1.2940104,1.931584,1.8976303,0.38480774,2.0485353,1.9768555,1.6260014,1.5430037,1.3845534,1.8070874,1.7844516,1.4600059,0.9507015,0.35085413,0.38103512,0.58098423,0.4678055,0.090543,0.018863125,0.05281675,0.2263575,0.65643674,1.2940104,1.9240388,2.3201644,2.263575,2.0862615,2.0787163,2.516341,3.561358,3.8858037,4.466788,5.3194013,5.5306683,4.738417,5.3646727,5.6778007,5.13077,4.323428,5.138315,5.7004366,5.956975,6.0248823,6.19465,5.956975,5.8966126,5.4174895,4.255521,2.5012503,2.3277097,2.305074,2.2899833,2.3126192,2.5917933,2.142851,1.8976303,1.6109109,1.2487389,1.0223814,1.1996948,1.0902886,0.935611,0.9016574,1.0676528,1.146878,1.0714256,1.0601076,1.1393328,1.1581959,1.1053791,1.2826926,1.3355093,1.2147852,1.1808317,1.0827434,1.2638294,1.5279131,1.7391801,1.8372684,1.6448646,1.4411428,1.3204187,1.3392819,1.5015048,1.5656394,1.5845025,1.7127718,2.0145817,2.4484336,2.6483827,3.519859,4.5422406,5.3458095,5.6853456,5.2665844,4.927048,4.29702,3.5424948,3.3425457,4.1800685,4.195159,3.8480775,3.4481792,3.1652324,3.0633714,2.969056,2.837014,2.727608,2.8219235,3.218049,3.8405323,4.3649273,4.7912335,5.413717,6.375736,7.84706,8.854351,9.363655,10.27663,9.665465,9.718282,10.084227,10.321902,9.880505,9.831461,9.95973,9.661693,9.137298,9.420244,10.699164,11.921495,12.54775,12.796744,13.619176,12.800517,11.77059,11.18206,11.114153,11.057564,10.695392,10.49167,10.469034,10.650121,11.065109,10.435081,10.18986,10.223814,10.31813,10.152134,10.216269,10.427535,10.79348,11.038701,10.593531,9.718282,9.22784,8.914713,8.771353,8.9788475,9.390063,9.861642,10.359629,10.970794,11.895086,13.230596,14.196388,14.811326,14.9358225,14.264296,13.275867,12.725064,12.291212,12.106354,12.743927,13.147598,12.400619,11.446144,10.506761,9.092027,9.612649,10.438853,10.801025,10.201178,8.394091,6.749226,5.372218,4.496969,4.1083884,3.942393,3.4330888,3.0897799,3.0331905,3.1727777,3.2067313,3.2746384,3.2557755,2.8747404,2.372981,2.5125682,2.7389257,2.9351022,3.3048196,3.8443048,4.357382,4.4177437,4.4705606,4.466788,4.3083377,3.8593953,4.025391,4.274384,4.429062,4.5761943,5.0779533,4.9534564,4.4101987,3.92353,3.4557245,2.4786146,2.474842,2.4069347,2.1353056,1.9730829,2.6672459,3.682082,3.572676,3.138824,2.7804246,2.505023,1.6675003,1.3091009,1.3392819,1.5316857,1.5467763,2.1051247,2.516341,2.7804246,3.108643,3.9197574,4.2894745,4.436607,4.859141,5.553304,6.043745,6.6662283,7.4471617,8.461998,9.473062,9.9257765,10.552032,11.080199,11.563096,11.864905,11.634775,12.076173,12.291212,11.759273,10.529396,9.239159,8.635539,8.420499,8.235641,8.171506,8.782671,10.03141,11.2801485,11.944131,11.604594,10.020092,9.57115,10.220041,10.714255,10.612394,10.284176,10.095545,9.880505,10.253995,11.3820095,13.008011,13.513543,13.807808,14.075664,14.543469,15.471535,17.28994,19.289433,21.553007,23.55627,24.17121,22.986605,21.507734,19.65915,17.595524,15.712983,15.377219,14.70192,14.335975,14.754736,16.28265,17.818108,19.093256,19.742147,19.54597,18.41041,18.293459,19.006485,20.183544,21.409647,22.22076,3.127506,2.9841464,3.108643,3.9763467,5.089271,5.0062733,4.014073,3.5538127,3.3010468,3.0822346,2.8709676,3.029418,3.029418,2.9464202,2.7653341,2.4031622,2.4861598,2.584248,2.674791,2.9011486,3.5764484,3.9612563,4.244203,4.5988297,5.149633,5.9796104,6.907676,7.9225125,8.654402,9.110889,9.650374,9.280658,8.8618965,8.397863,7.7678347,6.730363,5.119452,3.5387223,2.4823873,2.1390784,2.3880715,3.0935526,2.795515,2.2258487,1.8070874,1.6335466,1.7467253,2.474842,3.4481792,4.353609,4.927048,4.8327327,4.983638,4.3309736,3.199186,3.2482302,3.904667,4.606375,5.093044,5.3458095,5.560849,6.33801,6.519096,6.5530496,6.990674,8.518587,8.537451,8.107371,8.371455,9.22784,9.325929,8.544995,8.103599,7.443389,6.2625575,4.4894238,4.5950575,4.961002,6.4474163,8.201687,7.6810646,7.3453007,7.6923823,7.5905213,6.858632,6.300284,6.9454026,7.413208,7.1000805,5.9418845,4.402653,4.52715,5.492942,5.8702044,5.300538,4.52715,4.1989317,3.742444,3.5387223,3.5123138,3.127506,3.772625,4.61392,4.9459114,4.798779,4.957229,4.1536603,3.0331905,2.2107582,1.9353566,2.0975795,2.5125682,2.372981,1.8787673,1.2789198,0.8865669,0.9808825,1.4637785,1.6410918,1.6675003,2.535204,2.5691576,2.6823363,2.5238862,2.1353056,1.9542197,2.5767028,4.4516973,6.579458,8.186596,8.703445,9.073163,8.986393,8.590267,8.243186,8.503497,7.9225125,5.8588867,3.7575345,2.4974778,2.372981,1.9089483,1.8825399,2.6068838,4.0480266,5.8513412,3.6330378,4.08198,5.66271,7.0057645,6.8737226,6.937857,7.0359454,6.6247296,6.198423,7.3000293,7.1793056,6.0814714,5.3382645,5.2099953,4.881777,4.606375,4.3611546,4.564876,5.5570765,7.5603404,8.869441,11.336739,12.208215,10.740664,8.209232,6.643593,7.907422,11.544232,15.203679,14.622695,12.272349,11.25374,12.276122,14.698147,16.505234,17.667202,19.640285,20.145817,19.7761,21.983086,22.115128,22.986605,25.020048,28.223007,32.21067,38.186512,42.234535,44.99987,48.40278,55.642445,57.317493,59.811195,63.614002,68.73723,74.68666,76.82574,74.034,66.19825,54.963375,43.739815,37.707386,36.36056,41.842182,56.43847,82.58653,88.1172,70.959305,50.677673,36.67746,28.1966,23.895807,24.141027,26.812046,29.781101,30.909117,36.08516,44.411343,52.6583,56.098934,48.54614,38.450596,35.677715,36.307743,37.82811,39.14853,36.775547,37.6093,37.273537,34.602516,31.659868,38.684498,40.808483,37.560253,33.078377,36.092705,32.459667,19.817598,9.465516,6.7039547,10.789707,11.955449,20.500444,28.660633,31.893772,28.853037,24.435291,17.08999,12.193124,10.736891,9.333474,8.89585,9.0957985,7.937603,6.4134626,8.511042,5.485397,4.3083377,4.6629643,6.2663302,8.858124,10.084227,9.144843,7.0812173,6.013564,9.125979,10.057818,9.224068,7.7037,6.3342376,5.715527,7.194396,6.2323766,4.447925,3.2105038,3.6594462,3.9801195,3.6934,3.180323,2.7615614,2.6936543,3.1237335,4.6742826,8.480861,11.566868,6.8397694,9.906913,12.294985,12.845788,12.174261,12.683565,16.509007,22.254715,27.792929,32.489845,37.186764,36.156837,33.48582,29.652832,25.8123,23.805264,19.964731,17.769064,16.0827,14.664193,14.147344,12.989148,12.340257,11.6008215,10.770844,10.446399,9.009028,10.03141,11.812089,12.917468,12.162943,10.438853,8.937348,7.2396674,5.511805,4.538468,5.247721,5.1043615,5.093044,5.798525,7.4169807,4.032936,3.2218218,2.8936033,2.191895,1.4901869,1.3468271,1.1959221,1.0110635,0.7582976,0.4074435,0.20749438,0.2678564,0.35085413,0.3470815,0.2867195,0.63002837,0.935611,1.1808317,1.3732355,1.539231,1.8561316,1.1921495,0.41876137,0.003772625,0.018863125,0.06413463,0.10186087,0.07922512,0.030181,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24899325,0.5319401,0.7582976,0.9507015,1.116697,1.1242423,1.2751472,1.5430037,1.569412,2.2748928,2.1541688,1.7052265,1.2751472,1.0374719,0.5696664,0.38480774,0.39989826,0.44516975,0.2565385,0.47912338,1.0714256,1.5279131,1.3807807,0.20372175,0.63002837,0.58475685,0.482896,0.5357128,0.7432071,1.8297231,1.4939595,0.84884065,0.39989826,0.0754525,0.09808825,0.13958712,0.10186087,0.011317875,0.00754525,0.033953626,0.20749438,0.52439487,1.0072908,1.6712729,1.8146327,1.961765,2.0108092,2.1088974,2.6597006,3.531177,3.6066296,3.99521,4.9459114,5.855114,5.2250857,5.643847,6.1795597,6.2021956,5.3910813,5.349582,5.6363015,5.6023483,5.2665844,5.3571277,5.281675,5.198677,4.749735,3.7763977,2.293756,2.1956677,2.093807,2.0258996,2.11267,2.535204,2.305074,2.1353056,1.780679,1.2789198,0.94315624,1.2261031,1.1393328,0.9620194,0.875249,0.9507015,1.056335,1.0223814,1.026154,1.0902886,1.0978339,1.1053791,1.1317875,1.1657411,1.1657411,1.0902886,1.0072908,1.2110126,1.4600059,1.6410918,1.7919968,1.7580433,1.6524098,1.5543215,1.5241405,1.599593,1.539231,1.5731846,1.6712729,1.9127209,2.4823873,2.7238352,3.4670424,4.395108,5.1647234,5.4401255,5.7570257,5.4778514,4.7572803,3.8065786,2.897376,3.8669407,4.0291634,3.8443048,3.5274043,3.048281,2.8106055,2.6446102,2.6144292,2.848332,3.5538127,3.591539,3.6066296,3.9650288,4.6931453,5.485397,7.069899,8.182823,8.892077,9.476834,10.438853,10.103089,9.676784,9.676784,10.012547,9.982366,10.170997,10.529396,10.242677,9.612649,10.042727,10.834979,11.593277,12.2270775,12.687338,12.936331,12.068627,11.480098,11.359374,11.623458,11.9064045,11.815862,11.631002,11.438599,11.249968,11.034928,10.095545,9.616421,9.567377,9.703192,9.556059,9.537196,9.718282,9.922004,9.955957,9.590013,8.7600355,8.488406,8.492179,8.601585,8.782671,9.359882,9.797507,10.03141,10.423763,11.740409,13.170234,14.022847,14.407655,14.27184,13.358865,12.283667,11.793225,11.355601,11.114153,11.898859,12.079946,11.400873,10.54826,9.737145,8.729855,9.190115,9.737145,9.654147,8.654402,6.8699503,5.5495315,4.666737,4.164978,3.8707132,3.500996,3.3651814,3.1652324,3.1161883,3.2369123,3.3425457,3.0822346,2.6408374,2.2258487,2.0673985,2.4182527,2.6446102,2.8521044,3.0181,3.2746384,3.9386206,4.2064767,4.085753,3.9008942,3.7084904,3.2972744,3.6368105,3.9989824,4.293247,4.5535583,4.927048,4.5120597,3.9273026,3.350091,2.8256962,2.2862108,2.1503963,2.1843498,2.203213,2.2673476,2.6974268,3.3274553,3.3651814,2.9615107,2.323937,1.7127718,1.5467763,1.5128226,1.5203679,1.6448646,2.0862615,2.3956168,2.6031113,2.916239,3.410453,4.032936,4.3422914,4.689373,5.3080835,5.9984736,6.115425,6.537959,7.352846,8.699674,10.163452,10.801025,11.257513,12.083718,13.13628,13.853079,13.290957,12.857106,12.204442,11.144334,9.8239155,8.722309,8.013056,7.466025,7.5263867,8.246958,9.273112,9.952185,10.510533,10.461489,9.865415,9.318384,9.688101,10.480352,10.623712,9.963503,9.261794,9.876732,10.47658,11.261286,12.155397,12.83447,13.430545,13.705947,13.845533,14.335975,15.988385,18.184053,20.02132,21.734093,22.99415,22.89606,21.417192,19.998686,18.5085,16.825907,14.864142,14.494425,14.358611,14.524607,15.290449,17.191853,18.568861,19.097027,19.206434,19.036665,18.417955,18.010511,18.651857,19.719511,20.764528,21.51528,3.2935016,3.3312278,3.3689542,3.682082,4.1310244,4.1612053,3.7688525,3.5877664,3.5085413,3.3953626,3.108643,3.0105548,2.8181508,2.6672459,2.6068838,2.5993385,2.565385,2.7841973,2.9615107,3.0671442,3.3312278,3.7273536,4.0782075,4.4705606,4.98741,5.726845,6.696409,7.61693,8.597813,9.635284,10.61994,10.197406,9.563604,9.001483,8.492179,7.699928,6.4511886,4.8365054,3.3350005,2.354118,2.233394,2.535204,2.11267,1.569412,1.2789198,1.3807807,1.5203679,2.5880208,3.5500402,3.9386206,3.8556228,3.0671442,2.8709676,2.7615614,2.6068838,2.6672459,3.3538637,3.9499383,4.3196554,4.6742826,5.564622,6.5643673,6.9944468,7.8131065,9.378746,11.476325,11.706455,11.076427,10.574668,10.401127,9.989911,8.816625,7.798016,7.039718,6.300284,5.0025005,5.040227,5.6815734,6.903904,8.182823,8.511042,8.416726,9.016574,9.224068,8.688355,7.7942433,7.4396167,7.7716074,7.175533,5.3156285,3.1312788,3.1576872,4.1310244,4.768598,4.395108,2.9464202,2.7841973,2.7992878,2.9916916,3.2369123,3.2935016,3.9876647,5.0062733,5.4401255,5.2175403,5.0854983,3.451952,2.3428001,1.7618159,1.6071383,1.6825907,1.9504471,1.7240896,1.2826926,0.8526133,0.6187105,0.7092535,0.87147635,1.1619685,1.6260014,2.2862108,2.6785638,2.795515,2.5389767,2.1881225,2.3805263,3.1312788,4.9459114,6.609639,7.5112963,7.6282477,7.8734684,7.5905213,7.213259,6.903904,6.5228686,5.6023483,4.52715,3.6443558,3.138824,2.9916916,2.7125173,2.6710186,3.078462,3.7386713,4.025391,3.078462,3.5575855,4.4441524,4.9647746,4.5912848,4.236658,4.568649,4.919503,5.3873086,6.8246784,6.300284,5.191132,4.878004,5.3986263,5.43258,4.647874,4.395108,5.27413,7.020855,8.52236,10.438853,10.518079,9.152389,7.183078,5.8890676,6.3644185,7.4735703,9.408927,11.415963,11.781908,11.608367,12.102581,13.264549,15.267814,18.448135,19.968504,21.160654,21.636003,21.613369,21.915178,21.726547,23.880716,27.302486,31.199608,35.06278,42.830612,50.353226,55.77826,61.188206,72.60417,75.83731,75.245,76.489975,80.50404,83.50328,83.68814,81.447205,73.40396,59.739517,44.192528,35.726757,33.448093,36.696323,48.648,76.34284,99.94438,85.73668,59.105717,36.900043,27.426983,23.054512,23.246916,26.58946,30.584671,31.678732,34.870373,43.82281,57.219402,69.454025,70.653725,53.197784,43.600227,40.004917,40.065277,40.925434,37.786613,36.243607,34.15735,31.47501,30.218727,39.963417,46.044888,46.418377,42.185493,37.635708,27.49489,15.079182,7.201941,5.7909794,7.914967,9.0957985,17.003222,25.133228,29.279343,27.5213,24.265524,18.03692,13.211733,10.853842,8.744945,8.620448,8.771353,7.356619,5.515578,7.352846,5.3873086,4.429062,5.2892203,7.5490227,9.529651,9.175024,6.7643166,4.459243,4.2404304,7.911195,9.374973,9.307066,7.986647,6.085244,4.659192,10.076681,9.276885,6.4738245,4.236658,3.500996,3.7499893,3.8480775,3.712263,3.470815,3.440634,3.62172,4.983638,8.337502,11.038701,6.990674,8.60913,13.373956,14.607604,12.095036,12.102581,17.712475,23.80149,29.13221,33.74236,38.937263,39.46543,37.941288,34.98355,31.184519,27.110083,23.888262,20.311813,17.123945,14.999957,14.592513,13.43809,13.045737,12.37421,11.227332,10.238904,8.7600355,8.975075,10.174769,11.449917,11.69891,10.574668,9.710737,8.265821,6.3417826,4.9534564,5.9230213,4.9421387,4.557331,5.4967146,6.6850915,4.006528,3.361409,2.837014,1.8900851,1.3430545,1.2638294,1.1506506,0.9922004,0.7507524,0.3734899,0.14713238,0.15845025,0.59230214,1.1544232,1.0789708,1.7731338,1.5241405,1.297783,1.3770081,1.3732355,1.7844516,1.4071891,0.66020936,0.0150905,0.0,0.018863125,0.071679875,0.071679875,0.03772625,0.071679875,0.05281675,0.030181,0.011317875,0.026408374,0.1358145,0.026408374,0.0,0.0,0.10940613,0.55080324,0.10940613,0.27917424,0.724344,1.1317875,1.20724,1.5165952,1.5807298,1.5467763,1.5958204,1.9466745,2.4559789,2.6634734,2.4031622,1.8599042,1.569412,1.026154,0.72811663,0.58475685,0.52439487,0.5055317,0.58475685,0.9393836,1.2713746,1.2449663,0.52062225,0.29426476,0.40367088,0.52439487,0.80356914,1.8674494,2.7125173,2.474842,1.6939086,0.87902164,0.5093044,0.2867195,0.12826926,0.03772625,0.003772625,0.0,0.02263575,0.18863125,0.45648763,0.84884065,1.4637785,1.6184561,1.9844007,2.2711203,2.463524,2.7879698,3.6745367,4.13857,4.4931965,4.9044123,5.3759904,5.583485,6.247467,6.9454026,7.2623034,6.7756343,5.802297,5.5570765,5.20245,4.6252384,4.429062,4.52715,4.4743333,4.1272516,3.4368613,2.4371157,2.233394,2.1579416,2.1051247,2.1654868,2.6219745,2.4182527,2.3428001,1.9579924,1.3166461,0.935611,1.1808317,1.0978339,0.9695646,0.90543,0.8601585,0.8941121,0.90543,0.97333723,1.0638802,1.0450171,1.1619685,1.1091517,1.1053791,1.2034674,1.2600567,0.94315624,1.0638802,1.2751472,1.448688,1.7052265,1.841041,1.8674494,1.7957695,1.6788181,1.599593,1.5316857,1.5769572,1.7014539,1.9429018,2.3880715,2.5578396,3.2821836,4.0895257,4.738417,5.20245,6.043745,5.9984736,5.372218,4.429062,3.4029078,3.8443048,4.2027044,4.236658,3.8820312,3.2633207,2.837014,2.6974268,2.8143783,3.2218218,4.002755,3.9122121,3.5274043,3.7160356,4.640329,5.783434,7.141579,8.14887,8.869441,9.556059,10.627484,10.18986,9.937095,9.978593,10.231359,10.438853,10.982111,11.306557,10.872705,10.11818,10.435081,10.544487,10.846297,11.491416,12.185578,12.178034,11.774363,11.563096,11.717773,12.117672,12.340257,12.136535,11.6875925,11.216014,10.7557535,10.144588,9.193887,8.511042,8.280911,8.382772,8.379,8.390318,8.552541,8.718536,8.692128,8.2507305,7.665974,7.5829763,7.84706,8.27714,8.68081,9.073163,9.457971,9.627739,9.948412,11.3669195,12.687338,13.343775,13.407909,12.96274,12.106354,11.306557,11.016065,10.782163,10.604849,10.933067,10.552032,10.091772,9.488152,8.797762,8.186596,8.390318,8.329956,7.748972,6.628502,5.191132,4.557331,4.2404304,3.9574835,3.5839937,3.1350515,3.2218218,3.218049,3.2067313,3.2218218,3.2444575,2.7841973,2.2711203,1.9957186,2.0447628,2.305074,2.5087957,2.655928,2.7728794,3.0181,3.6934,4.08198,3.9989824,3.7914882,3.5651307,3.187868,3.519859,3.8593953,4.164978,4.406426,4.5912848,3.9008942,3.240685,2.7426984,2.463524,2.3880715,1.9730829,2.0258996,2.335255,2.6408374,2.637065,2.9652832,2.9766011,2.6106565,1.9655377,1.3015556,1.7693611,1.8221779,1.7882242,1.9391292,2.5012503,2.5012503,2.746471,3.0558262,3.440634,4.0970707,4.5988297,5.2665844,6.0022464,6.6322746,6.9227667,7.0170827,7.8395147,9.118435,10.495442,11.502733,11.615912,12.3289385,13.698401,14.947141,14.48688,13.030646,11.7894535,10.435081,9.122208,8.52236,7.8696957,7.326438,7.6018395,8.597813,9.416472,9.552286,9.631512,9.265567,8.82417,9.408927,9.971047,10.469034,10.34831,9.623966,8.888305,9.601331,10.95193,12.049765,12.58925,12.842015,13.034419,13.389046,13.70972,14.373701,16.31283,18.640541,20.111864,21.066338,21.42851,20.70794,19.734602,18.376457,17.063583,15.758255,13.981348,13.441863,13.898351,14.777372,15.973294,17.810562,18.742401,18.715992,18.429274,18.150099,17.72002,17.493662,18.429274,19.595015,20.455173,20.88148,3.3123648,3.5274043,3.610402,3.6858547,3.7575345,3.731126,3.470815,3.4594972,3.5651307,3.6254926,3.4255435,3.2520027,2.897376,2.584248,2.463524,2.595566,2.3767538,2.7917426,3.1840954,3.1954134,2.7615614,3.31991,3.7952607,4.187614,4.587512,5.198677,5.794752,6.8058157,8.043237,9.167479,9.665465,9.533423,9.016574,8.258276,7.5037513,7.1076255,6.4511886,5.587258,4.2328854,2.6182017,1.4864142,1.116697,0.7922512,0.58475685,0.55457586,0.7432071,0.79602385,1.9164935,2.9992368,3.5274043,3.5424948,2.7502437,2.4672968,2.3578906,2.3578906,2.6898816,3.3878171,4.191386,4.949684,5.723072,6.790725,7.250985,6.692637,7.413208,9.476834,10.740664,12.019584,12.381755,12.898605,13.204187,11.491416,9.167479,7.2057137,5.987156,5.726845,6.458734,6.356873,6.515323,6.126743,5.8173876,7.6697464,8.439363,8.892077,9.058073,8.926031,8.431817,6.7039547,6.439871,6.3644185,5.6589375,3.9725742,4.0895257,3.9008942,3.85185,3.7160356,2.637065,2.4408884,2.71629,3.0407357,3.350091,3.9159849,4.825187,5.6287565,5.956975,5.8588867,5.783434,3.3878171,2.305074,1.841041,1.6222287,1.6184561,1.5807298,1.2826926,0.94692886,0.72811663,0.7167987,0.79602385,0.95824677,1.1091517,1.3128735,1.7957695,2.123988,2.2975287,1.9844007,1.6109109,2.335255,3.6707642,4.745962,5.4967146,5.772116,5.342037,5.3080835,5.2590394,5.2099953,5.062863,4.606375,3.8971217,3.9197574,3.651901,2.9841464,2.7426984,2.9766011,2.9086938,3.1237335,3.500996,3.2218218,2.8256962,3.31991,3.783943,3.8178966,3.5274043,3.0671442,2.9124665,3.138824,3.7462165,4.67051,4.357382,4.406426,5.194905,6.3342376,6.6662283,5.1081343,4.376245,5.8400235,8.431817,8.616675,9.993684,8.7600355,6.719045,5.1760416,4.961002,6.598321,7.0849895,6.85486,6.8699503,8.612903,12.0233555,14.70192,15.905387,16.520325,19.04421,20.477808,20.432537,21.68505,23.458181,21.420965,20.590988,23.552498,29.305752,36.066296,41.27252,50.46263,60.810944,71.147934,82.82421,99.702934,104.22631,97.726074,90.96931,88.09457,86.623245,81.33402,77.79153,71.34411,60.0451,44.66411,33.542408,30.463947,32.440804,40.219955,58.275738,95.47382,95.93785,71.1668,39.92569,28.234325,23.809036,23.722265,26.815819,31.007204,33.27078,35.338177,41.381924,55.2765,74.83756,91.84078,73.60014,54.54084,42.940018,40.020004,39.933235,35.55322,32.950108,31.765503,31.22979,30.177227,40.81603,52.337627,56.562965,50.40227,35.84371,19.538425,9.107117,4.949684,5.3948536,6.7152724,7.6848373,13.977575,21.41342,26.525326,26.536644,22.42071,17.614386,13.494679,10.314357,7.194396,7.5792036,7.4735703,6.3644185,5.243949,6.6247296,4.878004,4.0706625,5.2779026,7.745199,8.8769865,8.096053,5.2288585,3.108643,3.4594972,6.8925858,8.763808,9.593785,8.722309,6.6247296,4.8855495,12.245941,11.3669195,8.303548,5.926794,3.9159849,3.904667,4.1536603,4.3007927,4.3611546,4.719554,4.636556,5.2552667,6.7869525,8.031919,6.3908267,6.6813188,14.030393,15.992157,11.962994,13.185325,19.647831,23.94485,28.166418,33.410366,39.78233,42.732525,43.5625,41.72523,37.141495,30.173454,27.476028,22.194353,16.957949,13.543724,12.849561,12.249713,12.261031,11.936585,11.027383,9.952185,9.352338,8.944894,9.231613,10.246449,11.566868,11.140562,10.691619,9.510788,7.5565677,5.451443,6.1606965,5.4401255,5.409944,6.3455553,6.673774,4.191386,3.3727267,2.6295197,1.6260014,1.237421,1.026154,0.84884065,0.7469798,0.6526641,0.41121614,0.27540162,0.47535074,1.3128735,2.2711203,2.0258996,3.6934,3.5877664,3.3576362,3.0633714,1.1732863,1.599593,1.2826926,0.65643674,0.11317875,0.0,0.0452715,0.0754525,0.1056335,0.11317875,0.056589376,0.09808825,0.0754525,0.060362,0.124496624,0.34330887,0.5394854,0.66775465,0.56589377,0.5998474,1.6524098,0.8262049,1.1204696,1.7316349,2.0900342,1.8146327,2.2560298,2.3503454,2.3428001,2.4031622,2.6219745,2.293756,2.8747404,3.0331905,2.546522,2.282438,1.6712729,1.1619685,0.7884786,0.66020936,0.97333723,0.8941121,0.98465514,1.2713746,1.4826416,1.056335,0.4376245,0.42630664,0.6752999,1.5279131,4.0216184,4.014073,4.055572,3.429316,2.2107582,1.2864652,0.7696155,0.331991,0.08299775,0.0150905,0.0,0.033953626,0.21881226,0.47535074,0.77716076,1.1732863,1.5920477,2.0145817,2.4559789,2.8445592,3.029418,3.8480775,4.9760923,5.6476197,5.5382137,4.776143,5.50426,6.6662283,7.6018395,7.9262853,7.5037513,6.2889657,5.7683434,5.2779026,4.606375,4.0103,4.172523,4.0291634,3.7047176,3.2821836,2.8181508,2.4522061,2.516341,2.6031113,2.6332922,2.8521044,2.444661,2.4333432,2.0900342,1.3996439,1.0336993,1.1808317,1.1053791,1.0186088,0.965792,0.8224323,0.7884786,0.84884065,0.97333723,1.0638802,0.9808825,1.177059,1.1091517,1.0450171,1.1355602,1.3845534,0.9280658,0.97710985,1.1732863,1.358145,1.5882751,1.7278622,1.9164935,1.9466745,1.7655885,1.478869,1.539231,1.5316857,1.690136,1.991946,2.191895,2.2711203,3.0860074,3.8593953,4.4403796,5.281675,5.9418845,6.2889657,6.047518,5.2892203,4.4403796,4.236658,4.7610526,4.738417,3.9574835,3.2557755,2.867195,3.0143273,3.3764994,3.7047176,3.8405323,3.8858037,3.5764484,3.7084904,4.587512,5.994701,6.598321,7.7414265,8.899622,9.918231,11.027383,10.306811,10.650121,11.09529,11.249968,11.32542,12.15917,12.079946,11.351829,10.593531,10.774617,10.469034,10.431308,10.8576145,11.559323,11.962994,12.178034,12.061082,12.057309,12.121444,11.717773,11.185833,10.412445,9.688101,9.137298,8.729855,8.13378,7.4773426,7.1076255,7.0585814,7.0246277,7.0849895,7.3415284,7.647111,7.7301087,7.2094865,7.066127,7.0057645,7.232122,7.809334,8.684583,8.793989,9.0807085,9.42779,10.023865,11.378237,12.445889,12.875969,12.630749,11.925267,11.261286,10.785934,10.56335,10.47658,10.359629,10.005001,9.186342,8.714764,8.262049,7.699928,7.0963078,6.990674,6.5266414,5.8173876,4.9723196,4.112161,3.7914882,3.7990334,3.6066296,3.1727777,2.969056,2.8822856,2.9803739,3.0671442,3.0407357,2.867195,2.3163917,2.0372176,1.9806281,2.04099,2.0673985,2.3578906,2.4899325,2.71629,3.1312788,3.663219,3.9688015,4.0103,3.893349,3.651901,3.259548,3.5387223,3.8292143,4.0706625,4.1762958,4.0178456,3.1614597,2.6144292,2.41448,2.4371157,2.4031622,1.9655377,2.003264,2.3956168,2.7728794,2.4974778,2.8785129,2.546522,2.0183544,1.7316349,2.0296721,2.5540671,2.2786655,2.0636258,2.2069857,2.4107075,2.4974778,2.837014,3.1048703,3.4330888,4.4177437,4.957229,5.5004873,6.1720147,7.0774446,8.341274,8.367682,8.98262,9.748463,10.525623,11.4838705,11.287694,11.638548,12.96274,14.532151,14.471789,12.453435,11.080199,9.703192,8.439363,8.182823,8.043237,7.9526935,8.390318,9.1825695,9.495697,9.307066,9.144843,8.846806,8.809079,10.016319,10.072908,9.997457,9.786189,9.507015,9.276885,9.556059,11.18206,12.347801,12.596795,12.815607,12.445889,12.951422,13.826671,14.977322,16.70141,18.621677,19.591242,19.91946,19.757236,19.104572,18.395319,17.014538,15.75071,14.747191,13.536179,13.226823,14.211478,15.599804,16.905132,18.040693,18.372684,18.142553,17.674747,17.169216,16.697638,17.127718,18.414183,19.666695,20.406128,20.557034,2.9464202,2.8596497,2.8030603,3.138824,3.6179473,3.3878171,3.85185,3.7198083,3.5236318,3.4481792,3.3274553,3.289729,2.969056,2.6332922,2.4220252,2.3503454,2.4823873,2.5993385,2.9954643,3.3727267,2.8219235,2.8219235,3.199186,3.6368105,4.0782075,4.7006907,5.0779533,5.6778007,6.700182,7.6886096,7.492433,7.466025,7.7829256,7.3377557,6.217286,5.692891,5.534441,5.300538,4.2630663,2.4861598,0.83752275,0.46026024,0.2565385,0.21881226,0.30181,0.41121614,0.39989826,0.4979865,1.3505998,2.6031113,2.8822856,1.750498,1.5656394,1.5279131,1.4600059,1.7995421,2.1541688,2.2786655,3.2859564,5.142088,6.6662283,7.254758,5.80607,5.1534057,6.300284,8.424272,7.1906233,6.398372,8.888305,13.238141,13.762536,12.445889,10.842525,9.590013,9.525878,11.672502,10.280403,7.84706,5.6476197,4.5799665,5.142088,6.4134626,7.032173,8.326183,9.933322,9.812597,10.506761,10.121953,9.608876,8.6732645,5.7683434,5.9984736,5.2062225,4.13857,3.31991,3.0520537,3.2482302,3.7462165,4.006528,3.953711,3.953711,5.2326307,6.1229706,6.8925858,7.1981683,6.089017,4.074435,3.0935526,2.323937,1.8259505,2.5314314,1.2751472,1.0148361,1.1204696,1.2411937,1.327964,1.2902378,1.50905,1.5241405,1.3694628,1.6033657,1.871222,1.8749946,1.3656902,0.8563859,1.6033657,3.8367596,4.4403796,4.8440504,5.281675,4.8063245,4.9647746,5.0213637,5.0477724,4.9723196,4.5912848,3.7877154,3.3463185,2.7011995,1.8900851,1.5731846,2.0108092,1.9278114,2.5314314,3.5538127,3.2331395,2.516341,2.4823873,2.493705,2.3578906,2.3201644,1.6373192,2.0673985,3.3123648,4.7912335,5.643847,6.9152217,6.5568223,6.696409,7.3981175,6.651138,4.4441524,3.5538127,4.7044635,7.175533,8.7751255,7.699928,6.2851934,4.817642,3.7613072,3.7990334,5.2628117,5.4212623,5.7079816,7.1604424,10.4049,15.214996,17.176762,17.904879,18.651857,20.323132,18.504726,17.354074,19.278114,22.337713,20.247679,19.515789,23.948624,29.984823,37.37917,49.19503,56.189476,69.44648,91.716286,120.73909,149.22618,152.31596,127.884445,101.951416,88.29829,88.45674,70.24251,61.158024,56.098934,51.06248,43.151283,32.50871,29.011486,31.309015,37.145267,43.396507,71.55915,91.37675,82.06214,50.46263,31.067568,26.672459,25.63876,28.09851,32.61057,36.164383,39.325844,41.461147,50.08537,68.35242,95.06261,91.410706,65.572,45.147003,39.042896,37.42821,29.69056,29.192572,32.520027,35.032597,30.882708,34.474247,48.399006,55.710354,48.368824,27.238352,12.113899,5.832478,4.323428,5.028909,6.8963585,7.2623034,13.389046,20.206179,24.525835,25.02382,19.470518,15.501716,12.46098,9.805053,7.0963078,6.6322746,5.873977,5.1043615,4.8440504,5.8437963,4.146115,3.31991,3.8141239,5.191132,6.119198,6.0701537,4.3007927,3.1954134,3.7462165,5.5382137,9.031664,10.570895,10.235131,8.439363,5.934339,7.5226145,8.284684,8.311093,7.454707,5.3571277,4.2706113,4.1989317,4.6214657,5.342037,6.515323,5.5985756,5.764571,6.3644185,6.6360474,5.7079816,7.5490227,11.370691,13.807808,14.249205,14.84528,17.225805,20.92675,25.770802,31.799456,39.246616,43.01924,45.69026,44.101986,38.15633,30.807257,27.094994,22.379211,17.20317,12.996693,12.068627,11.16697,11.627231,12.0724,11.808316,10.819888,10.7557535,10.733118,10.525623,10.687846,12.543978,12.702429,12.098808,10.989656,9.137298,5.828706,6.937857,7.273621,8.126234,9.480607,9.993684,4.9534564,3.2821836,2.4861598,1.6033657,1.1732863,0.8563859,0.63002837,0.5281675,0.5583485,0.7167987,0.76584285,1.5015048,1.8297231,1.5505489,1.3430545,2.7351532,4.9119577,6.700182,6.187105,0.73188925,3.4557245,2.203213,0.76207024,0.42630664,0.0,0.02263575,0.06790725,0.26408374,0.46026024,0.23013012,0.094315626,0.071679875,0.18485862,0.35462674,0.36594462,2.4295704,3.338773,2.837014,1.9089483,2.7615614,3.0407357,2.8106055,2.927557,3.4632697,3.7084904,4.4894238,4.610148,5.4363527,6.2097406,4.074435,2.7804246,3.199186,3.361409,2.686109,1.9542197,1.5241405,1.327964,1.237421,1.2789198,1.6335466,1.0336993,1.1506506,1.6071383,1.9466745,1.6184561,1.0186088,0.63002837,1.1883769,2.7540162,4.7308717,5.1835866,4.8553686,4.274384,3.4745877,1.9844007,1.3958713,0.70170826,0.21503963,0.02263575,0.0,0.071679875,0.32067314,0.5885295,0.7582976,0.73188925,1.3656902,1.6184561,2.0636258,2.897376,3.9197574,3.8593953,4.3309736,5.4401255,6.4474163,5.753253,5.692891,6.307829,7.0170827,7.383027,7.1264887,6.466279,6.319147,5.8626595,4.9760923,4.2404304,4.3649273,4.146115,3.7688525,3.380272,3.1124156,2.8332415,3.108643,3.3764994,3.3764994,3.1576872,2.6332922,2.546522,2.2560298,1.6222287,1.0223814,1.2185578,1.2223305,1.1280149,0.9922004,0.80734175,0.88279426,0.9997456,1.1242423,1.177059,1.0676528,1.0676528,0.98465514,0.8526133,0.7507524,0.8224323,0.9695646,1.1431054,1.4600059,1.7618159,1.6033657,1.2110126,1.5543215,1.901403,1.8787673,1.4637785,1.4298248,1.2449663,1.3355093,1.7769064,2.2899833,2.595566,3.4481792,4.0782075,4.5497856,5.783434,6.0022464,6.4134626,6.428553,5.855114,4.927048,4.9760923,5.2364035,4.5460134,3.1350515,2.6106565,2.7087448,3.1614597,3.6481283,3.904667,3.7084904,3.682082,3.6783094,3.9876647,4.7120085,5.7381625,6.9567204,7.7225633,8.66572,9.903141,11.000975,11.208468,10.9594755,11.050018,11.4838705,11.457462,12.838243,12.332711,11.404645,11.106608,12.068627,11.996947,11.189606,10.642575,10.789707,11.536687,12.121444,12.147853,11.7894535,11.072655,9.88805,9.424017,8.922258,8.2507305,7.61693,7.567886,7.5792036,7.1981683,6.8699503,6.647365,6.19465,5.855114,6.25124,6.6549106,6.7454534,6.620957,6.937857,6.7152724,6.587003,6.9755836,8.088508,8.722309,9.125979,9.854096,11.027383,12.344029,12.97783,13.057055,12.721292,12.140307,11.506506,10.540714,9.95973,9.771099,9.752235,9.446653,9.2995205,8.265821,7.564113,7.2057137,5.9984736,5.617439,4.957229,4.2064767,3.6971724,3.904667,3.4179983,3.1576872,2.848332,2.5804756,2.8219235,2.384299,2.354118,2.5804756,2.7691069,2.4861598,1.9881734,1.7429527,1.7957695,2.0447628,2.2296214,2.6446102,2.9011486,3.1161883,3.3689542,3.7235808,3.6481283,3.6330378,3.7235808,3.7235808,3.1727777,3.4066803,3.6745367,3.9386206,3.9688015,3.3727267,2.505023,2.5540671,2.674791,2.425798,1.7542707,1.9127209,2.1353056,2.4031622,2.6898816,2.9615107,2.7653341,2.1956677,1.5430037,1.81086,4.715781,4.6554193,3.5500402,2.463524,1.9844007,2.2296214,2.6182017,2.6144292,3.218049,4.406426,5.1269975,4.8327327,4.7346444,5.4174895,6.960493,8.926031,10.084227,10.604849,11.038701,11.434827,11.336739,11.042474,11.393328,12.611885,13.8719425,13.275867,11.529142,10.453944,9.4013815,8.390318,8.073418,8.303548,8.262049,8.52236,9.21275,9.993684,9.797507,9.574923,9.435335,9.431562,9.552286,9.639057,9.465516,9.156161,8.948667,9.216523,10.069136,11.299012,11.978085,11.951676,11.84227,12.377983,12.604341,13.475817,15.079182,16.618414,18.448135,19.270569,19.270569,18.983849,19.28566,18.13878,16.376965,15.022593,14.377474,14.022847,15.218769,16.644821,17.803017,18.470772,18.678267,18.629223,18.029375,17.346529,16.920223,16.969267,17.640795,18.840488,19.61765,19.787418,19.957186,2.6031113,2.7125173,2.8294687,3.0256453,3.1765501,2.9351022,3.0105548,3.350091,3.4179983,3.0671442,2.546522,3.229367,3.1652324,2.8106055,2.6446102,3.1539145,3.1350515,2.938875,2.71629,2.6106565,2.7728794,3.1954134,3.2784111,3.4934506,3.9725742,4.515832,4.8553686,5.342037,6.1908774,7.17176,7.6018395,7.488661,6.9755836,6.258785,5.4891696,4.7874613,4.406426,4.3083377,3.9989824,3.097325,1.3505998,0.6111652,0.36971724,0.29803738,0.2565385,0.27917424,0.392353,0.573439,1.1732863,2.1466236,3.0407357,2.5314314,2.233394,2.3201644,2.5540671,2.2899833,2.0258996,2.4522061,3.1765501,4.085753,5.3382645,4.919503,4.587512,4.919503,5.583485,5.383536,5.010046,4.7006907,5.4476705,7.0284004,8.001738,9.476834,8.952439,7.8810134,7.1076255,6.862405,6.4210076,6.300284,6.760544,7.4282985,7.3151197,7.8810134,8.597813,9.80128,11.246195,12.079946,11.59705,10.227587,7.8244243,5.2665844,4.4630156,4.6629643,4.4139714,4.3913355,4.779916,5.27413,5.7607985,4.983638,4.3686996,4.29702,4.112161,5.0515447,7.0472636,9.242931,9.914458,6.4926877,4.82896,3.731126,2.9615107,2.3805263,1.9466745,1.1091517,0.9393836,0.97710985,0.97710985,0.9242931,0.8601585,1.2185578,1.2789198,0.995973,0.9922004,1.1129243,1.086516,0.8978847,0.87147635,1.6750455,3.440634,4.353609,5.194905,5.9532022,5.80607,6.006019,5.723072,5.3080835,4.9232755,4.557331,3.9574835,3.3123648,2.5729303,2.0372176,2.3654358,2.41448,2.203213,2.4031622,2.7691069,2.1503963,1.2826926,1.2789198,1.3430545,1.1581959,0.87902164,1.1506506,2.7125173,4.4101987,5.4363527,5.3156285,5.111907,4.961002,4.666737,4.349837,4.4441524,3.531177,3.85185,4.9760923,6.858632,9.835234,9.133525,7.01331,5.1873593,4.432834,4.617693,5.66271,6.900131,7.624475,8.348819,10.785934,15.8676605,18.557543,19.768555,19.983595,19.263023,18.919714,19.50447,19.945868,19.945868,20.017548,21.752956,25.080412,31.376923,40.374634,50.17214,55.74808,65.97944,82.616714,102.879486,119.44885,127.79012,114.45013,97.145096,85.43109,80.66627,70.36323,60.252594,49.877876,40.14073,33.31228,29.788647,30.233816,34.798695,40.91412,43.287098,55.9518,79.17608,83.28824,63.00284,37.42444,31.048704,28.890762,30.07914,33.27078,36.628418,40.695305,44.577335,50.07405,63.859222,97.44313,95.168236,68.26565,46.889957,39.774784,34.20639,28.724768,27.977787,30.73935,33.595226,30.95816,31.569326,39.36357,41.5781,32.942562,15.690348,13.962485,11.363147,8.013056,5.247721,5.59103,8.484633,10.850069,13.819125,17.482344,20.862616,15.739391,12.54775,10.7557535,9.567377,7.9489207,7.7678347,5.9418845,4.647874,4.406426,4.0480266,2.927557,2.7011995,2.938875,3.4179983,4.093298,4.032936,3.361409,3.0860074,3.5274043,4.304565,8.246958,10.265312,10.329447,8.869441,6.7643166,6.4964604,6.0362,5.8400235,5.956975,6.013564,4.7044635,4.817642,5.583485,6.832224,9.031664,7.8998766,7.4169807,7.4018903,7.5905213,7.647111,8.669493,9.510788,11.027383,12.653384,12.381755,14.966003,17.165443,21.503962,26.800728,28.173964,33.606544,35.639988,34.587425,31.497646,28.17019,26.940315,22.447119,17.923742,14.841507,12.898605,11.449917,11.34051,11.879996,12.355347,12.049765,10.691619,10.502988,10.163452,9.948412,11.725319,12.253486,11.898859,13.298503,14.071891,6.828451,7.4999785,7.0849895,7.405663,8.016829,6.2361493,4.485651,3.3727267,2.4710693,1.6410918,1.0299267,0.7997965,0.6526641,0.55457586,0.59230214,0.98465514,1.4939595,1.4373702,4.1272516,7.1378064,2.282438,2.1881225,4.5233774,5.4363527,4.0103,2.293756,1.5618668,2.8709676,2.4408884,0.25276586,0.060362,0.094315626,0.482896,2.3163917,5.0968165,6.760544,6.138061,5.938112,7.0359454,8.537451,7.786698,6.043745,16.750456,24.56356,25.25018,25.68403,32.712433,34.542156,29.724512,20.368402,12.106354,14.252977,11.936585,9.137298,7.3075747,5.3684454,3.682082,3.2784111,2.897376,2.3277097,2.4182527,1.7731338,1.2751472,1.3392819,1.7655885,1.7316349,1.4071891,1.3694628,1.4373702,1.4600059,1.3241913,1.2826926,1.0035182,1.7165444,3.3236825,4.4139714,5.9682927,5.6551647,4.06689,2.0372176,0.6149379,1.2223305,0.9393836,0.452715,0.14713238,0.120724,0.32067314,0.49044126,0.90543,1.3807807,1.2713746,1.5430037,1.841041,2.1994405,2.8747404,4.3611546,5.753253,5.5570765,5.281675,5.4363527,5.534441,7.3075747,7.8998766,7.7037,7.3717093,7.809334,8.0206,7.673519,6.379509,4.776143,4.5233774,4.7120085,4.644101,4.29702,3.8895764,3.893349,3.572676,3.4745877,3.482133,3.4481792,3.2067313,2.9766011,2.6332922,2.1315331,1.5656394,1.1808317,1.1506506,1.20724,1.1016065,0.87147635,0.8337501,0.90543,0.9393836,1.026154,1.1129243,0.9808825,1.0601076,1.086516,1.0110635,0.875249,0.8111144,0.8978847,1.0751982,1.4675511,1.8184053,1.4449154,1.3845534,1.4939595,1.6033657,1.5543215,1.20724,1.3958713,1.4600059,1.5128226,1.690136,2.1541688,2.214531,2.505023,3.0143273,3.9499383,5.7079816,6.9152217,7.352846,7.322665,6.9755836,6.330465,5.745708,5.5683947,5.3910813,4.7950063,3.3538637,3.127506,3.531177,3.893349,3.8820312,3.5123138,4.014073,4.45547,4.9987283,5.5080323,5.564622,6.319147,7.3000293,8.050782,8.624221,9.58624,10.095545,9.944639,10.250222,11.016065,11.129244,11.668729,11.744182,11.910177,12.0724,11.4838705,10.921749,10.435081,10.344538,10.540714,10.484125,11.004747,10.902886,10.412445,9.684328,8.812852,8.341274,8.231868,7.907422,7.4396167,7.5565677,7.0812173,6.417235,6.138061,6.1078796,5.451443,5.2250857,5.5306683,5.8588867,5.9607477,5.828706,5.794752,5.836251,6.405917,7.3113475,7.707473,8.488406,9.2844305,10.231359,11.246195,12.027128,12.181807,12.585477,12.464753,11.872451,11.676274,10.789707,9.774872,9.307066,9.439108,9.590013,9.231613,8.873214,7.964011,6.5643673,5.3759904,4.164978,3.4481792,3.1539145,2.9916916,2.4672968,2.6332922,2.5804756,2.41448,2.2598023,2.2484846,2.0145817,2.003264,2.233394,2.4559789,2.1466236,1.9579924,2.0108092,2.142851,2.1994405,2.033445,2.233394,2.5540671,2.7653341,2.8822856,3.199186,3.350091,3.270866,3.0633714,2.9237845,3.1237335,3.1237335,3.150142,3.350091,3.4179983,2.6144292,2.2258487,2.191895,2.2447119,2.1805773,1.8523588,1.9994912,2.4107075,2.7540162,2.7691069,2.2748928,1.991946,1.5845025,1.991946,3.651901,6.4964604,6.398372,4.1762958,2.6710186,2.6672459,2.9124665,2.8822856,3.029418,3.561358,4.508287,5.726845,5.5306683,5.7381625,6.4436436,7.677292,9.439108,9.533423,10.103089,11.257513,12.449662,12.46098,11.6875925,12.702429,13.570132,13.494679,12.800517,11.034928,9.725827,8.631766,7.907422,8.107371,8.182823,8.337502,8.52236,8.733627,9.016574,9.631512,9.688101,9.627739,9.593785,9.393836,9.291975,9.529651,9.559832,9.484379,10.0465,11.729091,12.045992,11.46878,10.902886,11.68382,12.668475,13.8719425,15.211224,16.576914,17.814335,18.94235,19.289433,19.48561,19.53088,18.810308,16.98813,15.418718,14.890551,15.369675,16.01102,16.886269,17.784155,18.991394,20.213724,20.557034,20.017548,19.83269,19.319613,18.406637,17.625704,18.297232,18.885761,19.349794,19.696875,19.994913,2.372981,2.3390274,2.3465726,2.516341,2.8106055,3.0407357,3.2218218,3.6481283,3.7235808,3.3878171,3.1010978,3.1614597,3.2633207,3.1463692,2.9766011,3.3576362,3.199186,3.0218725,2.7389257,2.4031622,2.203213,2.6182017,2.867195,3.2218218,3.7763977,4.432834,4.7120085,4.9421387,5.6325293,6.63982,7.1906233,7.1302614,6.1795597,5.2137675,4.659192,4.508287,4.0517993,3.9461658,4.036709,3.7084904,1.901403,0.7696155,0.40367088,0.35085413,0.331991,0.23390275,0.44139713,0.633801,0.8941121,1.3505998,2.1956677,2.916239,2.6408374,2.6597006,3.2746384,3.783943,2.6672459,2.9841464,3.6556737,4.055572,4.025391,3.5651307,3.9273026,4.7346444,5.5306683,5.7683434,4.9723196,4.3611546,4.191386,4.6856003,6.058836,6.3908267,5.5382137,5.062863,5.4665337,6.145606,6.1720147,8.473316,9.748463,9.167479,8.345046,9.465516,10.114408,10.578441,10.702937,9.865415,8.639311,7.6810646,6.1531515,4.236658,3.138824,3.7047176,3.610402,3.62172,3.8971217,3.9801195,4.8327327,4.4177437,3.9574835,3.9197574,4.002755,4.6818275,7.4282985,8.82417,7.5565677,4.4403796,3.5236318,2.8445592,2.2748928,1.7580433,1.2789198,0.9922004,0.84884065,0.8224323,0.8978847,1.0525624,1.1619685,1.1808317,0.98465514,0.7092535,0.72811663,0.72811663,0.62625575,0.482896,0.482896,0.94315624,2.1881225,3.229367,4.1498876,4.8025517,4.821415,5.2628117,5.292993,5.149633,4.90064,4.45547,3.9574835,3.2482302,2.4295704,1.8448136,2.0673985,2.0145817,1.7957695,1.841041,2.0447628,1.7957695,0.98465514,0.754525,0.68661773,0.68661773,0.95824677,1.8297231,2.9539654,3.8820312,4.357382,4.2894745,3.9574835,3.7499893,3.5575855,3.4330888,3.6066296,3.2331395,3.3764994,3.783943,4.6252384,6.4926877,6.930312,6.40969,5.824933,5.281675,4.08198,5.2250857,6.722818,8.390318,9.952185,11.042474,14.203933,16.939087,18.104828,18.202915,19.379974,20.334448,20.228815,19.662922,20.096773,23.850534,23.356321,24.27307,28.438047,36.194565,46.414604,50.854984,57.989017,67.2244,77.78398,88.7095,97.66949,94.21754,85.72536,77.38409,72.211815,67.167816,60.70908,51.56424,41.00089,32.81052,30.633715,32.716206,38.322327,45.033825,48.74986,52.779022,74.294304,86.86469,77.04077,44.373615,33.851765,30.577126,31.278833,33.94608,37.79416,41.483784,45.520493,51.975456,64.98347,90.74295,94.662704,75.74299,55.672626,42.890972,32.55021,28.611588,26.012249,26.819592,29.607561,29.437794,30.02255,33.323597,32.9652,26.283878,14.351066,20.828663,15.882751,8.518587,4.327201,5.485397,7.7829256,8.182823,9.439108,12.498707,16.490145,14.071891,12.030901,10.623712,9.450426,7.4509344,6.7454534,5.062863,4.036709,3.742444,2.6936543,2.625747,2.5917933,3.2670932,4.164978,3.640583,3.6443558,3.4783602,3.2670932,3.3350005,4.191386,6.937857,8.416726,8.612903,7.8621507,6.862405,6.4738245,6.043745,5.915476,5.987156,5.7117543,5.8626595,6.417235,7.2660756,8.733627,11.581959,10.220041,9.529651,9.110889,8.710991,8.186596,8.771353,9.06939,9.590013,10.216269,10.216269,13.211733,14.943368,18.648085,23.518545,24.69183,31.358059,32.052223,30.479038,28.864353,27.958923,26.24238,23.231825,20.643805,18.640541,15.833707,13.822898,11.815862,11.11038,11.91395,13.309821,11.114153,10.846297,10.442626,9.665465,10.084227,10.887795,11.7894535,14.011529,15.120681,9.039209,8.326183,6.8397694,6.387054,6.851087,6.2097406,4.3083377,3.531177,2.8936033,2.0485353,1.3015556,1.0374719,0.76584285,1.1657411,1.9051756,1.6486372,1.448688,1.3845534,2.9237845,4.859141,3.2859564,3.519859,4.266839,4.817642,4.727099,3.783943,1.6712729,2.4371157,3.029418,2.3277097,1.146878,0.59230214,2.1164427,6.749226,13.094781,17.316349,17.810562,17.72002,17.512526,17.708702,18.87067,15.411173,23.16769,32.659615,37.545162,34.632698,39.948326,40.81603,37.239582,30.505445,23.186554,20.455173,15.807299,11.306557,7.8621507,5.2250857,3.3048196,2.4484336,2.1466236,2.1353056,2.4031622,2.0598533,1.7844516,1.9730829,2.354118,1.9844007,2.8634224,3.0218725,2.4974778,1.81086,1.9844007,1.297783,1.3468271,2.2748928,4.1762958,7.0812173,8.126234,7.624475,4.82896,1.2600567,0.7130261,1.3958713,1.1280149,0.5772116,0.211267,0.29049212,0.3961256,0.47912338,0.70170826,1.0487897,1.3015556,1.5430037,2.1013522,2.7540162,3.5123138,4.5988297,6.4964604,6.7680893,6.888813,7.1000805,6.4021444,7.8017883,8.514814,8.529905,8.14887,7.99042,8.3525915,8.469543,7.4773426,5.907931,5.692891,5.160951,5.1345425,4.9421387,4.5309224,4.5120597,3.9612563,3.5990841,3.531177,3.62172,3.4934506,3.4142256,2.957738,2.2975287,1.6561824,1.3128735,1.1317875,1.1016065,1.0186088,0.88279426,0.91297525,0.9922004,0.95824677,0.98465514,1.0638802,1.026154,0.9922004,0.9280658,0.86770374,0.8186596,0.7809334,0.76584285,1.1317875,1.5052774,1.6260014,1.3770081,1.3505998,1.2562841,1.1959221,1.1657411,1.0638802,1.3505998,1.4750963,1.5316857,1.6524098,1.991946,2.1692593,2.6332922,3.3236825,4.3422914,5.956975,7.0887623,7.326438,6.9793563,6.304056,5.50426,5.379763,5.511805,5.621211,5.1798143,3.410453,3.4859054,3.874486,4.123479,4.074435,3.8480775,4.22534,4.6214657,5.0515447,5.3759904,5.292993,5.270357,6.0814714,7.118943,8.175279,9.461743,10.03141,10.31813,10.729345,11.242422,11.404645,11.3820095,11.00852,11.52537,12.37421,11.200924,10.831206,10.412445,10.257768,10.359629,10.397354,10.269085,9.914458,9.442881,8.89585,8.231868,7.7942433,7.3868,6.8661776,6.3644185,6.2814207,6.2399216,5.753253,5.349582,5.1081343,4.640329,4.7044635,4.9723196,5.2628117,5.4174895,5.281675,5.270357,5.3156285,5.983383,7.0585814,7.541477,8.028146,8.646856,9.461743,10.480352,11.646093,12.012038,12.215759,12.053536,11.623458,11.32542,10.699164,9.593785,8.956212,9.061845,9.491924,9.156161,8.643084,7.488661,5.8400235,4.459243,3.3727267,2.757789,2.584248,2.5616124,2.123988,2.0862615,2.1051247,2.082489,2.04099,2.1164427,1.931584,1.9127209,1.9579924,1.9466745,1.7316349,1.7882242,2.0070364,2.0636258,1.8900851,1.7014539,1.6939086,1.7995421,1.9994912,2.2560298,2.516341,2.5917933,2.3503454,2.1466236,2.1956677,2.565385,2.6785638,2.8219235,2.9916916,2.9766011,2.335255,2.4031622,2.4069347,2.214531,1.9051756,1.7957695,1.8297231,1.9542197,2.0862615,2.0900342,1.7580433,1.4147344,1.5580941,2.444661,3.9159849,5.413717,5.2326307,3.7914882,2.7992878,2.7841973,3.0633714,2.9237845,3.2935016,3.7613072,4.3913355,5.726845,6.1342883,6.1041074,6.692637,8.080963,9.58624,9.574923,10.4049,11.932813,13.302276,12.951422,12.506252,12.928786,13.019329,12.393073,11.491416,10.650121,9.273112,8.22055,7.865923,8.107371,8.167733,8.122461,7.960239,8.039464,9.076936,9.880505,9.839006,9.390063,8.812852,8.209232,8.371455,9.024119,9.476834,9.733373,10.499215,11.778135,11.774363,11.1782875,10.8576145,11.853588,12.928786,14.607604,16.365646,17.886015,19.04421,19.289433,19.153618,18.97253,18.617905,17.512526,16.260014,15.07541,15.135772,16.429781,17.784155,18.09351,18.519815,19.515789,20.832436,21.503962,21.296469,20.99843,20.315586,19.391293,18.791445,18.780127,18.76881,18.893307,19.032892,18.806536,2.2673476,2.2484846,2.1881225,2.4484336,3.1199608,4.006528,4.1008434,4.4215164,4.508287,4.1574326,3.440634,2.8181508,2.7841973,2.8030603,2.7728794,3.0256453,2.8747404,2.7540162,2.5012503,2.1051247,1.7278622,2.04099,2.4182527,2.8445592,3.338773,3.9763467,4.504514,4.7044635,5.379763,6.4474163,6.9265394,6.8133607,5.9796104,5.0515447,4.4894238,4.561104,4.195159,4.164978,4.3422914,4.0706625,2.1692593,0.8186596,0.3734899,0.31312788,0.30935526,0.19994913,0.3734899,0.482896,0.6149379,0.9620194,1.8221779,3.2067313,3.3010468,3.380272,3.9612563,4.7836885,4.1008434,4.2328854,4.236658,3.7575345,3.0256453,2.848332,3.6066296,4.6554193,5.583485,6.19465,4.768598,3.8858037,3.4632697,3.5953116,4.561104,4.0706625,3.8292143,4.195159,5.2364035,6.7379084,7.8508325,9.578695,9.58624,8.194141,8.356364,10.080454,11.314102,11.404645,9.978593,6.9491754,5.5985756,5.342037,4.983638,4.1272516,3.199186,3.6028569,3.6292653,3.4029078,3.0558262,2.7351532,3.9348478,3.7877154,3.6141748,3.9499383,4.534695,4.561104,7.0812173,7.4584794,4.9534564,2.7691069,2.293756,1.8863125,1.4637785,1.0676528,0.8639311,0.84129536,0.72811663,0.7167987,0.8526133,1.0450171,1.2147852,1.1506506,0.98465514,0.9318384,1.2713746,1.4373702,1.1355602,0.8262049,0.7696155,1.0336993,1.5656394,2.1956677,2.7653341,3.259548,3.8141239,4.5120597,4.821415,4.825187,4.5120597,3.772625,3.3878171,2.7917426,2.1466236,1.6825907,1.720317,1.6410918,1.4713237,1.3807807,1.3694628,1.2562841,0.724344,0.41498876,0.3169005,0.5470306,1.3430545,2.2786655,2.8407867,3.138824,3.31991,3.5689032,3.2331395,2.8143783,2.674791,2.9011486,3.31991,3.3236825,3.0860074,2.9615107,3.1765501,3.8405323,4.3686996,4.776143,4.983638,4.7044635,3.4632697,4.719554,6.405917,8.186596,9.593785,10.03141,11.98563,15.124454,17.022083,17.976559,21.028612,21.696367,21.511507,20.081682,19.553514,24.631468,22.39053,22.560297,25.744392,32.138992,41.551693,47.07104,51.903774,56.81196,63.232967,73.28324,79.4628,79.54957,75.77317,70.43868,65.9304,61.39947,58.068245,53.122334,45.622353,36.485058,34.07435,36.179474,41.310246,47.674664,53.22042,54.352207,72.0345,90.648636,91.75778,54.088123,36.50769,31.859818,32.4823,34.40634,37.345215,40.793396,45.705353,53.846676,66.05866,82.228134,90.414734,79.62502,62.08609,45.407314,32.561527,29.366114,25.619896,25.276588,27.758974,27.95515,27.181763,27.415667,26.574371,23.499681,17.961468,23.876944,17.818108,9.820143,5.330719,5.240176,6.296511,6.3644185,7.111398,9.35611,13.057055,13.166461,12.249713,10.933067,9.25425,6.6813188,5.4174895,4.2404304,3.482133,2.9803739,2.0673985,2.8407867,2.806833,3.6594462,4.9760923,4.195159,4.255521,4.236658,3.85185,3.4632697,4.093298,5.560849,6.6322746,7.001992,6.960493,7.383027,7.145352,6.730363,6.719045,7.0170827,6.858632,8.224322,8.684583,9.325929,11.038701,14.48688,13.087236,11.996947,10.963248,10.012547,9.431562,8.620448,8.669493,8.892077,9.035437,9.2844305,11.3820095,13.2607765,17.04472,21.681276,22.941332,31.120384,30.731804,28.230553,27.038403,27.570343,27.053493,25.318087,23.643042,22.066084,19.379974,16.052519,12.2119875,10.325675,11.231105,14.128481,11.830952,11.065109,10.646348,10.001229,9.178797,9.88805,11.223559,13.385274,14.596286,11.102836,9.061845,6.862405,5.8702044,6.1908774,6.692637,4.5497856,3.7990334,3.2670932,2.4672968,1.5769572,1.2449663,1.2147852,1.7165444,2.3088465,1.9051756,1.6071383,1.9730829,2.2484846,2.5201135,3.7009451,3.9688015,3.7198083,3.9763467,4.5761943,4.187614,2.5502944,2.9464202,3.7990334,4.29702,4.3686996,2.7389257,5.80607,12.253486,20.126955,26.827137,29.27557,29.328386,27.559025,25.985842,28.057013,26.883726,30.686531,35.534355,37.50744,32.735065,38.295918,40.521767,38.20537,32.316307,26.00093,20.975796,15.811071,11.314102,7.8621507,5.4438977,3.6556737,2.7653341,2.5012503,2.546522,2.5389767,2.3163917,2.3692086,2.795515,3.199186,2.7087448,3.9273026,4.183841,3.8103511,3.3274553,3.429316,1.5241405,1.569412,2.8294687,5.05909,8.507269,9.175024,7.9036493,4.6026025,1.1204696,1.2261031,1.4901869,1.297783,0.8224323,0.3734899,0.39989826,0.58098423,0.7394345,0.995973,1.4147344,2.0296721,2.2409391,2.9086938,3.9310753,5.0779533,5.983383,7.383027,7.8395147,8.412953,8.843033,7.5603404,7.745199,8.329956,8.744945,8.75249,8.439363,8.68081,8.944894,8.186596,6.7152724,6.198423,5.5683947,5.6363015,5.5797124,5.2326307,5.1081343,4.5196047,3.8367596,3.5764484,3.7462165,3.8405323,3.7047176,3.2784111,2.5389767,1.7429527,1.4298248,1.1581959,1.0223814,0.9393836,0.8865669,0.90543,1.0072908,1.0035182,0.98842776,0.9922004,1.0072908,0.9808825,0.86770374,0.80356914,0.8262049,0.86770374,0.80734175,1.1732863,1.4411428,1.4600059,1.4449154,1.2638294,1.0487897,0.9280658,0.9280658,0.97710985,1.2751472,1.4411428,1.569412,1.7580433,2.1164427,2.384299,3.0143273,3.874486,4.930821,6.224831,7.092535,7.092535,6.598321,5.8702044,5.070408,5.379763,5.881522,5.926794,5.142088,3.440634,3.5085413,3.8480775,4.13857,4.2592936,4.323428,4.398881,4.5422406,4.7572803,4.9647746,5.0251365,4.6252384,5.3344917,6.79827,8.439363,9.454198,10.080454,10.631257,11.117926,11.566868,12.015811,11.408418,10.54826,10.842525,11.815862,11.144334,11.0613365,10.665211,10.525623,10.763299,11.050018,10.397354,9.650374,9.065618,8.707218,8.439363,8.062099,7.1906233,6.2814207,5.613666,5.311856,5.4288073,5.081726,4.5912848,4.1800685,3.953711,4.112161,4.395108,4.6327834,4.727099,4.666737,4.7610526,4.90064,5.4250345,6.2814207,7.0284004,7.496206,8.054554,8.763808,9.703192,10.948157,11.393328,11.627231,11.680047,11.502733,10.978339,10.306811,9.310839,8.748717,8.733627,8.733627,8.507269,7.8131065,6.8246784,5.6098933,4.134797,3.429316,2.8521044,2.4861598,2.3201644,2.2409391,1.9240388,1.8184053,1.8636768,1.9693103,1.9994912,1.9051756,1.8900851,1.8146327,1.6675003,1.5731846,1.6939086,1.8523588,1.7957695,1.5467763,1.3958713,1.3053282,1.2713746,1.3732355,1.599593,1.841041,1.780679,1.5580941,1.50905,1.7240896,2.033445,2.173032,2.3918443,2.5427492,2.5012503,2.1956677,2.5540671,2.5238862,2.1692593,1.8070874,1.9768555,1.8184053,1.5316857,1.388326,1.3920987,1.2449663,1.1242423,1.5128226,2.4899325,3.772625,4.7120085,4.025391,3.2972744,2.8106055,2.6974268,2.9351022,2.7540162,3.2859564,3.9876647,4.7233267,5.7419353,6.205968,6.4247804,7.1981683,8.560086,9.786189,10.114408,11.16697,12.645839,13.754991,13.20796,12.872196,12.694883,12.178034,11.268831,10.359629,10.174769,9.276885,8.416726,7.9262853,7.7225633,7.7829256,7.5188417,7.2057137,7.405663,8.937348,9.846551,9.597558,8.907167,8.239413,7.8131065,7.8923316,8.190369,8.405409,8.677037,9.556059,10.593531,10.657665,10.544487,10.887795,12.132762,13.181552,14.618922,16.275105,17.969013,19.508244,19.821371,19.353567,18.76881,18.13878,16.969267,16.109108,15.471535,15.897841,17.206944,18.199142,18.1086,18.474545,19.549744,20.915434,21.477554,21.375692,20.889025,20.334448,19.885506,19.613878,19.149845,18.715992,18.391546,18.131235,17.761518,2.3578906,2.637065,2.7653341,3.31991,4.3686996,5.455216,5.4703064,5.6513925,5.6023483,4.938366,3.2972744,2.5691576,2.1315331,1.9164935,1.9693103,2.4371157,2.3918443,2.2183034,1.9202662,1.6109109,1.5128226,1.7391801,2.0296721,2.335255,2.6785638,3.1312788,4.0970707,4.5422406,5.27413,6.300284,6.8473144,6.485142,6.187105,5.5683947,4.817642,4.7006907,4.4177437,4.4215164,4.4743333,4.044254,2.2862108,0.8601585,0.35839936,0.23013012,0.18485862,0.16222288,0.23767537,0.271629,0.513077,1.1091517,2.0900342,3.7273536,4.568649,4.7950063,4.779916,5.100589,5.80607,5.553304,4.4441524,3.0709167,2.5012503,2.463524,3.2255943,4.191386,4.919503,5.1534057,3.7763977,3.0897799,2.7992878,2.7615614,2.9615107,3.2972744,4.4630156,5.5004873,6.3116016,7.6508837,9.81637,9.152389,7.4999785,6.741681,8.790216,10.423763,11.732863,11.25374,8.718536,5.0741806,4.406426,4.4403796,4.376245,4.1008434,4.22534,4.429062,4.402653,3.8895764,3.0935526,2.6785638,3.7160356,3.5047686,3.519859,4.2706113,5.311856,5.010046,6.085244,5.7683434,3.7877154,2.3880715,1.8561316,1.5015048,1.1657411,0.87147635,0.7884786,0.72811663,0.724344,0.79602385,0.90543,0.9507015,0.9997456,1.1431054,1.2789198,1.539231,2.3126192,2.8256962,2.282438,1.7731338,1.7919968,2.2258487,2.082489,2.0636258,2.1315331,2.5087957,3.6745367,4.349837,4.5422406,4.315883,3.7009451,2.7389257,2.444661,2.082489,1.81086,1.7014539,1.7655885,1.6410918,1.5279131,1.2751472,0.87902164,0.47912338,0.29426476,0.13958712,0.15845025,0.5470306,1.5430037,2.1579416,2.5427492,2.71629,2.8332415,3.199186,2.6295197,2.003264,1.7014539,1.9202662,2.6898816,3.2067313,3.1010978,3.0105548,3.150142,3.3048196,3.0218725,3.259548,3.4444065,3.4330888,3.5123138,4.6516466,6.4549613,7.575431,7.907422,8.601585,10.650121,14.249205,17.37671,19.723284,22.703657,22.398075,23.126192,21.19838,18.433046,22.137764,21.104065,22.137764,25.661396,31.282606,37.805473,44.803696,48.625362,53.197784,60.731716,71.721375,74.8602,75.11674,72.95125,68.907,63.63664,56.396973,53.57882,52.49608,49.874104,41.861046,39.57861,40.94807,44.645245,49.651516,55.26141,56.03857,69.55212,92.716034,104.99216,68.390144,41.06502,33.708405,34.36484,36.14552,37.254673,40.408585,46.184475,54.55593,64.82879,75.663765,84.65016,78.37251,62.99152,45.45636,33.489594,29.79242,25.966978,25.608578,27.672205,26.464964,23.548725,22.515026,22.424482,22.239624,20.817345,20.255224,16.576914,12.283667,8.469543,4.8100967,4.8553686,5.4250345,6.043745,7.17176,10.201178,11.551778,11.317875,10.106862,8.280911,5.987156,4.5950575,3.783943,3.0897799,2.4408884,2.1353056,2.957738,3.0181,4.172523,5.907931,5.3344917,5.198677,4.8327327,4.395108,4.0480266,3.9688015,4.6629643,5.73439,6.349328,6.760544,8.311093,8.167733,7.5792036,7.5603404,8.29223,9.125979,10.480352,10.650121,11.351829,13.656902,17.99542,16.72782,15.520579,13.819125,12.185578,12.30253,9.378746,8.820397,9.4127,10.140816,10.178542,9.933322,12.215759,16.731592,20.96825,20.217497,28.041922,27.615616,25.348267,24.740875,26.393284,29.622652,28.841719,26.612097,24.235344,21.768045,16.761772,12.140307,9.933322,10.7557535,13.7851715,12.174261,10.989656,10.718028,10.691619,9.107117,9.431562,10.140816,11.879996,13.588995,12.50248,9.948412,7.624475,6.360646,6.1833324,6.319147,5.028909,4.0895257,3.3689542,2.6521554,1.6637276,1.297783,1.7316349,1.9240388,1.7769064,2.1541688,3.0558262,3.8556228,3.7084904,2.9652832,3.187868,2.7389257,2.7502437,2.6974268,2.6936543,3.4745877,3.470815,5.300538,5.8966126,5.6325293,8.322411,6.1606965,10.076681,16.35433,23.258234,31.041159,35.209908,35.345722,32.976517,31.02984,33.80649,35.775803,37.967697,35.922935,30.275316,26.725275,35.911617,40.699078,37.31126,27.777838,19.960958,17.01831,13.283413,9.906913,7.5037513,6.138061,4.7421894,4.085753,3.8405323,3.7235808,3.470815,3.0558262,3.2029586,3.8443048,4.5007415,4.274384,5.010046,5.13077,5.3646727,5.666483,5.2288585,1.8485862,1.6637276,3.5160866,6.1305156,8.122461,8.59404,5.9682927,3.0256453,1.3996439,1.5731846,1.4524606,1.5731846,1.388326,0.8639311,0.49421388,1.0374719,1.5015048,2.161714,3.0633714,4.014073,4.2064767,4.678055,5.772116,7.2887115,8.469543,9.208978,9.21275,9.522105,9.88805,8.744945,8.054554,8.031919,8.416726,8.903395,9.152389,9.114662,9.031664,8.182823,6.809588,6.1003346,6.058836,6.217286,6.19465,5.9494295,5.802297,5.3382645,4.293247,3.682082,3.7650797,4.0782075,3.832987,3.4632697,2.7313805,1.8599042,1.5316857,1.2147852,1.0223814,0.94315624,0.9242931,0.8941121,0.965792,1.0223814,0.9997456,0.9318384,0.9205205,1.0299267,0.98842776,0.94692886,0.9620194,0.98465514,0.97333723,1.1883769,1.3355093,1.358145,1.4524606,1.1393328,0.9318384,0.8186596,0.80356914,0.8941121,1.2411937,1.4901869,1.7052265,1.9693103,2.3880715,2.655928,3.1765501,4.025391,5.13077,6.2663302,7.111398,6.900131,6.3908267,5.926794,5.4438977,5.8437963,6.4511886,6.2625575,5.1345425,3.7763977,3.4142256,3.62172,3.9348478,4.191386,4.534695,4.504514,4.5460134,4.640329,4.749735,4.7950063,4.6252384,5.523123,7.303802,9.110889,9.4127,10.11818,10.650121,11.133017,11.664956,12.336484,11.408418,10.601076,10.529396,11.038701,11.200924,11.136789,10.782163,10.827434,11.34051,11.778135,10.895341,9.718282,8.907167,8.688355,8.843033,8.567632,7.4811153,6.296511,5.451443,5.081726,4.878004,4.4516973,3.9499383,3.5538127,3.440634,3.4330888,3.6896272,3.8820312,3.9273026,3.9688015,4.0895257,4.4215164,4.7950063,5.2665844,6.1078796,6.888813,7.6584287,8.461998,9.25425,9.895596,10.0276375,10.397354,10.868933,11.133017,10.733118,9.812597,8.9788475,8.529905,8.265821,7.4697976,7.4207535,6.862405,6.330465,5.7381625,4.3875628,3.9688015,3.4670424,2.8747404,2.3918443,2.4220252,2.0598533,1.7391801,1.7429527,1.9655377,1.9051756,1.9542197,1.9693103,1.8825399,1.7278622,1.6486372,1.6939086,1.659955,1.5241405,1.3241913,1.1317875,1.0676528,1.0751982,1.0525624,1.0525624,1.3015556,1.2298758,1.2487389,1.3619176,1.5543215,1.7844516,1.7919968,1.8825399,1.961765,1.9957186,2.003264,2.3126192,2.173032,1.9127209,1.8259505,2.1466236,1.8070874,1.327964,1.086516,1.0789708,0.91674787,1.0525624,1.3732355,2.1579416,3.3463185,4.5309224,3.572676,2.9766011,2.6408374,2.5201135,2.6483827,2.5691576,3.1614597,4.266839,5.481624,6.1606965,6.096562,6.9454026,8.0206,8.99771,9.910686,10.774617,12.113899,13.324911,13.822898,13.057055,12.50248,12.166716,11.480098,10.453944,9.688101,9.6051035,9.416472,8.741172,7.707473,6.94163,6.9944468,6.7831798,6.6586833,6.9755836,8.107371,9.065618,8.7600355,8.307321,8.213005,8.3525915,7.835742,7.1906233,6.6850915,6.6586833,7.5565677,8.8618965,9.246704,9.684328,10.665211,12.181807,13.181552,14.083209,15.343266,17.086218,19.108345,20.311813,19.798737,18.987621,18.28214,17.108854,16.207197,16.165699,16.795727,17.557796,17.550251,17.41821,18.184053,19.54597,20.760756,20.632486,20.270313,19.91946,19.87419,19.994913,19.715738,19.04421,18.470772,17.870924,17.425755,17.60684,2.7615614,3.3727267,4.074435,5.2628117,6.466279,6.330465,7.394345,7.484888,6.5945487,5.081726,3.6783094,3.3953626,2.6031113,1.6071383,1.0789708,2.0447628,2.022127,1.6373192,1.3958713,1.3807807,1.2826926,1.3430545,1.4222796,1.6373192,1.9844007,2.3503454,3.361409,4.063117,4.61392,5.2628117,6.349328,5.6023483,5.847569,5.485397,4.5535583,4.7006907,4.1762958,3.6669915,3.5764484,3.6179473,2.8219235,1.2110126,0.51684964,0.25276586,0.16222288,0.19994913,0.28294688,0.48666862,0.8224323,1.2864652,1.8448136,4.8138695,6.617184,6.688864,5.7570257,5.8437963,6.6850915,5.304311,3.821669,3.048281,2.4861598,2.1579416,2.203213,2.3088465,2.4672968,3.006782,3.0558262,3.1048703,2.9313297,2.8181508,3.5236318,4.7572803,5.451443,6.3719635,7.8319697,9.688101,10.506761,11.057564,10.978339,10.887795,12.3893,12.989148,10.684074,7.3075747,4.5497856,3.953711,4.9534564,4.5724216,4.063117,3.942393,3.9688015,5.8702044,4.9760923,3.8254418,3.289729,2.5314314,1.9957186,2.6295197,3.1916409,3.5424948,4.6554193,6.2663302,4.772371,3.180323,2.6068838,2.2899833,1.5430037,1.5241405,1.4675511,1.1544232,0.8865669,0.8865669,1.1242423,1.2864652,1.3392819,1.50905,1.4750963,1.4298248,1.50905,1.8863125,2.776652,3.338773,2.7653341,2.3201644,2.5804756,3.4481792,3.2520027,3.3425457,3.3915899,3.5047686,4.2102494,4.2102494,3.874486,3.3350005,2.7653341,2.3503454,1.9466745,1.7655885,1.7316349,1.8297231,2.0598533,1.8636768,1.8146327,1.4864142,0.845068,0.26031113,0.22258487,0.21503963,0.27917424,0.663982,1.7995421,2.1805773,2.3390274,2.2748928,2.1466236,2.2598023,1.7580433,1.1204696,0.6752999,0.56589377,0.7469798,1.9202662,2.6898816,3.097325,3.1237335,2.6710186,2.7691069,3.8254418,4.534695,4.538468,4.4403796,5.247721,6.379509,7.5112963,8.541223,9.627739,11.32542,13.781399,16.784409,19.61765,21.058792,22.303759,22.613113,21.35683,20.183544,23.039421,25.933023,26.34424,28.306005,32.444576,36.009705,39.3183,43.543636,48.74986,55.49909,64.851425,69.74452,77.89716,80.46255,75.12051,66.10017,58.079563,54.189987,53.60523,53.51846,49.149757,47.059723,47.931202,50.670128,54.431435,58.59264,56.287563,65.8738,91.33148,113.22779,88.72837,50.179684,36.900043,37.492348,42.381668,43.82281,44.799923,47.68221,53.75236,62.44449,71.32147,81.330246,77.285995,61.520195,42.279808,33.723495,27.49489,23.028103,22.284895,23.914669,23.254461,22.77911,23.228052,23.831673,22.684793,16.739138,13.102326,12.54775,12.672247,11.083972,5.43258,3.953711,4.436607,4.5950575,4.3913355,6.0286546,7.5905213,7.1566696,6.149379,5.3646727,4.9760923,4.0706625,3.3161373,2.8332415,2.625747,2.5616124,2.1353056,2.7615614,6.043745,9.544742,6.7756343,5.798525,4.044254,3.8782585,5.0779533,4.821415,4.881777,5.7570257,6.4134626,6.9227667,8.484633,9.178797,9.14107,8.873214,8.831716,9.431562,9.514561,10.718028,12.883514,16.422237,22.29244,21.073883,21.598278,19.934551,16.58446,16.524097,12.608112,11.936585,12.706201,13.475817,13.181552,10.38981,13.023102,17.96524,21.036158,16.984358,17.580433,18.7839,20.424992,22.63575,25.834936,32.41062,33.508453,30.652578,25.721758,20.949387,15.456445,11.649866,10.212496,10.661438,11.306557,11.012292,10.9594755,11.257513,11.046246,8.484633,8.59404,8.986393,10.159679,11.955449,13.5663595,11.819634,9.733373,8.080963,6.9189944,5.5985756,5.247721,4.2064767,3.229367,2.493705,1.6033657,1.297783,1.5316857,1.8749946,2.4597516,3.9989824,6.9869013,7.7187905,6.4926877,4.0782075,1.7089992,0.98842776,1.4939595,1.4524606,1.0789708,2.595566,4.2404304,9.276885,10.325675,7.6395655,9.0807085,8.869441,11.136789,15.422491,20.934296,26.551735,30.837437,31.026068,29.422703,30.033867,38.60527,36.394512,34.213936,30.882708,27.396803,26.93277,35.564537,36.51901,31.169428,22.439573,14.849052,13.113645,11.306557,9.25425,7.1868505,5.723072,4.5497856,4.074435,4.5497856,5.534441,5.873977,5.3609,5.142088,5.5683947,6.458734,7.0963078,8.424272,8.36391,8.114917,7.8432875,6.6850915,1.5920477,1.6750455,4.636556,7.9753294,8.986393,7.8395147,3.6443558,1.3053282,1.6939086,1.6335466,1.6222287,2.1579416,2.4182527,1.9730829,0.76207024,1.8259505,2.7313805,3.9348478,5.515578,7.1868505,7.7112455,7.7225633,8.175279,9.2995205,10.604849,12.264804,11.902632,11.431054,11.246195,10.208723,9.989911,8.816625,8.412953,9.005256,9.322156,8.650629,8.36391,7.786698,7.039718,7.066127,7.001992,6.9982195,6.8699503,6.6662283,6.6662283,6.058836,4.825187,3.9273026,3.7348988,4.0291634,4.0291634,3.5160866,2.8558772,2.2296214,1.6184561,1.2525115,1.0789708,1.1091517,1.2223305,1.1732863,1.0525624,0.97710985,0.9695646,0.995973,0.94692886,0.995973,1.1091517,1.1732863,1.1091517,0.83752275,0.9242931,1.3128735,1.4034165,1.1355602,0.97710985,0.8186596,0.79602385,0.65643674,0.49044126,0.7469798,1.4071891,1.7165444,1.9127209,2.093807,2.2296214,2.655928,3.0105548,3.6179473,4.606375,5.873977,6.9227667,6.4738245,5.583485,4.930821,4.821415,5.455216,5.945657,5.8588867,5.20245,4.4101987,3.9348478,3.8593953,3.712263,3.5689032,4.0593443,4.398881,4.908185,5.1647234,5.0138187,4.561104,4.9421387,6.326692,8.126234,9.669238,10.193633,10.853842,11.363147,11.566868,11.491416,11.3820095,11.299012,11.204697,11.332966,11.517824,11.200924,10.785934,10.416218,10.367173,10.740664,11.476325,10.27663,8.8618965,8.058327,7.964011,7.964011,7.9036493,7.118943,6.0626082,5.1798143,4.8968673,4.666737,4.0782075,3.5085413,3.1614597,3.0520537,2.806833,2.7917426,3.078462,3.4670424,3.4783602,3.5047686,3.802806,4.13857,4.5233774,5.2175403,6.0362,6.9189944,7.956466,8.797762,8.650629,8.382772,8.024373,8.488406,9.635284,10.269085,9.574923,8.793989,7.9715567,7.152897,6.40969,6.7379084,6.507778,6.043745,5.3910813,4.304565,4.0593443,4.0970707,3.7990334,3.1048703,2.5314314,2.191895,1.8221779,1.6675003,1.8297231,2.2598023,2.354118,2.4069347,2.2371666,1.8787673,1.5882751,1.6222287,1.5505489,1.3656902,1.0940613,0.77716076,0.7054809,0.80734175,0.8299775,0.80356914,1.0223814,1.1921495,1.4637785,1.5920477,1.6033657,1.7844516,1.81086,1.6071383,1.5203679,1.6222287,1.7089992,1.4034165,1.3015556,1.4524606,1.6448646,1.388326,1.0714256,0.95447415,1.0412445,1.2223305,1.297783,0.9922004,1.6109109,1.8976303,1.6863633,1.9089483,2.5804756,2.4710693,2.1956677,2.0862615,2.1956677,2.7351532,3.361409,4.485651,5.9796104,7.1868505,6.9680386,7.5716586,8.262049,8.763808,9.276885,10.899114,13.057055,14.245432,13.777626,11.763044,11.472552,11.076427,10.570895,9.910686,9.016574,9.14107,8.869441,7.9828744,6.7831798,6.089017,6.198423,6.537959,6.7379084,6.749226,6.8359966,7.2887115,7.3453007,7.6810646,8.254503,8.314865,7.145352,6.1078796,5.451443,5.406172,6.224831,7.5792036,8.469543,9.390063,10.484125,11.536687,12.427027,13.528633,15.01882,16.788181,18.448135,19.972277,19.813826,18.821627,17.53516,16.203424,15.754482,16.15438,16.91645,17.550251,17.56157,17.72002,19.089483,20.247679,20.387266,19.300749,19.108345,19.553514,19.957186,19.889278,19.180025,17.667202,17.278622,17.240896,17.448391,18.463226,2.516341,4.436607,5.5457587,5.975838,6.096562,6.5266414,6.9567204,7.364164,6.749226,5.1043615,3.3953626,2.4333432,1.4373702,0.80356914,0.66775465,0.90920264,0.935611,1.3694628,1.4826416,1.2147852,1.1846043,1.177059,1.1355602,1.1996948,1.4222796,1.7882242,2.565385,3.399135,4.3347464,5.160951,5.406172,5.0741806,5.553304,5.353355,4.4177437,4.1272516,3.6707642,3.2029586,3.0331905,2.9954643,2.444661,1.6260014,0.80356914,0.33953625,0.30935526,0.5017591,0.5394854,0.6375736,0.91297525,1.4864142,2.4672968,3.6179473,6.066381,6.5568223,5.0062733,4.52715,4.402653,4.353609,3.9386206,3.169005,2.5012503,1.9466745,3.3350005,4.659192,5.4438977,6.741681,5.9305663,5.7796617,6.903904,8.7600355,9.654147,10.152134,11.359374,13.909668,16.890041,17.818108,18.41041,17.765291,16.791954,15.297995,11.974312,10.718028,9.261794,7.77538,6.9189944,7.8319697,8.024373,7.141579,6.368191,5.8136153,4.478106,4.538468,4.3724723,4.164978,3.92353,3.5085413,3.2369123,3.6858547,4.3913355,4.515832,2.8822856,3.6858547,3.8065786,3.5651307,3.3651814,3.6934,2.4408884,1.7429527,1.388326,1.2261031,1.1544232,1.2298758,1.1732863,1.1581959,1.1959221,1.1317875,1.0751982,1.0412445,1.1053791,1.3920987,2.0560806,2.1692593,1.5052774,1.0072908,1.3505998,2.9464202,3.6896272,3.9122121,4.104616,4.3913355,4.4931965,4.266839,4.29702,3.783943,2.6597006,1.5807298,1.4901869,1.8749946,2.2899833,2.4974778,2.4861598,2.173032,2.0673985,1.6410918,0.875249,0.271629,0.24522063,0.4376245,0.724344,1.1204696,1.7882242,1.659955,1.4411428,1.2110126,1.0412445,1.026154,0.8865669,0.6187105,0.43007925,0.56589377,1.2864652,1.9202662,2.4597516,2.9200118,2.9049213,1.5845025,2.9501927,4.2027044,4.564876,4.3196554,4.8063245,6.0211096,7.069899,8.394091,10.359629,13.253232,17.048492,18.406637,19.527107,21.368149,23.620405,21.09652,21.09652,21.503962,22.382984,25.97075,30.377176,29.086939,28.200373,30.105547,33.48582,36.18702,39.159847,42.589165,47.576572,56.14798,66.22843,76.73897,82.922295,81.45097,70.44623,60.56195,56.578056,58.717136,62.625576,59.388664,54.918102,54.52575,54.86151,55.73299,60.120552,60.497814,69.02772,91.41825,113.506966,101.25348,63.602684,45.44127,44.464157,54.073032,63.35369,57.317493,51.518967,49.662834,55.21614,71.39316,91.478615,88.822685,68.81268,43.73227,32.746384,25.514263,20.319359,17.938831,17.516298,16.565596,21.371922,24.597515,24.299479,20.145817,13.430545,10.34831,8.756263,8.620448,8.733627,6.7152724,4.6516466,3.5349495,3.0445085,3.2331395,4.52715,6.5455046,6.647365,6.1418333,5.881522,6.2436943,6.1606965,5.5570765,4.6856003,3.9876647,4.112161,2.11267,2.2748928,4.644101,7.7301087,8.484633,5.50426,3.3878171,3.2633207,4.6214657,5.323174,4.349837,5.05909,6.039973,7.24344,9.997457,10.47658,10.367173,10.287949,10.631257,11.54046,10.729345,12.966512,16.195879,18.429274,17.727566,20.519308,21.209698,19.727057,16.946632,14.671739,16.143063,14.264296,12.0082655,11.053791,11.815862,9.49947,11.944131,14.966003,16.361876,15.920478,15.328176,16.437326,19.093256,22.235851,23.892035,30.66767,34.59497,34.71192,30.860073,23.68454,17.7917,13.290957,11.695138,12.121444,11.295239,10.465261,10.099318,9.982366,9.601331,8.141325,8.507269,9.125979,10.325675,12.049765,13.845533,14.883006,14.196388,11.246195,7.2660756,5.292993,4.659192,3.8593953,3.1954134,2.6295197,1.7957695,5.4665337,4.006528,3.7575345,6.4210076,9.061845,13.215506,10.970794,6.7114997,3.5387223,3.270866,1.1921495,1.3468271,1.720317,1.5430037,1.2864652,3.0331905,5.975838,11.246195,17.048492,18.685812,14.992412,12.830698,14.679284,19.700647,23.741129,26.219744,25.910389,23.503454,22.488617,29.143528,26.604551,26.593233,26.698868,25.257725,21.379465,21.941587,23.190327,23.560043,21.383238,14.883006,13.88326,12.434572,10.495442,8.461998,7.164215,6.851087,6.934085,7.118943,7.066127,6.3644185,5.402399,5.040227,5.836251,7.7829256,10.291721,9.857869,8.688355,7.752744,7.7640624,9.175024,2.8709676,2.191895,5.43258,9.514561,9.952185,9.488152,7.937603,7.3377557,7.2283497,4.647874,3.229367,3.5764484,3.731126,3.169005,2.7879698,3.9574835,5.587258,7.1076255,8.420499,9.895596,11.710228,12.257258,12.449662,12.683565,12.838243,15.07541,15.128226,13.754991,12.242168,12.404391,12.830698,12.0082655,10.861387,9.87296,9.114662,8.688355,8.827943,8.511042,7.9489207,8.578949,7.756517,7.24344,7.322665,7.5603404,6.828451,5.775889,4.7421894,4.123479,3.99521,4.1008434,4.0216184,3.5424948,2.9011486,2.1956677,1.3619176,1.1016065,0.95447415,0.94315624,1.0035182,1.0035182,0.88279426,0.80734175,0.8299775,0.90543,0.8978847,0.8978847,0.8526133,0.8601585,0.9280658,0.97333723,0.94315624,1.0638802,1.146878,1.116697,1.0374719,0.8903395,0.8186596,0.7130261,0.66020936,0.95447415,1.3317367,1.6222287,1.7165444,1.6976813,1.8599042,2.2899833,2.8558772,3.5236318,4.398881,5.726845,5.4401255,4.8365054,4.2517486,3.8820312,3.772625,4.564876,4.4403796,4.285702,4.2781568,3.8858037,3.399135,3.1463692,2.8822856,2.8181508,3.6179473,4.5196047,4.9723196,5.198677,5.138315,4.4516973,4.7421894,5.87775,7.232122,8.431817,9.374973,10.035183,10.899114,11.778135,12.408164,12.445889,11.2650585,10.386037,9.771099,9.695646,10.736891,9.989911,9.910686,9.710737,9.57115,10.646348,10.042727,9.156161,8.303548,7.7602897,7.7716074,7.405663,6.428553,5.304311,4.4403796,4.1762958,3.99521,3.651901,3.2859564,2.9803739,2.7841973,2.5012503,2.5767028,2.9049213,3.229367,3.1727777,3.0143273,3.1425967,3.2369123,3.4255435,4.266839,4.7120085,5.7004366,6.560595,6.8774953,6.466279,6.7152724,6.771862,6.930312,7.375482,8.145098,8.190369,7.7904706,7.1906233,6.63982,6.3832817,5.824933,5.485397,5.3382645,5.243949,4.949684,4.4818783,4.244203,4.0593443,3.6707642,2.7653341,2.2862108,1.9429018,1.7014539,1.6146835,1.8184053,2.757789,2.6219745,2.093807,1.6146835,1.3920987,1.4562333,1.297783,1.0223814,0.77716076,0.7432071,0.5998474,0.6526641,0.7167987,0.79602385,1.0827434,1.2826926,1.8334957,2.1654868,2.0862615,1.7618159,1.659955,1.5467763,1.4109617,1.2713746,1.1732863,1.0827434,1.0751982,1.1506506,1.1959221,0.9997456,0.7205714,0.9205205,1.1959221,1.358145,1.4298248,1.1053791,1.4373702,1.9957186,2.5616124,3.1048703,3.3463185,3.1312788,2.8106055,2.7426984,3.270866,3.270866,3.610402,4.3800178,5.13077,4.9044123,5.613666,6.8133607,8.054554,9.103344,9.937095,12.283667,14.037937,14.019074,12.14408,9.457971,10.442626,10.853842,10.235131,8.922258,8.043237,7.665974,7.175533,6.4436436,5.5797124,4.9044123,5.111907,5.4665337,5.87775,6.145606,5.956975,5.6476197,6.3644185,7.4471617,8.14887,7.6320205,5.80607,4.8930945,4.727099,5.240176,6.470052,7.413208,8.194141,9.06939,10.238904,11.815862,13.13628,14.075664,15.32063,16.946632,18.41041,19.300749,19.217752,18.463226,17.395575,16.42601,15.814844,15.196134,14.86037,15.079182,16.086473,16.614641,18.26705,19.806282,20.23636,18.791445,18.614132,19.436563,19.938324,19.493153,18.18028,18.070873,17.508753,17.63325,18.644312,19.794964,5.20245,4.9232755,4.9459114,4.9534564,4.957229,5.304311,4.979865,5.3646727,4.979865,3.6141748,2.293756,1.539231,0.8526133,0.48666862,0.452715,0.5357128,0.43007925,0.724344,0.94315624,0.9997456,1.1695137,0.86770374,0.80356914,0.90920264,1.116697,1.3732355,1.9768555,3.0935526,3.8593953,4.036709,4.036709,4.346064,4.7610526,4.8440504,4.6214657,4.5761943,4.0706625,3.4179983,3.1048703,3.0105548,2.4031622,1.6788181,0.8639311,0.452715,0.4979865,0.5998474,0.6526641,0.8224323,1.2600567,2.1353056,3.6330378,4.4743333,6.047518,6.628502,6.058836,5.753253,5.0553174,4.093298,3.229367,2.6332922,2.2748928,2.093807,2.9615107,4.0216184,5.7192993,9.782416,7.466025,7.375482,9.510788,12.574159,13.977575,12.355347,13.543724,15.728074,17.580433,18.26705,18.97253,16.84477,15.184815,14.456699,12.291212,10.616167,9.374973,8.643084,8.228095,7.6697464,7.1302614,6.560595,6.0022464,5.2892203,4.0404816,3.682082,3.5802212,3.6443558,3.6481283,3.2218218,3.0369632,3.3651814,4.055572,4.5535583,3.8895764,3.5274043,3.2784111,3.0331905,2.9237845,3.3463185,2.8747404,2.565385,2.3578906,2.203213,2.052308,1.659955,1.3845534,1.0978339,0.8111144,0.6790725,0.62625575,0.6111652,0.6375736,0.76584285,1.1355602,1.4864142,1.0601076,0.663982,0.87902164,2.052308,2.4974778,3.0256453,3.7877154,4.5309224,4.636556,3.8065786,3.3274553,2.7879698,2.0975795,1.4977322,1.5882751,2.1579416,2.6672459,2.746471,2.191895,1.8146327,1.5882751,1.1317875,0.49421388,0.15467763,0.181086,0.36594462,0.7394345,1.1883769,1.4298248,1.1996948,1.2525115,1.2110126,0.97710985,0.754525,0.8526133,0.5093044,0.392353,0.7884786,1.5920477,1.8599042,1.9655377,2.0447628,1.9693103,1.3317367,2.1202152,3.4029078,4.285702,4.8440504,6.115425,7.748972,7.8131065,8.27714,10.020092,12.860879,15.988385,16.803272,17.852062,19.711966,20.994658,18.814081,18.980076,20.892797,23.748674,26.547962,32.41062,31.429739,29.8641,30.66767,33.493366,38.337414,41.944046,44.61129,48.10474,55.66508,66.96032,74.85642,79.213806,79.11572,72.853165,63.217876,59.479206,61.463608,65.43996,64.11199,58.370052,57.411808,56.63842,55.408543,57.04209,59.218895,69.9407,94.99847,120.82209,114.46522,74.11699,54.55216,54.133396,65.428635,75.22237,64.3308,52.895977,46.380653,48.9234,63.35369,95.23992,99.140816,77.85189,47.335125,36.711414,30.181,25.872662,24.016531,23.103556,19.87419,23.805264,22.813063,19.568605,15.69412,11.7894535,9.748463,7.141579,6.4134626,7.224577,6.458734,4.5422406,3.1765501,2.4522061,2.4710693,3.361409,5.383536,6.379509,6.790725,6.700182,5.8664317,6.228604,6.258785,6.0739264,5.8437963,5.772116,3.7763977,3.3727267,4.647874,6.5945487,7.115171,5.0439997,3.682082,3.561358,4.349837,4.878004,4.195159,4.7421894,5.8211603,7.2057137,9.122208,11.329193,11.083972,10.899114,11.717773,12.902377,11.944131,14.117163,17.64834,19.930779,17.527617,21.375692,20.549488,18.09351,15.335721,11.891314,13.977575,13.487134,12.034674,10.842525,10.759526,8.98262,11.25374,13.245687,13.389046,12.864652,14.335975,17.712475,20.69662,22.020813,21.42851,24.914415,28.339958,29.332159,27.061039,22.235851,17.640795,14.841507,13.505998,12.989148,12.325166,10.718028,9.476834,8.605357,7.956466,7.24344,8.620448,10.220041,11.216014,11.853588,13.441863,15.467763,15.614895,12.792972,8.167733,5.1835866,5.0439997,4.4403796,3.6330378,2.8030603,2.0673985,3.92353,3.0935526,3.8103511,7.0585814,10.567122,11.993175,8.36391,4.304565,2.1843498,2.123988,0.98842776,0.84129536,1.0978339,1.3656902,1.4373702,3.361409,4.285702,10.393582,20.956932,28.347504,25.325632,20.647577,18.734856,20.790936,24.76351,23.741129,22.503708,20.994658,20.04773,21.394556,20.904116,21.322876,20.511763,18.063328,15.32063,17.029629,17.814335,19.134754,19.787418,15.890297,14.517061,13.053283,11.721546,10.299266,8.126234,8.145098,9.133525,9.574923,8.918486,7.575431,6.579458,6.379509,8.096053,10.714255,11.091517,10.212496,9.0543,8.27714,8.29223,9.239159,2.8521044,2.0258996,4.5837393,7.9526935,9.14107,9.997457,10.725573,9.703192,7.224577,5.492942,5.3571277,7.273621,8.405409,8.224322,8.484633,9.186342,10.170997,11.114153,11.898859,12.653384,14.120935,14.279386,14.000212,13.7700815,13.671993,15.267814,14.916959,14.022847,13.513543,13.822898,13.736128,13.253232,12.283667,11.072655,10.208723,9.997457,9.869187,9.386291,8.903395,9.590013,8.544995,7.8508325,7.435844,7.2358947,7.2057137,6.0512905,4.919503,4.1310244,3.8254418,3.983892,3.6858547,3.2746384,2.795515,2.2220762,1.4260522,1.0827434,1.0525624,1.0412445,0.9620194,0.91674787,0.8224323,0.7809334,0.7696155,0.76584285,0.7205714,0.84884065,0.77338815,0.7469798,0.84129536,0.9695646,0.87902164,0.95824677,1.0487897,1.0827434,1.0714256,0.90920264,0.7582976,0.66020936,0.7092535,1.0450171,1.2600567,1.5580941,1.6033657,1.4675511,1.6222287,1.8033148,2.3314822,2.8558772,3.308592,3.9348478,3.6254926,3.4255435,3.2218218,3.1048703,3.380272,3.953711,3.9989824,4.025391,4.063117,3.651901,3.048281,2.704972,2.5201135,2.625747,3.4179983,3.7801702,4.055572,4.557331,5.05909,4.7912335,5.2779026,5.9305663,6.7341356,7.7301087,9.005256,9.578695,10.231359,10.9594755,11.52537,11.476325,10.49167,9.74469,9.261794,9.107117,9.4127,8.990166,9.242931,9.480607,9.65792,10.3634,9.869187,9.107117,8.367682,7.8734684,7.8206515,7.24344,6.349328,5.3344917,4.4101987,3.7877154,3.4557245,3.519859,3.5274043,3.3576362,3.2105038,2.806833,2.584248,2.7313805,3.1010978,3.2255943,3.0256453,2.867195,2.6974268,2.655928,3.0671442,3.7650797,4.644101,5.4174895,5.802297,5.5193505,5.624984,5.824933,5.9532022,6.058836,6.432326,7.1793056,7.1906233,6.9152217,6.4964604,5.7909794,5.119452,4.5799665,4.2291126,4.115934,4.29702,4.0593443,3.8141239,3.4859054,3.1048703,2.795515,2.584248,2.3616633,2.2711203,2.2371666,2.003264,2.9426475,2.8822856,2.354118,1.7995421,1.5731846,1.4411428,1.2147852,0.9242931,0.6790725,0.6790725,0.58475685,0.62248313,0.77338815,1.0035182,1.2713746,1.4222796,1.8938577,2.1692593,2.1315331,2.0749438,1.6109109,1.2940104,1.0110635,0.77716076,0.7167987,0.95824677,1.0902886,1.0110635,0.7922512,0.69793564,0.5696664,0.8941121,1.1619685,1.20724,1.237421,1.3958713,1.6448646,2.3201644,3.199186,3.4745877,3.7047176,3.9725742,3.8178966,3.4481792,3.731126,3.8178966,4.191386,4.768598,5.311856,5.413717,6.126743,7.0170827,8.009283,9.027891,9.97482,11.744182,13.43809,13.4644985,11.706455,9.540969,10.106862,10.612394,10.095545,8.733627,7.8696957,7.3981175,6.6134114,5.783434,5.1269975,4.7912335,4.8968673,4.919503,5.1043615,5.3873086,5.372218,5.062863,5.643847,6.6549106,7.326438,6.6020937,5.0439997,4.5535583,4.7346444,5.2628117,5.9003854,6.888813,7.9225125,9.178797,10.729345,12.562841,13.6833105,14.547242,15.384765,16.388283,17.716248,18.991394,18.983849,18.157644,17.071129,16.395828,15.290449,14.252977,13.513543,13.422999,14.464244,15.845025,18.297232,20.266542,20.723028,19.15739,18.912169,18.761265,18.772581,18.719765,18.112373,17.784155,17.60684,18.02183,19.051756,20.30804,5.9117036,4.5120597,3.863168,3.802806,4.1197066,4.5422406,3.7386713,3.7235808,3.3161373,2.263575,1.2600567,0.8639311,0.56589377,0.40367088,0.36971724,0.41121614,0.30935526,0.35839936,0.60362,1.0035182,1.4260522,0.9318384,0.7469798,0.7582976,0.8978847,1.146878,1.7391801,2.8106055,3.380272,3.338773,3.4594972,3.9197574,4.1612053,4.4894238,4.919503,5.1835866,4.561104,3.712263,3.2784111,3.1237335,2.3390274,1.6712729,0.94315624,0.6073926,0.66020936,0.62248313,0.80356914,0.98842776,1.3468271,2.0447628,3.229367,4.06689,5.2326307,6.617184,8.024373,9.175024,7.405663,4.90064,3.361409,3.350091,4.304565,4.3875628,5.2590394,6.477597,8.039464,10.397354,8.194141,8.835487,11.604594,15.399856,18.742401,17.467255,18.433046,19.68933,20.217497,19.968504,19.327158,16.91645,14.78869,13.328684,11.2801485,9.454198,7.8734684,7.0963078,6.79827,5.73439,5.040227,5.070408,5.0553174,4.6327834,3.832987,3.0331905,2.6483827,2.6785638,2.9049213,2.8558772,2.625747,2.927557,3.4481792,3.8707132,3.8443048,3.5764484,3.2859564,3.0746894,3.006782,3.1048703,3.0633714,2.9313297,2.7125173,2.4371157,2.1692593,1.5958204,1.2223305,0.84129536,0.49044126,0.45648763,0.41121614,0.35839936,0.31312788,0.3169005,0.44516975,0.80734175,0.6752999,0.55080324,0.724344,1.2789198,1.4675511,2.0598533,2.7615614,3.2557755,3.187868,2.282438,1.6788181,1.7580433,2.3126192,2.565385,2.1881225,2.2258487,2.3013012,2.1390784,1.5807298,1.3015556,1.0940613,0.724344,0.28294688,0.19994913,0.26408374,0.35085413,0.60362,0.90543,0.8563859,0.9507015,1.2826926,1.2940104,1.0072908,1.0148361,0.8903395,0.5319401,0.52439487,1.0299267,1.7995421,2.142851,1.871222,1.5015048,1.2600567,1.0638802,1.4562333,2.8445592,4.4215164,5.881522,7.3905725,8.858124,8.495952,8.303548,9.314611,11.608367,13.234368,14.347293,16.309057,18.429274,17.972786,17.316349,18.018057,20.028866,23.39782,28.287142,33.021786,32.629433,31.852272,32.5653,33.78763,40.25391,45.060234,47.689754,49.877876,55.597176,64.851425,70.29532,73.31719,74.38862,73.05311,65.96435,63.059425,63.632866,65.31923,64.11199,59.84515,59.283028,57.77398,54.574795,52.81675,54.740788,65.511635,91.09003,120.425964,125.45864,81.97537,61.15425,62.180405,75.29405,81.79428,67.695984,53.42414,44.543385,44.818787,56.212112,94.711754,105.38451,84.50303,49.345936,38.197826,33.738586,30.075367,29.049213,29.430248,26.868635,25.948114,20.074137,13.962485,13.087236,23.69963,14.071891,7.541477,5.142088,5.6551647,5.5797124,4.8138695,3.5575855,2.8898308,2.957738,2.9464202,4.4101987,5.6589375,6.3229194,6.2097406,5.3156285,5.553304,5.783434,5.8890676,5.855114,5.7796617,4.5837393,4.3913355,5.6400743,7.3415284,7.092535,5.987156,5.5080323,5.3571277,5.2062225,4.719554,4.644101,4.9459114,5.8098426,7.066127,8.20546,11.23865,11.374464,11.378237,12.291212,13.407909,12.966512,15.328176,18.327412,19.828917,17.753973,20.673985,19.383747,16.840998,14.120935,10.423763,12.170488,13.083464,12.800517,11.574413,10.272858,9.35611,10.601076,12.611885,14.652876,16.641048,15.214996,17.753973,20.349539,20.870161,18.983849,20.455173,22.50748,23.141281,21.711456,18.908396,16.18456,15.916705,15.539442,14.339747,13.430545,11.446144,9.710737,8.2507305,7.224577,6.94163,8.669493,10.125726,10.676529,10.804798,12.0724,14.075664,15.079182,13.622949,9.918231,5.8211603,5.9796104,5.111907,4.376245,3.9386206,2.987919,2.6182017,2.2447119,3.6028569,7.0170827,11.393328,7.6810646,4.2894745,2.2069857,1.4411428,1.0299267,0.72811663,0.48666862,0.6375736,1.2034674,1.8938577,3.7084904,4.0291634,9.329701,19.94964,30.101774,30.090458,27.170444,23.8279,22.349031,24.812555,22.428255,21.579414,21.100292,20.066593,17.787928,16.644821,16.086473,14.977322,13.200415,11.634775,14.6302395,16.094019,17.908651,19.500698,17.87847,15.569623,14.083209,13.385274,12.777881,10.902886,10.167224,10.408672,10.412445,9.756008,8.793989,8.544995,7.779153,9.042982,11.559323,11.208468,10.197406,9.895596,9.725827,9.631512,10.054046,4.164978,2.4371157,4.5460134,8.397863,10.121953,12.117672,12.012038,10.125726,8.039464,8.59404,8.548768,10.065364,11.649866,12.808062,14.045483,14.188843,14.441608,14.377474,14.177525,14.600059,15.520579,15.230087,14.219024,13.2607765,13.415455,14.524607,14.0983,13.675766,13.758763,13.822898,14.128481,14.015302,13.2607765,12.045992,10.982111,11.231105,10.842525,10.303039,10.125726,10.850069,9.325929,8.318638,7.496206,6.952948,7.2170315,6.205968,5.093044,4.29702,3.9688015,3.9876647,3.6292653,3.2255943,2.8294687,2.3428001,1.5467763,1.1808317,1.1959221,1.1581959,0.9808825,0.91674787,0.84129536,0.7809334,0.73188925,0.70170826,0.6828451,0.8111144,0.724344,0.68661773,0.79602385,0.95824677,0.7997965,0.94692886,1.0676528,1.0751982,1.1431054,0.95824677,0.7432071,0.6375736,0.7205714,0.995973,1.1846043,1.4373702,1.4373702,1.267602,1.4034165,1.5618668,2.0296721,2.4031622,2.5427492,2.5729303,2.5087957,2.5125682,2.5087957,2.595566,3.0331905,3.5236318,3.802806,3.8820312,3.7348988,3.2746384,2.6408374,2.4522061,2.493705,2.7087448,3.218049,3.0030096,3.3312278,4.002755,4.640329,4.6742826,5.3458095,5.907931,6.5756855,7.5603404,9.092027,9.857869,10.386037,10.751981,10.884023,10.56335,9.846551,9.246704,8.918486,8.7751255,8.473316,8.345046,8.692128,9.235386,9.752235,10.106862,9.665465,9.024119,8.424272,8.001738,7.8017883,7.3453007,6.4926877,5.458988,4.45547,3.6669915,3.3425457,3.6179473,3.821669,3.7009451,3.4255435,2.9237845,2.5578396,2.6295197,2.9652832,2.916239,2.7125173,2.4333432,2.233394,2.203213,2.3578906,3.2029586,4.1612053,4.8629136,5.1232247,4.930821,4.8402777,5.028909,5.142088,5.1571784,5.383536,6.1116524,6.398372,6.296511,5.8400235,5.040227,4.3800178,3.7613072,3.361409,3.2557755,3.4179983,3.3236825,3.2142766,2.8936033,2.4823873,2.4371157,2.4220252,2.4522061,2.5880208,2.6823363,2.372981,2.867195,2.8181508,2.4107075,1.901403,1.6071383,1.4260522,1.1016065,0.80356914,0.63002837,0.58475685,0.58475685,0.6187105,0.8337501,1.177059,1.3656902,1.4562333,1.6863633,1.9127209,2.0447628,2.033445,1.3392819,0.94692886,0.7092535,0.56212115,0.5281675,0.7469798,0.8563859,0.7432071,0.52062225,0.5281675,0.6752999,1.1317875,1.4901869,1.6750455,1.9240388,2.022127,2.142851,2.5314314,3.1161883,3.500996,3.9122121,4.2592936,4.13857,3.7462165,3.874486,4.191386,4.5460134,5.0666356,5.7004366,6.2135134,6.7341356,7.352846,8.054554,8.899622,10.035183,11.302785,12.766563,12.777881,11.2801485,9.80128,9.6051035,9.778644,9.390063,8.394091,7.6320205,7.141579,6.175787,5.323174,4.8629136,4.749735,4.6252384,4.466788,4.5196047,4.7874613,5.0213637,5.036454,5.4703064,6.1041074,6.398372,5.4703064,4.376245,4.3611546,4.7233267,5.119452,5.5570765,6.643593,8.009283,9.495697,11.042474,12.679792,13.604086,14.434063,15.192361,15.961976,16.886269,18.082191,18.361366,17.927513,17.093763,16.263786,14.588741,13.317367,12.438345,12.272349,13.460726,15.701665,18.55377,20.519308,20.802254,19.338476,18.991394,18.150099,17.731337,17.870924,17.946377,18.014284,18.052011,18.414183,19.149845,20.017548,3.9989824,3.640583,3.180323,3.2067313,3.8103511,4.5988297,3.6707642,3.0897799,2.474842,1.6750455,0.7582976,0.51684964,0.41876137,0.36971724,0.32444575,0.28294688,0.32067314,0.3734899,0.6111652,1.0789708,1.6675003,1.2713746,0.9280658,0.7092535,0.7130261,1.0638802,1.7278622,2.425798,2.9652832,3.3425457,3.731126,3.7499893,3.8443048,4.266839,4.889322,5.1873593,4.5196047,3.7650797,3.4557245,3.3915899,2.655928,2.0560806,1.327964,0.94315624,0.9205205,0.84884065,1.0902886,1.1808317,1.2336484,1.3355093,1.5580941,2.1843498,3.7499893,6.1908774,9.110889,11.7894535,9.2995205,6.1078796,4.3649273,4.908185,7.2585306,7.7678347,9.699419,12.287439,13.822898,11.649866,10.801025,12.562841,15.101818,18.240643,23.450638,24.842735,25.627441,26.106565,25.917934,24.031622,21.994404,20.689075,18.233097,14.264296,9.937095,7.6886096,5.534441,4.2781568,4.025391,4.183841,3.821669,4.1612053,4.5196047,4.515832,4.0895257,2.9086938,2.2296214,2.142851,2.4786146,2.8332415,2.5276587,2.9351022,3.229367,3.0218725,2.3126192,3.127506,3.5085413,3.6971724,3.7235808,3.3878171,2.897376,2.5578396,2.1768045,1.720317,1.3166461,1.0072908,0.69793564,0.44516975,0.32444575,0.40367088,0.36971724,0.27540162,0.19240387,0.15467763,0.15467763,0.22258487,0.28294688,0.41498876,0.6187105,0.79602385,1.1280149,1.5203679,1.6222287,1.3543724,0.90920264,0.4376245,0.30181,1.327964,3.0218725,3.5689032,2.546522,1.8636768,1.3996439,1.1280149,1.1317875,0.9808825,0.8186596,0.56212115,0.31312788,0.362172,0.5055317,0.5885295,0.6413463,0.63002837,0.44516975,0.88279426,1.2298758,1.1091517,0.79602385,1.2147852,0.72811663,0.573439,0.7167987,1.146878,1.8749946,2.6295197,2.214531,1.5430037,1.026154,0.59607476,1.2600567,2.7351532,4.727099,6.673774,7.7376537,8.511042,8.560086,8.465771,8.990166,11.083972,12.057309,13.973803,16.67123,18.708447,17.338985,18.044466,19.119663,20.391039,23.424229,31.569326,32.440804,32.097492,32.716206,34.127167,33.81781,40.12187,45.595947,48.8819,50.96439,55.163322,60.316727,64.48925,67.97516,70.502815,71.230934,67.29608,64.700516,63.546097,63.074516,61.68619,60.026237,59.637657,57.091133,52.45458,49.274254,50.36077,58.241783,79.4628,109.02509,130.38193,87.56263,64.530754,66.33029,82.08478,85.016106,71.93264,59.596157,49.892967,46.210884,53.4166,92.06337,107.331184,87.64185,49.100716,35.504173,32.67848,28.720995,27.491117,29.196344,30.377176,24.329659,16.62973,9.533423,11.344283,36.402058,17.886015,8.141325,4.719554,4.719554,4.798779,5.5495315,4.432834,3.7235808,3.7688525,2.969056,3.7688525,4.568649,4.772371,4.5912848,5.0175915,4.938366,4.8666863,4.5950575,4.2517486,4.3196554,3.9876647,4.5233774,6.428553,8.677037,8.699674,8.145098,8.507269,8.654402,7.8696957,5.847569,5.8702044,5.798525,6.1908774,7.0887623,8.0206,10.38981,11.189606,11.570641,12.162943,13.117417,13.664448,16.667458,18.749947,18.629223,17.112627,18.323639,17.829426,16.505234,14.483108,11.140562,13.030646,14.000212,13.562587,11.917723,9.955957,10.484125,10.31813,12.385528,17.350302,23.593996,17.180534,16.675003,18.387774,19.451654,17.833199,19.368656,20.470263,20.458946,19.112118,16.663685,15.211224,16.52787,17.135263,16.146835,15.290449,12.917468,11.034928,9.525878,8.443134,8.00551,8.669493,8.692128,8.744945,9.239159,10.31813,11.838497,13.626721,13.93985,11.895086,7.432071,6.790725,5.323174,5.2892203,6.1908774,4.8025517,3.5274043,4.3611546,5.7306175,8.099826,13.962485,4.9949555,3.240685,2.8030603,1.5882751,1.297783,5.6815734,4.8855495,2.776652,1.6524098,2.2484846,3.2859564,3.9574835,7.865923,15.437581,23.922215,27.359077,28.404093,25.978296,22.164171,22.213217,21.560553,22.137764,22.005722,20.43631,17.946377,13.513543,11.68382,12.0082655,12.664702,10.438853,11.959221,14.841507,17.742655,19.406384,18.659403,15.818617,14.841507,14.8339615,15.045229,14.875461,13.385274,11.819634,10.567122,9.906913,10.03141,10.582213,8.865668,8.831716,10.838752,11.657412,9.680555,10.525623,10.955703,10.589758,11.883769,6.937857,3.7537618,5.613666,10.831206,12.755245,15.094273,12.332711,10.325675,11.25374,13.649357,11.623458,10.79348,11.634775,13.611631,15.192361,16.59955,17.437073,16.51278,14.879233,15.826162,16.603323,16.086473,14.407655,12.717519,13.170234,13.781399,13.830443,13.5663595,13.230596,13.068373,14.475562,15.098045,14.7170105,13.407909,11.54046,12.061082,11.570641,11.283921,11.657412,12.393073,10.065364,8.846806,8.043237,7.4207535,7.1868505,6.2436943,5.240176,4.644101,4.4516973,4.1612053,3.8971217,3.4670424,3.0181,2.4786146,1.5769572,1.2789198,1.2336484,1.1581959,1.0035182,0.9922004,0.8941121,0.754525,0.70170826,0.7469798,0.79602385,0.7507524,0.6488915,0.6375736,0.7507524,0.9318384,0.7205714,0.94692886,1.1129243,1.1016065,1.1959221,1.0072908,0.7884786,0.69039035,0.7469798,0.88279426,1.1129243,1.2487389,1.2110126,1.1053791,1.237421,1.5769572,2.0108092,2.2975287,2.3503454,2.1956677,2.1541688,2.093807,2.1579416,2.3880715,2.7238352,3.3878171,3.7084904,3.6179473,3.187868,2.6219745,2.2069857,2.3465726,2.6068838,2.7728794,2.8521044,2.6295197,3.1840954,3.7499893,3.99521,4.0480266,4.8365054,5.7004366,6.549277,7.5112963,8.937348,10.182315,10.933067,11.09529,10.748209,10.148361,9.484379,8.82417,8.431817,8.29223,8.103599,8.043237,8.314865,8.820397,9.34102,9.552286,9.405154,9.0807085,8.5563135,7.967784,7.586749,7.5037513,6.647365,5.4703064,4.3649273,3.6669915,3.4444065,3.6066296,3.7650797,3.663219,3.187868,2.6332922,2.41448,2.5729303,2.7728794,2.293756,2.0975795,1.961765,1.9542197,2.0900342,2.3616633,3.0860074,4.1536603,4.7120085,4.6026025,4.3875628,4.236658,4.304565,4.3422914,4.3686996,4.6516466,4.7874613,5.036454,4.8855495,4.3649273,4.0593443,3.399135,2.9652832,2.886058,3.029418,2.9841464,2.8558772,2.9049213,2.7992878,2.4786146,2.161714,2.1466236,2.3767538,2.625747,2.7691069,2.7917426,2.867195,2.6823363,2.2975287,1.8184053,1.3958713,1.2713746,0.8903395,0.6187105,0.543258,0.4678055,0.55080324,0.62625575,0.8526133,1.1657411,1.2864652,1.3128735,1.3807807,1.6410918,1.8636768,1.448688,0.8903395,0.66775465,0.6073926,0.59230214,0.5281675,0.46026024,0.47912338,0.513077,0.5583485,0.69793564,1.1544232,1.690136,2.2258487,2.7200627,3.199186,2.8030603,2.7389257,2.6710186,2.7653341,3.6707642,4.134797,4.104616,3.8971217,3.7952607,4.006528,4.3686996,4.6026025,5.138315,5.8928404,6.247467,6.677546,7.4169807,8.111144,8.8618965,10.246449,11.457462,12.30253,11.853588,10.419991,9.537196,9.005256,8.646856,8.235641,7.6923823,7.0849895,6.462507,5.458988,4.738417,4.45547,4.2404304,3.9612563,3.9574835,4.1197066,4.398881,4.779916,5.1232247,5.511805,5.73439,5.4967146,4.4177437,3.6669915,3.9801195,4.45547,4.9119577,5.8513412,6.8850408,8.390318,9.74469,10.782163,11.793225,12.630749,13.490907,14.543469,15.573396,15.984612,16.501461,17.16167,17.440845,17.006994,15.746937,13.947394,12.513797,11.551778,11.514051,13.174006,15.652621,18.21046,19.783646,19.896824,18.693357,18.33873,17.640795,17.165443,17.154125,17.501207,18.644312,18.761265,18.915941,19.334703,19.410156,3.0822346,3.4859054,3.1010978,2.9351022,3.4029078,4.3196554,3.3915899,2.5087957,1.8787673,1.4298248,0.80734175,0.5772116,0.362172,0.23390275,0.18485862,0.1358145,0.17354076,0.32067314,0.44894236,0.63002837,1.1280149,1.1657411,0.935611,0.694163,0.6488915,0.9922004,1.5279131,2.003264,2.5314314,3.1463692,3.7688525,3.2821836,3.3048196,3.6179473,3.942393,3.9688015,3.5538127,3.519859,3.92353,4.4743333,4.5460134,3.4481792,2.3390274,1.7052265,1.6033657,1.6788181,1.5203679,1.5618668,1.5580941,1.4335974,1.3128735,1.7165444,3.187868,4.991183,6.6360474,7.91874,7.6886096,6.017337,4.6516466,4.561104,5.9494295,8.356364,11.053791,15.916705,21.171972,21.390783,20.123182,22.424482,23.016785,21.998177,24.842735,27.07613,27.872154,27.725021,26.55928,23.726038,24.872917,24.940825,22.133991,16.980585,12.3289385,9.435335,7.092535,5.304311,4.402653,5.0515447,4.8553686,4.5761943,4.255521,4.0178456,4.0895257,4.187614,3.5877664,3.3689542,3.4896781,2.806833,2.5616124,3.2520027,3.4745877,2.886058,2.2296214,2.9841464,3.2105038,3.399135,3.5575855,3.2029586,1.9844007,1.9429018,1.8636768,1.2902378,0.5357128,0.41121614,0.34330887,0.26408374,0.16976812,0.120724,0.09808825,0.1358145,0.18485862,0.20372175,0.1659955,0.41121614,0.5017591,0.5055317,0.47912338,0.44139713,0.73566186,1.0751982,1.2147852,1.0789708,0.76207024,0.29803738,0.40367088,1.3845534,2.4371157,1.6184561,1.2261031,1.0110635,0.9620194,1.0827434,1.388326,1.0223814,0.5281675,0.19994913,0.14335975,0.29049212,0.7054809,1.1204696,1.2223305,1.0186088,0.8224323,0.8111144,0.9997456,0.9393836,0.6413463,0.58098423,0.58098423,0.6451189,0.77716076,1.0601076,1.6335466,2.6106565,2.41448,1.6335466,0.80356914,0.41121614,0.9507015,2.0636258,3.9725742,5.956975,6.349328,6.590776,7.0359454,7.6093845,8.729855,11.291467,13.917213,16.15438,17.908651,19.134754,19.866644,22.013268,22.379211,24.44661,28.909626,33.644268,30.143274,29.384975,30.98457,33.565044,34.760967,39.81251,44.56602,49.42516,54.69929,60.60722,61.278748,62.282265,64.72315,67.643166,68.00911,64.296844,58.977448,56.05366,56.974182,60.62231,57.841885,54.782288,50.455086,46.380653,46.599464,50.383408,56.219658,70.6424,94.80229,124.451355,91.40693,66.33784,66.33784,83.79378,86.39689,84.22008,82.7978,73.275696,58.468143,52.839386,89.535706,107.41418,89.16599,49.006397,32.686024,27.740112,23.016785,19.70442,19.051756,22.371666,16.109108,10.770844,6.0814714,4.745962,12.438345,7.5188417,5.5080323,5.873977,6.688864,4.640329,5.7117543,5.13077,3.5990841,2.1994405,2.3956168,3.410453,3.9914372,3.9989824,3.8103511,4.3347464,4.7120085,4.5950575,4.236658,3.8292143,3.5236318,3.440634,3.821669,5.0553174,6.820906,8.103599,9.578695,11.385782,12.879742,12.755245,9.031664,8.0206,7.383027,7.2660756,7.5301595,7.752744,9.631512,10.34831,10.457717,10.748209,12.238396,14.007756,17.097536,18.840488,18.444365,16.969267,17.101309,16.33924,16.33924,16.414692,13.536179,15.120681,14.675511,12.826925,10.469034,8.7600355,11.555551,11.41219,11.427281,13.35132,17.56157,18.063328,19.542198,20.368402,20.202406,20.017548,20.519308,21.232334,21.296469,20.470263,19.104572,17.112627,17.120173,17.071129,17.240896,20.232588,15.99593,13.27964,12.525115,12.593022,10.785934,8.933576,7.7904706,7.643338,8.401636,9.597558,10.514306,12.242168,13.238141,12.559069,9.87296,6.5643673,4.821415,6.25124,8.929804,7.4169807,4.644101,11.77059,13.7851715,11.242422,20.26277,9.009028,9.80128,7.914967,1.7354075,2.7615614,26.065065,22.7527,11.344283,3.2633207,2.8219235,2.04099,1.7542707,4.063117,9.64283,17.746428,23.069601,23.748674,20.98334,17.674747,18.417955,20.662666,21.424738,20.8513,19.572378,18.693357,13.517315,12.019584,12.7477,13.04951,9.0957985,9.669238,11.962994,14.366156,15.422491,13.826671,12.276122,13.041965,14.290704,15.316857,16.524097,17.025856,15.769572,13.400364,11.385782,12.0082655,11.642321,10.287949,11.042474,13.306048,12.755245,7.7037,9.14107,9.639057,8.563859,12.053536,8.820397,5.3646727,5.8966126,10.106862,13.185325,14.66042,12.740154,11.996947,13.664448,15.641303,11.649866,10.329447,9.525878,8.345046,7.17176,14.996184,19.304522,18.297232,15.022593,17.365393,18.168962,17.346529,15.79598,14.562332,14.830189,13.245687,13.58145,13.958713,13.739901,13.521088,14.313339,16.633503,17.923742,16.923996,13.702174,13.177779,12.359119,12.457208,13.332457,13.502225,10.7557535,10.31813,9.846551,8.786444,8.345046,6.858632,5.6061206,4.878004,4.5912848,4.2706113,3.9801195,3.62172,3.1237335,2.4182527,1.478869,1.1506506,1.0487897,1.026154,1.0299267,1.1129243,0.91674787,0.7432071,0.7167987,0.80734175,0.80734175,0.62625575,0.6073926,0.6451189,0.68661773,0.7469798,0.62625575,0.8224323,1.0299267,1.0978339,1.0374719,0.9280658,0.80734175,0.77338815,0.8224323,0.87147635,1.1016065,1.0789708,1.0525624,1.1393328,1.297783,1.4939595,1.8070874,2.0070364,2.003264,1.8297231,1.659955,1.8938577,2.214531,2.5502944,3.0520537,3.893349,4.2517486,3.9461658,3.048281,1.8787673,2.0598533,2.3880715,2.5917933,2.5314314,2.2296214,2.7389257,3.2067313,3.4330888,3.4896781,3.7084904,4.7572803,5.6513925,6.3116016,6.7643166,7.141579,8.778898,10.001229,10.227587,9.601331,9.001483,8.843033,8.394091,8.043237,7.835742,7.432071,7.515069,7.9225125,8.367682,8.635539,8.575176,9.110889,9.303293,8.741172,7.7225633,7.232122,7.356619,6.7643166,5.6325293,4.3649273,3.5689032,3.0445085,2.867195,2.9728284,3.1237335,2.9313297,2.3201644,2.2409391,2.4182527,2.5276587,2.1956677,2.0372176,2.2371666,2.354118,2.3880715,2.776652,3.5085413,4.0404816,4.2592936,4.217795,4.1197066,3.85185,3.6481283,3.6292653,3.6481283,3.2972744,3.199186,2.927557,2.6106565,2.3616633,2.2899833,2.022127,2.1013522,2.4408884,2.897376,3.2670932,3.2520027,3.361409,3.4217708,3.3463185,3.1124156,3.0897799,3.127506,3.127506,3.1463692,3.4029078,3.682082,3.361409,2.6823363,1.8938577,1.237421,0.8224323,0.67152727,0.56212115,0.41876137,0.32067314,0.45648763,0.7092535,0.8601585,0.91674787,1.1129243,1.0035182,1.297783,1.5241405,1.3656902,0.65643674,0.694163,0.6451189,0.5055317,0.35839936,0.38103512,0.44139713,0.66775465,0.9242931,1.1996948,1.6033657,2.1654868,2.4522061,2.8709676,3.3312278,3.2331395,3.2105038,3.1237335,3.1576872,3.5387223,4.5007415,4.478106,4.4630156,4.4177437,4.38379,4.4705606,4.4705606,4.745962,5.311856,5.8928404,5.904158,6.198423,7.2057137,8.103599,8.854351,10.208723,11.197151,11.106608,10.280403,9.416472,9.537196,9.280658,8.409182,7.643338,7.1566696,6.6058664,5.704209,4.67051,4.055572,3.7877154,3.187868,3.1765501,3.5236318,3.802806,3.983892,4.425289,4.927048,4.8402777,4.606375,4.2819295,3.5236318,3.108643,3.4745877,4.2291126,5.2288585,6.560595,7.3679366,8.575176,9.57115,10.095545,10.253995,10.695392,11.736636,13.041965,14.177525,14.618922,15.056546,15.773345,15.98084,15.380992,14.158662,13.415455,12.113899,11.148107,11.257513,13.015556,14.369928,16.237377,17.599297,17.886015,16.984358,16.935314,16.675003,16.505234,16.682549,17.440845,18.221779,19.078165,19.73083,19.934551,19.470518,2.6785638,2.927557,2.8822856,2.837014,2.9501927,3.2670932,2.3201644,1.5958204,1.2449663,1.1355602,0.845068,0.48666862,0.3055826,0.28294688,0.30935526,0.22258487,0.23013012,0.23013012,0.3734899,0.65643674,0.935611,0.7167987,0.79602385,0.76207024,0.59230214,0.663982,1.4826416,2.1353056,2.3993895,2.5125682,3.1954134,3.3915899,3.2482302,3.1840954,3.229367,3.0407357,3.5047686,4.3007927,5.323174,6.398372,7.281166,6.952948,4.719554,2.806833,2.0560806,1.9240388,2.3201644,2.4672968,2.3465726,2.0673985,1.8372684,1.2525115,1.9466745,2.848332,3.259548,2.8407867,3.9688015,4.3007927,4.7572803,5.2288585,4.5724216,7.0170827,9.06939,10.921749,12.755245,14.750964,18.4255,22.020813,23.533634,23.046967,22.718748,21.620914,22.186808,22.869654,22.869654,22.115128,24.503199,24.024076,21.066338,17.455936,16.467508,11.827179,8.643084,6.628502,5.7607985,6.270103,5.723072,5.2552667,5.3759904,5.6551647,4.7233267,4.636556,3.4557245,2.5201135,2.3088465,2.4672968,2.203213,2.4484336,2.8822856,3.240685,3.3123648,3.591539,3.3915899,3.4594972,3.5990841,2.6785638,1.6750455,1.6071383,1.7995421,1.7919968,1.3392819,0.77716076,0.46026024,0.38858038,0.4074435,0.23013012,0.16976812,0.17731337,0.2678564,0.3470815,0.20372175,0.33953625,0.4979865,0.52439487,0.41876137,0.34330887,0.5017591,0.8337501,1.2449663,1.6071383,1.7882242,1.5279131,1.1921495,1.1544232,1.2525115,0.77338815,0.7054809,0.52062225,0.49421388,0.6790725,0.875249,0.41121614,0.20749438,0.1659955,0.25276586,0.4979865,0.5319401,0.9922004,1.3317367,1.3128735,0.9808825,0.8941121,1.1280149,1.116697,0.80734175,0.6790725,1.1053791,0.9280658,0.935611,1.5052774,2.595566,6.1116524,5.13077,2.9501927,1.3505998,0.6073926,0.65643674,1.3053282,2.8785129,4.798779,5.5797124,5.304311,6.3455553,8.303548,11.295239,15.965749,16.4826,18.8254,22.024584,24.838963,25.72553,26.51778,25.895298,26.857317,30.116865,34.123394,34.945824,33.436775,31.471237,30.584671,31.97677,37.22449,42.649525,51.402016,62.221905,69.40875,67.337585,64.49303,61.86728,60.42991,61.135387,59.00763,53.767452,49.84015,50.722942,58.962357,56.706326,52.28858,46.806957,41.9365,39.9106,46.127888,55.140686,70.536766,92.21427,116.40812,92.97257,69.148445,65.089096,78.19143,83.088295,106.214485,148.72443,156.3904,118.532104,68.0242,89.6338,101.596794,85.89513,50.492813,29.328386,23.650587,19.806282,16.735365,14.709465,15.328176,9.835234,5.5759397,4.3083377,6.8737226,13.204187,6.9755836,5.0062733,6.515323,8.575176,6.1041074,4.346064,3.338773,2.5691576,2.11267,2.6408374,3.078462,3.5538127,3.5764484,3.2444575,3.2218218,3.5123138,3.5349495,3.410453,3.2105038,2.9766011,3.2331395,3.7198083,4.9157305,6.470052,7.224577,7.8206515,12.249713,15.863888,16.060064,12.279895,10.269085,8.262049,7.61693,8.050782,7.654656,9.827688,9.144843,8.643084,9.699419,12.019584,13.981348,17.742655,19.606333,19.383747,20.398582,19.436563,17.787928,16.867407,16.35433,14.158662,14.600059,13.008011,10.70671,8.495952,6.609639,9.650374,10.767072,10.782163,11.359374,15.022593,19.21398,20.270313,20.458946,19.889278,16.505234,17.77661,19.059301,19.58747,19.700647,20.873934,20.281631,21.647322,20.617395,17.18808,15.705438,14.252977,13.35132,12.966512,12.1252165,8.922258,7.5716586,6.771862,7.5565677,9.491924,10.646348,11.446144,12.811834,14.181297,14.452927,11.98563,8.371455,5.8098426,6.085244,7.537705,5.0477724,18.342503,12.864652,5.6589375,5.7306175,14.037937,6.2097406,5.3873086,4.3875628,4.5912848,15.90916,9.280658,8.624221,7.7150183,4.6516466,1.8599042,3.187868,2.5201135,3.180323,6.541732,12.019584,13.505998,14.532151,15.433809,17.425755,22.60557,22.975286,19.527107,17.04472,16.59955,15.554533,12.223305,9.491924,8.76758,9.49947,9.167479,8.326183,7.967784,8.182823,8.341274,7.073672,6.7454534,9.001483,12.313848,14.498198,12.717519,12.181807,13.045737,13.245687,11.951676,9.567377,11.974312,12.287439,13.45318,14.641558,11.242422,10.525623,10.080454,9.242931,7.967784,6.828451,5.956975,4.719554,6.643593,11.544232,15.539442,14.1926155,13.860624,13.396591,12.860879,13.528633,10.31813,9.808825,9.484379,9.133525,10.868933,12.045992,14.48688,15.135772,14.068119,14.494425,16.444872,18.233097,17.006994,14.037937,14.747191,15.973294,15.494171,14.93205,14.739646,14.226569,14.237886,14.713238,16.931541,19.319613,17.425755,16.810818,15.056546,13.996439,13.856852,13.234368,12.1101265,11.974312,11.257513,9.831461,8.98262,8.07719,6.673774,5.696664,5.221313,4.45547,4.112161,3.7462165,3.1124156,2.2786655,1.6033657,1.4373702,1.2411937,1.1959221,1.2487389,1.0902886,0.88279426,0.72811663,0.7130261,0.8337501,0.9922004,0.95447415,0.8186596,0.6187105,0.47912338,0.6375736,0.7507524,0.77338815,0.90543,1.0487897,0.7922512,0.7696155,0.7092535,0.7054809,0.7809334,0.91674787,1.2562841,1.20724,1.1732863,1.3204187,1.5769572,1.3430545,1.6146835,1.7580433,1.6071383,1.478869,1.4637785,1.7052265,2.0900342,2.5729303,3.1614597,4.247976,4.52715,3.9159849,2.757789,1.841041,1.9240388,2.4220252,2.4974778,2.2296214,2.6182017,3.2105038,3.832987,4.357382,4.6818275,4.745962,5.3080835,7.0585814,8.812852,9.876732,10.069136,10.680302,11.604594,11.7894535,10.944386,9.514561,8.643084,8.073418,7.752744,7.6093845,7.5301595,7.4396167,7.6093845,7.8395147,8.00551,8.062099,8.103599,8.284684,8.265821,7.8734684,7.122716,7.3717093,7.220804,6.3644185,4.9723196,3.682082,2.8709676,2.565385,2.674791,2.9313297,2.8822856,2.4069347,2.3767538,2.444661,2.372981,2.0145817,2.2447119,2.3013012,2.2711203,2.41448,3.169005,3.2935016,3.2935016,3.3123648,3.399135,3.4972234,2.9954643,2.5691576,2.6408374,3.0558262,3.1010978,2.9237845,2.4371157,1.9806281,1.7052265,1.5430037,1.267602,1.2562841,1.3958713,1.6109109,1.8599042,2.6597006,2.7804246,2.7426984,2.7426984,2.637065,3.3727267,3.8669407,4.0782075,4.134797,4.3422914,4.2894745,3.482133,2.5691576,1.8787673,1.3958713,0.8639311,0.55080324,0.41121614,0.38103512,0.38103512,0.42630664,0.56212115,0.70170826,0.8337501,1.0412445,1.2223305,1.2034674,1.0336993,0.7809334,0.52062225,0.47157812,0.41876137,0.35085413,0.3169005,0.41876137,0.663982,0.7394345,0.8299775,0.9997456,1.1883769,2.1013522,2.1390784,2.4522061,3.350091,4.29702,3.0218725,2.5767028,2.71629,3.2557755,4.074435,3.6594462,4.3385186,4.9987283,5.0854983,4.606375,4.6931453,5.010046,5.3948536,5.7004366,5.8211603,6.387054,6.832224,7.5226145,8.43559,9.144843,10.231359,10.502988,9.7069645,8.473316,8.29223,7.8696957,7.303802,6.7341356,6.0324273,4.798779,4.4630156,3.6556737,2.987919,2.71629,2.7238352,3.0558262,3.772625,4.496969,5.0062733,5.2288585,4.98741,4.3875628,3.7801702,3.3236825,2.9766011,2.6597006,3.229367,4.1989317,5.270357,6.330465,7.164215,7.8395147,8.424272,8.835487,8.83926,9.246704,10.352083,11.514051,12.449662,13.200415,14.558559,15.384765,15.592259,15.105591,13.856852,12.223305,10.967021,10.340765,10.63503,12.196897,13.249459,14.84528,16.097792,16.731592,17.067356,17.527617,17.957695,18.433046,18.881989,19.1008,18.406637,18.285913,18.62545,18.934805,18.334957,2.897376,2.5125682,2.2484846,2.1994405,2.305074,2.3277097,1.7995421,1.4675511,1.3204187,1.2185578,0.9016574,0.67152727,0.51684964,0.40367088,0.29049212,0.14335975,0.15845025,0.124496624,0.17731337,0.3470815,0.573439,0.46026024,0.63002837,0.6790725,0.58475685,0.67152727,1.5128226,2.3088465,2.6182017,2.516341,2.5767028,2.9803739,3.2067313,3.1199608,2.8143783,2.6068838,2.9954643,3.289729,3.8103511,4.6554193,5.704209,5.2326307,3.8593953,2.9501927,2.8030603,2.6332922,2.546522,2.474842,2.1051247,1.4977322,1.0714256,0.62248313,1.0487897,1.6750455,2.2409391,2.897376,3.6896272,4.4441524,5.2062225,6.156924,7.6131573,11.200924,12.777881,12.355347,11.415963,12.879742,19.772327,23.243143,23.145054,20.194862,15.988385,14.777372,15.150862,16.969267,19.278114,20.311813,21.90386,20.900343,17.991648,14.603831,12.90615,10.70671,9.646602,8.458225,7.043491,6.4926877,6.417235,5.4778514,5.2967653,5.7796617,5.13077,3.8367596,2.7313805,2.1956677,2.323937,2.9011486,3.3651814,3.138824,3.1916409,3.572676,3.410453,4.08198,4.3800178,4.2781568,3.7198083,2.6219745,2.1654868,1.9429018,1.6712729,1.3468271,1.237421,1.1544232,0.73566186,0.4074435,0.29803738,0.21503963,0.20749438,0.17731337,0.17731337,0.1961765,0.1961765,0.23767537,0.38103512,0.4376245,0.38480774,0.35839936,0.3470815,0.46026024,0.6752999,0.965792,1.2864652,1.569412,1.3166461,0.94692886,0.6451189,0.362172,0.35462674,0.23767537,0.211267,0.2867195,0.32821837,0.15467763,0.116951376,0.20372175,0.3470815,0.44894236,0.36594462,0.6752999,0.935611,0.94692886,0.7582976,0.86770374,1.0374719,1.2034674,1.146878,0.52062225,0.9016574,0.7054809,0.80356914,1.4449154,2.233394,4.5837393,3.640583,2.2748928,1.7278622,1.6184561,0.965792,1.1695137,2.173032,3.482133,4.187614,4.4516973,4.8742313,6.187105,8.6581745,12.098808,14.856597,19.395065,25.914162,31.286379,29.06053,28.215462,26.464964,25.291677,25.657623,28.007969,32.88597,34.900555,32.72752,28.389004,27.253443,34.138485,39.684242,47.003136,55.985756,63.28956,61.203297,59.501842,56.578056,53.759907,55.306683,60.3205,56.762917,51.17566,49.27048,55.9103,58.268192,54.03531,48.20283,42.54012,35.609806,39.835148,49.926918,66.11148,86.64588,107.840485,92.82921,70.483955,63.806408,74.309395,82.05082,123.77228,190.48361,221.46819,190.08371,103.78869,100.06511,99.344536,82.54126,51.228474,27.645796,20.798481,20.77962,19.263023,14.811326,12.898605,6.1418333,10.080454,12.185578,9.665465,9.480607,6.1078796,4.0782075,5.138315,7.466025,5.6815734,3.4670424,2.625747,2.1277604,1.7844516,2.2711203,2.8256962,3.150142,3.1425967,2.837014,2.3767538,2.595566,2.5691576,2.5314314,2.5314314,2.444661,2.8898308,3.500996,4.715781,6.2814207,7.277394,7.3415284,11.302785,15.513034,16.976812,13.358865,11.317875,9.024119,8.126234,8.397863,7.7376537,9.597558,8.458225,7.696155,8.809079,11.431054,13.196642,16.58446,18.866898,19.719511,21.209698,19.221525,18.033148,17.36162,16.67123,15.165953,12.966512,10.740664,8.941121,7.496206,5.80607,6.881268,8.537451,9.87296,10.925522,12.694883,16.18456,18.044466,18.312323,17.033401,14.252977,18.549997,19.417702,19.059301,18.900852,19.58747,21.013521,22.537663,21.779364,18.587723,15.030138,14.618922,13.460726,12.653384,11.898859,9.533423,8.137552,8.201687,8.6732645,9.205205,10.140816,10.465261,11.834724,13.88326,15.022593,12.438345,8.993938,7.4697976,6.700182,5.7872066,4.1083884,13.902123,8.688355,5.9682927,10.823661,15.912932,7.2283497,4.1612053,2.6068838,4.3347464,16.98813,7.2057137,14.743419,15.214996,5.723072,4.82896,5.168496,4.104616,4.534695,6.934085,9.352338,10.612394,14.460471,18.802763,23.307278,29.381203,22.326395,16.28265,13.170234,12.332711,10.559577,9.21275,6.6850915,5.8098426,6.937857,7.914967,6.006019,4.9647746,4.247976,3.5877664,2.9954643,2.9954643,4.961002,8.07719,10.974566,11.736636,10.967021,10.801025,11.34051,12.174261,12.400619,12.510024,11.69891,12.064855,12.955194,10.929295,10.091772,9.137298,8.050782,7.0548086,6.56814,5.772116,3.5953116,4.3309736,8.835487,14.517061,16.003475,16.124199,14.634012,12.242168,10.593531,10.087999,9.480607,8.922258,8.597813,8.692128,10.518079,13.664448,16.625957,17.614386,14.558559,14.754736,16.62973,16.392056,14.449154,15.418718,17.01831,16.535416,15.792209,15.584714,15.686575,15.584714,16.146835,18.097282,20.206179,19.270569,18.014284,16.078928,14.498198,13.641812,13.196642,12.366665,12.540206,12.076173,10.710483,9.559832,8.473316,6.952948,5.96452,5.560849,4.8855495,4.327201,3.7990334,3.059599,2.2409391,1.8334957,1.5128226,1.2902378,1.2411937,1.2751472,1.1280149,0.8941121,0.72811663,0.7205714,0.845068,0.935611,1.0110635,0.9507015,0.73188925,0.5055317,0.5998474,0.77338815,0.7997965,0.8639311,0.9242931,0.724344,0.68661773,0.6752999,0.694163,0.73566186,0.7922512,1.1732863,1.2864652,1.2110126,1.1053791,1.20724,1.2261031,1.5543215,1.6637276,1.4637785,1.3355093,1.3505998,1.5279131,1.9391292,2.5201135,3.0331905,3.572676,3.380272,2.7879698,2.1503963,1.8297231,1.6071383,1.9957186,2.2220762,2.1843498,2.4597516,2.8936033,3.8895764,4.738417,4.9987283,4.4630156,5.138315,6.752999,8.926031,10.816116,11.133017,10.770844,11.427281,12.321393,12.408164,10.386037,8.477088,7.7904706,7.707473,7.752744,7.564113,7.7301087,7.9262853,7.9753294,7.907422,7.960239,7.816879,7.7301087,7.673519,7.5527954,7.2057137,7.281166,7.01331,6.368191,5.383536,4.1574326,3.0709167,2.516341,2.4899325,2.727608,2.7238352,2.3993895,2.4786146,2.5125682,2.3163917,1.9504471,2.191895,2.323937,2.4069347,2.6182017,3.2557755,3.5462675,3.4632697,3.2972744,3.2331395,3.3425457,2.8521044,2.6446102,2.7200627,2.9086938,2.886058,2.3692086,1.8599042,1.5316857,1.3845534,1.2751472,1.1846043,1.1242423,1.0714256,1.0601076,1.1544232,1.6486372,1.9429018,2.263575,2.4861598,2.1051247,2.6144292,3.6028569,4.3083377,4.4215164,4.08198,3.7650797,2.867195,1.9806281,1.3958713,1.086516,0.7092535,0.513077,0.43385187,0.44139713,0.55080324,0.6149379,0.6149379,0.6413463,0.724344,0.8224323,0.95447415,0.90920264,0.7507524,0.55457586,0.41498876,0.36971724,0.3961256,0.41121614,0.41498876,0.45648763,0.73188925,0.8601585,0.94692886,1.0714256,1.2562841,2.0372176,2.1013522,2.493705,3.3840446,4.0480266,3.3915899,2.9200118,2.6219745,2.5691576,2.9426475,2.9426475,3.4179983,4.327201,5.13077,4.7950063,4.8968673,5.1081343,5.413717,5.7306175,5.926794,5.8211603,5.783434,6.3455553,7.432071,8.329956,9.333474,9.4013815,8.714764,7.7942433,7.484888,7.2924843,6.8850408,6.462507,5.87775,4.640329,3.9122121,3.1840954,2.6408374,2.4031622,2.5276587,2.9728284,3.8254418,4.7006907,5.2137675,4.983638,4.45547,4.104616,3.6896272,3.127506,2.516341,2.5087957,3.5123138,4.5196047,5.240176,6.096562,6.6850915,6.9491754,7.2887115,7.8017883,8.29223,9.046755,10.167224,11.02361,11.563096,12.325166,13.494679,14.4114275,14.898096,14.7321005,13.604086,11.653639,10.367173,10.072908,10.804798,12.294985,13.490907,15.131999,16.67123,17.882242,18.866898,18.991394,19.032892,19.240387,19.47429,19.21398,18.92726,18.685812,18.463226,18.289686,18.233097,2.7728794,2.1353056,1.8523588,1.9051756,2.0560806,1.841041,1.6260014,1.5580941,1.5316857,1.4071891,1.0223814,0.9997456,0.8526133,0.5772116,0.3055826,0.30181,0.21881226,0.124496624,0.071679875,0.09808825,0.23767537,0.2678564,0.40367088,0.47912338,0.482896,0.58098423,1.2864652,2.0296721,2.4408884,2.4597516,2.3201644,2.546522,2.9200118,2.8822856,2.4333432,2.1353056,2.0787163,1.8674494,1.9127209,2.3503454,3.048281,2.584248,2.2711203,2.4823873,2.9916916,2.9615107,2.4031622,2.1843498,1.7542707,1.0487897,0.4678055,0.65643674,1.2902378,1.8674494,2.565385,4.2291126,5.3910813,6.63982,8.039464,9.865415,12.593022,14.713238,14.879233,13.487134,12.340257,14.68683,22.688566,25.646305,23.488363,17.810562,11.876224,10.653893,10.827434,13.36641,17.584206,21.122927,20.847527,18.12369,14.815099,12.012038,10.023865,9.623966,9.899368,8.76758,6.432326,5.3910813,5.4476705,4.779916,4.772371,5.3873086,5.172269,4.2328854,3.4368613,2.9539654,3.0181,3.9084394,5.0968165,4.5120597,4.123479,4.3309736,3.9801195,4.323428,4.7648253,4.6516466,3.7952607,2.4672968,2.3428001,2.0447628,1.5656394,1.1053791,1.0751982,1.0751982,0.72811663,0.48666862,0.51684964,0.6790725,0.724344,0.5470306,0.331991,0.19994913,0.19994913,0.211267,0.2565385,0.27917424,0.28294688,0.32067314,0.29426476,0.2678564,0.28294688,0.38103512,0.59607476,1.1996948,1.2902378,1.1091517,0.8262049,0.5357128,0.29049212,0.14335975,0.10940613,0.1358145,0.08677038,0.124496624,0.116951376,0.181086,0.29803738,0.29426476,0.35839936,0.73188925,0.8224323,0.59230214,0.573439,0.9242931,1.0223814,1.1657411,1.1921495,0.4640329,0.6752999,0.5885295,0.72811663,1.1393328,1.3845534,2.04099,1.5807298,1.418507,1.8787673,2.173032,2.41448,2.203213,2.2975287,2.8407867,3.3463185,3.7952607,3.942393,4.5988297,6.047518,8.043237,12.491161,17.844517,24.586197,30.731804,31.810774,29.856554,27.34776,24.7786,23.092237,23.661903,27.260988,31.293924,30.731804,26.498919,25.487854,31.667414,36.466194,41.646008,47.127632,51.013435,49.096943,49.34971,49.05167,47.829338,47.67089,57.015682,58.079563,54.95583,51.945274,53.537323,56.42715,52.967655,47.51244,41.513966,33.516,35.639988,45.40354,60.297867,77.51613,93.94214,89.3018,71.2083,64.040306,73.581276,87.02314,132.20033,202.41643,65535.0,231.29964,134.34695,111.97528,102.23437,83.510826,53.382645,28.622906,21.896315,22.356575,20.104319,13.792717,10.612394,5.523123,12.830698,14.490653,7.816879,5.451443,4.7120085,3.4142256,4.085753,5.96452,4.979865,3.1727777,2.7011995,2.214531,1.7014539,2.4823873,2.7087448,2.7691069,2.848332,2.8407867,2.3578906,2.1315331,1.9466745,1.8787673,1.8938577,1.8599042,2.4069347,3.380272,4.821415,6.405917,7.462252,7.3113475,10.220041,14.234114,16.663685,14.071891,12.1101265,9.937095,8.8769865,8.89585,8.616675,9.684328,8.590267,7.699928,8.284684,10.510533,12.279895,14.966003,17.225805,18.878216,20.904116,19.089483,19.047983,19.342249,18.908396,17.04472,12.577931,10.121953,8.963757,8.209232,6.7643166,5.692891,6.9869013,9.514561,11.800771,12.034674,13.038192,14.649103,14.852824,13.513543,12.370438,16.218515,17.278622,17.414436,18.161417,20.756983,21.620914,22.484844,22.14531,20.225042,17.172989,16.825907,14.777372,14.094527,14.739646,13.562587,11.004747,10.8576145,10.329447,9.235386,9.963503,9.408927,10.412445,12.657157,14.449154,12.706201,9.507015,8.412953,7.1906233,6.006019,7.4207535,7.699928,5.2665844,7.273621,13.358865,15.645076,8.831716,4.436607,3.6934,7.0548086,14.188843,9.771099,19.210207,17.803017,5.6853456,7.84706,8.3525915,8.22055,8.741172,9.835234,10.072908,14.958458,18.980076,22.156626,24.99364,28.487091,17.825653,11.604594,8.643084,7.4811153,6.3531003,5.6815734,4.115934,3.7462165,4.727099,5.2590394,3.8103511,2.7917426,2.0296721,1.4713237,1.1846043,1.1053791,2.0749438,3.904667,6.2021956,8.367682,8.511042,8.333729,9.103344,10.79348,12.113899,11.076427,10.306811,10.834979,11.778135,10.336992,9.34102,8.816625,8.00551,7.122716,7.3717093,5.5193505,3.3161373,3.078462,5.9682927,12.027128,17.056038,17.086218,14.769827,11.827179,9.073163,9.582467,9.163706,8.771353,8.495952,7.575431,11.057564,13.807808,15.803526,16.524097,14.924504,14.2944765,14.554788,14.709465,14.747191,15.614895,15.641303,16.052519,16.531643,16.716501,16.180788,17.293713,18.033148,18.840488,19.519562,19.210207,17.70493,16.071383,14.671739,13.822898,13.800262,12.83447,13.117417,12.823153,11.517824,10.182315,8.922258,7.2358947,6.1418333,5.7607985,5.330719,4.7233267,4.115934,3.240685,2.3088465,2.0372176,1.6033657,1.448688,1.3732355,1.2826926,1.1581959,0.8941121,0.7922512,0.83752275,0.935611,0.875249,0.8941121,0.91297525,0.784706,0.58475685,0.5998474,0.7130261,0.784706,0.8639311,0.90543,0.784706,0.6828451,0.69039035,0.6828451,0.633801,0.62248313,0.95824677,1.2261031,1.1996948,0.9695646,0.9507015,1.116697,1.3430545,1.3920987,1.2751472,1.2713746,1.3053282,1.4335974,1.7957695,2.305074,2.6483827,2.7238352,2.3767538,2.022127,1.8334957,1.7580433,1.4600059,1.6260014,1.8184053,1.8561316,1.8146327,2.1315331,2.9237845,3.5462675,3.6481283,3.1840954,3.7047176,4.821415,7.1000805,9.850324,11.09529,10.687846,11.057564,12.223305,13.196642,11.970539,9.831461,8.586494,7.9828744,7.6584287,7.115171,7.8508325,8.27714,8.273367,7.9300575,7.564113,7.5037513,7.462252,7.3453007,7.175533,7.0887623,7.066127,6.8058157,6.360646,5.6400743,4.395108,3.270866,2.6068838,2.4484336,2.6144292,2.704972,2.3578906,2.4107075,2.5012503,2.4408884,2.2069857,2.3993895,2.565385,2.7841973,3.1161883,3.5839937,3.8178966,3.7914882,3.5689032,3.308592,3.2369123,2.8822856,2.806833,2.8407867,2.837014,2.655928,1.9466745,1.50905,1.3204187,1.2713746,1.1732863,1.1883769,1.2562841,1.2223305,1.1016065,1.086516,1.0751982,1.3091009,1.6825907,1.9542197,1.7693611,1.9806281,3.078462,3.9008942,3.9008942,3.1199608,2.6295197,2.0070364,1.4675511,1.0902886,0.80734175,0.59230214,0.52062225,0.5055317,0.5319401,0.6488915,0.66775465,0.63002837,0.633801,0.6828451,0.7167987,0.80356914,0.7582976,0.62625575,0.4979865,0.49421388,0.43007925,0.41498876,0.4376245,0.47912338,0.4979865,0.7922512,0.95824677,1.1091517,1.2713746,1.3732355,1.9089483,1.9844007,2.2975287,2.938875,3.410453,3.2369123,2.776652,2.3918443,2.2748928,2.4899325,2.5087957,2.637065,3.3840446,4.4441524,4.67051,4.7610526,5.0666356,5.5004873,5.8136153,5.59103,5.330719,5.243949,5.7004366,6.647365,7.6093845,7.9526935,7.835742,7.5263867,7.2094865,6.9793563,6.952948,6.620957,6.1531515,5.4778514,4.2517486,3.3953626,2.8030603,2.4031622,2.1956677,2.263575,3.0105548,3.9763467,4.8025517,5.1081343,4.4630156,3.7499893,3.5877664,3.350091,2.8256962,2.2484846,2.474842,3.6179473,4.6214657,5.2099953,5.8664317,6.25124,6.3531003,6.6322746,7.2472124,8.035691,8.771353,9.593785,10.159679,10.578441,11.415963,12.649611,13.702174,14.283158,14.177525,13.230596,11.593277,10.336992,10.1294985,11.00852,12.370438,13.981348,15.988385,17.897333,19.346022,20.130728,19.493153,18.723537,18.429274,18.591496,18.565088,19.051756,19.002712,18.715992,18.534906,18.844261,2.214531,1.8674494,1.8334957,1.9881734,2.0749438,1.6976813,1.5618668,1.5807298,1.6033657,1.50905,1.20724,1.2261031,1.0676528,0.7092535,0.38103512,0.58475685,0.35839936,0.18863125,0.090543,0.049044125,0.0452715,0.1056335,0.17731337,0.24899325,0.30935526,0.3772625,0.9318384,1.5430037,1.9844007,2.2183034,2.3918443,2.3428001,2.3993895,2.282438,1.9429018,1.5430037,1.2298758,1.0374719,1.0035182,1.0978339,1.1996948,1.0714256,1.1808317,1.6335466,2.2069857,2.3616633,1.8334957,1.6712729,1.4335974,0.9808825,0.48666862,1.20724,2.3126192,3.0331905,3.5689032,5.0854983,6.8661776,8.529905,10.691619,13.109872,14.698147,13.426772,12.347801,11.751727,12.717519,17.112627,24.405111,26.763002,23.609087,17.195625,12.623203,11.491416,12.37421,15.433809,20.013775,24.623924,22.062311,16.705183,12.536433,10.804798,10.038955,9.578695,9.7069645,7.9941926,4.9044123,3.7990334,3.5689032,3.8707132,4.5422406,5.1345425,4.9421387,5.485397,4.9723196,4.1762958,3.953711,5.2326307,6.360646,5.621211,5.2099953,5.5985756,5.534441,4.2328854,4.1310244,4.244203,3.8782585,2.637065,2.3880715,2.0485353,1.8976303,1.8636768,1.5015048,0.8262049,0.5055317,0.56212115,0.87902164,1.20724,1.3053282,1.0223814,0.66020936,0.38480774,0.24522063,0.23390275,0.17354076,0.14713238,0.17354076,0.21881226,0.2867195,0.26408374,0.24522063,0.26408374,0.29426476,0.8186596,1.2185578,1.4335974,1.3770081,0.965792,0.39989826,0.14713238,0.11317875,0.181086,0.20749438,0.18863125,0.15467763,0.13204187,0.14335975,0.181086,0.452715,0.9620194,0.935611,0.47535074,0.5357128,0.95824677,1.0638802,1.0827434,1.0299267,0.69793564,0.7205714,0.7167987,0.73566186,0.7469798,0.62625575,0.5696664,0.63002837,1.1657411,2.1466236,3.1576872,5.036454,4.4931965,3.731126,3.5764484,3.4745877,3.4934506,3.9197574,4.696918,5.8173876,7.3377557,11.45369,16.248695,20.587215,25.269043,32.995377,31.550463,28.732311,25.574625,23.145054,22.56407,21.107838,24.257978,25.865116,25.208681,26.993132,30.282862,33.65936,36.6171,38.37514,37.880928,36.658596,37.805473,40.978252,43.72095,41.44983,49.225212,53.81272,55.208595,53.974945,51.23979,49.859013,47.15027,42.664616,37.15658,32.59548,34.67797,43.558727,55.23123,66.74151,76.203255,81.71129,71.01589,66.01339,75.38459,94.59103,131.26094,188.49544,230.60925,225.56525,145.0197,118.67169,107.165184,87.40795,56.347927,30.969479,25.276588,22.141537,16.859861,9.982366,7.326438,6.9491754,11.506506,10.427535,4.183841,4.2781568,3.519859,3.2859564,4.2706113,5.624984,4.957229,3.5424948,3.1463692,2.516341,1.8938577,3.0181,2.704972,2.5238862,2.7728794,3.2067313,3.0558262,2.1843498,1.780679,1.5920477,1.4713237,1.3732355,1.8485862,3.187868,4.9044123,6.4549613,7.250985,7.092535,9.310839,12.551523,15.026365,14.539697,13.158916,11.189606,10.223814,10.378491,10.306811,10.442626,9.691874,9.001483,9.0543,10.26154,12.166716,14.490653,16.290195,17.84829,20.692848,19.681786,20.22127,21.138018,21.130472,18.761265,14.019074,11.793225,10.827434,10.106862,8.865668,6.7567716,7.062354,9.80128,12.913695,12.276122,11.276376,11.744182,11.744182,11.016065,10.948157,11.744182,15.369675,17.542706,18.968758,25.318087,23.967487,25.00496,25.25018,23.85808,22.315077,20.53817,17.308804,17.20317,19.851553,19.964731,16.097792,14.169979,12.045992,9.895596,10.178542,9.190115,9.525878,11.133017,13.008011,13.166461,10.442626,8.75249,7.6320205,8.00551,12.196897,6.2663302,5.7004366,8.43559,11.480098,10.917976,8.52236,5.0515447,8.099826,15.011275,12.879742,10.812344,14.667966,12.479843,5.9192486,10.295494,11.615912,13.011784,13.879487,13.917213,13.117417,22.601797,23.552498,21.956678,20.787165,19.99114,11.544232,6.9189944,4.4743333,3.4896781,4.1498876,2.8219235,2.2711203,2.5012503,2.9049213,2.263575,2.142851,1.3543724,1.0186088,1.1808317,0.80734175,0.58475685,0.69039035,1.1921495,1.991946,2.8106055,4.104616,5.3571277,6.7869525,7.9338303,7.6395655,8.186596,9.288202,10.876478,11.68382,9.25425,9.107117,9.5183325,9.25425,8.318638,7.9262853,4.9723196,4.123479,3.9348478,4.979865,9.831461,16.075155,16.014793,13.649357,11.136789,8.790216,8.541223,8.812852,9.050528,9.016574,8.7600355,11.589504,12.811834,11.876224,10.585986,13.075918,13.936077,12.857106,13.143826,14.875461,14.909414,13.472044,15.094273,16.663685,16.84477,16.06761,18.542452,18.881989,18.949896,19.002712,17.689838,16.505234,15.490398,14.762281,14.43029,14.637785,13.513543,13.630494,13.324911,12.106354,10.638803,9.574923,7.7640624,6.4436436,5.934339,5.666483,5.304311,4.6742826,3.6066296,2.4786146,2.2069857,1.7844516,1.7089992,1.5807298,1.3166461,1.1544232,0.8903395,0.8903395,1.0072908,1.0714256,0.88279426,0.7582976,0.80356914,0.77338815,0.6526641,0.6413463,0.6790725,0.7696155,0.91297525,1.0110635,0.8865669,0.73566186,0.72811663,0.66775465,0.543258,0.52062225,0.7469798,1.0525624,1.1355602,1.0035182,1.0110635,1.0110635,1.0072908,1.0110635,1.0601076,1.2487389,1.2826926,1.3845534,1.6373192,1.9579924,2.1013522,2.1503963,2.161714,2.1353056,2.0183544,1.7391801,1.5203679,1.4713237,1.4335974,1.3015556,1.0072908,1.2751472,1.3694628,1.3619176,1.3732355,1.5354583,1.6373192,2.3956168,4.779916,8.254503,10.785934,10.978339,11.106608,11.691365,12.679792,13.426772,12.174261,10.20495,8.503497,7.4018903,6.5945487,7.7112455,8.186596,8.190369,7.8017883,7.0057645,7.009537,7.2623034,7.2472124,6.9265394,6.730363,6.7831798,6.820906,6.560595,5.7872066,4.3196554,3.4217708,2.7992878,2.5767028,2.6936543,2.927557,2.4069347,2.2899833,2.474842,2.727608,2.6898816,2.8445592,2.938875,3.1425967,3.4934506,3.8895764,3.8593953,3.9461658,3.7952607,3.3953626,3.0709167,2.8747404,2.7615614,2.7653341,2.757789,2.4408884,1.7580433,1.418507,1.2902378,1.2562841,1.20724,1.1808317,1.4449154,1.5467763,1.4034165,1.3241913,1.1129243,1.0676528,1.086516,1.1959221,1.5430037,1.7995421,2.6483827,3.150142,2.8936033,1.9957186,1.4864142,1.2713746,1.177059,1.0412445,0.73188925,0.60362,0.56589377,0.573439,0.5998474,0.62248313,0.5470306,0.5885295,0.67152727,0.72811663,0.7167987,0.84129536,0.7469798,0.56589377,0.46026024,0.6149379,0.52439487,0.422534,0.4074435,0.49044126,0.58098423,0.8941121,1.0412445,1.2411937,1.448688,1.3505998,1.7089992,1.7882242,1.8825399,2.173032,2.7313805,2.4069347,2.1202152,2.2183034,2.637065,2.9200118,2.6144292,2.6295197,3.0256453,3.7047176,4.395108,4.4931965,5.0213637,5.560849,5.6589375,4.817642,5.081726,5.323174,5.7192993,6.3229194,7.0849895,6.5530496,6.3908267,6.4926877,6.6813188,6.700182,6.6586833,6.258785,5.5495315,4.5460134,3.2670932,2.727608,2.384299,2.11267,1.9164935,1.9164935,2.9237845,3.9650288,4.7233267,4.881777,4.0970707,3.2670932,3.0407357,2.7917426,2.3880715,2.1956677,2.5616124,3.4972234,4.4516973,5.172269,5.7117543,6.119198,6.304056,6.609639,7.1378064,7.7640624,8.13378,8.544995,9.001483,9.590013,10.533169,12.185578,13.313594,13.751218,13.426772,12.381755,11.268831,10.295494,10.084227,10.774617,12.019584,14.060574,16.42601,18.500954,19.783646,19.87796,18.700903,17.421982,16.825907,17.082445,17.73511,18.43682,18.648085,18.923487,19.364883,19.61765,2.0447628,1.9730829,1.7957695,1.6448646,1.5241405,1.3430545,1.3543724,1.5430037,1.5543215,1.388326,1.388326,0.9997456,0.8262049,0.6451189,0.422534,0.35085413,0.20372175,0.120724,0.08677038,0.071679875,0.0452715,0.0452715,0.08299775,0.1358145,0.24522063,0.48666862,1.0148361,1.81086,2.2409391,2.233394,2.3201644,2.3692086,1.9127209,1.5052774,1.3241913,1.1883769,1.3732355,1.4373702,1.3015556,1.0035182,0.68661773,0.5394854,0.513077,0.49421388,0.482896,0.58098423,0.52062225,0.5017591,0.48666862,0.48666862,0.6111652,1.1355602,2.6219745,4.006528,4.949684,5.828706,5.168496,5.2062225,5.9532022,6.8473144,6.7756343,5.2967653,6.4021444,8.771353,11.706455,15.135772,20.873934,22.096264,19.91946,16.588232,15.501716,17.663431,22.04722,26.55928,29.215208,28.151327,23.258234,16.13929,11.25374,9.65792,8.986393,9.035437,9.891823,9.016574,6.2399216,3.7386713,3.7499893,4.6516466,5.342037,5.330719,4.745962,4.4894238,4.112161,4.063117,4.7572803,6.5756855,6.0512905,5.3986263,5.80607,7.0849895,7.6584287,3.7914882,3.097325,3.610402,4.187614,4.515832,3.8103511,3.1199608,3.4066803,4.0782075,2.9916916,1.4147344,0.63002837,0.3470815,0.32821837,0.36594462,0.6111652,0.67152727,0.56212115,0.3772625,0.3055826,0.15845025,0.13204187,0.18485862,0.24522063,0.18485862,0.18485862,0.1659955,0.1659955,0.18485862,0.18485862,0.41498876,0.80356914,1.1581959,1.2562841,0.8563859,0.32821837,0.116951376,0.041498873,0.09808825,0.42630664,0.1961765,0.26408374,0.23390275,0.094315626,0.23013012,0.3734899,0.41121614,0.38103512,0.35462674,0.42630664,0.58475685,0.845068,1.1317875,1.3204187,1.237421,0.90543,0.73188925,0.543258,0.331991,0.26031113,0.32067314,0.5281675,1.2713746,3.2821836,7.6131573,8.360137,7.7037,6.9944468,6.2663302,4.2404304,4.0970707,4.2328854,5.455216,7.435844,8.744945,12.4307995,18.761265,23.98635,26.868635,28.68704,30.735577,27.725021,23.133736,19.685556,19.319613,17.206944,19.527107,22.899834,25.589716,27.479801,29.826374,31.784365,29.06053,24.024076,25.695349,28.966215,30.343224,35.545673,43.415367,45.927937,48.43296,46.044888,45.086643,46.47874,45.74685,42.01195,39.778557,36.632187,32.765247,30.961933,35.074093,43.554955,52.24708,58.74732,62.410534,70.367004,68.43165,68.593864,77.05209,94.17604,125.17193,162.3285,186.66948,181.47081,132.26447,115.61209,106.36162,87.04578,56.762917,31.12793,24.87669,18.931032,11.879996,5.594803,5.20245,7.8508325,12.955194,13.645585,9.808825,8.088508,4.2064767,3.5462675,5.1458607,6.971811,5.9192486,4.61392,3.410453,2.4559789,1.9579924,2.1503963,2.7238352,2.6597006,2.927557,3.5689032,3.6783094,2.7011995,2.0372176,1.6750455,1.5203679,1.3732355,1.3505998,2.3692086,3.942393,5.50426,6.40969,6.25124,7.54525,9.110889,10.729345,13.185325,14.539697,12.872196,12.792972,14.188843,12.238396,11.834724,11.77059,12.204442,12.789199,12.679792,14.094527,17.033401,18.693357,19.180025,21.50019,19.670467,18.368912,17.874697,17.931286,17.761518,16.063837,14.796235,13.185325,11.378237,10.453944,8.937348,8.367682,10.095545,12.385528,10.4049,9.820143,10.86516,11.408418,11.034928,11.046246,13.70972,24.178753,27.551481,24.17121,29.600016,29.441565,34.42143,36.598236,34.251663,31.859818,25.318087,19.908142,19.274342,22.820608,25.72553,22.90738,18.218006,13.513543,10.152134,9.016574,9.797507,10.038955,10.272858,11.080199,13.106099,11.778135,10.106862,9.06939,9.084481,10.023865,6.300284,10.178542,14.618922,14.652876,7.3415284,4.5460134,5.3910813,15.603577,26.627188,15.641303,8.073418,8.314865,9.337247,9.967276,14.86037,12.370438,13.04951,15.490398,17.48989,16.03743,25.069094,23.631723,20.07791,17.621931,14.313339,8.514814,5.1798143,3.2633207,2.565385,3.7235808,1.8184053,1.599593,2.0372176,2.1805773,1.1280149,0.7130261,0.63002837,0.7092535,0.7696155,0.6111652,0.3772625,0.32821837,0.40367088,0.5394854,0.68661773,1.1996948,1.9768555,3.4745877,5.100589,5.2326307,7.039718,9.205205,10.480352,10.291721,8.729855,8.141325,9.495697,10.167224,9.635284,9.476834,6.436098,5.1458607,4.889322,5.938112,9.552286,13.570132,13.86817,11.925267,9.205205,7.141579,7.8508325,8.484633,8.880759,8.771353,7.7829256,7.33021,9.495697,10.231359,8.5563135,6.590776,10.216269,11.216014,13.283413,15.773345,13.687083,14.517061,16.418465,15.214996,12.928786,17.77661,18.72731,18.636768,20.583443,22.194353,15.641303,14.735873,14.592513,14.524607,14.366156,14.464244,13.098554,12.838243,12.736382,12.079946,10.4049,9.869187,8.243186,6.832224,6.1418333,5.873977,5.9720654,5.089271,3.8103511,2.7313805,2.4861598,1.9881734,1.8334957,1.6335466,1.3128735,1.1280149,0.935611,0.9205205,1.026154,1.0902886,0.87147635,0.79602385,0.935611,0.935611,0.77338815,0.76207024,0.84884065,0.9620194,1.0827434,1.1204696,0.9016574,0.77716076,0.7469798,0.7167987,0.6526641,0.58098423,0.69039035,0.90920264,0.9695646,0.9016574,1.0223814,0.9242931,0.8903395,0.9695646,1.1393328,1.297783,1.2223305,1.2411937,1.3996439,1.6033657,1.6033657,1.8825399,2.4371157,2.7125173,2.5314314,2.1051247,1.4939595,1.3355093,1.327964,1.1883769,0.6413463,0.7130261,0.5319401,0.4074435,0.4376245,0.47157812,0.7432071,1.659955,4.402653,8.345046,11.076427,11.065109,11.208468,10.7218,10.412445,12.694883,12.96274,11.099063,9.035437,7.7414265,7.2170315,7.6697464,7.2962565,7.149124,7.3868,7.2623034,6.7869525,6.858632,6.937857,6.779407,6.439871,6.549277,6.8435416,6.700182,5.8588867,4.395108,3.8103511,3.138824,2.867195,3.048281,3.3425457,2.7426984,2.4823873,2.6672459,3.0445085,3.0218725,2.9615107,3.0369632,2.9615107,2.8256962,3.0822346,3.6330378,4.0517993,3.953711,3.4255435,3.0218725,2.9728284,2.9954643,3.0218725,2.8822856,2.3201644,1.5882751,1.3770081,1.2713746,1.2449663,1.6486372,1.5618668,1.7240896,1.6863633,1.4109617,1.2525115,1.2751472,1.1242423,0.9808825,0.935611,1.0072908,1.5580941,2.2899833,2.546522,2.1315331,1.3128735,1.0072908,0.9016574,0.84129536,0.7696155,0.73188925,0.67152727,0.663982,0.6413463,0.58475685,0.55080324,0.513077,0.66775465,0.80734175,0.7922512,0.5357128,0.5696664,0.5357128,0.4376245,0.33576363,0.33576363,0.3734899,0.482896,0.5357128,0.56589377,0.76207024,1.0186088,1.1921495,1.3656902,1.4600059,1.267602,1.4977322,1.8599042,2.0108092,1.9127209,1.8146327,1.7052265,2.263575,2.9652832,3.3953626,3.2482302,3.5802212,3.7160356,3.9688015,4.357382,4.640329,4.847823,5.2099953,5.247721,4.8440504,4.255521,4.587512,5.0439997,5.534441,6.1342883,7.111398,6.598321,6.2135134,6.115425,6.3116016,6.651138,6.628502,5.8626595,4.7950063,3.731126,2.837014,2.203213,2.1353056,2.0749438,1.8674494,1.7693611,2.123988,2.9992368,3.9461658,4.447925,3.9386206,3.350091,3.2670932,3.0746894,2.6332922,2.305074,2.9766011,3.7650797,4.45547,5.0553174,5.798525,6.458734,6.907676,7.0812173,7.141579,7.4471617,7.8734684,8.458225,9.084481,9.714509,10.359629,11.653639,12.510024,12.928786,12.528888,10.514306,9.25425,9.050528,9.288202,9.906913,11.3820095,13.543724,15.596032,17.37671,18.51227,18.402864,17.7917,17.097536,16.58446,16.505234,17.08999,17.112627,17.716248,18.71222,19.640285,19.7761,1.2261031,1.1129243,1.0110635,1.0035182,1.0374719,0.9016574,1.1016065,1.2826926,1.3807807,1.4600059,1.6939086,1.1959221,0.8601585,0.5772116,0.331991,0.181086,0.4640329,0.38480774,0.1961765,0.060362,0.0452715,0.08299775,0.29803738,0.35839936,0.29426476,0.5017591,1.0336993,1.6750455,2.0749438,2.1541688,2.123988,2.191895,2.1956677,1.9994912,1.6637276,1.4713237,1.50905,1.388326,1.1619685,0.94315624,0.91674787,0.7130261,0.59230214,0.44894236,0.30935526,0.29803738,0.40367088,0.4074435,0.39989826,0.3961256,0.34330887,0.45648763,0.95447415,1.4713237,1.8674494,2.2296214,2.3993895,3.2520027,4.187614,4.6252384,4.002755,6.2097406,9.310839,11.336739,12.064855,13.011784,15.430037,16.21097,14.762281,12.215759,11.461235,15.965749,20.768301,25.227543,27.936289,26.736593,23.363867,15.924251,10.472807,9.608876,12.453435,14.260523,13.890805,11.249968,7.4207535,4.6554193,4.5196047,4.798779,4.979865,4.7421894,3.953711,5.406172,5.5080323,5.3080835,5.541986,6.6360474,7.322665,5.9607477,5.6551647,6.8774953,7.4999785,3.942393,2.8030603,2.4559789,2.5276587,3.8820312,3.6443558,2.9464202,2.7313805,3.1237335,3.4557245,2.0258996,1.1883769,0.7884786,0.7884786,1.2449663,1.9957186,1.6486372,1.0336993,0.5772116,0.3169005,0.23013012,0.17354076,0.19994913,0.271629,0.2678564,0.211267,0.241448,0.31312788,0.34330887,0.2565385,0.29426476,0.6828451,0.86770374,0.73566186,0.633801,0.34330887,0.27540162,0.20749438,0.11317875,0.16976812,0.1056335,0.090543,0.13958712,0.241448,0.3734899,0.3055826,0.26031113,0.32444575,0.43385187,0.392353,0.46026024,0.7130261,0.73566186,0.573439,0.7092535,0.6828451,0.5696664,0.3961256,0.26031113,0.34330887,0.30935526,0.44139713,0.98842776,2.1956677,4.2819295,6.960493,8.646856,9.310839,8.710991,6.3908267,5.6778007,7.115171,9.903141,12.845788,14.358611,15.505488,20.360857,28.207916,34.42143,30.46772,31.531599,31.290152,27.634478,21.583187,17.28994,16.4411,14.750964,15.999702,20.202406,23.635496,25.589716,23.299732,19.83269,18.13878,21.021067,24.63524,26.197107,28.966215,33.644268,38.38646,43.69077,40.502903,37.36785,37.22072,37.382942,33.77631,32.59925,31.433512,30.158363,30.946842,38.12615,43.294643,49.960873,56.7931,57.623074,61.90123,64.345894,67.85443,75.71658,91.60311,121.91992,143.49179,155.70378,152.52345,122.48582,111.205666,101.830696,82.27341,53.62032,30.113092,22.72252,17.410664,10.797253,4.7308717,6.300284,15.064092,19.862871,17.520071,9.88805,3.85185,2.6936543,3.5085413,5.534441,7.326438,6.72659,7.1076255,4.5007415,2.7917426,2.9313297,2.9200118,2.584248,2.4295704,2.493705,2.8256962,3.482133,3.2557755,2.282438,1.4600059,1.1016065,0.935611,0.8526133,1.2261031,2.3918443,3.942393,4.749735,5.342037,6.620957,7.9489207,9.74469,13.475817,16.59955,14.064346,11.717773,11.495189,11.408418,12.479843,12.3289385,12.947649,14.498198,15.30554,15.920478,17.7917,19.11589,19.58747,20.413673,18.700903,16.784409,15.07541,14.460471,16.320375,16.520325,13.615403,11.00852,10.065364,10.121953,10.484125,10.38981,9.861642,9.016574,8.062099,7.164215,8.635539,10.4049,11.736636,13.230596,15.365902,23.126192,26.117884,24.525835,29.139755,29.769783,35.172184,39.20512,38.899536,34.447838,29.72074,24.937052,22.764019,23.94485,27.302486,30.995888,26.24238,18.848034,12.698656,9.774872,12.234623,12.543978,13.124963,14.9358225,17.48989,15.46399,12.559069,12.325166,13.875714,11.917723,13.807808,20.583443,20.938068,13.777626,8.194141,3.4934506,5.292993,8.692128,10.906659,11.306557,15.399856,18.127462,17.071129,13.038192,10.103089,10.921749,14.102073,16.38451,16.0827,13.106099,22.503708,24.789919,22.990377,19.425245,15.716756,11.781908,7.54525,5.0854983,4.817642,5.4703064,2.6936543,2.5427492,3.62172,4.06689,1.5316857,1.3317367,0.8111144,0.7092535,1.0789708,1.2826926,1.146878,0.7997965,0.51684964,0.42630664,0.5017591,0.65643674,1.146878,2.0787163,3.3123648,4.4516973,7.224577,10.106862,12.2119875,12.400619,9.276885,9.295748,9.163706,9.857869,11.050018,11.087745,9.491924,8.511042,7.0774446,5.8890676,7.3905725,11.574413,14.045483,13.8719425,11.332966,7.9225125,7.322665,8.273367,8.98262,8.756263,8.001738,8.858124,11.763044,13.52486,13.155144,11.853588,10.672756,11.52537,12.132762,11.947904,12.136535,11.785681,12.864652,13.283413,13.468271,16.373192,17.206944,17.652113,18.51227,19.938324,21.402102,16.21097,16.131744,16.848543,16.399601,15.147089,13.65313,13.181552,13.226823,13.226823,12.528888,10.782163,8.597813,7.0057645,6.228604,5.666483,5.492942,4.8855495,3.9008942,2.9464202,2.7804246,2.3880715,2.0485353,1.8033148,1.6222287,1.4109617,1.0676528,0.9695646,0.98465514,0.965792,0.7469798,0.7432071,0.9280658,1.0525624,1.0186088,0.8601585,0.8299775,0.9280658,1.0412445,1.116697,1.1808317,0.9016574,0.76584285,0.77716076,0.83752275,0.76207024,0.8224323,0.9280658,0.9016574,0.77338815,0.77716076,0.90543,0.965792,1.0336993,1.1016065,1.0638802,0.9922004,1.1431054,1.4713237,1.8259505,1.931584,2.5729303,2.8898308,2.7653341,2.305074,1.8372684,1.3241913,0.95824677,0.8865669,0.87902164,0.3470815,0.44894236,0.44894236,0.38103512,0.32067314,0.3734899,0.633801,1.6222287,4.485651,8.605357,11.615912,9.982366,9.691874,9.001483,8.058327,8.873214,9.378746,9.563604,8.9788475,7.7829256,6.741681,6.7152724,6.6020937,6.617184,6.911449,7.5792036,6.9982195,6.4436436,6.405917,6.688864,6.428553,6.0286546,6.0776987,6.2097406,5.824933,4.0782075,3.2369123,3.1576872,3.1614597,3.1463692,3.5839937,3.006782,2.6483827,2.6446102,2.8106055,2.6672459,2.625747,2.6332922,2.4672968,2.3088465,2.7389257,3.0746894,3.5085413,3.6707642,3.4632697,3.0709167,3.059599,3.0860074,2.927557,2.5502944,2.1353056,1.5618668,1.2864652,1.1657411,1.1732863,1.3920987,1.4147344,1.5279131,1.5656394,1.4562333,1.237421,1.1355602,0.9922004,0.8941121,0.84129536,0.7394345,1.0940613,1.6222287,1.750498,1.4260522,1.1053791,0.83752275,0.70170826,0.62625575,0.56589377,0.5017591,0.46026024,0.48666862,0.5357128,0.58475685,0.633801,0.62625575,0.6790725,0.94692886,1.2902378,1.267602,0.8337501,0.7469798,0.70170826,0.58098423,0.44516975,0.5394854,0.5696664,0.5998474,0.663982,0.7507524,0.94692886,1.1808317,1.3732355,1.4147344,1.1808317,1.20724,1.8448136,2.3616633,2.5087957,2.546522,2.535204,2.335255,2.625747,3.4142256,4.0178456,3.9688015,3.8178966,4.1574326,4.859141,5.1043615,4.9987283,4.878004,4.5497856,4.13857,4.112161,4.606375,5.4438977,5.915476,6.149379,7.0849895,6.221059,5.413717,5.191132,5.621211,6.2851934,5.726845,4.8742313,3.783943,2.71629,2.1654868,1.9994912,2.0372176,1.9768555,1.81086,1.8184053,2.0070364,2.746471,3.5424948,4.06689,4.168751,3.9914372,3.7877154,3.4896781,3.078462,2.5729303,2.8634224,3.5236318,4.3083377,5.119452,5.9796104,6.2097406,6.6624556,6.94163,6.9869013,7.066127,7.515069,8.386545,9.076936,9.514561,10.18986,11.23865,11.257513,10.555805,9.367428,7.8508325,7.277394,7.3415284,7.877241,8.8618965,10.4049,12.792972,14.592513,15.746937,16.42601,16.999449,17.071129,16.995676,16.848543,16.897587,17.603067,17.772837,18.127462,18.87067,19.711966,19.836462,0.6375736,0.633801,0.62248313,0.6413463,0.6488915,0.5281675,0.76584285,0.8601585,0.91297525,0.98842776,1.1280149,0.8224323,0.543258,0.331991,0.20372175,0.1659955,0.32067314,0.23390275,0.11317875,0.060362,0.090543,0.15467763,0.44516975,0.5017591,0.362172,0.55080324,0.7922512,1.116697,1.4260522,1.6410918,1.7278622,1.5656394,1.5656394,1.5958204,1.6033657,1.6146835,1.5279131,1.5543215,1.4713237,1.2864652,1.2223305,1.1280149,0.875249,0.6111652,0.44139713,0.44894236,0.513077,0.482896,0.42630664,0.38103512,0.31312788,0.23013012,0.46026024,1.1581959,2.0296721,2.3428001,2.6031113,3.6254926,4.7421894,5.553304,5.9494295,11.314102,18.368912,21.75673,21.190834,21.462463,20.772074,18.991394,16.022339,13.234368,13.45318,17.240896,20.179771,22.04722,22.847017,22.820608,19.478064,15.022593,12.400619,13.162688,17.45971,18.591496,16.67123,12.90615,8.586494,5.1043615,5.4665337,5.4212623,4.7874613,4.104616,4.6327834,5.8400235,6.25124,6.126743,5.7796617,5.583485,8.314865,8.3525915,7.24344,6.0550632,5.402399,3.6292653,3.3840446,2.8407867,2.263575,3.9989824,4.7044635,3.6330378,3.0709167,4.991183,11.087745,10.419991,5.5495315,2.0372176,1.8674494,3.4330888,3.7537618,3.470815,2.6597006,1.5015048,0.26408374,0.331991,0.2678564,0.26031113,0.30181,0.19994913,0.17731337,0.24522063,0.30935526,0.331991,0.3470815,0.34330887,0.6790725,0.91674787,1.0412445,1.4864142,1.2034674,0.73566186,0.33576363,0.14335975,0.18863125,0.20749438,0.14713238,0.14713238,0.21503963,0.23767537,0.14713238,0.116951376,0.15467763,0.21503963,0.20749438,0.271629,0.42630664,0.5017591,0.47912338,0.4979865,0.6790725,0.56212115,0.41121614,0.3772625,0.52062225,0.4376245,0.7054809,1.7278622,3.591539,6.039973,8.7751255,7.8734684,6.9265394,6.934085,6.3153744,5.8928404,7.3075747,10.450171,13.845533,14.652876,15.973294,22.303759,30.203636,36.024796,35.90407,33.16892,32.36535,30.05273,25.35204,19.934551,16.071383,13.804035,15.030138,19.478064,24.688059,23.394047,18.666948,14.66042,14.030393,17.912424,20.75321,20.975796,23.031876,27.577888,31.456148,34.926964,34.447838,33.881947,33.953625,32.26349,28.905853,28.094738,27.857063,28.596497,33.06706,39.974735,43.37387,47.387943,52.439487,55.265182,57.362762,60.618538,64.51189,70.22742,80.67759,110.67373,127.36759,135.62587,133.57733,112.61663,103.75096,93.678055,75.9203,51.12284,27.061039,21.31533,19.217752,13.238141,5.3458095,7.0057645,21.779364,22.005722,16.70141,11.529142,8.805306,3.832987,3.440634,4.293247,4.798779,5.1232247,6.8359966,4.8440504,3.127506,3.108643,3.6330378,3.1237335,2.5691576,2.595566,3.199186,3.7462165,3.3651814,2.3578906,1.5769572,1.267602,1.0525624,0.91297525,0.9695646,1.5845025,2.7313805,3.99521,4.61392,5.96452,7.1076255,8.254503,10.785934,12.46098,11.031156,10.144588,10.668983,10.695392,13.396591,12.992921,13.004238,14.407655,15.611122,15.199906,16.82968,18.097282,18.055782,17.210714,16.991903,15.886524,14.222796,13.226823,15.045229,15.524352,12.619431,9.812597,8.771353,9.325929,10.567122,10.012547,9.058073,8.843033,10.242677,8.612903,8.68081,9.522105,10.744436,12.487389,16.109108,21.013521,22.552752,21.477554,23.952396,24.801237,28.483318,31.931498,33.165146,31.248653,30.346996,28.185282,24.925734,21.85859,21.405874,27.913652,27.645796,22.152855,14.905642,11.272603,12.00072,13.81158,15.588487,17.025856,18.614132,16.275105,12.494934,10.310584,10.589758,12.034674,15.98084,19.395065,18.293459,12.449662,5.3948536,4.5497856,8.959985,8.729855,5.1760416,10.808571,17.693611,19.99114,19.61765,18.572634,18.97253,19.161163,20.866388,20.987112,18.61036,14.984866,19.1008,22.590479,23.069601,20.65135,17.935059,15.931795,11.619685,8.2507305,6.881268,6.379509,3.9763467,3.5047686,4.0895257,4.236658,1.8448136,1.4713237,1.0487897,1.2411937,1.8297231,1.7429527,1.177059,0.72811663,0.46026024,0.4074435,0.5394854,0.4979865,0.94692886,1.7580433,2.6785638,3.3161373,6.628502,10.008774,12.521342,12.89106,9.469289,9.310839,8.484633,8.654402,9.623966,9.367428,9.005256,9.344792,8.397863,6.700182,7.3188925,9.937095,11.5857315,12.3289385,11.902632,9.703192,8.620448,10.152134,10.657665,9.352338,8.303548,6.851087,8.001738,9.918231,11.2650585,11.189606,11.050018,10.484125,9.544742,8.82417,9.442881,9.623966,10.148361,10.461489,10.733118,11.846043,13.355092,14.584969,16.309057,17.980331,17.73511,16.592005,16.761772,17.123945,16.663685,14.5132885,14.219024,13.585222,13.592768,13.849306,12.611885,11.2801485,9.495697,7.8508325,6.63982,5.8702044,5.772116,5.1647234,4.1272516,3.1199608,2.9803739,2.9237845,2.6332922,2.2220762,1.8184053,1.5543215,1.2638294,1.0902886,1.1355602,1.2487389,1.0299267,0.9242931,0.87902164,0.9242931,0.95824677,0.7582976,0.80734175,0.95447415,0.9922004,0.935611,1.0299267,0.91297525,0.814887,0.8262049,0.875249,0.7432071,0.77716076,0.90543,0.94692886,0.875249,0.83752275,0.8563859,0.9280658,1.0186088,1.0902886,1.1091517,0.8865669,1.0827434,1.4977322,1.8938577,2.003264,2.4522061,2.6106565,2.3956168,2.0258996,2.0258996,1.6712729,1.2940104,1.0601076,0.8903395,0.4678055,0.47535074,0.482896,0.44139713,0.38858038,0.43385187,0.49044126,1.2411937,3.4670424,6.9755836,10.578441,9.314611,9.06939,8.228095,6.858632,6.7379084,7.7338815,8.028146,7.9451485,7.605612,6.9227667,6.7567716,6.4964604,6.066381,5.9305663,7.073672,6.63982,6.224831,6.4247804,6.960493,6.670001,6.6058664,6.832224,6.9152217,6.356873,4.5837393,3.7235808,3.3236825,3.029418,2.8332415,3.097325,2.8030603,2.4182527,2.3126192,2.4597516,2.4522061,2.493705,2.7917426,2.8785129,2.7389257,2.7841973,2.8822856,3.0558262,3.2029586,3.2331395,3.1010978,3.0633714,3.0105548,2.7879698,2.3503454,1.750498,1.3392819,1.1129243,1.1016065,1.2185578,1.2638294,1.3770081,1.4034165,1.3204187,1.1808317,1.1242423,1.1317875,1.0978339,1.0072908,0.90920264,0.935611,1.116697,1.3015556,1.2826926,1.1053791,1.0638802,0.77716076,0.66020936,0.6073926,0.5470306,0.452715,0.4678055,0.58098423,0.6828451,0.784706,1.0412445,1.3392819,1.2562841,1.2525115,1.3656902,1.2110126,0.83752275,0.62625575,0.52439487,0.4678055,0.39989826,0.47157812,0.5772116,0.6828451,0.79602385,0.965792,1.1204696,1.0374719,0.91297525,0.8337501,0.76584285,1.2110126,1.9429018,2.655928,3.0746894,2.9501927,2.9841464,2.886058,3.0445085,3.6330378,4.5950575,4.2064767,4.146115,4.4403796,4.7836885,4.5309224,5.0439997,5.040227,4.727099,4.398881,4.447925,5.4703064,6.149379,6.326692,6.228604,6.477597,5.5382137,5.0477724,5.1232247,5.564622,5.885295,4.82896,3.7763977,2.8407867,2.161714,1.8787673,1.991946,1.9655377,1.8636768,1.7429527,1.6863633,1.7655885,2.3277097,3.0558262,3.731126,4.236658,4.353609,4.0895257,3.821669,3.5877664,3.0897799,3.0860074,3.399135,3.983892,4.82896,5.96452,5.907931,5.96452,6.066381,6.2625575,6.72659,7.1906233,7.956466,8.812852,9.552286,9.97482,10.38981,9.8239155,8.612903,7.273621,6.519096,6.7831798,7.3151197,8.111144,9.163706,10.465261,11.902632,12.981603,13.841762,14.543469,15.0905,15.731846,16.007248,16.320375,16.840998,17.527617,17.882242,18.02183,18.274595,18.693357,19.063074,0.41876137,0.41876137,0.39989826,0.41121614,0.44516975,0.45648763,0.5357128,0.52439487,0.52062225,0.543258,0.55080324,0.482896,0.31312788,0.21503963,0.22258487,0.2263575,0.26408374,0.27540162,0.22258487,0.14713238,0.16976812,0.23013012,0.513077,0.56212115,0.392353,0.47535074,0.5772116,0.7582976,0.9620194,1.1355602,1.2147852,1.0525624,1.1016065,1.3317367,1.6184561,1.750498,1.81086,1.9127209,2.0070364,1.9806281,1.6825907,1.5807298,1.4071891,1.0676528,0.7130261,0.754525,0.7922512,0.6828451,0.58098423,0.51684964,0.4376245,0.5017591,0.98465514,1.9391292,3.006782,3.3953626,4.183841,5.9305663,7.798016,9.318384,10.416218,15.645076,23.22428,27.211945,27.215717,28.39655,27.845745,25.619896,22.009495,18.666948,18.614132,19.33093,19.519562,20.100546,21.254969,22.443346,18.576405,16.229834,16.286423,18.595268,21.983086,21.4436,19.232841,15.309312,10.170997,4.82896,5.624984,5.715527,4.930821,4.195159,5.50426,5.372218,5.764571,5.96452,5.50426,4.1536603,7.1793056,7.6207023,6.48137,4.8666863,3.9914372,3.399135,3.863168,3.5575855,2.9766011,4.949684,8.75249,11.529142,13.072145,14.551015,18.516043,16.414692,8.167733,2.6672459,2.637065,4.647874,3.7198083,4.8666863,5.251494,3.7613072,0.9808825,0.5319401,0.33953625,0.331991,0.35462674,0.1659955,0.14713238,0.2678564,0.34330887,0.331991,0.33576363,0.5357128,0.9205205,1.20724,1.4449154,2.0183544,1.5845025,0.8526133,0.32821837,0.18485862,0.27917424,0.21881226,0.150905,0.14335975,0.17731337,0.14713238,0.09808825,0.12826926,0.116951376,0.060362,0.09808825,0.14335975,0.21503963,0.30181,0.35839936,0.32067314,0.4979865,0.482896,0.45648763,0.52062225,0.694163,0.845068,1.2034674,2.7011995,5.032682,6.6322746,9.035437,7.6886096,6.307829,6.228604,6.398372,6.2361493,7.7716074,10.567122,13.290957,13.70972,15.875206,21.967995,29.13221,35.42495,39.80874,36.51901,34.40634,31.286379,26.883726,22.847017,17.006994,14.920732,16.463736,20.36463,24.193844,19.859098,14.569878,11.148107,11.00852,14.181297,15.535669,15.743164,18.485863,23.692085,27.525072,28.547453,28.475773,28.532362,28.58518,27.136492,24.940825,24.812555,25.887753,28.536135,34.379932,39.672924,42.898518,47.750114,54.3258,59.128353,58.728455,59.086853,60.44877,63.63664,70.031235,97.47708,111.831924,120.0487,121.19935,106.501205,96.066124,84.18236,68.2317,47.565254,23.503454,17.516298,16.848543,12.668475,5.8513412,6.9567204,23.854307,21.707684,15.23386,11.729091,11.072655,4.5988297,4.9232755,4.919503,3.029418,3.2520027,5.138315,4.168751,3.0445085,2.9086938,3.3350005,3.0897799,2.5201135,2.4597516,2.9803739,3.3727267,3.048281,2.3314822,1.8749946,1.7089992,1.267602,1.3845534,1.3732355,1.6939086,2.6634734,4.447925,4.6742826,5.798525,6.700182,7.405663,9.046755,9.046755,8.209232,8.246958,9.175024,9.329701,12.585477,12.464753,12.287439,13.143826,13.86817,13.328684,14.1926155,14.86037,14.720782,14.154889,14.916959,14.943368,14.124708,13.287186,14.177525,14.84528,12.823153,10.284176,8.6581745,8.631766,9.978593,9.4127,8.971302,9.910686,12.73261,10.63503,9.303293,8.7600355,9.042982,10.223814,15.656394,18.893307,19.523335,18.632996,18.840488,19.87796,21.790682,23.348776,24.065575,24.20139,25.110592,25.800982,23.990122,20.123182,17.357847,23.465727,26.34424,24.933279,19.859098,13.404137,13.106099,17.04472,19.278114,18.900852,20.059048,16.859861,12.347801,9.125979,8.431817,10.159679,13.830443,13.996439,11.898859,10.31813,13.585222,22.582933,16.569368,7.9828744,5.1269975,12.151625,17.829426,19.56106,21.058792,24.593742,31.007204,26.295197,24.58997,24.046711,22.665932,18.304777,16.233604,17.765291,19.25925,19.346022,18.919714,17.50498,14.1058445,10.710483,8.224322,6.4738245,5.0062733,4.3347464,4.6856003,4.8666863,2.2447119,1.4562333,1.1242423,1.5015048,2.1881225,2.1202152,1.3920987,0.8526133,0.5470306,0.4640329,0.5394854,0.5017591,0.965792,1.6863633,2.3993895,2.8256962,5.9720654,9.0957985,11.604594,12.408164,9.944639,9.937095,8.6732645,8.307321,8.695901,7.405663,7.4396167,8.280911,8.367682,7.7678347,8.167733,9.148616,9.688101,10.144588,10.378491,9.733373,10.529396,12.3289385,12.068627,9.6201935,7.798016,5.73439,4.9119577,5.5004873,7.0170827,8.314865,9.827688,9.314611,8.122461,7.2396674,7.3000293,8.612903,9.405154,9.397609,8.8769865,8.722309,9.967276,11.080199,13.20796,15.158407,13.381501,15.520579,16.897587,17.723793,17.429527,14.667966,14.094527,13.739901,13.928532,14.166207,13.13628,11.419736,10.265312,8.710991,6.832224,5.7419353,5.798525,5.20245,4.183841,3.2331395,3.1048703,3.2142766,3.127506,2.7200627,2.123988,1.7542707,1.4260522,1.2223305,1.2298758,1.3392819,1.237421,1.0035182,0.845068,0.8224323,0.84129536,0.66020936,0.7167987,0.87902164,0.90920264,0.814887,0.84884065,0.8978847,0.87147635,0.8865669,0.9016574,0.72811663,0.7167987,0.80356914,0.8563859,0.8337501,0.7809334,0.7507524,0.7809334,0.8601585,0.95824677,1.0223814,0.935611,1.146878,1.4524606,1.720317,1.8938577,2.2258487,2.2673476,2.1164427,1.991946,2.2447119,1.9127209,1.8334957,1.7919968,1.599593,1.0714256,0.60362,0.63002837,0.68661773,0.77338815,1.3430545,0.97710985,1.0601076,2.305074,5.2137675,10.057818,9.186342,8.801534,8.096053,6.85486,5.451443,6.5568223,6.760544,6.8661776,7.032173,6.7643166,6.5040054,6.3153744,5.9117036,5.666483,6.620957,6.462507,6.3153744,6.6058664,7.092535,6.8737226,7.281166,7.6282477,7.4282985,6.462507,4.7836885,3.8820312,3.451952,3.0331905,2.595566,2.5427492,2.4899325,2.1390784,1.961765,2.0560806,2.1315331,2.191895,2.704972,2.9803739,2.848332,2.6446102,2.7200627,2.7200627,2.7917426,2.938875,3.0407357,2.9916916,2.757789,2.4069347,1.961765,1.3958713,1.1431054,1.0374719,1.146878,1.327964,1.2562841,1.2940104,1.3091009,1.1619685,0.935611,0.91674787,1.0412445,1.0827434,1.0601076,1.056335,1.2185578,1.4675511,1.3996439,1.146878,0.9016574,0.9280658,0.66020936,0.56589377,0.5319401,0.4979865,0.45648763,0.4979865,0.6375736,0.7997965,0.95824677,1.1242423,1.4109617,1.4222796,1.3505998,1.2147852,0.88279426,0.69793564,0.52062225,0.4376245,0.44516975,0.43007925,0.42630664,0.5470306,0.6828451,0.7922512,0.91674787,0.98842776,0.79602385,0.6073926,0.55080324,0.62625575,1.1393328,1.6184561,2.2183034,2.7917426,2.9086938,2.7992878,2.9464202,3.127506,3.451952,4.3649273,4.006528,4.255521,4.666737,4.889322,4.696918,5.2250857,5.172269,4.776143,4.402653,4.564876,5.794752,6.1531515,6.2135134,6.168242,5.836251,4.8553686,4.8402777,5.1534057,5.3269467,5.070408,3.7914882,2.8407867,2.2560298,1.991946,1.9240388,1.991946,1.8938577,1.8070874,1.7693611,1.6712729,1.6863633,2.1541688,2.8445592,3.5500402,4.08198,4.221567,4.025391,3.8820312,3.8443048,3.6481283,3.663219,3.9310753,4.357382,4.9534564,5.8400235,5.6400743,5.462761,5.515578,5.824933,6.2436943,6.7454534,7.5226145,8.431817,9.186342,9.35611,9.424017,8.726082,7.594294,6.5040054,6.0626082,6.7114997,7.533932,8.492179,9.537196,10.627484,11.408418,12.030901,12.683565,13.355092,13.807808,14.230342,14.5132885,15.23386,16.395828,17.463482,17.942604,18.006739,17.938831,17.976559,18.312323,0.47912338,0.35839936,0.26408374,0.2678564,0.3734899,0.51684964,0.40367088,0.36971724,0.36594462,0.35085413,0.29426476,0.33953625,0.24899325,0.23013012,0.30181,0.29049212,0.38858038,0.5017591,0.44894236,0.27540162,0.2678564,0.30181,0.482896,0.49421388,0.32444575,0.27540162,0.43007925,0.6187105,0.73188925,0.7394345,0.70170826,0.80734175,1.0299267,1.3392819,1.6373192,1.7580433,2.161714,2.2598023,2.4710693,2.6823363,2.2673476,2.214531,2.1541688,1.6561824,0.965792,0.98842776,1.1317875,1.026154,0.875249,0.754525,0.6187105,0.94315624,1.7014539,2.546522,3.259548,3.7537618,5.560849,8.567632,11.6875925,14.064346,15.060319,17.301258,21.217243,24.152346,25.729303,27.819336,29.803738,29.532108,26.849771,23.246916,21.85859,19.338476,17.765291,19.002712,22.235851,23.959942,20.089228,18.923487,20.375948,23.107328,24.51829,23.446865,21.941587,17.904879,11.385782,4.5912848,5.2137675,5.8400235,5.59103,4.930821,5.6778007,4.447925,4.6252384,5.05909,4.8100967,3.169005,5.010046,4.6629643,4.164978,4.2630663,4.4177437,3.651901,4.2328854,4.244203,4.1197066,6.617184,14.381247,22.967741,26.879953,24.680513,19.002712,14.996184,8.024373,4.991183,6.9227667,8.975075,4.4177437,6.3908267,8.160188,6.63982,2.372981,0.80356914,0.3734899,0.36594462,0.35839936,0.211267,0.20749438,0.362172,0.482896,0.4979865,0.45648763,0.8526133,1.388326,1.6750455,1.7127718,1.8787673,1.2336484,0.6149379,0.2867195,0.27917424,0.36971724,0.23390275,0.211267,0.21503963,0.241448,0.3734899,0.41121614,0.52062225,0.43385187,0.19240387,0.150905,0.150905,0.19240387,0.16976812,0.10940613,0.17731337,0.2678564,0.41498876,0.59607476,0.79602385,1.0299267,1.5430037,1.9051756,3.4066803,5.349582,5.040227,7.0887623,8.126234,8.235641,7.7716074,7.356619,7.424526,9.665465,12.049765,13.562587,14.1926155,16.784409,20.492899,26.68755,34.496883,40.84621,39.88419,36.983044,31.776821,26.1707,24.310795,19.647831,17.184307,17.953922,20.394812,20.33822,14.679284,10.378491,8.718536,9.450426,10.79348,10.831206,12.166716,15.603577,20.685303,25.706667,26.087702,24.35984,22.616886,22.043447,22.948877,22.013268,22.945105,25.431265,28.996395,33.01424,36.79441,41.20838,50.390953,62.57653,70.099144,67.97138,61.85219,57.355217,57.55894,63.029247,86.370476,97.605354,106.20316,111.69988,103.694374,89.54703,74.509346,58.95104,41.615826,19.625195,11.717773,10.231359,8.469543,5.511805,6.221059,20.160908,19.508244,14.6151495,10.770844,8.194141,4.315883,7.696155,7.8923316,3.4972234,2.1315331,3.3651814,2.897376,2.5427492,2.7540162,2.637065,2.6408374,2.354118,2.1579416,2.2560298,2.6521554,2.4899325,2.2107582,2.11267,2.052308,1.4373702,1.9164935,2.0673985,2.41448,3.3878171,5.2967653,5.587258,6.6813188,7.3490734,7.726336,9.318384,8.8618965,8.054554,7.413208,7.254758,7.699928,10.453944,10.827434,11.000975,11.574413,11.563096,11.932813,11.400873,10.86516,11.027383,12.377983,13.558814,13.947394,13.864397,13.63804,13.607859,15.056546,14.683057,12.909923,10.555805,8.843033,9.408927,9.314611,9.405154,10.344538,12.604341,10.650121,8.797762,7.8244243,7.8319697,8.262049,13.619176,16.414692,17.384256,17.150352,16.222288,17.37671,18.270823,18.153872,17.448391,17.742655,17.637022,19.76101,21.051247,20.421219,18.738628,22.03213,25.793438,28.573862,27.615616,18.848034,17.410664,21.651094,23.428001,21.579414,21.90386,17.569115,13.185325,10.495442,9.522105,8.567632,9.771099,8.805306,6.9189944,9.835234,27.755201,41.64978,23.420456,8.43559,8.59404,12.347801,16.82968,19.851553,22.805517,27.374166,35.579628,27.174217,24.012758,24.367384,24.989868,21.088974,15.833707,14.151116,14.694374,16.335466,18.135008,16.309057,13.577678,10.982111,8.763808,6.3644185,5.2552667,4.689373,5.3759904,6.0362,3.4066803,2.0787163,1.4713237,1.5543215,2.0673985,2.516341,2.1013522,1.5165952,1.0412445,0.8299775,0.90543,0.7507524,1.0336993,1.5618668,2.214531,2.9237845,5.330719,7.835742,9.993684,11.197151,10.668983,10.544487,8.933576,8.360137,8.567632,6.5530496,5.987156,6.1644692,7.201941,8.484633,8.66572,9.21275,9.680555,9.431562,8.646856,8.345046,11.423509,12.955194,12.098808,9.337247,6.4926877,5.926794,4.4403796,3.4972234,3.7763977,5.194905,6.983129,7.9715567,7.91874,7.1604424,6.63982,9.088254,10.121953,9.80128,8.797762,8.401636,8.371455,8.541223,10.103089,12.306303,12.453435,14.324657,16.81459,18.448135,18.285913,15.916705,13.411682,13.536179,14.034165,14.117163,14.460471,11.480098,10.453944,8.990166,6.722818,5.300538,5.2364035,4.7950063,4.063117,3.3576362,3.1954134,3.2331395,3.2972744,3.0181,2.444661,2.0749438,1.6033657,1.3845534,1.2713746,1.2034674,1.2298758,0.97710985,0.87147635,0.83752275,0.7997965,0.6828451,0.6187105,0.7469798,0.83752275,0.8224323,0.77338815,0.8601585,0.875249,0.91297525,0.9393836,0.7884786,0.7092535,0.69039035,0.6828451,0.6451189,0.5583485,0.5885295,0.58098423,0.63002837,0.73566186,0.77716076,0.9997456,1.1996948,1.3091009,1.3845534,1.6184561,2.0258996,2.0296721,2.003264,2.1013522,2.2711203,2.0447628,2.354118,2.5578396,2.335255,1.7014539,0.7130261,0.86770374,1.1091517,1.4222796,2.8106055,2.5427492,1.4373702,1.4109617,3.8178966,9.465516,8.729855,8.009283,7.6697464,7.0849895,4.6290107,5.251494,5.6589375,5.934339,6.1116524,6.1908774,5.8136153,5.9682927,6.1229706,6.156924,6.3531003,6.428553,6.319147,6.488915,6.8397694,6.741681,7.303802,7.6395655,7.2698483,6.1229706,4.5761943,3.5462675,3.4368613,3.1954134,2.6144292,2.323937,2.2786655,1.9579924,1.7014539,1.6335466,1.6712729,1.7089992,2.2069857,2.493705,2.41448,2.3013012,2.4597516,2.444661,2.4899325,2.6446102,2.7804246,2.7238352,2.3163917,1.8259505,1.4222796,1.1732863,1.0223814,1.0601076,1.2336484,1.3920987,1.2864652,1.1808317,1.1959221,1.0940613,0.8639311,0.73566186,0.8903395,0.965792,1.1016065,1.2940104,1.3958713,1.7316349,1.5958204,1.146878,0.68661773,0.6526641,0.4640329,0.38858038,0.3772625,0.41121614,0.47535074,0.56212115,0.68661773,0.8941121,1.0902886,1.026154,0.90920264,1.086516,1.177059,1.0186088,0.66775465,0.62625575,0.5470306,0.52062225,0.5394854,0.52062225,0.49044126,0.56589377,0.65643674,0.69039035,0.62248313,0.5696664,0.5319401,0.5470306,0.63002837,0.754525,0.91674787,0.995973,1.3204187,1.9391292,2.6483827,2.3163917,2.5540671,2.7728794,2.9049213,3.3953626,3.338773,3.9197574,4.6214657,5.1835866,5.572167,5.409944,4.9534564,4.349837,3.9499383,4.315883,5.1647234,5.292993,5.4891696,5.753253,5.27413,4.376245,4.610148,4.82896,4.5535583,3.9688015,2.897376,2.2786655,2.022127,1.9994912,2.0372176,1.9466745,1.8334957,1.7731338,1.7693611,1.7165444,1.7240896,2.2296214,2.9086938,3.500996,3.7914882,3.772625,3.712263,3.7273536,3.863168,4.1008434,4.357382,4.7912335,5.142088,5.3458095,5.5495315,5.3194013,5.240176,5.458988,5.8136153,5.836251,6.3832817,7.284939,8.043237,8.431817,8.465771,8.537451,8.065872,7.394345,6.749226,6.2135134,6.752999,7.4999785,8.405409,9.4013815,10.408672,11.129244,11.706455,12.181807,12.593022,12.992921,12.81938,12.902377,13.747445,15.297995,16.965494,17.652113,17.976559,17.991648,17.859608,17.825653,0.5017591,0.34330887,0.27917424,0.271629,0.26031113,0.1358145,0.16222288,0.32444575,0.3961256,0.32067314,0.19994913,0.124496624,0.071679875,0.05281675,0.1056335,0.29049212,0.39989826,0.3169005,0.23767537,0.2565385,0.36594462,0.3772625,0.33576363,0.21881226,0.090543,0.090543,0.12826926,0.12826926,0.150905,0.2263575,0.33576363,0.56589377,0.72811663,0.8563859,1.0148361,1.2826926,1.780679,2.1994405,2.516341,2.7313805,2.8521044,3.5123138,2.9992368,1.961765,1.0638802,0.97710985,1.3920987,1.569412,1.3505998,0.9016574,0.7167987,0.8262049,1.1280149,1.569412,2.1541688,2.9615107,5.2062225,8.726082,12.879742,16.403374,17.380484,17.452164,17.399347,18.312323,19.7761,19.836462,21.986858,22.386757,20.474035,17.380484,15.916705,13.607859,13.626721,14.913187,16.610868,18.052011,15.890297,19.047983,21.918951,22.831926,24.076893,26.434784,24.53338,18.214233,10.220041,6.1795597,5.6287565,6.930312,6.9491754,5.3609,4.6554193,4.349837,4.557331,4.4215164,3.8556228,3.5236318,5.832478,6.224831,5.9796104,5.907931,6.349328,4.61392,5.4363527,5.406172,5.0175915,8.66572,17.029629,24.291933,24.114618,16.229834,6.439871,6.3417826,8.616675,15.052773,23.303505,26.868635,13.075918,10.416218,10.26154,8.084735,3.4330888,1.0148361,0.43007925,0.32821837,0.16222288,0.19994913,0.47912338,0.5583485,0.69793564,0.9808825,1.297783,1.2864652,1.9240388,2.282438,2.1013522,1.7693611,0.98842776,0.65643674,0.5357128,0.49044126,0.5017591,0.7582976,0.84129536,0.633801,0.47157812,1.1431054,1.3656902,1.6033657,1.3468271,0.68661773,0.32067314,0.32067314,0.35839936,0.29426476,0.19994913,0.33576363,0.6413463,0.76207024,1.0676528,1.5807298,1.9844007,2.4484336,2.8936033,3.6368105,4.636556,5.4778514,6.405917,6.9491754,7.786698,8.627994,8.224322,9.397609,12.344029,15.011275,16.561823,17.380484,19.783646,22.775337,27.094994,33.255688,41.51774,39.00517,35.749393,31.531599,27.325123,25.299223,23.918442,20.50799,18.327412,17.689838,15.931795,10.631257,8.145098,8.631766,10.79348,11.857361,12.147853,12.506252,14.177525,17.493662,21.851044,24.182526,25.07664,24.8201,24.269297,24.842735,22.839472,24.299479,26.32915,27.570343,28.166418,31.441057,37.888474,50.771988,68.80514,86.151665,87.04201,71.30639,56.721416,52.190495,57.755116,79.39867,88.25301,94.93433,101.10635,99.45771,84.1484,64.70429,47.308716,32.32008,14.268067,7.835742,6.7379084,5.956975,4.4743333,5.2779026,12.577931,14.158662,13.792717,12.223305,7.1566696,4.666737,9.673011,10.650121,5.5268955,1.6939086,2.8785129,2.1503963,2.052308,3.0897799,3.7235808,3.3576362,2.7691069,2.6068838,2.9313297,3.2482302,2.003264,1.9240388,1.9957186,1.8523588,1.7542707,1.961765,2.5540671,2.9803739,3.3953626,4.640329,6.858632,9.522105,10.148361,9.148616,9.797507,9.989911,11.057564,10.269085,7.9300575,7.3717093,9.812597,9.544742,9.635284,10.804798,11.427281,12.894833,11.446144,9.8239155,9.740918,11.902632,14.720782,13.630494,12.777881,13.204187,12.864652,15.562078,18.101055,17.999193,14.984866,11.016065,9.454198,8.971302,8.695901,8.345046,8.209232,7.0359454,5.455216,6.1418333,8.541223,8.835487,9.507015,11.827179,14.200161,15.70921,16.11288,16.697638,16.810818,17.180534,17.987877,18.829172,17.278622,17.889788,20.051502,22.511253,23.375185,22.560297,29.000168,34.36107,35.217453,33.078377,24.631468,23.209188,24.899324,25.544443,20.723028,16.475054,14.698147,11.766817,8.873214,12.0082655,7.6395655,5.292993,8.477088,16.25624,23.23937,14.966003,19.934551,21.813318,15.558306,7.4169807,13.849306,21.251196,23.601542,21.4436,21.896315,22.299986,25.329405,24.842735,21.492645,22.733839,20.402355,18.685812,16.720274,15.241405,16.569368,15.411173,10.472807,8.137552,8.888305,7.277394,4.323428,4.044254,4.817642,5.7117543,6.470052,4.5761943,3.187868,2.3088465,2.1277604,3.006782,3.029418,2.6332922,2.1390784,1.9806281,2.7011995,1.6373192,1.20724,1.6071383,2.3880715,2.4710693,4.1574326,6.9491754,8.567632,9.0807085,10.925522,8.103599,6.466279,6.126743,6.515323,6.3945994,4.5497856,4.0706625,5.8098426,8.239413,7.4471617,9.631512,11.000975,11.563096,11.053791,8.941121,9.246704,10.103089,10.33322,8.98262,5.311856,3.832987,3.783943,4.2592936,4.1310244,2.0447628,4.0103,5.1232247,6.405917,7.6886096,7.6282477,11.121698,10.125726,8.473316,8.122461,9.171251,8.424272,8.14887,9.540969,12.257258,14.418973,16.007248,16.667458,16.516552,16.173243,16.784409,13.13628,13.091009,13.392818,13.340002,14.815099,11.959221,9.846551,8.14887,6.6662283,5.3269467,4.459243,4.2404304,4.0404816,3.6594462,3.3425457,3.2821836,3.108643,2.7313805,2.3428001,2.4408884,1.9881734,1.7014539,1.5128226,1.3656902,1.20724,1.1581959,1.0148361,0.8941121,0.84129536,0.8526133,0.6828451,0.80734175,0.8978847,0.83752275,0.70170826,0.69039035,0.724344,0.8224323,0.9205205,0.8865669,0.7394345,0.7469798,0.7469798,0.65643674,0.47157812,0.4376245,0.45648763,0.5357128,0.6451189,0.7167987,0.7922512,0.88279426,1.0110635,1.1280149,1.1280149,1.4109617,1.5430037,1.6788181,1.8674494,2.0749438,2.6597006,2.916239,2.3390274,1.3619176,1.3732355,0.72811663,1.1317875,1.5958204,2.0900342,3.5538127,5.4363527,2.5540671,0.63002837,1.9844007,5.523123,6.085244,5.485397,5.349582,5.583485,4.349837,4.093298,4.266839,4.610148,5.119452,6.058836,5.6778007,5.915476,6.2323766,6.2323766,5.6476197,5.7192993,5.3269467,5.534441,6.205968,5.9984736,6.168242,6.6850915,6.8774953,6.319147,4.8666863,3.7801702,3.2520027,2.9803739,2.776652,2.595566,2.214531,1.8184053,1.4600059,1.2223305,1.2223305,1.4034165,1.7618159,2.0862615,2.263575,2.2899833,2.1541688,2.11267,2.191895,2.293756,2.1805773,1.9994912,1.6675003,1.3392819,1.1091517,1.0374719,0.86770374,0.98842776,1.146878,1.2147852,1.1883769,1.237421,1.0223814,0.9016574,0.91674787,0.80734175,0.95447415,1.1657411,1.4713237,1.7014539,1.4939595,1.2525115,1.1732863,0.8865669,0.45648763,0.3961256,0.2867195,0.2867195,0.35839936,0.4640329,0.55080324,0.8903395,1.1129243,1.2525115,1.3920987,1.6486372,1.2223305,1.0412445,0.97333723,0.9242931,0.83752275,0.9242931,0.6073926,0.36971724,0.35839936,0.3961256,0.59230214,0.7582976,0.8224323,0.7582976,0.6111652,0.4376245,0.35085413,0.31312788,0.35085413,0.5357128,0.754525,0.83752275,1.177059,1.8787673,2.746471,2.4522061,2.727608,2.8747404,2.6898816,2.4559789,2.4672968,3.1312788,4.0593443,4.90064,5.342037,5.1081343,4.255521,3.7462165,3.85185,4.1197066,4.1197066,4.2404304,4.5196047,4.749735,4.45547,4.2102494,4.2894745,3.9688015,3.3236825,3.187868,2.8596497,2.2183034,1.841041,1.8146327,1.7542707,1.9504471,1.8599042,1.6222287,1.3958713,1.3732355,1.5203679,2.161714,2.897376,3.440634,3.5839937,3.5839937,3.5689032,3.682082,3.9688015,4.3347464,4.689373,4.7950063,4.878004,4.961002,4.851596,4.6818275,4.8327327,5.198677,5.66271,6.1041074,6.700182,7.254758,7.7112455,7.9791017,7.9036493,7.816879,7.5490227,7.3075747,7.1302614,6.8963585,7.3490734,7.635793,8.130007,8.907167,9.752235,10.167224,10.699164,11.091517,11.234878,11.200924,11.54046,11.570641,11.932813,12.936331,14.57365,15.916705,17.112627,17.659658,17.546478,17.225805,0.8941121,0.52062225,0.32067314,0.21881226,0.16976812,0.1358145,0.150905,0.21503963,0.211267,0.1358145,0.11317875,0.116951376,0.09808825,0.08299775,0.08677038,0.094315626,0.15467763,0.35462674,0.47535074,0.47157812,0.4640329,0.30181,0.24899325,0.2263575,0.19240387,0.150905,0.120724,0.1056335,0.10940613,0.150905,0.26408374,0.5055317,0.58475685,0.59607476,0.6488915,0.86770374,1.0751982,1.3317367,1.9164935,2.7351532,3.3048196,3.240685,2.4295704,1.5845025,1.1242423,1.1959221,1.6033657,1.7769064,1.5580941,1.1016065,0.8865669,1.3996439,2.033445,2.8407867,3.4670424,3.169005,4.9949555,8.348819,12.774108,16.946632,18.674494,16.607096,15.724301,16.252468,17.803017,19.398838,19.621422,18.251959,17.112627,16.991903,17.637022,16.0412,16.222288,17.222033,17.554024,15.196134,14.4114275,15.23386,16.233604,16.98813,18.085964,15.792209,12.875969,9.714509,7.0963078,6.228604,6.0324273,6.304056,5.726845,4.3649273,3.6783094,3.380272,3.2633207,3.0407357,3.059599,4.2819295,4.889322,4.3611546,3.5387223,3.2520027,4.29702,4.6516466,4.870459,5.349582,6.330465,7.8621507,10.657665,13.36641,12.525115,9.159933,8.782671,11.710228,15.69412,23.179008,30.169682,26.234835,12.608112,7.4169807,5.7419353,4.406426,1.9806281,1.1544232,1.0110635,1.0299267,0.8526133,0.28294688,0.35839936,0.5772116,0.9393836,1.3204187,1.4939595,1.569412,2.2560298,2.5880208,2.1994405,1.3430545,0.8941121,0.59230214,0.5394854,0.66775465,0.7582976,1.1544232,1.5052774,1.5015048,1.2449663,1.2411937,1.5807298,1.9051756,1.9429018,1.6637276,1.297783,0.7997965,0.482896,0.422534,0.62248313,1.0299267,1.2185578,1.4071891,1.6675003,2.0145817,2.3880715,1.931584,2.3088465,3.1048703,4.0216184,4.9044123,6.1531515,7.9489207,10.370946,12.909923,14.449154,13.815352,13.947394,14.758509,15.916705,16.82968,17.301258,19.032892,22.718748,27.49489,30.935526,31.984314,31.143019,27.683523,23.443092,22.831926,23.035648,20.032639,18.516043,18.531134,15.516807,10.608622,7.647111,6.7944975,8.035691,11.197151,13.50977,16.403374,18.836716,20.357084,21.092747,24.439064,26.834682,27.540163,26.480055,24.231571,22.424482,23.578907,23.805264,23.292187,26.31406,29.59247,33.780083,43.25692,58.33233,75.23746,92.78017,79.41376,59.079308,47.157814,50.481495,70.00483,74.9432,81.281204,92.169,97.94489,79.07045,56.71387,38.107285,24.925734,13.264549,7.254758,5.6098933,4.961002,4.564876,6.3153744,10.393582,10.457717,11.189606,12.245941,8.243186,4.9723196,10.099318,11.261286,5.938112,1.4600059,2.4031622,2.1013522,2.0372176,2.6106565,3.138824,3.0143273,3.6330378,4.0593443,3.9348478,3.482133,2.8822856,2.3013012,2.0636258,2.1202152,2.0598533,2.2069857,3.3274553,3.731126,3.470815,4.346064,6.156924,7.91874,8.6581745,8.405409,8.186596,10.020092,9.839006,9.891823,10.321902,9.163706,10.178542,8.582722,7.6923823,8.605357,10.182315,10.702937,12.1101265,12.272349,11.370691,11.891314,14.475562,12.740154,12.091263,13.332457,12.679792,14.34352,16.912678,18.293459,17.23335,13.324911,10.570895,9.673011,9.027891,8.035691,7.111398,5.3156285,3.500996,4.06689,6.228604,6.0022464,7.484888,9.371201,11.197151,13.124963,15.931795,16.750456,16.837225,16.991903,17.844517,19.866644,17.897333,17.112627,18.168962,20.406128,21.839725,30.003687,29.550972,31.437284,38.21669,44.06803,35.364586,28.611588,23.431774,20.360857,20.832436,22.258488,17.071129,11.6008215,9.295748,10.763299,5.4250345,12.491161,17.67852,15.256495,8.043237,15.75071,16.67123,14.4152,11.370691,8.695901,13.656902,18.055782,18.991394,18.082191,21.4436,24.963459,23.58645,20.643805,18.791445,20.025093,17.908651,15.878979,15.535669,15.712983,12.483616,15.599804,14.9358225,14.030393,13.849306,12.781653,10.804798,9.295748,7.2698483,5.3156285,5.613666,4.9647746,4.508287,4.346064,4.4403796,4.606375,4.4818783,4.0404816,3.0746894,2.1277604,2.505023,1.4222796,1.1996948,1.6222287,2.282438,2.5804756,5.5080323,8.073418,8.397863,7.575431,9.691874,8.4544525,7.33021,6.628502,6.304056,5.9192486,5.0515447,4.821415,5.413717,6.428553,6.8850408,8.073418,11.947904,14.637785,13.475817,6.9869013,6.326692,7.77538,9.092027,8.7751255,6.0776987,5.5570765,6.115425,6.7077274,5.847569,1.5807298,2.2560298,2.8445592,4.346064,6.7567716,9.058073,9.220296,7.6848373,7.884786,9.7069645,9.488152,8.469543,8.477088,9.450426,10.861387,11.672502,14.335975,14.743419,14.25675,13.962485,14.709465,13.102326,13.238141,13.332457,12.626976,11.3971,9.118435,9.2844305,8.511042,6.375736,5.4363527,4.247976,3.8971217,3.9197574,3.863168,3.2821836,3.3576362,3.270866,3.1350515,3.0331905,3.0030096,2.5993385,2.214531,1.8448136,1.50905,1.2525115,1.177059,1.116697,1.0374719,0.94315624,0.87902164,0.80734175,0.8865669,0.9242931,0.88279426,0.8865669,0.77338815,0.77716076,0.8601585,0.95447415,0.94692886,0.8299775,0.7922512,0.76584285,0.6752999,0.47157812,0.38858038,0.34330887,0.38103512,0.513077,0.7054809,0.66020936,0.7167987,0.9016574,1.1846043,1.4600059,1.4675511,1.3619176,1.5203679,1.8523588,1.8070874,2.2069857,2.372981,1.9504471,1.3845534,1.9353566,1.4335974,1.5241405,2.5691576,4.187614,5.251494,6.9944468,3.3350005,0.8299775,1.4524606,2.5691576,3.9725742,3.2784111,3.410453,4.432834,3.5802212,3.6179473,3.3010468,3.240685,3.7198083,4.678055,4.9459114,5.2250857,5.8173876,6.304056,5.523123,5.353355,4.8629136,4.9760923,5.541986,5.3269467,5.583485,6.126743,6.017337,5.2552667,4.768598,4.376245,3.7575345,3.1237335,2.6332922,2.4107075,2.003264,1.5769572,1.2223305,0.9997456,0.9393836,1.1242423,1.3468271,1.5015048,1.5656394,1.6184561,1.7467253,1.8372684,1.8674494,1.7995421,1.5731846,1.3392819,1.3053282,1.2261031,1.056335,0.9507015,0.87902164,0.9808825,1.086516,1.1393328,1.2034674,1.2110126,1.0751982,1.0450171,1.1317875,1.1016065,1.5015048,1.3656902,1.1544232,1.0186088,0.8111144,0.76207024,0.724344,0.60362,0.39989826,0.21503963,0.211267,0.24522063,0.331991,0.46026024,0.58475685,0.8111144,1.026154,1.0751982,0.965792,0.8903395,0.80734175,0.8337501,0.98465514,1.116697,0.97333723,0.784706,0.5470306,0.41498876,0.422534,0.47157812,0.52062225,0.5998474,0.66775465,0.68661773,0.6111652,0.43007925,0.3470815,0.32821837,0.35462674,0.41121614,0.58475685,0.66775465,0.91297525,1.3996439,2.052308,1.7882242,1.9655377,2.093807,2.003264,1.871222,1.9994912,2.8294687,3.7047176,4.346064,4.8629136,4.2517486,3.5349495,3.180323,3.180323,3.059599,3.6141748,4.1800685,4.466788,4.398881,4.112161,3.7801702,3.651901,3.4632697,3.1463692,2.8332415,2.3767538,2.1088974,1.9466745,1.8070874,1.6222287,1.5618668,1.629774,1.5203679,1.2525115,1.1883769,1.3543724,1.7089992,2.2069857,2.6785638,2.8030603,3.078462,3.6028569,4.112161,4.4931965,4.8100967,4.98741,5.0213637,4.9459114,4.870459,4.9760923,5.292993,5.270357,5.2552667,5.5570765,6.4436436,6.858632,7.3717093,7.673519,7.707473,7.673519,7.4584794,7.062354,6.730363,6.5530496,6.458734,6.4021444,6.620957,7.3188925,8.409182,9.495697,10.544487,10.751981,10.744436,10.7557535,10.650121,10.525623,10.657665,11.080199,11.781908,12.706201,14.049255,14.973549,15.380992,15.441354,15.592259,0.8639311,0.633801,0.5696664,0.4074435,0.1659955,0.1358145,0.1659955,0.150905,0.13204187,0.116951376,0.10940613,0.11317875,0.094315626,0.09808825,0.10940613,0.06413463,0.1056335,0.20749438,0.27917424,0.29049212,0.2678564,0.23767537,0.3055826,0.3470815,0.29803738,0.17731337,0.14335975,0.08677038,0.06413463,0.09808825,0.181086,0.41121614,0.55457586,0.5885295,0.56212115,0.6149379,0.60362,0.7507524,1.1657411,1.8485862,2.6936543,2.3126192,1.6222287,1.146878,1.0902886,1.3241913,1.6335466,1.720317,1.599593,1.5920477,2.3390274,2.795515,3.731126,4.5309224,5.270357,6.7152724,10.574668,14.947141,18.79899,20.764528,19.153618,15.716756,14.679284,14.720782,15.011275,15.196134,15.9695215,16.459963,16.493916,16.607096,18.029375,18.274595,19.40261,19.779873,18.71222,16.467508,14.886778,14.369928,14.377474,13.845533,11.204697,11.249968,9.073163,6.749226,5.4476705,5.462761,5.5080323,5.7494807,5.3948536,4.534695,4.1762958,3.5236318,2.9954643,2.4786146,2.2786655,3.108643,3.6556737,3.9914372,4.1083884,4.032936,3.8405323,3.6179473,3.802806,4.4818783,5.3910813,5.938112,6.5455046,7.062354,6.7454534,6.4511886,8.616675,10.853842,11.759273,13.634267,15.192361,11.548005,6.903904,4.8553686,3.4557245,2.0598533,1.3430545,0.9016574,0.8526133,0.814887,0.6111652,0.27917424,0.2867195,0.49421388,0.9808825,1.6184561,2.052308,1.7354075,1.9542197,2.0183544,1.659955,1.0148361,0.633801,0.8601585,1.2185578,1.5279131,1.8863125,2.282438,2.8709676,2.6483827,1.659955,0.9808825,1.4600059,1.7467253,2.0447628,2.4295704,2.8407867,2.2711203,1.5505489,1.2525115,1.6410918,2.6785638,3.6292653,4.168751,4.22534,4.002755,3.9801195,3.0671442,2.9728284,3.4972234,4.4177437,5.455216,8.677037,11.404645,13.528633,14.928277,15.467763,15.294222,14.128481,13.234368,13.008011,12.958967,15.105591,21.043703,26.438557,29.13221,29.13221,28.728539,28.879444,28.245644,26.468737,24.148573,23.371412,22.684793,21.130472,18.602814,15.8676605,12.875969,10.79348,8.688355,7.5037513,10.069136,17.029629,20.956932,22.232079,22.341486,23.861853,26.604551,29.37366,29.754694,27.343987,23.741129,20.972023,19.998686,18.889534,18.55377,22.737612,28.449366,31.807001,37.386715,47.878384,64.089355,92.11241,80.922806,57.78907,41.56301,42.67216,60.96562,64.91556,70.06519,80.771904,90.1846,74.64139,51.45106,31.939043,20.183544,12.996693,6.6850915,4.689373,4.534695,5.7419353,9.827688,12.264804,13.81158,15.082954,14.792462,9.767326,6.0512905,11.423509,13.732355,9.065618,1.7240896,2.3918443,2.173032,2.0296721,2.3805263,3.1010978,3.3048196,4.689373,5.2779026,4.5724216,3.5689032,3.7084904,2.7728794,2.1881225,2.305074,2.4031622,2.9916916,4.5422406,4.878004,3.9612563,3.8707132,4.7572803,6.0211096,7.043491,7.7414265,8.567632,11.204697,10.770844,11.038701,11.864905,9.220296,8.831716,7.8998766,7.594294,8.43559,10.321902,10.352083,12.162943,12.917468,12.596795,14.000212,14.66042,12.419481,11.498961,12.385528,11.827179,13.656902,16.4826,18.116146,17.308804,13.743673,11.02361,10.303039,9.699419,8.571404,7.5226145,5.194905,3.2821836,2.7502437,3.2369123,3.0520537,4.3121104,5.624984,7.5829763,10.26154,13.230596,13.822898,14.592513,14.78869,14.498198,14.641558,13.422999,13.736128,15.131999,18.361366,25.35204,33.01424,32.972744,33.821583,38.793903,45.780804,36.76423,27.132719,22.526344,23.465727,25.35204,23.31105,20.613623,16.41092,11.087745,6.2399216,7.6622014,14.475562,14.818871,9.122208,10.11818,14.743419,12.860879,10.763299,10.544487,10.11818,11.031156,15.211224,16.893814,16.622187,21.277605,22.53389,24.710693,21.639776,15.411173,16.380737,13.079691,12.985375,13.479589,12.668475,9.382519,17.7502,19.508244,18.26705,15.878979,12.449662,10.7218,9.480607,8.643084,8.160188,7.9828744,7.605612,6.221059,5.4174895,5.6778007,6.368191,6.48137,6.537959,5.247721,3.3274553,3.4745877,1.720317,1.3770081,1.750498,2.3578906,2.9464202,6.3455553,9.42779,10.054046,9.020347,10.069136,9.639057,8.360137,6.952948,5.9003854,5.451443,5.2967653,5.3269467,5.1156793,5.13077,6.7341356,7.8131065,12.098808,16.459963,16.837225,8.231868,7.4282985,8.710991,8.933576,7.6207023,6.9755836,6.0286546,7.4282985,8.499724,7.5226145,3.7160356,3.7348988,2.535204,2.5125682,4.376245,7.152897,8.892077,8.952439,9.97482,11.457462,9.740918,9.65792,9.733373,10.133271,10.623712,10.56335,13.026875,12.868423,12.702429,13.445636,14.302021,12.570387,12.555296,12.691111,12.3893,12.0082655,10.201178,9.906913,8.956212,7.001992,5.5080323,4.0404816,3.9386206,4.402653,4.606375,3.7047176,3.712263,3.6179473,3.7499893,3.9763467,3.712263,3.350091,2.8143783,2.2862108,1.8636768,1.5580941,1.3996439,1.2487389,1.1355602,1.0412445,0.91297525,0.8337501,0.84884065,0.8639311,0.8865669,0.995973,0.95447415,0.91674787,0.9393836,1.0110635,1.0638802,0.95824677,0.8224323,0.73566186,0.68661773,0.58475685,0.40367088,0.3169005,0.32444575,0.422534,0.6187105,0.633801,0.87902164,1.0714256,1.146878,1.2487389,1.1883769,1.2185578,1.3770081,1.5505489,1.4826416,1.9844007,2.3654358,1.901403,1.1280149,1.8636768,1.6863633,1.5128226,2.8898308,4.9723196,4.5233774,9.525878,5.070408,1.3091009,1.5015048,2.003264,3.8669407,2.5767028,2.535204,4.08198,3.5236318,3.4670424,2.7879698,2.4861598,2.927557,3.8480775,4.1272516,4.323428,4.6026025,4.851596,4.659192,5.3873086,5.1345425,4.881777,4.949684,4.991183,5.1345425,5.6476197,5.5985756,4.930821,4.4441524,4.466788,3.561358,2.71629,2.3314822,2.1994405,1.8523588,1.4524606,1.1619685,1.0450171,1.0450171,0.9205205,0.9620194,1.0487897,1.1204696,1.2110126,1.3543724,1.4524606,1.448688,1.3166461,1.0638802,0.8903395,0.9393836,0.97710985,0.94315624,0.91297525,0.9016574,1.0186088,1.0978339,1.0978339,1.086516,1.2826926,1.2638294,1.3015556,1.3920987,1.2487389,1.3958713,1.146878,0.814887,0.56589377,0.392353,0.39989826,0.38103512,0.362172,0.32821837,0.20372175,0.24522063,0.32821837,0.55457586,0.87147635,1.0789708,1.0412445,1.0299267,0.8903395,0.65643674,0.55457586,0.56212115,0.66775465,0.77716076,0.80734175,0.6790725,0.6790725,0.58098423,0.5017591,0.5017591,0.62625575,0.7394345,0.69793564,0.62625575,0.59607476,0.59230214,0.49044126,0.39989826,0.35462674,0.35085413,0.35462674,0.4678055,0.5885295,0.79602385,1.1280149,1.5656394,1.448688,1.4524606,1.4864142,1.5543215,1.7618159,1.9844007,2.727608,3.3463185,3.6783094,4.0404816,3.640583,3.3236825,3.1576872,3.0520537,2.7389257,3.0897799,3.731126,4.3309736,4.5233774,3.9008942,3.4594972,3.289729,2.957738,2.4597516,2.2069857,2.0975795,2.0108092,1.7844516,1.478869,1.3845534,1.327964,1.4675511,1.478869,1.3656902,1.4750963,1.7467253,1.9429018,2.1088974,2.2673476,2.425798,2.7540162,3.2255943,3.6481283,4.0178456,4.496969,4.587512,4.4894238,4.3913355,4.3686996,4.38379,4.5233774,4.459243,4.5950575,5.1043615,5.934339,6.405917,6.971811,7.4509344,7.699928,7.6320205,7.152897,6.617184,6.1795597,5.881522,5.6513925,5.704209,6.1833324,6.94163,7.9036493,9.073163,9.989911,10.246449,10.137043,9.80128,9.239159,9.114662,9.390063,9.899368,10.393582,10.544487,11.593277,12.989148,13.947394,14.27184,14.358611,1.8448136,1.0940613,0.80356914,0.59230214,0.331991,0.15467763,0.15845025,0.13958712,0.12826926,0.12826926,0.10940613,0.1358145,0.116951376,0.09808825,0.090543,0.0754525,0.07922512,0.071679875,0.08299775,0.120724,0.16976812,0.2263575,0.2867195,0.32444575,0.30935526,0.18485862,0.22258487,0.13204187,0.056589376,0.05281675,0.08677038,0.26408374,0.46026024,0.58098423,0.6375736,0.7394345,0.633801,0.6149379,0.80356914,1.2411937,1.8749946,1.5128226,1.0751982,0.8865669,1.0601076,1.4901869,1.7240896,1.7089992,1.4713237,1.4750963,2.6521554,3.4859054,4.557331,6.085244,8.409182,11.996947,15.871433,18.500954,19.862871,19.319613,15.656394,12.966512,12.079946,12.619431,13.800262,14.445381,15.648849,20.066593,23.163918,24.148573,25.940569,29.17371,31.048704,29.566063,25.574625,22.771564,19.059301,15.961976,13.754991,11.7026825,8.07719,9.016574,8.265821,6.888813,5.9192486,6.330465,5.560849,5.3910813,5.1269975,4.67051,4.496969,3.6179473,2.6332922,1.8485862,1.5618668,2.0560806,2.6974268,3.3274553,3.802806,3.821669,2.9237845,2.2975287,2.7426984,3.500996,4.115934,4.395108,4.515832,4.52715,4.7044635,5.462761,7.360391,8.963757,8.00551,6.6247296,5.1647234,2.173032,2.8407867,3.2331395,2.3654358,0.8337501,0.8299775,0.6526641,0.62248313,0.5055317,0.29803738,0.211267,0.24899325,0.41121614,0.8941121,1.569412,1.991946,1.5845025,1.5618668,1.5958204,1.5618668,1.5279131,1.2600567,1.478869,1.81086,2.203213,2.9539654,3.3123648,3.772625,3.410453,2.3503454,1.7580433,1.8523588,1.9391292,2.3993895,3.218049,3.9650288,3.8669407,3.3576362,3.1840954,3.904667,5.885295,7.3717093,7.273621,6.722818,6.258785,5.847569,5.3646727,5.413717,5.666483,6.1116524,7.0359454,12.136535,14.558559,15.079182,14.803781,15.184815,17.701157,17.565342,14.66042,11.272603,12.0724,16.38451,23.416683,28.472,30.25268,30.852528,26.44233,25.665169,26.868635,27.442074,23.824127,23.09601,23.420456,22.160398,19.104572,16.467508,13.856852,13.241914,11.370691,8.918486,10.499215,18.75372,24.024076,24.695602,22.975286,24.90687,28.109829,30.811028,30.690304,27.415667,22.647068,19.496925,17.286167,15.754482,15.939341,20.16468,26.604551,30.965706,35.06278,42.102493,56.68369,80.247505,71.2347,50.983253,35.606033,35.983295,52.654526,56.13666,60.554405,70.58204,81.43211,70.182144,46.999363,27.29494,17.135263,13.223051,8.197914,5.323174,4.568649,6.149379,10.54826,11.570641,13.404137,14.807553,14.385019,10.593531,8.91094,14.011529,16.32792,11.819634,1.9693103,2.7426984,2.3918443,2.263575,2.8181508,3.6330378,3.6292653,5.353355,5.855114,4.636556,3.6707642,3.8103511,2.9954643,2.2899833,2.1051247,2.1881225,3.4859054,5.594803,6.628502,6.25124,5.6589375,4.8855495,5.2364035,6.006019,6.9454026,8.2507305,10.729345,10.691619,11.672502,12.974057,9.635284,8.126234,7.333983,6.9944468,7.3188925,8.986393,9.152389,10.616167,11.740409,12.925014,16.618414,15.30554,12.679792,11.544232,12.404391,13.434318,14.102073,16.01102,17.169216,16.467508,13.713491,11.16697,10.057818,9.439108,8.76758,7.914967,5.7683434,3.9688015,2.7351532,2.0636258,1.7278622,2.4069347,3.259548,4.745962,6.8774953,9.208978,10.246449,12.608112,13.241914,11.830952,10.808571,11.046246,12.672247,14.498198,17.7917,26.280106,33.47073,36.84723,38.016743,40.05396,47.519985,44.62261,32.791656,24.544699,23.84299,26.07261,22.647068,20.323132,16.429781,11.106608,7.3151197,8.529905,13.257004,12.936331,8.869441,12.189351,12.58925,9.74469,8.541223,9.786189,10.18986,8.299775,10.940613,16.101564,20.519308,19.666695,21.005976,25.329405,22.005722,12.951422,12.623203,9.578695,10.38981,10.506761,9.273112,9.906913,18.474545,22.039675,20.790936,16.101564,10.518079,8.695901,8.175279,9.110889,10.469034,10.038955,8.348819,6.3945994,5.406172,5.6400743,6.379509,6.571913,6.752999,6.1531515,5.05909,4.821415,2.493705,2.04099,2.2409391,2.867195,4.7120085,8.360137,10.355856,10.529396,9.891823,10.61994,11.09529,10.510533,8.843033,6.79827,5.798525,5.6589375,5.66271,5.2250857,4.817642,5.9796104,6.741681,10.33322,15.128226,17.003222,9.322156,9.88805,11.174516,9.827688,6.8133607,7.4094353,7.149124,8.533678,9.242931,8.43559,6.749226,5.975838,3.6745367,2.6597006,3.9008942,6.530414,8.797762,9.310839,9.58624,9.922004,9.405154,9.190115,9.88805,10.280403,10.080454,9.929549,11.027383,10.672756,10.710483,11.672502,12.774108,11.774363,12.385528,13.219278,13.389046,12.491161,13.302276,11.4838705,9.190115,7.405663,5.934339,4.063117,4.006528,4.689373,5.070408,4.1574326,4.06689,4.032936,4.557331,5.119452,4.2064767,3.6858547,3.2444575,2.7879698,2.3390274,2.0108092,1.5731846,1.3505998,1.237421,1.1506506,1.0110635,0.935611,0.935611,0.9507015,0.97710985,1.086516,1.0827434,1.0374719,1.0186088,1.0638802,1.20724,1.1053791,0.87147635,0.754525,0.76207024,0.63002837,0.3961256,0.331991,0.33953625,0.392353,0.5394854,0.6149379,0.9016574,1.0487897,1.026154,1.1242423,1.026154,1.1091517,1.2940104,1.4675511,1.4600059,1.8825399,2.6634734,2.2598023,1.1431054,1.7919968,1.7354075,1.4562333,2.9086938,4.9723196,3.4557245,9.710737,6.5643673,2.4522061,1.2185578,2.1315331,4.6516466,2.6446102,1.9089483,3.3953626,3.2369123,2.7728794,2.4823873,2.2371666,2.3692086,3.6594462,3.4859054,3.7650797,3.9273026,3.783943,3.5424948,4.515832,4.610148,4.5233774,4.6214657,4.961002,4.504514,4.851596,4.9760923,4.508287,3.7348988,3.7386713,2.938875,2.2296214,1.9278114,1.7844516,1.6260014,1.4147344,1.1959221,1.0638802,1.1355602,0.8639311,0.79602385,0.8299775,0.9016574,0.97333723,1.116697,1.1808317,1.1204696,0.9695646,0.80734175,0.7130261,0.7696155,0.8941121,0.9997456,0.9922004,0.97333723,1.0638802,1.1846043,1.2487389,1.1959221,1.4335974,1.4411428,1.5165952,1.5958204,1.2411937,1.1280149,0.8111144,0.4979865,0.29426476,0.19240387,0.21503963,0.19994913,0.211267,0.24522063,0.24899325,0.33953625,0.44894236,0.66020936,0.9808825,1.3166461,1.1053791,0.88279426,0.663982,0.52062225,0.56212115,0.58475685,0.6375736,0.67152727,0.65643674,0.58098423,0.6149379,0.5583485,0.482896,0.47535074,0.6073926,0.8111144,0.76207024,0.6413463,0.56589377,0.60362,0.5357128,0.42630664,0.3734899,0.41121614,0.47535074,0.59230214,0.62248313,0.7205714,0.91674787,1.1242423,1.1317875,1.2261031,1.3128735,1.4298248,1.7655885,2.0975795,2.5540671,2.938875,3.2444575,3.6556737,3.610402,3.6066296,3.482133,3.187868,2.7879698,3.048281,3.482133,4.063117,4.425289,3.863168,3.4594972,3.1614597,2.7011995,2.1390784,1.8636768,1.9579924,1.8863125,1.6071383,1.2826926,1.2940104,1.2487389,1.3166461,1.3468271,1.3543724,1.5241405,1.871222,1.9429018,1.9164935,1.9579924,2.1994405,2.595566,2.927557,3.169005,3.410453,3.8556228,4.0103,3.9763467,4.063117,4.247976,4.1574326,4.074435,4.1272516,4.4516973,5.0062733,5.5495315,6.058836,6.6360474,7.213259,7.6093845,7.533932,6.888813,6.360646,5.938112,5.594803,5.2665844,5.4665337,6.043745,6.790725,7.665974,8.805306,9.435335,9.57115,9.288202,8.7600355,8.258276,8.224322,8.416726,8.748717,9.027891,8.937348,10.321902,11.978085,13.151371,13.536179,13.27964,2.9766011,1.5807298,0.91297525,0.7167987,0.6488915,0.27540162,0.20749438,0.20372175,0.181086,0.124496624,0.1056335,0.1659955,0.14713238,0.08677038,0.041498873,0.0754525,0.026408374,0.018863125,0.0452715,0.11317875,0.26408374,0.24522063,0.16976812,0.17731337,0.23767537,0.17354076,0.29803738,0.20749438,0.08677038,0.02263575,0.02263575,0.10940613,0.27540162,0.47157812,0.68661773,0.9507015,0.875249,0.69793564,0.7582976,1.0487897,1.2185578,1.0487897,0.8262049,0.7922512,1.0638802,1.6637276,1.8033148,1.6410918,1.1808317,0.90543,1.7769064,3.1765501,4.221567,6.628502,10.521852,14.449154,16.026112,15.124454,13.505998,11.714001,9.065618,8.544995,7.9489207,9.431562,13.079691,16.908905,18.968758,27.1629,33.71595,36.107796,37.06604,41.28761,43.143738,40.193546,33.90835,29.679241,24.133482,18.734856,14.449154,11.46878,9.22784,7.5490227,7.7904706,7.9489207,7.6131573,7.9753294,6.085244,5.1345425,4.636556,4.323428,4.146115,3.4142256,2.0749438,1.3204187,1.4713237,1.9768555,2.3428001,2.4295704,2.41448,2.233394,1.5882751,1.5543215,2.384299,3.2520027,3.7877154,4.0782075,4.006528,4.1612053,4.425289,4.9987283,6.417235,8.031919,7.6810646,7.1038527,6.1342883,2.7313805,2.7540162,2.704972,1.9429018,0.87147635,0.94315624,0.80734175,0.76584285,0.7092535,0.58475685,0.42630664,0.49421388,0.66775465,1.0827434,1.5203679,1.4147344,1.3355093,1.5203679,1.7769064,2.0560806,2.4672968,2.4182527,2.1088974,1.9994912,2.4786146,3.8556228,4.349837,4.217795,3.9348478,3.8707132,4.304565,3.4934506,2.9841464,3.1161883,3.7462165,4.221567,4.930821,5.270357,5.745708,6.9491754,9.574923,10.367173,9.088254,8.179051,8.152642,7.6131573,7.726336,8.503497,8.922258,8.990166,9.759781,14.966003,15.731846,14.581196,13.970031,16.28265,21.847271,24.307022,20.330677,14.188843,17.77661,21.854816,24.250433,25.559534,27.01954,30.494127,24.435291,22.556524,23.348776,24.012758,20.4514,21.439827,21.09652,20.647577,19.647831,15.99593,12.306303,12.777881,12.400619,10.842525,12.449662,17.818108,24.435291,25.921707,23.046967,23.737356,28.075874,30.41113,29.913143,26.427238,20.458946,18.12369,16.87118,16.158154,16.580687,19.87419,24.291933,30.562035,35.496628,40.47272,51.42088,60.56195,53.601456,40.333134,29.928234,30.935526,45.44504,48.22169,52.20936,62.116272,74.41503,65.4475,42.4873,23.23937,14.551015,12.404391,9.812597,6.56814,4.979865,5.975838,9.084481,8.575176,8.733627,10.287949,12.257258,11.978085,13.766309,17.63325,18.059555,12.698656,2.3767538,3.5764484,2.9124665,2.837014,3.8669407,4.557331,3.9914372,5.5759397,5.8664317,4.395108,3.6669915,3.2105038,2.9011486,2.3767538,1.7316349,1.4826416,3.1237335,5.4363527,7.3075747,8.137552,7.8206515,5.553304,4.7950063,4.9119577,5.4967146,6.3832817,8.058327,8.590267,10.597303,12.913695,10.597303,8.197914,6.56814,5.523123,5.2137675,6.126743,6.560595,7.8131065,9.374973,11.947904,17.437073,15.301767,12.958967,12.366665,13.88326,16.263786,15.165953,15.343266,15.531898,15.045229,13.754991,11.261286,9.291975,8.439363,8.394091,7.9451485,6.7756343,5.7381625,4.564876,3.3651814,2.637065,2.9766011,3.3161373,3.5462675,4.115934,5.9984736,7.726336,11.363147,12.566614,11.208468,11.344283,12.702429,14.154889,15.814844,18.387774,23.182781,32.361576,38.280827,40.24259,42.15154,52.488533,60.958076,47.719933,30.863846,21.353058,23.005466,21.760502,16.422237,11.321648,9.291975,11.672502,6.907676,10.801025,14.656648,14.030393,8.741172,10.827434,8.062099,6.428553,7.5490227,8.669493,7.0548086,7.1000805,15.026365,24.586197,17.063583,20.892797,23.141281,19.56106,12.913695,12.958967,9.65792,8.718536,7.8131065,7.798016,12.725064,16.52787,20.33822,19.960958,15.256495,10.174769,8.13378,7.9753294,9.22784,10.570895,9.869187,6.5530496,5.0213637,4.564876,4.7308717,5.2967653,4.949684,4.8629136,5.7079816,6.8171334,6.2021956,3.5462675,3.180323,3.2482302,3.8895764,7.2358947,10.661438,10.729345,9.963503,9.895596,11.038701,12.181807,12.653384,11.348056,8.718536,6.802043,6.255012,5.8664317,5.5759397,5.323174,5.0515447,4.919503,7.424526,11.129244,13.008011,8.428044,12.106354,14.241659,12.049765,7.877241,9.193887,9.525878,9.046755,8.379,8.14887,8.99771,7.2396674,5.4401255,4.776143,5.6325293,7.6093845,8.371455,7.677292,6.466279,6.089017,8.307321,7.5829763,9.107117,9.812597,9.152389,9.0957985,8.922258,8.850578,8.7751255,9.031664,10.38981,10.967021,12.325166,13.6833105,13.905896,11.498961,14.992412,12.479843,8.963757,6.881268,6.1078796,4.085753,3.9008942,4.5196047,4.9421387,4.2102494,4.2517486,4.4441524,5.2364035,5.8966126,4.52715,3.742444,3.5990841,3.399135,2.9313297,2.4786146,1.7882242,1.478869,1.3920987,1.3694628,1.2487389,1.0789708,1.0638802,1.0827434,1.0978339,1.1280149,1.0902886,1.0978339,1.1016065,1.1506506,1.3732355,1.267602,0.94315624,0.7922512,0.814887,0.62625575,0.35462674,0.34330887,0.36594462,0.3772625,0.5017591,0.60362,0.73188925,0.8224323,0.9205205,1.1695137,1.1016065,1.0827434,1.2902378,1.599593,1.5731846,1.6373192,2.7200627,2.6144292,1.4449154,1.690136,1.6637276,1.5958204,2.9615107,4.745962,3.4217708,7.8923316,7.6282477,4.1008434,0.513077,1.7693611,4.8553686,2.938875,1.5958204,2.3692086,2.7992878,1.8448136,2.3126192,2.305074,1.961765,3.4896781,2.957738,3.4029078,3.7273536,3.429316,2.625747,2.9501927,3.3689542,3.863168,4.4139714,5.0175915,3.9348478,3.8858037,3.9876647,3.7084904,2.8785129,2.5729303,2.2183034,1.8900851,1.5958204,1.2864652,1.3053282,1.3317367,1.1883769,0.98465514,1.0827434,0.9205205,0.8299775,0.8186596,0.8639311,0.9016574,1.0336993,1.0487897,0.9620194,0.84129536,0.8111144,0.7394345,0.80356914,0.9808825,1.1506506,1.0902886,1.0336993,1.0714256,1.2411937,1.4562333,1.4939595,1.5618668,1.5316857,1.6071383,1.6373192,1.1242423,0.8978847,0.5357128,0.27540162,0.17731337,0.14335975,0.1659955,0.16222288,0.1659955,0.211267,0.32821837,0.47912338,0.59607476,0.6413463,0.72811663,1.1091517,0.90920264,0.62248313,0.47535074,0.5319401,0.6752999,0.7205714,0.69039035,0.70170826,0.754525,0.7469798,0.58475685,0.47912338,0.43007925,0.43007925,0.452715,0.6752999,0.7205714,0.663982,0.5885295,0.62625575,0.5394854,0.45648763,0.44894236,0.543258,0.72811663,0.84884065,0.7130261,0.65643674,0.7507524,0.79602385,0.90543,1.237421,1.4562333,1.539231,1.7580433,2.1768045,2.41448,2.757789,3.289729,3.8971217,4.0970707,4.1762958,3.874486,3.2935016,2.886058,3.3274553,3.4859054,3.682082,3.893349,3.742444,3.5160866,3.1124156,2.674791,2.2598023,1.8636768,1.8146327,1.7052265,1.5052774,1.3053282,1.3053282,1.2147852,1.1657411,1.1506506,1.1732863,1.2223305,1.5241405,1.539231,1.5656394,1.7467253,2.0673985,2.5012503,2.795515,2.9803739,3.108643,3.2557755,3.5236318,3.7198083,4.0970707,4.534695,4.5309224,4.425289,4.5799665,4.878004,5.2175403,5.4967146,5.9720654,6.4964604,6.9982195,7.3490734,7.375482,6.779407,6.3719635,6.0776987,5.824933,5.572167,5.726845,6.187105,6.8963585,7.7829256,8.729855,9.027891,8.786444,8.262049,7.7829256,7.748972,7.816879,7.809334,7.835742,7.9489207,8.171506,10.121953,11.46878,12.332711,12.67602,12.325166,1.0827434,1.0450171,0.9016574,0.9016574,0.95824677,0.6413463,0.49421388,0.38480774,0.2678564,0.1659955,0.1659955,0.120724,0.07922512,0.049044125,0.041498873,0.0754525,0.0150905,0.0,0.056589376,0.17731337,0.33576363,0.19994913,0.150905,0.17354076,0.211267,0.1358145,0.22258487,0.18863125,0.10940613,0.0452715,0.0452715,0.0452715,0.1358145,0.31312788,0.48666862,0.47157812,0.4979865,0.40367088,0.33576363,0.38858038,0.59607476,0.5357128,0.4640329,0.62248313,1.0638802,1.6637276,1.478869,1.0035182,0.784706,1.116697,2.0447628,2.8521044,3.8103511,4.9459114,6.0286546,6.5756855,7.432071,7.0585814,5.9230213,4.708236,4.3196554,4.636556,4.478106,5.2288585,8.254503,14.909414,21.926497,30.878935,36.798183,37.579117,33.964943,30.852528,31.769276,31.878681,29.76224,27.41944,22.733839,20.63626,19.24416,16.675003,11.046246,7.5301595,7.220804,7.9828744,8.096053,6.2399216,5.3382645,4.67051,4.1612053,3.8141239,3.7537618,3.5689032,2.2447119,2.1315331,3.1010978,2.5012503,2.674791,3.2369123,3.4255435,2.9464202,1.9693103,2.323937,3.6481283,4.689373,5.0553174,5.1873593,4.0517993,3.6141748,4.0480266,5.3194013,7.1868505,6.858632,6.089017,4.7535076,3.3651814,3.097325,4.429062,3.0671442,2.1654868,2.674791,3.3727267,1.7618159,1.5128226,1.780679,1.9391292,1.5882751,1.5241405,1.8297231,2.3201644,2.4861598,1.50905,1.6071383,2.1466236,2.444661,2.3578906,2.2748928,2.372981,2.0372176,1.9353566,2.7728794,5.3080835,6.458734,5.3910813,5.1647234,6.6850915,8.710991,7.001992,5.0666356,3.6858547,3.2444575,3.7084904,5.0138187,6.228604,7.5716586,9.159933,11.000975,8.963757,8.107371,8.624221,9.688101,9.446653,8.443134,9.457971,11.057564,12.543978,13.947394,15.863888,14.320885,13.347548,15.173498,20.202406,25.499172,29.76224,28.577635,25.284132,30.95816,29.773556,25.140774,20.972023,19.666695,22.096264,24.133482,24.944597,23.65813,20.462717,16.618414,18.693357,18.489635,18.678267,18.218006,12.359119,9.333474,9.325929,9.861642,10.702937,13.837989,16.414692,21.97554,24.989868,24.601288,24.627695,27.336441,28.581408,27.336441,23.303505,16.905132,16.063837,17.867151,19.429018,20.145817,21.681276,23.405365,30.214954,35.191048,37.239582,41.10652,44.61129,39.144756,31.060022,25.61235,26.93277,39.714424,42.42317,44.686745,52.722435,69.337074,60.63363,38.095966,19.425245,10.963248,7.6923823,5.5306683,5.1835866,5.7192993,7.4509344,11.917723,10.38981,9.654147,12.068627,16.361876,17.591751,20.032639,21.451145,18.69713,11.778135,3.8292143,5.2326307,4.0178456,3.731126,4.9949555,5.5080323,4.9723196,5.8173876,5.855114,4.5724216,3.1425967,2.6182017,2.7087448,2.565385,1.9089483,1.0072908,1.5920477,2.565385,3.3651814,3.8178966,4.134797,2.5616124,1.7655885,1.780679,2.565385,3.9688015,4.908185,5.6098933,7.4169807,9.80128,10.374719,6.934085,5.168496,4.798779,5.0251365,4.5007415,4.183841,5.43258,7.115171,9.344792,13.456953,12.396846,12.128989,13.694629,15.773345,14.724555,15.237633,14.954685,13.6833105,12.449662,13.472044,11.461235,9.49947,8.360137,8.179051,8.484633,8.631766,9.782416,8.7751255,5.9682927,5.247721,6.0286546,5.2099953,4.3196554,4.5309224,6.6662283,7.364164,9.26934,10.533169,11.465008,14.539697,15.079182,13.758763,14.6302395,18.078419,20.813572,29.750921,33.878174,36.44733,42.28358,57.785297,74.018906,62.165314,41.8535,26.71773,24.397566,20.662666,14.366156,10.212496,8.646856,5.8136153,6.4134626,9.050528,12.15917,12.672247,6.043745,11.891314,8.07719,4.085753,4.006528,6.5455046,8.13378,9.1976595,11.676274,14.999957,16.097792,17.23335,16.939087,15.792209,16.720274,25.008732,14.169979,8.869441,7.8508325,9.639057,12.543978,12.800517,12.196897,12.566614,13.739901,13.517315,11.223559,10.47658,9.940866,8.880759,7.17176,5.0854983,4.0216184,3.5349495,3.942393,6.349328,4.45547,4.5761943,6.255012,8.080963,7.6886096,4.515832,4.45547,4.821415,5.330719,8.103599,9.752235,10.940613,11.642321,11.966766,12.162943,12.162943,11.566868,10.789707,9.646602,7.3377557,6.9491754,5.926794,5.523123,5.8437963,5.8437963,4.610148,6.0248823,7.3113475,7.062354,5.2175403,13.543724,17.795471,16.165699,12.551523,16.55428,12.442118,7.3679366,5.1760416,6.507778,8.790216,6.507778,6.7152724,7.092535,6.828451,6.620957,7.8319697,6.5040054,5.2892203,5.402399,6.620957,8.661947,9.756008,9.865415,9.133525,7.888559,8.926031,9.148616,9.061845,9.265567,10.438853,10.450171,10.223814,9.857869,9.7296,10.499215,10.325675,10.072908,8.096053,5.1534057,4.4101987,3.4330888,3.5839937,4.1800685,4.4441524,3.4783602,4.2102494,4.8063245,5.1534057,5.2364035,5.1269975,4.3196554,4.349837,4.274384,3.712263,2.806833,2.4899325,1.8259505,1.629774,1.8825399,1.7240896,1.0148361,0.7922512,0.8563859,0.995973,1.0072908,1.0072908,1.1242423,1.2525115,1.3732355,1.5580941,1.4713237,1.0110635,0.66775465,0.62625575,0.7469798,0.36971724,0.29426476,0.26408374,0.2565385,0.48666862,0.7205714,0.73188925,0.84884065,1.0336993,0.9016574,1.20724,1.2185578,1.3091009,1.4373702,1.1431054,0.83752275,1.7052265,2.071171,1.5203679,0.8865669,1.3845534,2.04099,3.3651814,4.8742313,5.081726,8.107371,9.084481,5.5683947,0.10940613,0.24522063,2.625747,3.0897799,2.5427492,2.1390784,3.3123648,2.1503963,2.3654358,2.3880715,1.9391292,1.9994912,2.1692593,2.3692086,2.516341,2.5276587,2.3201644,2.4408884,3.0935526,3.5538127,3.8443048,4.7610526,4.22534,3.4481792,2.9539654,2.7804246,2.4861598,2.0372176,1.7844516,1.7052265,1.6033657,1.1129243,0.9808825,0.965792,0.965792,0.9620194,1.0223814,0.935611,0.8526133,0.8526133,0.9507015,1.0827434,0.9620194,0.9318384,0.9620194,0.995973,0.94692886,0.77338815,0.8526133,0.9620194,0.9922004,0.9318384,0.8941121,0.95824677,1.0789708,1.2638294,1.5580941,1.4939595,1.5430037,1.5580941,1.4071891,0.9922004,0.6375736,0.3772625,0.23390275,0.19240387,0.1659955,0.14335975,0.14713238,0.21503963,0.35462674,0.55080324,0.66020936,0.8224323,0.83752275,0.72811663,0.77716076,0.76584285,0.5998474,0.52439487,0.56589377,0.5017591,0.5885295,0.63002837,0.63002837,0.62625575,0.68661773,0.55080324,0.5281675,0.6073926,0.67152727,0.48666862,0.67152727,0.7167987,0.6375736,0.5281675,0.56589377,0.5281675,0.65643674,0.7092535,0.7054809,0.9016574,0.8639311,0.72811663,0.663982,0.73566186,0.87147635,1.2223305,1.3317367,1.4298248,1.6109109,1.8297231,2.2220762,2.757789,3.3764994,3.9574835,4.349837,4.617693,4.610148,3.9876647,3.059599,2.776652,3.0822346,3.240685,3.2972744,3.229367,2.9615107,2.8521044,2.8596497,2.5917933,2.071171,1.7542707,1.4600059,1.4524606,1.4298248,1.2826926,1.0978339,1.0374719,1.0676528,1.0978339,1.086516,1.0374719,1.146878,1.3392819,1.5882751,1.8749946,2.1654868,2.2748928,2.505023,2.8407867,3.108643,2.9766011,3.1350515,3.4217708,3.9197574,4.5196047,4.8968673,4.8138695,4.689373,4.719554,4.9345937,5.20245,5.726845,6.2361493,6.7114997,7.118943,7.4018903,7.0585814,6.670001,6.432326,6.3644185,6.3153744,6.3644185,6.85486,7.5301595,8.182823,8.620448,8.096053,7.6093845,7.164215,6.7831798,6.515323,6.907676,7.066127,7.1906233,7.4396167,7.964011,9.016574,9.7069645,10.386037,11.117926,11.7026825,0.9016574,0.68661773,0.68661773,0.7696155,0.8639311,0.94692886,1.0223814,0.76584285,0.4640329,0.2678564,0.181086,0.16976812,0.09808825,0.03772625,0.018863125,0.0150905,0.003772625,0.030181,0.22258487,0.47912338,0.482896,0.27917424,0.18863125,0.13958712,0.116951376,0.16222288,0.150905,0.14335975,0.116951376,0.071679875,0.02263575,0.07922512,0.23013012,0.35839936,0.38480774,0.26408374,0.24899325,0.2263575,0.21503963,0.22258487,0.26408374,0.26408374,0.33953625,0.5696664,0.97333723,1.5052774,0.9393836,0.5885295,0.70170826,1.3091009,2.2296214,3.180323,4.7572803,5.9192486,6.590776,7.6395655,7.6923823,6.907676,6.221059,6.0362,6.2097406,5.6287565,5.4363527,7.828197,13.128735,19.80251,25.42372,27.045948,28.728539,30.399813,27.849518,26.291424,24.408884,22.107582,20.489126,21.854816,20.281631,19.636513,19.1008,17.818108,14.905642,12.864652,11.332966,10.27663,9.295748,7.6093845,6.304056,6.2361493,5.9532022,5.0666356,4.255521,3.92353,3.0218725,2.4823873,2.516341,2.6106565,2.1881225,2.5389767,2.9426475,3.1124156,3.2029586,3.429316,4.0103,4.432834,4.587512,4.7610526,5.2062225,5.5382137,5.0779533,4.8100967,7.383027,9.239159,8.7600355,6.643593,3.92353,1.9881734,2.4861598,2.9464202,3.5047686,3.7273536,2.6144292,1.629774,1.4864142,1.5845025,2.0108092,3.5538127,3.0331905,2.686109,2.516341,2.293756,1.5731846,2.022127,2.2371666,2.203213,2.1579416,2.5917933,2.2484846,3.2142766,3.772625,3.7613072,4.5535583,4.3422914,3.3915899,3.6858547,5.9003854,9.371201,9.812597,8.805306,7.213259,5.5004873,3.7575345,5.5004873,7.118943,8.786444,10.397354,11.5857315,10.427535,8.816625,6.9454026,5.1798143,4.036709,5.6815734,9.408927,13.053283,16.124199,19.794964,20.274086,16.607096,15.531898,18.474545,21.519053,22.7942,25.842482,27.087448,26.359331,26.857317,23.488363,19.410156,18.293459,19.783646,19.519562,20.474035,24.031622,24.276842,20.972023,19.557287,23.635496,24.076893,21.915178,18.863125,17.338985,11.559323,10.27663,11.038701,12.536433,14.607604,17.067356,22.24717,26.321604,27.834427,27.702385,28.566317,26.78941,23.710949,19.753464,14.392565,15.531898,18.30855,20.470263,21.35683,21.877453,22.14531,27.34776,33.42923,37.299942,36.83591,33.425457,28.653088,24.291933,22.10381,23.84299,34.34975,36.285107,36.869865,43.2041,62.267174,54.97092,35.489082,18.731083,10.133271,5.6513925,5.0062733,4.134797,4.0291634,5.062863,7.020855,7.360391,11.879996,18.863125,24.510744,22.95265,29.426476,24.85028,16.65614,9.405154,4.768598,6.7114997,5.4476705,4.919503,5.836251,5.6551647,5.9682927,6.8925858,6.3908267,4.617693,3.9122121,3.4179983,3.1463692,2.7125173,1.9768555,1.056335,0.7922512,0.9507015,1.4449154,2.6974268,5.613666,2.9916916,1.3053282,0.86770374,1.659955,3.308592,4.5309224,8.797762,13.781399,15.784663,9.7296,8.922258,7.6018395,6.0362,4.5761943,3.6594462,3.380272,3.6707642,6.802043,10.868933,9.808825,11.627231,11.744182,12.823153,15.094273,16.361876,17.57666,15.762027,13.721037,12.706201,12.411936,10.533169,9.261794,8.578949,8.299775,8.069645,11.936585,11.59705,9.5032425,7.4471617,6.530414,7.7602897,8.963757,8.254503,6.330465,6.485142,7.816879,8.744945,10.416218,12.626976,13.807808,11.359374,11.1782875,14.5132885,19.625195,21.813318,23.767538,24.378702,25.472763,28.78513,35.949345,49.87033,49.764698,41.759186,32.659615,29.939552,26.476282,17.056038,8.9788475,5.3080835,4.847823,4.8138695,7.7187905,11.536687,12.811834,6.63982,6.579458,3.9348478,2.0787163,2.173032,3.187868,8.439363,8.98262,8.7751255,9.906913,12.608112,13.030646,17.421982,19.002712,17.16167,17.440845,13.045737,10.469034,8.699674,7.4584794,7.2094865,7.84706,7.594294,8.869441,11.291467,11.6875925,9.929549,7.9753294,6.971811,6.643593,5.304311,4.447925,3.7801702,3.7084904,4.8365054,7.9828744,5.7607985,6.326692,8.511042,10.514306,9.899368,6.1606965,4.402653,3.7650797,4.0517993,5.7570257,6.9189944,6.9454026,6.7680893,7.0585814,8.22055,8.929804,8.069645,7.6093845,8.14887,8.8769865,8.6732645,7.3151197,6.3417826,6.530414,7.907422,7.466025,8.314865,9.156161,8.714764,5.7192993,11.321648,12.89106,14.437836,17.056038,18.912169,11.114153,6.488915,5.191132,6.058836,6.590776,5.481624,5.372218,6.0739264,6.8850408,6.598321,7.492433,6.4474163,5.696664,6.0814714,7.0510364,8.971302,9.782416,9.420244,8.714764,9.367428,9.1825695,9.510788,9.559832,9.556059,10.718028,9.997457,10.578441,11.133017,11.16697,10.997202,9.918231,9.865415,9.442881,8.141325,6.3153744,4.4177437,4.3083377,4.557331,4.3121104,3.31991,3.3576362,3.591539,3.832987,4.134797,4.798779,3.953711,3.8593953,3.6443558,3.1237335,2.795515,2.5578396,2.0145817,1.6712729,1.5279131,1.0789708,0.70170826,0.663982,0.754525,0.87902164,1.0676528,1.0299267,1.056335,1.1808317,1.3920987,1.6524098,1.5505489,1.1695137,0.8601585,0.7469798,0.7582976,0.46026024,0.32821837,0.26408374,0.271629,0.4640329,0.5772116,0.5319401,0.6828451,0.9242931,0.694163,0.9393836,1.1846043,1.1883769,1.0940613,1.4260522,1.1091517,1.690136,1.9768555,1.6184561,1.0940613,1.7278622,2.8898308,4.0970707,5.1458607,6.1078796,6.5945487,10.314357,7.8131065,0.392353,0.09808825,1.3845534,3.2633207,2.9426475,1.237421,2.565385,2.1994405,2.2560298,2.3013012,2.0560806,1.4147344,1.8787673,2.022127,2.214531,2.4107075,2.173032,2.335255,2.8294687,3.199186,3.3576362,3.5877664,3.7348988,3.4029078,2.8143783,2.252257,2.0485353,1.6146835,1.3920987,1.3091009,1.2336484,0.9808825,0.77716076,0.80356914,0.83752275,0.8262049,0.875249,0.84884065,0.7507524,0.72811663,0.8186596,0.9242931,0.8601585,0.845068,0.9507015,1.1280149,1.2147852,1.0336993,0.9393836,0.8526133,0.7884786,0.845068,0.98465514,1.1016065,1.1393328,1.1695137,1.3845534,1.2185578,1.2185578,1.3204187,1.3166461,0.8337501,0.51684964,0.38858038,0.31312788,0.24522063,0.23013012,0.21503963,0.2263575,0.30935526,0.43385187,0.5017591,0.59230214,0.7054809,0.8224323,0.87902164,0.80356914,0.73188925,0.6149379,0.5772116,0.62248313,0.6375736,0.6752999,0.7394345,0.7432071,0.6752999,0.5998474,0.51684964,0.52439487,0.5998474,0.633801,0.4376245,0.6526641,0.7205714,0.6413463,0.5055317,0.5017591,0.51684964,0.52439487,0.5885295,0.7054809,0.80356914,0.9318384,0.845068,0.90543,1.1242423,1.1619685,1.2034674,1.6071383,1.9353566,2.142851,2.5767028,2.5767028,3.029418,3.5839937,4.134797,4.8365054,4.5988297,4.4630156,4.0706625,3.410453,2.837014,2.7426984,3.2105038,3.4859054,3.3538637,3.1539145,2.7804246,2.4597516,2.1579416,1.841041,1.4864142,1.2411937,1.1996948,1.2638294,1.3128735,1.1959221,1.056335,0.98842776,0.965792,0.98465514,1.0638802,1.2487389,1.388326,1.4939595,1.6260014,1.9089483,2.2069857,2.6634734,3.048281,3.2746384,3.4142256,3.3878171,3.2935016,3.3463185,3.6594462,4.2027044,4.3309736,4.447925,4.568649,4.715781,4.8855495,5.3344917,5.8400235,6.3342376,6.7152724,6.900131,6.802043,6.48137,6.2663302,6.1720147,5.938112,6.096562,6.6247296,7.1868505,7.598067,7.8508325,7.7678347,7.375482,6.8359966,6.356873,6.187105,6.3908267,6.5643673,6.7152724,6.9189944,7.3188925,8.047009,8.348819,8.582722,9.016574,9.835234,0.5696664,0.422534,0.44894236,0.56212115,0.7696155,1.1883769,1.327964,0.9808825,0.73188925,0.6413463,0.24899325,0.21881226,0.15467763,0.094315626,0.05281675,0.026408374,0.018863125,0.03772625,0.29426476,0.663982,0.694163,0.32821837,0.26031113,0.21881226,0.1358145,0.15845025,0.12826926,0.14335975,0.12826926,0.090543,0.08677038,0.16222288,0.18485862,0.211267,0.23390275,0.17731337,0.1659955,0.13204187,0.10186087,0.09808825,0.120724,0.181086,0.331991,0.5470306,0.7809334,0.94315624,0.51684964,0.44894236,0.7809334,1.4298248,2.1994405,2.9766011,4.285702,5.50426,6.507778,7.665974,6.94163,5.7117543,5.0138187,5.2062225,5.9796104,6.1833324,6.507778,8.582722,13.106099,19.855326,26.525326,27.947605,28.019285,28.045694,26.706413,29.39252,29.83769,28.626678,27.283625,28.260735,26.90259,22.40562,17.7917,14.48688,12.325166,12.257258,11.91395,11.77059,11.751727,11.25374,8.401636,7.001992,6.439871,6.1720147,5.7419353,5.553304,5.406172,4.825187,3.893349,3.2255943,3.0709167,2.7011995,2.6823363,3.180323,3.9688015,3.8782585,3.8895764,3.731126,3.429316,3.3350005,4.7874613,5.772116,6.349328,7.3792543,10.544487,10.193633,7.77538,5.4438977,3.783943,1.81086,2.263575,4.2517486,5.3269467,4.8100967,3.7914882,2.8634224,2.142851,1.7429527,2.0108092,3.5123138,3.4066803,2.8445592,2.2748928,1.8146327,1.267602,1.5015048,1.901403,2.0975795,2.0673985,2.1390784,2.0258996,2.8256962,3.4029078,3.8556228,5.5268955,5.247721,6.1720147,9.099571,12.943876,14.728328,14.049255,12.045992,9.163706,6.519096,5.8928404,8.07719,8.714764,8.75249,8.899622,9.601331,8.952439,7.3188925,5.5306683,4.432834,4.881777,9.386291,13.483362,16.576914,18.881989,21.420965,19.31584,14.698147,13.102326,15.411173,17.867151,18.75372,20.647577,21.737865,21.575642,21.092747,17.723793,15.143317,16.094019,18.814081,17.01831,16.146835,20.964478,23.544952,22.409393,22.526344,26.049976,25.578398,23.258234,20.345766,17.20317,14.049255,14.554788,15.113135,14.324657,12.996693,16.648594,21.217243,24.70692,26.63096,28.004196,28.158873,25.238861,20.685303,16.029884,12.864652,15.62244,18.542452,20.277859,20.938068,22.100037,22.590479,25.016277,27.970242,29.898052,29.10203,24.476791,20.511763,18.463226,18.7839,21.11161,29.788647,31.044931,31.59196,37.499893,54.2013,49.285572,32.49739,17.45971,9.49947,5.6363015,5.081726,4.5761943,4.447925,4.8930945,5.9796104,7.7829256,15.554533,23.65813,29.113348,31.614597,37.356533,27.800474,16.214743,8.914713,5.251494,5.994701,5.2099953,5.2288585,6.0248823,5.2137675,5.643847,6.771862,6.6322746,5.270357,4.7006907,4.285702,3.8593953,3.199186,2.3126192,1.4449154,0.9242931,0.8337501,0.94692886,1.4109617,2.7502437,1.5769572,0.9808825,1.2223305,2.2258487,3.591539,5.1345425,8.480861,15.920478,22.737612,17.222033,14.679284,12.789199,10.178542,7.0284004,5.070408,4.666737,4.7421894,7.0057645,9.703192,7.594294,10.186088,11.400873,12.54775,13.95494,14.992412,15.23386,14.015302,12.913695,12.355347,11.5857315,9.665465,11.000975,10.816116,8.537451,7.816879,12.359119,10.967021,8.563859,7.907422,9.578695,9.239159,11.332966,11.559323,9.590013,9.058073,8.137552,7.696155,9.922004,12.770335,9.963503,10.846297,13.015556,16.11288,19.866644,24.107073,21.802,18.746174,18.387774,20.975796,23.548725,34.225254,43.106014,41.57433,31.339195,24.431519,22.72252,15.912932,8.827943,4.315883,3.2331395,3.6971724,6.8473144,10.680302,11.92904,6.058836,3.5764484,2.1994405,1.720317,1.841041,2.1654868,6.0776987,7.5037513,9.291975,10.902886,8.439363,10.072908,14.260523,16.316603,14.962231,12.325166,11.087745,10.091772,8.443134,6.696409,6.85486,4.9647746,5.028909,6.488915,8.069645,7.7602897,7.805561,6.2323766,5.191132,5.100589,4.644101,3.5839937,3.187868,3.7914882,5.4288073,7.8621507,5.4665337,6.221059,8.677037,11.174516,11.84227,9.06939,6.307829,4.5799665,4.395108,5.7683434,6.0512905,5.458988,4.851596,4.8327327,5.723072,6.590776,5.983383,5.715527,6.3531003,7.220804,8.571404,7.5188417,6.6020937,6.8133607,7.5905213,6.8774953,7.8961043,9.718282,10.170997,5.824933,8.461998,9.322156,12.713746,17.440845,16.810818,9.725827,7.284939,7.7187905,8.654402,7.1038527,5.2250857,5.081726,5.59103,6.5341864,8.552541,7.6093845,6.56814,6.1078796,6.4926877,7.541477,9.703192,9.21275,8.812852,9.408927,10.091772,8.865668,9.593785,10.155907,10.038955,10.355856,9.820143,11.000975,12.494934,13.034419,11.480098,10.27663,9.544742,9.514561,9.137298,6.092789,4.447925,4.768598,4.7648253,3.8480775,3.1614597,2.969056,2.9615107,3.3651814,4.093298,4.749735,3.610402,3.3463185,3.0558262,2.5427492,2.3163917,2.2560298,1.9504471,1.6750455,1.5015048,1.3015556,0.8111144,0.68661773,0.65643674,0.65643674,0.845068,0.8262049,0.845068,0.9695646,1.2034674,1.478869,1.4562333,1.146878,0.9016574,0.845068,0.9016574,0.62625575,0.3961256,0.2565385,0.24522063,0.3734899,0.5696664,0.47157812,0.5281675,0.72811663,0.59607476,0.7469798,1.0525624,1.1016065,1.026154,1.5128226,1.6146835,1.6863633,1.9768555,2.1843498,1.4637785,2.071171,2.8709676,3.410453,3.9574835,5.5193505,4.561104,8.7600355,7.4735703,0.8941121,0.041498873,0.4979865,2.3201644,2.5578396,1.327964,1.8221779,2.704972,2.3880715,2.0975795,2.0372176,1.358145,1.629774,1.9089483,2.1013522,2.1277604,1.9089483,1.7693611,2.0183544,2.463524,2.8332415,2.746471,2.7351532,2.9237845,2.746471,2.1881225,1.7919968,1.2411937,1.0035182,0.935611,0.90920264,0.8186596,0.67152727,0.66775465,0.68661773,0.68661773,0.694163,0.70170826,0.66020936,0.6488915,0.69039035,0.7394345,0.8639311,0.9205205,0.9695646,1.0374719,1.116697,0.9922004,0.91297525,0.9318384,1.0336993,1.1242423,1.1393328,1.2110126,1.1808317,1.1431054,1.4335974,1.3053282,1.1280149,1.0374719,0.9393836,0.52062225,0.32444575,0.2678564,0.25276586,0.241448,0.23390275,0.2678564,0.33576363,0.44139713,0.5319401,0.52439487,0.62625575,0.77716076,0.9205205,0.97710985,0.83752275,0.7809334,0.6451189,0.5998474,0.70170826,0.8903395,0.76207024,0.7696155,0.784706,0.72811663,0.58098423,0.5357128,0.513077,0.5470306,0.58098423,0.4376245,0.5470306,0.543258,0.47912338,0.43007925,0.4979865,0.6111652,0.5772116,0.6375736,0.814887,0.935611,1.1431054,1.0412445,1.0336993,1.1883769,1.2449663,1.3241913,1.659955,2.0975795,2.4371157,2.4522061,2.214531,2.848332,3.5764484,4.1574326,4.8968673,4.696918,4.432834,4.183841,3.9008942,3.3953626,3.097325,3.1916409,3.308592,3.2482302,3.0218725,2.4295704,2.11267,1.7995421,1.4260522,1.1544232,1.1544232,1.1544232,1.2261031,1.3204187,1.267602,1.1431054,1.0525624,0.98465514,0.9997456,1.2411937,1.1204696,1.2298758,1.3920987,1.5845025,1.9466745,2.1654868,2.5276587,2.916239,3.2331395,3.3953626,3.2859564,3.1614597,3.1576872,3.3651814,3.8254418,4.266839,4.5535583,4.617693,4.564876,4.689373,5.1232247,5.7494807,6.1908774,6.356873,6.436098,6.247467,6.0324273,5.8966126,5.832478,5.73439,5.938112,6.2889657,6.6586833,6.9982195,7.33021,7.281166,7.141579,6.832224,6.4134626,6.0776987,5.9796104,6.2889657,6.458734,6.5002327,6.990674,7.5792036,7.8998766,7.964011,7.911195,8.013056,0.28294688,0.23390275,0.241448,0.34330887,0.6149379,1.1506506,1.3053282,0.995973,0.7922512,0.7582976,0.4074435,0.39989826,0.35839936,0.24522063,0.094315626,0.041498873,0.041498873,0.05281675,0.3734899,0.9205205,1.2223305,0.55457586,0.46026024,0.47535074,0.38480774,0.23013012,0.14713238,0.13958712,0.120724,0.08299775,0.120724,0.16222288,0.124496624,0.10186087,0.124496624,0.12826926,0.124496624,0.08299775,0.056589376,0.071679875,0.13204187,0.24522063,0.3961256,0.543258,0.6073926,0.47912338,0.33576363,0.5055317,0.97710985,1.539231,1.7844516,2.142851,2.837014,3.7386713,4.689373,5.50426,4.8930945,3.7763977,3.1161883,3.259548,3.953711,5.0854983,7.7414265,9.714509,11.299012,15.294222,21.571869,24.254206,24.646559,24.042938,23.722265,27.732567,30.181,30.388494,29.369886,29.826374,29.882963,24.899324,18.4255,12.83447,9.318384,10.035183,10.578441,11.133017,11.925267,13.219278,9.861642,7.424526,6.620957,6.9680386,6.7869525,6.1833324,6.119198,5.7192993,4.825187,3.9876647,4.285702,3.904667,3.8858037,4.6290107,5.8664317,5.0439997,4.3121104,3.9197574,3.8971217,4.063117,4.9647746,5.587258,6.5643673,8.179051,10.38981,9.020347,6.360646,4.4403796,3.4368613,1.6637276,1.8938577,4.496969,5.9909286,5.455216,4.515832,3.5877664,2.3654358,1.8070874,2.2447119,3.3840446,4.2894745,3.682082,2.6182017,1.7882242,1.539231,1.2411937,1.6222287,1.9806281,1.9655377,1.5845025,2.1768045,3.4481792,4.938366,7.1076255,11.32542,13.373956,16.867407,20.025093,20.741892,16.58446,13.849306,11.593277,9.0807085,6.9152217,7.0472636,8.66572,9.450426,8.552541,7.3905725,9.639057,8.805306,6.79827,5.081726,4.6818275,6.1720147,10.718028,13.9888935,15.377219,15.845025,17.886015,15.01882,11.721546,10.767072,12.332711,13.992666,14.264296,14.966003,16.120426,17.320122,17.727566,15.671484,14.034165,14.784918,16.463736,14.2077055,13.555041,17.927513,21.58696,22.620659,22.967741,26.506464,26.09902,23.41291,19.817598,16.392056,17.320122,19.293203,19.372429,16.950403,13.736128,16.305285,19.123436,21.371922,22.97906,24.631468,24.861599,23.08092,18.931032,14.120935,12.419481,15.660167,18.923487,19.934551,19.364883,20.85507,22.296213,22.65084,22.616886,22.367893,21.583187,18.395319,15.731846,14.369928,14.969776,18.070873,24.352295,25.027594,27.015768,34.270527,47.776524,44.373615,29.094484,15.384765,8.624221,6.1116524,5.6400743,5.3344917,5.27413,6.006019,8.537451,11.287694,18.957441,26.14429,33.399048,47.24081,48.629135,32.674706,17.206944,9.408927,5.7909794,4.447925,3.8141239,4.315883,5.304311,5.0553174,5.492942,6.7454534,7.220804,6.462507,5.1760416,5.0251365,4.496969,3.7877154,3.006782,2.1994405,1.6788181,1.6410918,1.6976813,1.6863633,1.6863633,7.54525,7.33021,4.8327327,2.8521044,3.2331395,5.0175915,7.364164,15.614895,25.861345,24.94837,21.319103,18.516043,14.988639,10.925522,8.262049,7.032173,6.326692,7.6320205,9.703192,8.567632,10.521852,12.034674,13.573905,14.939595,15.279131,13.377728,13.290957,13.087236,12.061082,10.714255,8.379,10.38981,10.578441,8.175279,7.786698,13.52486,11.155652,8.111144,8.326183,12.253486,9.80128,11.2801485,12.792972,12.362892,9.955957,7.7225633,6.2399216,8.899622,12.668475,8.114917,13.35132,14.864142,16.03743,18.033148,19.779873,17.40689,14.830189,14.867915,17.652113,20.658894,25.902843,35.217453,36.711414,28.35505,18.018057,16.007248,12.264804,7.7225633,3.832987,2.5578396,3.7235808,5.7909794,7.635793,7.6207023,3.6028569,1.7542707,1.7429527,1.9579924,1.8448136,1.9051756,4.104616,7.635793,10.680302,10.925522,5.564622,6.851087,8.75249,9.81637,9.337247,7.3453007,7.805561,7.5716586,6.277648,4.8855495,5.6589375,3.640583,4.08198,5.1873593,5.7306175,5.0553174,6.7152724,6.722818,6.273875,5.802297,4.9685473,3.187868,2.9426475,4.1272516,5.987156,7.0849895,7.4735703,7.492433,8.201687,10.03141,12.770335,11.529142,8.66572,6.9152217,7.0812173,8.031919,7.333983,5.9984736,5.0213637,4.878004,5.5382137,6.8133607,6.9567204,6.1041074,5.100589,5.492942,7.145352,6.398372,6.119198,7.01331,7.5905213,6.6850915,7.111398,8.639311,9.639057,7.0887623,6.809588,7.2698483,10.352083,14.136025,12.909923,10.087999,11.185833,12.427027,11.521597,7.654656,5.5683947,5.643847,6.1003346,6.7643166,9.088254,8.967529,7.5829763,7.360391,8.439363,8.66572,9.461743,8.707218,8.688355,9.669238,9.914458,9.25425,9.952185,10.725573,10.740664,9.639057,10.03141,11.268831,12.1252165,11.846043,10.163452,9.2844305,8.526133,8.390318,7.997965,5.0553174,4.112161,4.768598,4.859141,3.893349,3.059599,3.3274553,2.9237845,3.059599,3.802806,4.074435,2.9011486,2.7125173,2.6521554,2.3277097,1.8297231,1.9127209,1.8146327,1.6373192,1.5052774,1.5882751,1.0525624,0.875249,0.69793564,0.513077,0.65643674,0.6526641,0.58475685,0.6413463,0.8601585,1.1544232,1.2826926,1.0940613,0.88279426,0.8262049,0.965792,0.77338815,0.49044126,0.29803738,0.24522063,0.23013012,0.46026024,0.38103512,0.3734899,0.4979865,0.5281675,0.5281675,0.77716076,0.9318384,1.0336993,1.5241405,1.81086,1.6524098,1.9994912,2.6219745,2.093807,2.1503963,2.7125173,2.9652832,3.218049,4.9157305,3.5387223,5.832478,5.323174,1.5467763,0.049044125,0.090543,1.327964,1.9881734,1.629774,1.1732863,2.4408884,2.0636258,1.7429527,1.8372684,1.3656902,1.358145,1.7127718,1.9278114,1.8523588,1.6939086,1.4637785,1.5165952,1.8297231,2.2069857,2.263575,2.0862615,2.2786655,2.354118,2.0975795,1.5656394,1.056335,0.9016574,0.8601585,0.8224323,0.8186596,0.7054809,0.6488915,0.62248313,0.6073926,0.6073926,0.62248313,0.66020936,0.70170826,0.73188925,0.7394345,0.8563859,0.9620194,1.0035182,0.98842776,0.995973,0.935611,0.935611,1.0751982,1.267602,1.3015556,1.1657411,1.1883769,1.1959221,1.1959221,1.3807807,1.2789198,1.0450171,0.8111144,0.5998474,0.27917424,0.1961765,0.16976812,0.18485862,0.211267,0.22258487,0.35085413,0.42630664,0.49044126,0.5583485,0.6111652,0.73566186,0.8186596,0.91674787,0.9997456,0.9507015,1.0035182,0.9242931,0.8111144,0.784706,0.98842776,0.8337501,0.784706,0.77338815,0.73188925,0.58475685,0.59230214,0.56212115,0.5394854,0.51684964,0.44139713,0.49044126,0.49044126,0.47912338,0.4678055,0.47912338,0.6828451,0.7167987,0.7130261,0.754525,0.84129536,1.026154,1.0902886,1.1506506,1.2298758,1.2826926,1.5882751,1.7844516,2.033445,2.3163917,2.4559789,2.2107582,2.6823363,3.2859564,3.874486,4.7233267,4.644101,4.3347464,4.0970707,3.9650288,3.7047176,3.6028569,3.7009451,3.6443558,3.3350005,2.916239,2.0900342,1.7354075,1.4449154,1.1242423,0.995973,1.0714256,1.0978339,1.146878,1.20724,1.1921495,1.1544232,1.0450171,0.9280658,0.8978847,1.0789708,0.98842776,1.1242423,1.327964,1.5618668,1.9164935,2.0749438,2.3654358,2.71629,3.0181,3.127506,2.957738,2.8898308,2.969056,3.2369123,3.731126,4.2404304,4.5007415,4.5120597,4.436607,4.5837393,5.0439997,5.564622,5.8437963,5.885295,6.0211096,5.9230213,5.715527,5.5382137,5.4703064,5.5080323,5.723072,5.9532022,6.255012,6.549277,6.617184,6.40969,6.477597,6.48137,6.2399216,5.726845,5.6363015,6.0022464,6.2021956,6.258785,6.858632,7.0849895,7.3792543,7.454707,7.2396674,6.8774953,0.1358145,0.124496624,0.116951376,0.181086,0.38480774,0.784706,0.95447415,0.8186596,0.6526641,0.573439,0.55080324,0.56212115,0.5281675,0.362172,0.150905,0.13958712,0.14335975,0.15467763,0.49044126,1.1581959,1.8561316,0.935611,0.754525,0.77338815,0.6752999,0.35839936,0.28294688,0.24522063,0.18485862,0.120724,0.15845025,0.14335975,0.12826926,0.11317875,0.10186087,0.10940613,0.090543,0.0754525,0.10186087,0.17354076,0.27917424,0.36971724,0.4640329,0.52062225,0.49421388,0.32821837,0.3961256,0.73188925,1.2185578,1.5203679,1.1016065,1.0412445,1.2261031,1.5580941,1.9278114,2.1994405,2.4597516,1.9429018,1.5052774,1.5467763,2.0372176,2.9992368,7.677292,10.321902,9.937095,10.303039,14.060574,16.675003,17.863379,17.91997,17.701157,19.636513,22.239624,23.544952,23.72981,25.140774,25.717985,23.616632,19.18757,13.52486,8.424272,8.126234,8.307321,8.639311,9.442881,11.68382,9.793735,7.647111,6.8963585,7.352846,6.971811,5.587258,5.2137675,5.093044,4.908185,4.7950063,5.270357,5.4212623,5.8437963,6.752999,7.9791017,6.4549613,5.093044,4.8402777,5.6891184,6.6850915,6.3229194,5.7381625,5.7419353,6.326692,6.673774,7.066127,6.387054,5.1081343,3.519859,1.7429527,1.2336484,3.4029078,5.0854983,5.0968165,4.247976,4.1272516,3.0218725,2.7087448,3.712263,5.2779026,7.2623034,5.8513412,3.8367596,2.7351532,2.7615614,2.022127,2.0145817,2.2598023,2.41448,2.2711203,3.8820312,5.2590394,7.541477,11.7026825,18.55377,22.85079,26.51778,26.423466,21.420965,12.332711,9.435335,8.439363,7.8961043,7.2623034,6.907676,7.0510364,8.484633,8.065872,6.9869013,10.774617,9.7220545,7.4584794,5.7192993,5.4778514,6.952948,9.118435,11.378237,11.664956,10.812344,12.559069,11.099063,9.906913,10.159679,11.506506,12.049765,10.899114,10.589758,12.679792,16.078928,17.04472,16.4826,15.365902,14.603831,13.890805,11.732863,13.494679,16.188334,19.15739,21.304014,21.088974,26.15561,26.86109,23.54118,18.704676,17.025856,20.296722,22.232079,22.028357,19.934551,17.267305,16.490145,17.520071,19.119663,20.225042,19.972277,20.074137,20.104319,17.689838,13.70972,12.276122,15.00373,18.48209,19.01403,17.293713,18.376457,20.225042,19.693102,18.49718,17.380484,16.11288,14.388792,13.098554,11.634775,11.219787,14.905642,18.406637,18.62545,22.205671,31.12793,42.728752,39.144756,25.299223,13.030646,7.2283497,5.8211603,6.1116524,5.764571,5.723072,7.394345,12.642066,15.69412,21.851044,28.788902,40.51045,67.31495,60.34691,38.212917,19.274342,10.284176,6.3719635,3.4029078,2.463524,2.916239,4.08198,5.270357,5.915476,7.1076255,7.9036493,7.6093845,5.7570257,6.089017,5.4665337,4.6818275,4.002755,3.1727777,2.6332922,2.8332415,3.2331395,3.5387223,3.6971724,15.188588,14.479335,9.042982,4.3686996,3.9574835,5.6363015,7.6395655,13.95494,22.737612,26.325377,24.503199,21.405874,17.512526,13.702174,11.227332,9.0543,7.250985,8.27714,11.151879,11.446144,13.36641,13.196642,13.932304,16.452417,19.56106,14.275613,14.554788,15.724301,15.286676,12.894833,9.378746,8.692128,8.228095,7.435844,7.7829256,14.053028,11.740409,8.612903,8.75249,12.540206,9.016574,9.797507,12.234623,13.13628,8.771353,6.832224,6.33801,9.593785,13.679539,10.423763,16.373192,15.086727,13.909668,14.569878,13.185325,11.962994,11.363147,12.166716,15.041456,20.534397,20.1345,24.20139,27.53639,25.699121,15.026365,10.823661,8.495952,5.836251,3.1124156,3.029418,4.244203,4.187614,3.1840954,1.7542707,0.6073926,0.68661773,1.7693611,2.2786655,1.9391292,1.7844516,3.6443558,8.601585,10.446399,7.816879,4.1762958,3.6594462,3.4972234,3.3878171,3.1765501,2.8596497,3.983892,3.9763467,3.0633714,2.071171,2.425798,2.9464202,3.6481283,4.1574326,4.2592936,3.874486,5.9532022,7.4811153,7.99042,7.4094353,6.0550632,3.4557245,2.9992368,4.2894745,6.1531515,6.609639,10.868933,10.159679,8.627994,9.027891,12.736382,12.411936,9.808825,8.688355,9.639057,10.072908,9.125979,7.3868,6.307829,6.3455553,6.9567204,8.748717,9.450426,7.6923823,4.817642,4.878004,5.383536,4.6742826,5.160951,7.0246277,8.186596,7.5905213,7.0510364,7.0359454,7.7187905,9.001483,7.0963078,6.7152724,7.696155,9.405154,10.763299,13.751218,17.629477,17.308804,12.362892,7.0359454,6.2851934,6.72659,7.4169807,7.805561,7.752744,10.38981,8.858124,8.771353,10.702937,10.212496,9.261794,9.144843,9.144843,9.050528,9.137298,9.993684,10.47658,11.057564,11.102836,8.850578,9.9257765,10.955703,10.544487,9.073163,8.68081,7.564113,7.0057645,6.6247296,5.9003854,4.1574326,4.0593443,4.9987283,5.5306683,5.0025005,3.5764484,4.6818275,3.62172,2.8143783,2.927557,2.8898308,2.0183544,2.0749438,2.4069347,2.4522061,1.7316349,1.9768555,1.8900851,1.6524098,1.5165952,1.7655885,1.4071891,1.177059,0.8224323,0.46026024,0.5696664,0.5998474,0.40367088,0.34330887,0.5281675,0.7922512,1.0601076,1.0789708,0.8978847,0.7167987,0.9016574,0.8262049,0.5696664,0.40367088,0.331991,0.116951376,0.2565385,0.26031113,0.25276586,0.30181,0.4376245,0.30181,0.44516975,0.7054809,1.0148361,1.3958713,1.6146835,1.5920477,2.022127,2.727608,2.6521554,2.0598533,2.686109,3.1727777,3.4444065,4.708236,4.478106,3.9310753,3.3915899,2.4974778,0.18485862,0.08677038,0.69793564,1.6109109,2.0183544,0.694163,1.3505998,1.2864652,1.2751472,1.4411428,1.2525115,1.0751982,1.3694628,1.6071383,1.6222287,1.6033657,1.4750963,1.4109617,1.4034165,1.5241405,1.9240388,1.901403,1.7542707,1.7655885,1.8221779,1.3996439,1.086516,1.0336993,0.98465514,0.8978847,0.9242931,0.79602385,0.7054809,0.62625575,0.58098423,0.6149379,0.6149379,0.69039035,0.77338815,0.83752275,0.87147635,0.7997965,0.87902164,0.95824677,0.98465514,0.995973,1.0412445,1.1053791,1.20724,1.3053282,1.3091009,1.1732863,1.1355602,1.237421,1.3619176,1.2147852,1.0186088,0.87147635,0.68661773,0.44516975,0.18485862,0.1659955,0.14713238,0.15467763,0.19240387,0.23390275,0.44894236,0.49044126,0.51684964,0.60362,0.72811663,0.8526133,0.7997965,0.8262049,0.97333723,1.086516,1.1996948,1.237421,1.0789708,0.845068,0.9016574,0.8563859,0.784706,0.7394345,0.7054809,0.6149379,0.6149379,0.5998474,0.5394854,0.4640329,0.46026024,0.48666862,0.56589377,0.6111652,0.5885295,0.5017591,0.7092535,0.79602385,0.7054809,0.55080324,0.60362,0.77338815,1.0638802,1.267602,1.3091009,1.267602,1.7618159,1.9353566,1.9164935,2.033445,2.8143783,2.6219745,2.5502944,2.7615614,3.3538637,4.353609,4.3385186,4.1272516,3.863168,3.6707642,3.6179473,4.006528,4.5120597,4.3196554,3.429316,2.6597006,1.81086,1.3770081,1.1732863,1.1016065,1.1280149,1.0978339,1.056335,1.0299267,1.0223814,1.0072908,1.0450171,0.94315624,0.83752275,0.784706,0.7507524,0.98842776,1.1619685,1.3204187,1.5165952,1.7957695,1.9806281,2.2786655,2.5616124,2.7389257,2.7615614,2.5804756,2.5616124,2.7238352,3.1048703,3.7386713,4.115934,4.2291126,4.2517486,4.3083377,4.4818783,4.949684,5.2137675,5.3382645,5.4288073,5.613666,5.80607,5.560849,5.251494,5.100589,5.168496,5.3609,5.613666,5.983383,6.2323766,5.8098426,5.4967146,5.6061206,5.783434,5.7494807,5.2779026,5.3910813,5.6400743,5.828706,6.0626082,6.722818,6.477597,6.590776,6.752999,6.7341356,6.405917,0.1358145,0.11317875,0.124496624,0.120724,0.11317875,0.19994913,0.35839936,0.4979865,0.5696664,0.55080324,0.42630664,0.2565385,0.1961765,0.1961765,0.2867195,0.58098423,0.49421388,0.5017591,0.6149379,0.98842776,1.8938577,1.1959221,0.97710985,0.7884786,0.51684964,0.38103512,0.68661773,0.7167987,0.5583485,0.3772625,0.42630664,0.35462674,0.23390275,0.181086,0.1961765,0.18485862,0.1358145,0.150905,0.24899325,0.39989826,0.5357128,0.46026024,0.422534,0.41121614,0.41121614,0.41121614,0.5583485,1.1355602,1.3920987,1.1016065,0.56589377,0.5017591,0.6451189,0.80356914,0.90543,0.9922004,1.750498,1.5618668,1.2940104,1.7580433,3.7235808,2.4672968,3.3689542,6.3832817,10.352083,13.000465,14.66042,15.935568,16.192106,15.184815,13.060828,14.196388,17.501207,21.45869,25.140774,28.22678,20.1345,15.62244,13.3626375,11.721546,8.744945,6.0701537,5.485397,6.168242,7.0812173,6.9567204,8.167733,7.5263867,7.1000805,7.3000293,6.8963585,5.59103,6.0512905,6.247467,5.7570257,5.783434,5.915476,5.6287565,5.8928404,6.6586833,6.8661776,5.80607,4.8440504,4.8138695,5.881522,7.5527954,7.8319697,6.466279,5.2326307,4.8930945,5.172269,7.7225633,8.390318,7.115171,4.8063245,3.3425457,1.8636768,2.9237845,3.4481792,3.1010978,4.2706113,7.043491,6.9680386,6.779407,8.107371,11.487643,13.856852,9.258021,5.492942,4.9723196,4.715781,4.2404304,3.8254418,3.8820312,4.6516466,6.224831,9.009028,6.043745,5.3948536,9.937095,17.335213,17.712475,14.037937,9.567377,6.304056,4.961002,7.118943,7.7338815,7.9225125,8.088508,7.91874,6.8925858,5.704209,5.9720654,7.164215,6.5756855,6.930312,6.5341864,6.9680386,8.710991,11.136789,12.310076,14.268067,16.11288,16.392056,13.106099,12.936331,10.585986,9.835234,11.133017,11.59705,10.876478,10.295494,12.691111,16.459963,15.516807,15.24895,15.977067,15.626213,13.6833105,11.231105,15.16218,16.105335,17.670975,20.013775,19.866644,26.751684,27.200626,25.276588,22.714975,18.904623,20.323132,21.73032,22.209444,21.454918,19.74592,16.984358,19.270569,22.322622,23.084692,19.715738,17.84829,16.739138,14.7736,12.128989,10.789707,13.045737,14.909414,15.580941,15.558306,16.633503,16.731592,15.565851,14.056801,12.928786,12.694883,10.231359,9.156161,8.722309,9.352338,12.6345215,14.381247,14.313339,17.108854,24.623924,35.90407,30.629942,21.171972,11.668729,5.198677,3.783943,5.481624,5.7419353,5.9230213,7.9791017,14.449154,17.014538,25.499172,36.858547,53.473186,83.15997,61.897457,39.533337,21.87368,11.242422,6.470052,4.1762958,3.059599,2.8181508,3.4255435,5.172269,6.258785,7.1264887,7.5527954,7.598067,7.598067,8.575176,7.9413757,6.560595,5.100589,4.0291634,3.2331395,3.8971217,4.7950063,5.2590394,5.172269,3.8443048,4.1310244,6.56814,9.842778,10.816116,11.5857315,10.982111,11.332966,13.336229,16.0827,18.451908,16.927769,14.094527,11.653639,10.419991,8.933576,7.4999785,8.262049,10.763299,11.947904,17.73511,13.045737,8.944894,12.713746,27.860836,17.30503,16.13929,21.979313,28.336185,24.627695,18.523588,12.777881,8.98262,7.4773426,7.356619,7.564113,8.612903,8.869441,8.314865,8.560086,6.670001,9.884277,11.910177,10.834979,9.125979,6.609639,11.785681,16.648594,17.73511,16.11288,15.101818,14.818871,12.340257,11.11038,20.949387,14.68683,7.9413757,5.1269975,6.7869525,9.582467,8.571404,13.2607765,19.406384,21.741638,13.977575,9.57115,8.039464,5.541986,2.4823873,3.4934506,3.3123648,1.9391292,0.8337501,0.48666862,0.41121614,0.6187105,1.8070874,2.7087448,2.7728794,2.1503963,3.8858037,5.96452,6.1418333,4.349837,2.7011995,2.6031113,2.4031622,2.7087448,3.0558262,1.9089483,1.6750455,1.599593,1.3053282,0.8262049,0.59607476,1.5354583,1.9164935,2.033445,1.9429018,1.478869,2.2598023,3.108643,4.195159,5.6778007,7.6886096,4.0782075,2.5880208,3.0709167,4.949684,7.232122,9.918231,11.027383,11.566868,12.064855,12.58925,11.170743,7.8998766,6.0550632,6.375736,7.0359454,7.964011,7.707473,7.635793,7.9451485,7.673519,9.031664,8.763808,7.322665,5.5382137,4.6252384,4.7572803,3.9310753,4.4441524,6.307829,7.2472124,7.1378064,7.5490227,7.515069,7.413208,8.986393,8.937348,7.435844,6.0550632,7.3453007,14.815099,21.994404,24.07312,18.674494,9.34102,5.5080323,7.0849895,7.8432875,8.722309,9.144843,7.0359454,8.729855,8.431817,8.16396,9.027891,11.200924,12.566614,11.627231,9.703192,8.186596,8.514814,9.088254,10.386037,10.853842,9.986138,8.299775,7.9715567,9.408927,10.612394,11.133017,12.083718,8.458225,5.9682927,5.2175403,5.342037,3.9989824,4.98741,7.0472636,8.07719,7.4094353,5.798525,7.213259,5.372218,3.169005,2.1202152,2.3654358,1.7655885,1.7354075,2.1088974,2.5125682,2.3654358,3.059599,2.5578396,1.9240388,1.780679,2.305074,2.1088974,1.4750963,0.77716076,0.33953625,0.41121614,0.6073926,0.4376245,0.36971724,0.48666862,0.47157812,0.7432071,1.0940613,1.0374719,0.694163,0.7922512,0.7582976,0.58475685,0.5470306,0.56589377,0.21503963,0.23767537,0.271629,0.24899325,0.20372175,0.29049212,0.20372175,0.2565385,0.58098423,0.9695646,0.8865669,1.3845534,1.5580941,2.052308,2.674791,2.3956168,2.2258487,2.6031113,3.1765501,3.7198083,4.134797,7.7716074,6.477597,4.979865,4.0782075,0.6111652,0.21881226,0.18485862,1.5882751,2.987919,0.41121614,0.58475685,0.76207024,0.8299775,0.8639311,1.1431054,0.8865669,1.0450171,1.2336484,1.3619176,1.6184561,1.2147852,1.0299267,0.91674787,0.90920264,1.2525115,1.5430037,1.6637276,1.6222287,1.50905,1.50905,1.2185578,1.0072908,0.86770374,0.80356914,0.83752275,0.7432071,0.62625575,0.55080324,0.543258,0.58098423,0.58098423,0.543258,0.55457586,0.6488915,0.80734175,0.7582976,0.6752999,0.65643674,0.77338815,1.0676528,1.3958713,1.4524606,1.3166461,1.2110126,1.478869,1.5882751,1.3694628,1.4449154,1.690136,1.2525115,0.76207024,0.6488915,0.6073926,0.452715,0.120724,0.1358145,0.1358145,0.150905,0.19994913,0.32067314,0.4678055,0.58475685,0.7696155,0.935611,0.83752275,0.875249,0.86770374,0.8903395,0.965792,1.0374719,0.86770374,0.91674787,0.9280658,0.8526133,0.8526133,0.7696155,0.7394345,0.72811663,0.7092535,0.68661773,0.49044126,0.4074435,0.4074435,0.46026024,0.5357128,0.422534,0.46026024,0.4979865,0.5357128,0.73188925,0.7582976,0.633801,0.52439487,0.55457586,0.8224323,1.2261031,1.3355093,1.3166461,1.2298758,1.0223814,1.3996439,1.7429527,1.991946,2.2899833,2.9615107,2.4823873,2.0372176,2.1692593,2.8898308,3.6481283,3.8669407,3.893349,3.832987,3.731126,3.5689032,4.3385186,4.67051,4.063117,2.7238352,1.5241405,1.3656902,1.2185578,1.2110126,1.3619176,1.5580941,1.5920477,1.2826926,1.0299267,0.95824677,0.8865669,0.8865669,0.9507015,1.0336993,1.1053791,1.1280149,1.1431054,1.2449663,1.3845534,1.5769572,1.9089483,2.04099,2.1956677,2.41448,2.5804756,2.3956168,2.372981,2.4823873,2.6974268,3.029418,3.5538127,3.983892,4.134797,4.172523,4.191386,4.22534,4.606375,4.919503,5.2364035,5.4212623,5.1269975,5.2967653,5.2288585,4.938366,4.6290107,4.715781,4.8629136,5.1345425,5.5457587,5.847569,5.553304,5.455216,5.413717,5.4250345,5.458988,5.4476705,5.3382645,5.311856,5.3344917,5.564622,6.3342376,6.126743,6.119198,6.3153744,6.428553,5.904158,0.10186087,0.094315626,0.11317875,0.11317875,0.10186087,0.1358145,0.19994913,0.15467763,0.211267,0.392353,0.513077,0.5357128,0.51684964,0.58475685,0.69793564,0.6413463,0.38858038,0.33953625,0.5319401,0.84129536,0.965792,0.91297525,0.8978847,0.9242931,0.94692886,0.88279426,1.1280149,1.026154,0.9016574,0.87147635,0.84129536,0.66020936,0.60362,0.5696664,0.49421388,0.35462674,0.2867195,0.29426476,0.32444575,0.38858038,0.58475685,0.52062225,0.69039035,0.7432071,0.6451189,0.7054809,1.0940613,1.1996948,1.0299267,0.6790725,0.30935526,0.24899325,0.32067314,0.422534,0.5055317,0.5998474,1.2411937,1.5467763,1.5656394,1.8146327,3.2821836,4.214022,4.214022,5.036454,7.0472636,9.216523,11.140562,10.469034,10.061591,11.276376,13.977575,15.777118,19.700647,25.027594,29.66415,30.143274,22.628204,17.652113,15.165953,13.93985,11.52537,11.996947,12.585477,12.755245,11.536687,7.5075235,5.406172,5.692891,6.4474163,6.7756343,6.8246784,6.85486,6.9567204,7.01331,6.8774953,6.3455553,6.752999,7.405663,8.009283,8.179051,7.4396167,7.1000805,6.760544,6.085244,5.4665337,6.013564,7.0472636,7.1000805,6.964266,6.5455046,4.8553686,6.119198,6.138061,5.010046,3.5236318,3.169005,3.2444575,4.055572,4.6026025,4.851596,5.7494807,7.281166,7.4282985,8.00551,11.0613365,18.885761,17.142809,11.868678,8.145098,7.643338,8.60913,6.7643166,5.6891184,5.149633,5.2326307,6.349328,8.175279,6.2927384,5.2967653,6.590776,8.424272,5.824933,5.7796617,6.4549613,6.94163,7.277394,7.4169807,6.515323,6.4738245,7.2472124,6.820906,8.703445,10.008774,8.835487,5.6325293,3.1727777,4.3649273,6.930312,9.850324,12.219532,13.264549,12.909923,11.98563,11.419736,11.272603,10.714255,11.951676,12.442118,12.0724,11.268831,10.997202,11.7026825,13.396591,15.588487,17.357847,17.323895,18.587723,17.77661,15.950659,13.65313,10.876478,14.1058445,16.135517,17.663431,19.391293,22.028357,25.650078,26.449873,27.411894,28.02683,24.276842,20.391039,16.758,15.8676605,16.98813,16.16947,14.075664,16.810818,20.315586,21.749184,19.481836,16.754227,13.558814,11.16697,10.472807,11.970539,13.59654,12.974057,12.377983,12.536433,12.615658,13.094781,11.7894535,10.31813,9.405154,8.899622,7.3415284,6.1795597,5.692891,6.5832305,9.97482,11.446144,12.81938,16.120426,22.171717,30.56958,27.63825,19.568605,11.299012,5.73439,3.7235808,4.38379,4.678055,5.481624,7.8508325,13.023102,14.822643,22.183035,34.760967,52.420624,75.21482,56.13666,36.232292,21.918951,14.260523,8.971302,6.579458,4.285702,3.3312278,3.9725742,5.455216,6.4436436,7.1981683,7.5829763,7.756517,8.14887,9.2995205,9.382519,8.718536,7.424526,5.43258,4.187614,4.715781,5.492942,5.873977,6.1003346,6.488915,8.495952,10.740664,12.189351,12.162943,8.322411,7.7602897,8.126234,8.778898,10.774617,14.4114275,13.879487,10.895341,7.805561,7.5905213,7.322665,9.884277,10.929295,10.47658,12.913695,18.523588,15.562078,12.272349,14.947141,27.947605,18.26705,15.32063,17.595524,21.420965,21.002203,22.232079,25.299223,23.790173,17.074902,10.284176,8.273367,9.25425,8.488406,6.4964604,9.035437,8.831716,10.465261,12.151625,12.064855,8.345046,15.23386,15.47908,12.849561,12.261031,19.787418,18.26705,13.743673,12.027128,13.392818,12.58925,8.047009,7.383027,7.6923823,7.5263867,6.8850408,5.9305663,9.0957985,15.369675,20.492899,16.969267,11.133017,8.062099,5.221313,2.5880208,2.6144292,1.7580433,0.8601585,0.43007925,0.7696155,1.9730829,1.7995421,2.3277097,3.440634,3.9763467,1.7240896,3.4783602,5.3646727,6.1078796,5.4363527,4.093298,3.7688525,4.123479,3.3010468,1.4449154,0.69793564,0.7205714,0.65643674,0.60362,0.76207024,1.448688,1.0902886,0.935611,1.0186088,1.1393328,0.87147635,0.9280658,1.2487389,1.9504471,3.6481283,7.4584794,6.6662283,5.304311,5.349582,6.4511886,5.9494295,6.9755836,10.733118,13.513543,13.656902,11.574413,9.084481,5.7117543,3.893349,4.715781,7.914967,7.8734684,8.186596,8.469543,8.616675,8.786444,9.661693,9.005256,7.7112455,6.4021444,5.4174895,4.478106,4.2291126,5.2364035,7.254758,9.250477,9.325929,7.835742,6.688864,7.0359454,9.242931,10.042727,8.963757,9.103344,12.479843,20.028866,26.1707,21.998177,15.369675,10.831206,9.646602,9.627739,8.167733,7.424526,7.5490227,6.670001,7.4773426,8.07719,8.726082,9.522105,10.393582,11.879996,11.7894535,10.446399,8.669493,7.7716074,8.443134,8.963757,8.854351,7.9526935,6.432326,7.8696957,9.986138,10.718028,10.638803,12.928786,10.699164,7.643338,5.5570765,5.119452,5.8664317,4.979865,6.066381,6.643593,5.9720654,5.0553174,4.8402777,4.749735,3.863168,2.6182017,2.7917426,1.9504471,1.6033657,1.841041,2.3767538,2.5125682,2.7200627,2.5993385,2.3692086,2.3993895,3.2067313,2.5729303,1.7693611,1.1242423,0.77716076,0.7054809,0.754525,0.49421388,0.38480774,0.49421388,0.52062225,0.46026024,0.69793564,0.7696155,0.62625575,0.633801,0.65643674,0.4979865,0.4074435,0.39989826,0.26408374,0.19994913,0.23390275,0.20372175,0.124496624,0.19240387,0.17354076,0.24522063,0.60362,1.0110635,0.7997965,1.2789198,1.418507,1.6222287,1.9844007,2.2484846,1.8749946,1.8259505,2.3428001,3.150142,3.4745877,7.1038527,5.956975,5.7909794,8.001738,9.631512,2.1994405,0.20749438,1.0751982,2.282438,1.3770081,0.52062225,0.62248313,0.73188925,0.68661773,1.0827434,0.83752275,0.73188925,0.90920264,1.237421,1.3015556,1.2110126,1.0525624,0.9318384,0.90543,0.995973,1.1317875,1.2110126,1.2826926,1.3732355,1.4977322,1.2826926,1.1053791,1.0676528,1.1016065,0.97333723,0.845068,0.7092535,0.59230214,0.52062225,0.52062225,0.5093044,0.5055317,0.5394854,0.5998474,0.6488915,0.63002837,0.663982,0.784706,0.965792,1.0940613,1.1959221,1.1732863,1.146878,1.1959221,1.358145,1.5354583,1.2449663,1.0299267,1.0035182,0.84884065,0.633801,0.5885295,0.46026024,0.22258487,0.09808825,0.10186087,0.10940613,0.12826926,0.19240387,0.34330887,0.5319401,0.66020936,0.8337501,1.0186088,1.0450171,0.965792,0.8903395,0.875249,0.91674787,0.9393836,0.91674787,0.8978847,0.8601585,0.8186596,0.8299775,0.784706,0.80734175,0.8526133,0.8337501,0.6149379,0.58475685,0.65643674,0.663982,0.59607476,0.6187105,0.47912338,0.392353,0.33953625,0.36594462,0.56212115,0.56589377,0.59230214,0.633801,0.68661773,0.7507524,0.8224323,1.0299267,1.056335,0.88279426,0.80356914,1.1808317,1.3166461,1.4901869,1.8334957,2.3503454,2.6446102,2.2786655,2.2447119,2.7841973,3.4029078,3.663219,3.7801702,3.7688525,3.7235808,3.8254418,4.2819295,4.08198,3.270866,2.2560298,1.780679,1.6524098,1.5920477,1.448688,1.2449663,1.177059,1.146878,0.9997456,0.8941121,0.87902164,0.935611,0.95447415,1.0223814,1.1431054,1.2826926,1.3845534,1.418507,1.4524606,1.5430037,1.6825907,1.7957695,2.1164427,2.293756,2.3201644,2.323937,2.5804756,2.516341,2.4295704,2.5578396,2.9501927,3.4444065,3.531177,3.5990841,3.5839937,3.5462675,3.640583,3.8443048,4.093298,4.447925,4.798779,4.859141,4.696918,4.636556,4.4931965,4.293247,4.2517486,4.6214657,5.1345425,5.553304,5.80607,5.9796104,5.775889,5.7004366,5.66271,5.59103,5.4212623,5.2552667,5.1081343,5.089271,5.300538,5.8437963,5.8626595,5.9984736,6.1003346,6.013564,5.587258,0.06413463,0.07922512,0.13958712,0.15845025,0.116951376,0.0754525,0.09808825,0.041498873,0.08299775,0.21503963,0.24899325,0.47157812,0.5093044,0.47912338,0.47535074,0.56589377,0.56589377,0.6790725,0.79602385,0.8224323,0.6790725,0.9280658,1.0902886,1.2864652,1.4298248,1.237421,1.3430545,1.237421,1.1091517,1.0110635,0.87147635,0.7884786,0.7884786,0.8262049,0.8111144,0.6149379,0.45648763,0.5583485,0.62248313,0.6111652,0.7696155,0.98465514,1.3732355,1.4524606,1.2336484,1.1883769,1.056335,0.9393836,0.7469798,0.48666862,0.25276586,0.18485862,0.2678564,0.38858038,0.6526641,1.3996439,1.358145,1.8448136,1.9768555,1.8221779,2.3578906,2.6219745,3.712263,6.092789,8.669493,8.809079,9.525878,11.310329,14.581196,18.312323,20.036411,19.613878,19.628967,21.983086,24.997414,23.394047,19.900597,17.82188,15.954432,14.479335,14.939595,15.297995,15.686575,16.678776,16.927769,13.147598,7.6886096,5.8173876,5.5193505,5.8136153,6.741681,6.63982,6.8699503,7.1038527,7.092535,6.6850915,7.149124,7.8621507,8.152642,7.8696957,7.383027,6.8058157,6.670001,6.247467,5.587258,5.511805,6.247467,6.72659,7.284939,7.6622014,7.001992,7.84706,7.303802,5.6853456,4.217795,5.0213637,4.0593443,3.482133,3.5764484,3.92353,3.3915899,5.5495315,5.8664317,5.7570257,7.5792036,14.641558,13.713491,9.522105,6.752999,6.48137,6.175787,4.4516973,3.6179473,3.6556737,4.146115,4.244203,4.478106,3.5802212,3.1576872,3.4029078,3.0633714,2.252257,5.4288073,8.722309,9.963503,8.699674,7.5792036,7.5829763,9.012801,10.691619,9.971047,9.820143,10.514306,10.03141,8.231868,6.8397694,7.4697976,8.318638,10.435081,12.800517,12.340257,12.287439,11.7555,11.476325,11.200924,9.65792,9.525878,10.269085,11.400873,12.336484,12.396846,12.81938,13.570132,15.007503,17.01831,19.029121,18.38023,17.493662,16.546734,15.448899,13.845533,13.211733,13.494679,15.294222,18.651857,23.054512,24.657877,27.85329,30.777075,31.007204,25.563307,20.557034,15.863888,14.219024,15.482853,16.663685,16.0827,16.965494,18.112373,18.678267,18.150099,17.056038,14.950912,12.483616,10.868933,11.891314,12.830698,11.77059,10.872705,10.763299,10.540714,11.563096,11.080199,9.903141,8.703445,8.013056,5.8400235,4.52715,4.285702,5.304311,7.7716074,9.246704,11.544232,14.852824,19.549744,26.197107,25.19359,17.640795,10.544487,6.4926877,3.682082,3.7009451,3.8065786,4.5950575,6.7379084,10.963248,13.219278,19.806282,30.694077,45.478996,63.4216,45.369587,30.041412,20.57967,15.999702,11.208468,9.371201,6.8850408,5.2854476,5.0968165,5.855114,7.1038527,7.598067,8.126234,9.110889,10.612394,10.370946,10.3634,10.227587,9.397609,7.111398,5.3156285,5.8928404,6.971811,7.352846,6.5228686,7.1604424,8.465771,10.521852,12.845788,14.381247,13.72481,9.8239155,7.149124,7.183078,8.420499,11.98563,12.00072,9.590013,6.7680893,6.4247804,7.567886,11.431054,13.290957,12.974057,14.864142,18.599041,17.4333,15.928022,18.078419,27.317577,21.82841,17.591751,15.743164,15.841252,15.856343,19.953413,25.917934,27.804247,23.277096,13.588995,10.265312,12.347801,14.5132885,14.071891,10.967021,12.491161,14.18507,13.95494,12.0233555,10.914205,26.034885,21.1267,17.040947,18.874443,15.946886,15.9695215,14.347293,12.340257,10.616167,9.273112,11.955449,14.275613,13.140053,9.703192,9.348565,9.246704,8.76758,10.099318,12.47607,12.223305,9.159933,8.103599,6.3719635,3.8254418,2.8332415,2.1768045,1.3468271,0.86770374,1.3732355,3.610402,3.4972234,2.8596497,3.0520537,3.4745877,1.5882751,5.6023483,6.255012,5.621211,4.738417,3.6179473,2.886058,2.6295197,1.8184053,0.6073926,0.34330887,0.56589377,0.452715,0.36971724,0.52439487,0.9507015,0.6828451,0.5583485,0.724344,0.98842776,0.8262049,0.6526641,0.845068,1.5845025,3.4783602,7.5565677,8.099826,6.9265394,6.375736,6.5756855,5.4401255,7.1340337,12.728837,16.558052,16.320375,13.087236,8.98262,5.4401255,4.055572,5.481624,9.424017,7.7301087,7.8923316,8.567632,9.291975,10.510533,11.114153,10.023865,8.416726,6.911449,5.5985756,4.5950575,4.5837393,5.1156793,6.300284,8.809079,10.914205,9.5183325,7.8131065,7.9036493,10.801025,10.495442,9.34102,10.050273,14.000212,21.232334,23.643042,18.651857,14.049255,12.238396,10.197406,9.495697,8.126234,7.2396674,7.0548086,6.8699503,7.375482,8.627994,8.778898,8.201687,9.495697,10.902886,10.253995,9.26934,8.511042,7.3905725,8.6732645,8.75249,8.209232,7.5301595,7.1302614,7.6395655,8.986393,9.258021,8.89585,10.684074,11.559323,9.190115,6.7379084,5.59103,5.3910813,4.123479,4.5309224,5.2628117,5.2364035,3.6481283,4.074435,4.1574326,3.5839937,2.7087448,2.5502944,1.8221779,1.3128735,1.4298248,1.9466745,1.9994912,2.071171,2.2598023,2.4220252,2.565385,2.8747404,2.795515,2.1881225,1.4675511,0.98465514,1.0336993,1.1846043,0.80356914,0.56589377,0.65643674,0.7432071,0.51684964,0.59230214,0.6752999,0.6413463,0.5394854,0.5696664,0.49044126,0.4074435,0.35085413,0.26408374,0.21503963,0.2867195,0.24522063,0.11317875,0.15845025,0.181086,0.21503963,0.452715,0.72811663,0.52062225,0.8941121,1.1016065,1.267602,1.4901869,1.8636768,1.6410918,1.4260522,1.9466745,2.9011486,2.9351022,4.7836885,5.300538,5.5004873,8.318638,18.595268,4.217795,0.271629,0.452715,1.1317875,1.3619176,0.45648763,0.38858038,0.5319401,0.6375736,0.83752275,0.87902164,0.7167987,0.76584285,1.0336993,1.1091517,1.1129243,0.97710985,0.86770374,0.84884065,0.9016574,0.97333723,1.1129243,1.3241913,1.5656394,1.7618159,1.4109617,1.2223305,1.116697,1.0487897,0.9808825,0.88279426,0.7809334,0.663982,0.5583485,0.5394854,0.4979865,0.5319401,0.6111652,0.68661773,0.6752999,0.7432071,0.79602385,0.8865669,1.0072908,1.0978339,1.2147852,1.2298758,1.2638294,1.2902378,1.1431054,1.2147852,1.1242423,0.95447415,0.7809334,0.663982,0.58475685,0.44894236,0.27917424,0.1358145,0.090543,0.09808825,0.1056335,0.12826926,0.20749438,0.3961256,0.6488915,0.8337501,0.94315624,0.995973,1.0336993,1.0110635,0.91674787,0.8337501,0.7997965,0.79602385,0.845068,0.84884065,0.845068,0.8337501,0.7884786,0.69793564,0.68661773,0.73566186,0.76207024,0.60362,0.5885295,0.6149379,0.55080324,0.42630664,0.4376245,0.46026024,0.43385187,0.3734899,0.33953625,0.4074435,0.46026024,0.5093044,0.6073926,0.7394345,0.8224323,0.9808825,1.2185578,1.2261031,0.97333723,0.7092535,0.8978847,0.98465514,1.2449663,1.6976813,2.123988,2.2598023,2.0145817,1.9089483,2.1353056,2.546522,2.987919,3.482133,3.8593953,4.025391,3.953711,3.6594462,3.2859564,2.674791,1.961765,1.5807298,1.3770081,1.267602,1.1695137,1.0601076,0.9808825,0.935611,0.90543,0.90543,0.9280658,0.94692886,0.9393836,0.9997456,1.1053791,1.2336484,1.3392819,1.4637785,1.5807298,1.6976813,1.8146327,1.9240388,2.1654868,2.263575,2.2371666,2.2069857,2.4031622,2.4786146,2.4333432,2.6031113,3.048281,3.5387223,3.5877664,3.6783094,3.7386713,3.7499893,3.742444,3.6934,3.7877154,4.006528,4.217795,4.1612053,4.112161,4.0593443,4.032936,4.055572,4.1083884,4.564876,5.0968165,5.4778514,5.6853456,5.904158,5.704209,5.481624,5.3269467,5.160951,4.749735,4.485651,4.4101987,4.4818783,4.715781,5.1835866,5.481624,5.5985756,5.515578,5.3344917,5.2628117,0.05281675,0.0754525,0.12826926,0.1358145,0.094315626,0.05281675,0.094315626,0.056589376,0.049044125,0.071679875,0.03772625,0.35085413,0.392353,0.35839936,0.38858038,0.58475685,0.67152727,0.7092535,0.7130261,0.7130261,0.7582976,0.9997456,1.177059,1.4675511,1.7316349,1.4864142,1.5354583,1.4562333,1.2449663,0.98842776,0.8601585,0.9205205,0.90543,0.9280658,0.9205205,0.6526641,0.4376245,0.52439487,0.6488915,0.70170826,0.73188925,1.1204696,1.659955,1.8938577,1.7919968,1.750498,1.1431054,0.7997965,0.5772116,0.3961256,0.25276586,0.23013012,0.30181,0.43385187,0.7469798,1.50905,1.1921495,1.5354583,1.8448136,2.0183544,2.5616124,2.1277604,3.5538127,6.511551,9.14107,8.058327,9.623966,14.226569,19.112118,22.315077,22.639523,20.69662,18.285913,17.874697,19.01403,18.342503,18.28214,17.497435,15.441354,13.694629,15.965749,17.25976,16.195879,15.928022,16.840998,16.535416,10.612394,7.0849895,5.8136153,6.5040054,8.737399,8.575176,8.888305,8.926031,8.582722,8.394091,9.118435,9.540969,9.665465,9.680555,9.952185,8.348819,6.990674,6.0324273,5.2967653,4.2592936,4.1612053,4.7572803,5.753253,6.719045,7.073672,7.654656,7.0359454,6.0286546,5.455216,6.1342883,4.0970707,2.5389767,2.173032,2.6898816,2.7728794,4.9459114,5.191132,4.61392,4.821415,7.914967,7.33021,4.90064,3.6066296,3.7801702,3.1199608,2.04099,1.9391292,2.5691576,3.2520027,2.8709676,2.0636258,1.8448136,2.1541688,2.584248,2.354118,2.686109,6.7152724,10.412445,11.604594,9.982366,8.582722,8.835487,10.423763,12.147853,11.92904,10.978339,10.63503,10.601076,10.789707,11.321648,10.303039,9.435335,9.397609,10.178542,11.091517,11.091517,11.472552,12.0233555,12.264804,11.423509,9.676784,9.673011,10.729345,12.147853,13.245687,13.128735,12.875969,13.985121,16.177015,17.414436,15.920478,16.418465,16.833452,16.4826,16.105335,13.373956,12.909923,14.5132885,17.614386,21.281378,23.948624,29.022804,31.807001,30.26777,25.016277,21.032385,16.365646,14.015302,14.886778,17.77661,17.335213,16.659912,16.644821,17.297485,17.723793,17.014538,15.445127,13.321139,11.506506,11.423509,11.868678,12.287439,11.92904,10.861387,10.008774,10.751981,10.529396,9.733373,8.684583,7.647111,5.4212623,4.214022,3.983892,4.6026025,5.8173876,7.673519,9.808825,12.291212,16.014793,22.692339,22.858335,15.928022,9.725827,6.6322746,3.6028569,3.3312278,3.561358,4.002755,5.1458607,8.269594,11.219787,16.803272,26.483828,39.601246,53.371326,40.438766,30.041412,22.718748,17.859608,13.717264,13.472044,10.770844,7.432071,5.304311,6.2851934,7.062354,7.4697976,8.258276,9.899368,12.577931,13.309821,12.381755,11.61214,11.249968,9.97482,7.5829763,7.2660756,7.5716586,7.515069,6.590776,6.5530496,6.6360474,7.7829256,9.97482,12.2270775,14.581196,10.438853,7.3000293,7.3981175,7.699928,11.9064045,15.279131,14.132254,9.454198,6.9227667,9.87296,14.04171,16.29774,16.222288,16.078928,17.391802,17.21826,17.655886,19.719511,23.333685,22.560297,19.346022,17.214487,17.150352,17.60684,18.866898,23.26955,26.8045,26.140518,18.595268,15.728074,18.648085,26.864862,30.690304,11.25374,14.803781,17.267305,15.663939,12.264804,14.581196,28.35505,28.207916,24.205162,20.172226,13.656902,12.1252165,15.716756,14.1058445,8.692128,12.596795,13.917213,14.596286,13.781399,11.936585,10.808571,10.269085,7.8432875,5.8173876,5.27413,6.1003346,5.564622,6.205968,6.0739264,4.7874613,3.531177,4.293247,3.3727267,2.1805773,2.11267,4.5497856,6.2663302,5.50426,4.4139714,3.531177,1.7655885,5.5268955,5.2326307,3.8971217,2.9426475,2.1956677,1.5505489,1.0714256,0.7092535,0.4979865,0.543258,0.7205714,0.5394854,0.45648763,0.5583485,0.55080324,1.0827434,1.2487389,1.2449663,1.1996948,1.1581959,1.3505998,1.931584,2.8219235,4.5988297,8.488406,9.2995205,8.024373,6.9265394,6.48137,5.406172,7.99042,13.875714,17.833199,17.70493,14.381247,10.284176,6.3153744,4.8063245,6.428553,10.212496,8.179051,8.224322,9.231613,10.367173,11.072655,12.027128,10.880251,9.099571,7.3000293,5.2364035,4.002755,4.074435,4.142342,4.3800178,6.462507,10.197406,10.895341,9.839006,8.793989,10.001229,10.197406,9.420244,10.257768,13.826671,19.723284,17.410664,15.350811,13.951167,12.593022,9.639057,8.296002,7.8017883,7.6282477,7.586749,7.8508325,7.5263867,9.0957985,8.8769865,7.567886,10.212496,10.868933,9.465516,8.345046,8.16396,7.914967,9.242931,9.295748,8.854351,8.582722,9.050528,7.7829256,8.126234,8.16396,7.8017883,8.793989,11.796998,10.397354,8.269594,6.862405,5.3910813,4.4215164,4.406426,4.9760923,5.172269,3.4557245,4.2102494,4.3913355,3.731126,2.6031113,2.022127,1.5845025,1.20724,1.2525115,1.599593,1.6373192,1.4901869,1.7957695,2.2258487,2.4710693,2.2409391,2.795515,2.3277097,1.5505489,1.0412445,1.2223305,1.4600059,1.0450171,0.72811663,0.73188925,0.76207024,0.55080324,0.4979865,0.51684964,0.513077,0.392353,0.44894236,0.41876137,0.35085413,0.27917424,0.24899325,0.20372175,0.32821837,0.3169005,0.15467763,0.1358145,0.19994913,0.20372175,0.3169005,0.49044126,0.44894236,0.69039035,0.87147635,0.995973,1.1393328,1.4449154,1.5241405,1.267602,1.8599042,2.9652832,2.7087448,3.31991,4.696918,4.7950063,6.349328,16.87118,4.5535583,0.5885295,0.08677038,0.5772116,2.033445,0.663982,0.26031113,0.482896,0.8186596,0.58475685,0.86770374,0.845068,0.79602385,0.88279426,1.1355602,1.116697,0.935611,0.77338815,0.7205714,0.76207024,0.83752275,0.98465514,1.2600567,1.5807298,1.7316349,1.4977322,1.2826926,1.0789708,0.94315624,0.9997456,0.95447415,0.875249,0.76207024,0.6451189,0.5696664,0.55457586,0.6111652,0.694163,0.76584285,0.77716076,0.9280658,1.0186088,1.0336993,1.0148361,1.0487897,1.2713746,1.327964,1.3241913,1.2525115,0.9997456,0.88279426,0.87147635,0.8262049,0.724344,0.66020936,0.5357128,0.32067314,0.17354076,0.12826926,0.1056335,0.1056335,0.10940613,0.15467763,0.29049212,0.58098423,0.7394345,0.8978847,1.0035182,1.0110635,0.9016574,0.965792,0.90543,0.814887,0.754525,0.754525,0.72811663,0.7432071,0.7997965,0.84884065,0.7809334,0.6488915,0.5583485,0.5583485,0.6111652,0.58098423,0.573439,0.5583485,0.49044126,0.3961256,0.40367088,0.41121614,0.3961256,0.36971724,0.3470815,0.3734899,0.45648763,0.5772116,0.7054809,0.814887,0.8903395,1.0148361,1.1317875,1.1431054,0.9997456,0.7167987,0.83752275,0.90920264,1.116697,1.4411428,1.6863633,1.7127718,1.6071383,1.539231,1.6033657,1.8146327,2.2711203,2.7992878,3.31991,3.6330378,3.4368613,2.7540162,2.354118,1.9693103,1.569412,1.3355093,1.1695137,0.9620194,0.8526133,0.84884065,0.8111144,0.754525,0.7922512,0.8601585,0.9205205,0.9808825,1.1129243,1.1053791,1.1544232,1.2751472,1.2789198,1.4260522,1.5958204,1.7882242,1.9542197,1.9730829,2.093807,2.1390784,2.1390784,2.142851,2.203213,2.463524,2.637065,2.8558772,3.138824,3.3953626,3.519859,3.6669915,3.7613072,3.772625,3.7160356,3.5575855,3.4934506,3.5877664,3.742444,3.7009451,3.802806,3.8178966,3.8858037,4.006528,4.0517993,4.4894238,4.9760923,5.3609,5.6061206,5.775889,5.775889,5.5683947,5.342037,5.0439997,4.376245,3.9574835,3.802806,3.8820312,4.146115,4.564876,4.8025517,4.908185,4.7874613,4.568649,4.606375,0.08299775,0.08299775,0.071679875,0.05281675,0.03772625,0.060362,0.120724,0.08299775,0.030181,0.00754525,0.041498873,0.2678564,0.26031113,0.32444575,0.513077,0.6488915,0.7054809,0.5055317,0.41121614,0.5583485,0.87902164,0.97333723,1.1053791,1.4147344,1.7391801,1.6109109,1.6561824,1.5920477,1.3128735,0.9808825,1.0336993,1.1506506,1.1280149,1.1091517,1.0487897,0.73566186,0.43385187,0.29426476,0.392353,0.573439,0.45648763,0.7809334,1.2826926,1.6976813,1.9202662,1.9768555,1.3204187,0.79602385,0.47157812,0.32067314,0.241448,0.35462674,0.3772625,0.5281675,0.7696155,0.83752275,0.7130261,0.8224323,1.4675511,2.6672459,4.1310244,5.0025005,6.25124,7.907422,9.1825695,8.458225,11.514051,15.9695215,18.674494,18.983849,18.761265,17.444618,15.961976,15.0376835,15.377219,17.670975,18.983849,17.587978,14.698147,12.457208,13.913441,16.520325,14.298248,11.815862,11.691365,14.618922,11.091517,8.065872,7.0170827,8.401636,11.657412,11.77059,11.781908,11.23865,10.393582,10.212496,11.604594,11.944131,12.106354,12.445889,12.759018,10.352083,7.6395655,5.66271,4.353609,2.5314314,1.991946,2.8294687,3.85185,4.425289,4.459243,4.5497856,4.1800685,4.666737,5.7570257,5.6287565,3.8178966,2.2748928,1.629774,2.252257,4.255521,5.6400743,5.9494295,5.855114,5.402399,3.9914372,2.003264,0.94315624,0.8601585,1.3807807,1.7052265,1.3392819,1.8900851,2.6521554,3.150142,3.108643,2.1051247,2.0183544,2.5917933,3.5047686,4.3385186,3.742444,6.205968,8.763808,9.993684,10.008774,9.461743,9.125979,9.318384,10.057818,11.106608,12.645839,12.411936,11.936585,12.14408,13.340002,10.63503,9.7069645,8.14887,6.8359966,9.906913,10.208723,10.902886,11.638548,12.581704,14.403882,13.12119,12.721292,12.00072,11.302785,12.54775,12.147853,12.00072,13.226823,14.679284,12.947649,13.057055,15.23386,16.388283,15.897841,15.580941,13.762536,14.007756,14.913187,15.829934,16.856089,21.952906,27.577888,29.109575,26.431011,23.933533,21.171972,16.897587,14.083209,14.222796,17.335213,16.293968,15.75071,16.407146,17.523844,16.931541,15.30554,13.396591,12.045992,11.434827,11.0613365,11.502733,13.490907,13.656902,11.68382,10.295494,9.933322,9.175024,8.850578,8.612903,6.937857,5.6287565,4.9157305,4.4139714,4.093298,4.255521,6.4549613,7.745199,8.941121,11.834724,19.206434,19.538425,14.053028,8.83926,5.9796104,3.5462675,3.138824,3.772625,3.874486,3.712263,5.4250345,8.360137,12.362892,21.78691,35.28159,45.807213,43.00038,35.666397,26.864862,19.40261,15.829934,16.644821,15.256495,10.691619,5.6098933,6.326692,6.1908774,6.8661776,7.9489207,9.684328,12.97783,17.139036,15.754482,13.502225,12.619431,12.917468,10.457717,8.816625,7.779153,7.213259,7.032173,6.549277,6.228604,6.470052,7.2698483,8.20546,9.95973,8.797762,8.582722,9.552286,8.322411,12.46098,19.43279,20.168453,14.049255,8.933576,13.132507,17.425755,19.783646,19.447882,16.954176,16.248695,16.101564,18.8254,21.96045,18.297232,19.24416,18.119919,18.931032,22.04722,24.178753,20.704166,21.077656,23.08092,24.484337,23.073374,21.632233,23.876944,38.20537,47.855747,10.933067,15.505488,19.934551,17.80679,12.215759,15.769572,26.163155,33.334915,27.634478,14.596286,14.93205,10.801025,15.645076,14.754736,9.431562,16.98813,9.812597,7.8131065,10.050273,12.58925,8.480861,7.5527954,7.0548086,5.3344917,2.8596497,2.2409391,2.3692086,3.0445085,4.0178456,4.647874,3.9197574,5.828706,5.032682,3.5123138,2.8445592,4.2102494,8.590267,9.06939,7.4282985,4.8629136,2.022127,2.9539654,2.6710186,1.9164935,1.2147852,0.8563859,0.88279426,1.0450171,1.1280149,1.0374719,0.80734175,0.7884786,0.7696155,0.84884065,0.965792,0.90920264,2.1579416,2.4559789,2.093807,1.5618668,1.539231,2.5201135,3.8858037,5.3194013,7.2887115,11.019837,11.642321,10.33322,8.578949,7.020855,5.462761,7.798016,13.004238,16.950403,17.474798,14.392565,11.563096,7.4207535,5.492942,6.85486,10.125726,8.60913,8.703445,9.903141,11.02361,10.201178,11.721546,10.978339,9.469289,7.6622014,4.957229,2.957738,2.8596497,2.806833,2.5578396,3.4934506,7.533932,11.559323,12.562841,10.34831,7.5565677,9.544742,9.665465,10.56335,13.313594,17.425755,11.940358,13.151371,13.93985,11.978085,9.759781,8.080963,7.809334,8.246958,8.956212,9.793735,7.8734684,9.061845,9.092027,8.348819,11.857361,11.363147,9.691874,8.254503,7.888559,8.83926,9.49947,9.81637,9.997457,10.178542,10.435081,7.6508837,7.4018903,7.635793,7.6848373,8.303548,10.895341,10.114408,8.733627,7.7225633,6.2814207,5.9720654,5.4740787,5.311856,5.3458095,4.776143,4.772371,5.160951,4.504514,2.837014,1.6561824,1.4298248,1.297783,1.3091009,1.448688,1.6448646,1.2034674,1.4864142,1.9768555,2.2220762,1.8146327,2.5767028,2.1051247,1.4260522,1.1204696,1.3204187,1.5769572,1.2298758,0.8865669,0.76207024,0.6413463,0.4979865,0.3734899,0.31312788,0.29803738,0.2263575,0.30181,0.29049212,0.23013012,0.17731337,0.211267,0.14335975,0.28294688,0.32821837,0.211267,0.1056335,0.20749438,0.19994913,0.25276586,0.41121614,0.5998474,0.7167987,0.79602385,0.86770374,0.9620194,1.1204696,1.4449154,1.1921495,1.720317,2.8256962,2.7426984,3.1840954,3.9725742,3.8858037,3.821669,6.828451,3.6368105,1.1581959,0.049044125,0.6187105,2.8445592,1.0336993,0.31312788,0.58475685,1.1053791,0.48666862,0.784706,0.9620194,0.91674787,0.8563859,1.3317367,1.3204187,0.9808825,0.6790725,0.5583485,0.55080324,0.6488915,0.73188925,0.9620194,1.2562841,1.3166461,1.3958713,1.2411937,1.0450171,0.94692886,1.0299267,1.0299267,0.95824677,0.8526133,0.73188925,0.60362,0.6451189,0.7167987,0.784706,0.8526133,0.9507015,1.0450171,1.177059,1.177059,1.0412445,0.9318384,1.2110126,1.2751472,1.2185578,1.086516,0.90920264,0.663982,0.573439,0.5885295,0.6413463,0.66775465,0.43007925,0.23390275,0.14335975,0.14335975,0.124496624,0.116951376,0.14335975,0.24899325,0.4678055,0.8337501,0.8639311,0.86770374,0.95824677,1.0374719,0.814887,0.91297525,0.8903395,0.8186596,0.7582976,0.77716076,0.6149379,0.60362,0.68661773,0.77338815,0.7432071,0.633801,0.51684964,0.482896,0.52062225,0.52062225,0.5470306,0.55457586,0.543258,0.52439487,0.52062225,0.362172,0.29426476,0.30935526,0.3772625,0.452715,0.52062225,0.72811663,0.87147635,0.9016574,0.8941121,0.8111144,0.7884786,0.83752275,0.9205205,0.935611,1.0638802,1.056335,1.0223814,1.0299267,1.1016065,1.2864652,1.2789198,1.3053282,1.4222796,1.50905,1.7957695,2.0183544,2.3767538,2.727608,2.5767028,2.0975795,1.7014539,1.388326,1.1846043,1.177059,1.1544232,0.91674787,0.7469798,0.7205714,0.7092535,0.69039035,0.73566186,0.814887,0.9205205,1.0676528,1.3958713,1.3128735,1.3015556,1.4298248,1.3430545,1.3996439,1.5165952,1.7580433,1.9957186,1.8674494,1.8938577,1.931584,2.003264,2.1013522,2.1881225,2.5540671,2.897376,3.1048703,3.1652324,3.1614597,3.3651814,3.5085413,3.531177,3.4670424,3.451952,3.3538637,3.229367,3.270866,3.482133,3.663219,3.7801702,3.8895764,4.002755,4.08198,4.055572,4.3347464,4.678055,5.0553174,5.3948536,5.583485,5.873977,5.885295,5.6891184,5.281675,4.561104,3.9574835,3.5651307,3.531177,3.8141239,4.1762958,4.085753,4.2102494,4.195159,3.9876647,3.8292143,0.1659955,0.08299775,0.033953626,0.026408374,0.049044125,0.060362,0.011317875,0.0,0.0,0.041498873,0.19994913,0.11317875,0.071679875,0.116951376,0.24899325,0.44139713,1.0148361,1.0035182,0.814887,0.6828451,0.67152727,0.7582976,1.1619685,1.4373702,1.478869,1.5241405,1.4034165,1.3732355,1.2449663,1.1431054,1.50905,1.50905,1.6939086,1.8599042,1.8825399,1.7240896,1.0412445,0.48666862,0.31312788,0.4074435,0.26031113,0.43007925,0.5093044,0.814887,1.2223305,1.1581959,0.80734175,0.4979865,0.30181,0.23013012,0.23013012,0.59607476,0.59607476,0.8526133,1.2789198,1.0827434,0.80356914,1.0148361,2.1503963,4.0480266,5.9494295,11.321648,15.116908,16.546734,16.331694,16.724047,15.55076,14.298248,13.951167,13.70972,10.985884,11.717773,12.2119875,12.596795,13.555041,16.32792,18.1086,18.534906,16.161926,12.178034,10.423763,9.0543,8.959985,8.986393,8.744945,8.635539,7.3679366,6.6850915,7.0057645,8.507269,11.106608,10.789707,10.016319,9.156161,8.4544525,8.028146,10.453944,11.521597,11.246195,9.854096,7.7678347,6.620957,6.0286546,4.8402777,3.218049,2.655928,3.4255435,4.8063245,4.9723196,3.712263,2.4559789,1.7995421,1.2751472,1.9730829,3.6028569,4.5309224,4.3611546,3.4481792,2.637065,2.425798,2.9766011,4.8553686,6.3153744,7.443389,7.3717093,4.2706113,1.9881734,0.84129536,0.5319401,0.66775465,0.77716076,1.2411937,1.5958204,2.2673476,3.1840954,3.7688525,2.8030603,2.0145817,1.9164935,2.655928,3.9989824,2.9728284,3.2821836,4.2064767,5.1760416,5.798525,7.3000293,8.269594,8.0206,7.5905213,9.752235,15.011275,16.4826,15.769572,14.158662,12.619431,9.933322,9.242931,8.858124,8.001738,6.8058157,10.759526,11.68382,11.729091,12.268577,13.917213,17.25976,17.931286,16.199652,13.181552,10.850069,10.03141,10.284176,11.114153,11.4838705,9.812597,12.155397,14.003984,14.981093,14.577423,12.162943,11.868678,11.329193,11.732863,12.581704,11.7026825,15.365902,21.153109,23.43932,22.137764,22.673477,19.478064,17.414436,15.294222,13.600313,14.464244,15.565851,17.029629,17.448391,15.758255,11.231105,11.012292,10.982111,10.789707,10.56335,10.940613,12.223305,12.321393,11.419736,10.295494,10.344538,9.016574,7.9791017,8.428044,9.159933,6.5455046,5.873977,5.9984736,5.3269467,3.9386206,3.5839937,5.149633,6.2814207,6.8133607,8.318638,14.128481,13.483362,10.748209,7.564113,5.0213637,3.6934,2.9728284,3.663219,3.8141239,3.218049,3.3878171,4.6818275,6.4436436,14.053028,26.555508,36.65105,45.524265,36.685005,25.197363,18.357594,15.671484,13.498452,19.059301,18.127462,9.537196,5.20245,5.3986263,6.7643166,8.047009,9.337247,12.083718,18.395319,19.606333,16.614641,12.562841,12.83447,11.917723,10.642575,10.227587,10.352083,9.156161,10.20495,11.080199,12.611885,13.95494,12.58925,11.246195,10.057818,12.132762,15.082954,11.031156,9.507015,11.898859,15.030138,15.988385,12.128989,14.913187,19.123436,22.458437,23.156372,20.017548,18.433046,17.908651,24.442837,31.395784,19.470518,14.879233,12.551523,13.95494,18.391546,22.99415,21.726547,18.13878,15.4074,15.90916,21.254969,19.70442,18.723537,33.93476,48.90831,15.181043,16.890041,26.40083,23.111101,9.190115,9.567377,38.058243,30.260225,18.94235,16.45619,14.724555,16.188334,10.631257,8.307321,10.529396,9.673011,3.874486,6.8925858,10.502988,9.752235,2.9766011,6.4436436,12.31762,12.030901,5.583485,1.5580941,1.7165444,1.9391292,2.493705,3.1237335,3.0520537,2.5012503,2.546522,3.1161883,3.4670424,2.1956677,6.8473144,9.046755,8.98262,6.6586833,1.8599042,2.0447628,2.7238352,2.4182527,1.2110126,0.7469798,1.5052774,2.5917933,2.927557,2.1164427,0.44139713,0.47912338,1.3128735,1.6863633,1.50905,1.8599042,2.8747404,2.625747,2.1843498,1.9278114,1.5241405,3.270866,5.4476705,8.695901,12.691111,16.158154,16.976812,16.74291,13.72481,8.733627,5.0968165,5.4401255,10.925522,16.003475,17.320122,13.732355,10.521852,7.6697464,6.5530496,7.586749,10.223814,7.1340337,7.01331,8.171506,9.239159,9.14107,10.201178,10.072908,9.280658,7.9715567,5.9192486,3.0633714,2.1466236,2.0258996,2.0183544,1.9089483,5.3609,12.404391,16.603323,15.086727,8.544995,9.397609,10.152134,11.246195,13.249459,16.874952,13.189097,12.83447,12.513797,11.491416,11.627231,11.332966,9.303293,8.941121,10.853842,12.830698,9.193887,8.707218,9.005256,9.5032425,11.3820095,10.321902,9.012801,8.009283,7.7678347,8.620448,8.695901,9.208978,10.110635,10.593531,9.0807085,5.4174895,5.0968165,6.1531515,7.2924843,7.888559,7.069899,6.2889657,5.772116,5.670255,6.0739264,6.964266,5.3458095,4.2894745,4.9119577,6.3644185,5.5080323,5.0854983,4.908185,4.2819295,1.9994912,1.5467763,1.2789198,1.20724,1.327964,1.6335466,1.2789198,1.6561824,1.9429018,1.8636768,1.6939086,2.1202152,1.780679,1.4600059,1.4675511,1.6033657,2.003264,1.6863633,1.2751472,1.0450171,0.8865669,0.60362,0.422534,0.35085413,0.32444575,0.21503963,0.19994913,0.2263575,0.21503963,0.16222288,0.1358145,0.10186087,0.10186087,0.150905,0.19240387,0.1056335,0.1659955,0.17354076,0.22258487,0.36594462,0.6111652,0.62248313,0.76207024,0.9695646,1.1091517,0.9620194,1.267602,1.0299267,0.965792,1.4864142,2.7313805,2.7804246,2.5729303,2.493705,2.8521044,3.874486,4.08198,1.7655885,0.116951376,0.21881226,1.0374719,1.0751982,0.5055317,0.59230214,1.1846043,0.73188925,0.7432071,0.91297525,0.935611,0.95447415,1.5430037,1.7240896,1.1091517,0.59230214,0.4678055,0.44139713,0.47912338,0.543258,0.66020936,0.80734175,0.91674787,0.91674787,1.0638802,1.1280149,1.056335,0.94692886,0.94692886,0.95447415,0.8865669,0.76207024,0.70170826,0.7130261,0.7997965,0.94692886,1.1204696,1.267602,0.97333723,1.0299267,1.1204696,1.0525624,0.7469798,0.87147635,0.9997456,1.0676528,0.995973,0.70170826,0.543258,0.513077,0.482896,0.422534,0.41121614,0.25276586,0.13958712,0.1056335,0.124496624,0.1358145,0.1358145,0.2565385,0.49421388,0.77338815,0.9318384,1.237421,0.9997456,0.80734175,0.8639311,1.0223814,1.0714256,0.965792,0.7696155,0.6073926,0.65643674,0.52062225,0.4979865,0.4979865,0.48666862,0.48666862,0.513077,0.55457586,0.63002837,0.6526641,0.45648763,0.44516975,0.46026024,0.45648763,0.422534,0.3961256,0.3470815,0.34330887,0.41876137,0.52439487,0.55080324,0.56212115,0.6187105,0.73566186,0.8563859,0.87147635,0.845068,0.965792,1.0525624,1.1657411,1.6184561,1.4335974,1.1883769,0.94315624,0.845068,1.1129243,1.1619685,1.1204696,1.20724,1.4109617,1.4939595,1.7165444,1.9089483,2.2862108,2.674791,2.5012503,2.4522061,2.1315331,1.6976813,1.2751472,0.94692886,0.9695646,0.9205205,0.8526133,0.8337501,0.9318384,1.1129243,1.086516,1.116697,1.2261031,1.1883769,1.3619176,1.358145,1.3505998,1.4147344,1.5241405,1.4298248,1.4222796,1.5430037,1.720317,1.7693611,1.659955,1.6410918,1.8070874,2.1277604,2.4559789,2.7238352,2.7653341,2.897376,3.2105038,3.5387223,3.821669,3.8103511,3.6745367,3.5500402,3.5236318,3.5236318,3.5349495,3.5575855,3.6141748,3.7235808,3.821669,3.8895764,3.9574835,4.06689,4.2894745,4.164978,4.044254,4.195159,4.5799665,4.8365054,5.2288585,5.481624,5.413717,5.0968165,4.851596,4.1310244,3.6594462,3.5689032,3.8103511,4.164978,4.055572,4.063117,4.0593443,3.9386206,3.6481283,0.33953625,0.31312788,0.2565385,0.1358145,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0452715,0.22258487,0.21503963,0.3055826,0.35462674,0.35085413,0.43007925,0.6828451,0.7507524,0.6187105,0.45648763,0.6111652,0.8111144,1.0374719,1.2487389,1.4826416,1.8561316,1.7429527,1.5015048,1.2298758,1.0412445,1.0940613,1.3091009,2.191895,2.6219745,2.2447119,1.478869,0.94315624,0.44516975,0.211267,0.20749438,0.150905,0.36971724,0.47535074,0.56589377,0.6187105,0.5017591,0.5093044,0.422534,0.29049212,0.23013012,0.422534,0.87902164,0.7394345,0.6828451,0.845068,0.814887,0.845068,1.4977322,5.040227,10.099318,11.664956,12.336484,14.196388,15.109364,14.366156,12.706201,12.385528,10.801025,10.33322,11.69891,13.977575,14.84528,13.6682205,13.721037,15.482853,16.644821,17.712475,17.810562,15.626213,12.0233555,10.03141,9.533423,8.718536,7.3981175,5.87775,4.938366,4.4403796,5.20245,6.0286546,6.9454026,9.193887,8.533678,7.8319697,7.194396,6.7341356,6.609639,8.152642,8.714764,7.99042,6.571913,5.9607477,6.247467,6.0701537,5.5268955,5.0854983,5.5495315,5.194905,5.572167,5.726845,5.330719,4.689373,3.7952607,2.9086938,2.6295197,3.169005,4.3611546,3.99521,3.4670424,3.361409,3.682082,3.8405323,3.1539145,3.6556737,4.659192,5.1873593,3.9801195,2.7238352,1.961765,1.4939595,1.4260522,2.1692593,1.4600059,3.0030096,5.6061206,7.756517,7.5905213,5.6400743,4.2517486,3.802806,4.0706625,4.2404304,2.8558772,2.425798,3.4029078,4.9760923,5.040227,6.270103,7.997965,9.978593,12.162943,14.694374,15.705438,15.55076,15.211224,14.577423,12.472299,12.559069,13.317367,12.89106,11.551778,11.714001,11.672502,12.140307,13.155144,14.064346,13.52486,18.002966,20.357084,18.953669,15.181043,13.43809,15.188588,14.3095665,13.0646,12.332711,11.604594,11.487643,11.668729,11.193378,10.544487,11.61214,10.382264,10.140816,10.310584,10.604849,11.046246,13.702174,15.931795,18.02183,19.621422,19.757236,17.165443,16.475054,16.120426,16.06761,17.833199,19.312067,19.168707,17.957695,15.343266,10.084227,11.932813,13.690856,13.8870325,12.611885,11.514051,11.604594,11.495189,11.125471,10.401127,9.208978,8.563859,9.26934,10.797253,11.148107,6.8737226,5.119452,5.100589,4.7120085,3.6971724,3.6481283,3.9386206,4.659192,5.27413,6.228604,8.956212,10.31813,9.590013,6.760544,3.6179473,3.742444,2.6408374,3.029418,3.2255943,2.7615614,2.3880715,2.8030603,3.6971724,8.047009,17.580433,32.78411,37.95638,32.546436,26.668686,22.956423,16.561823,13.558814,15.788436,19.21398,18.516043,7.0963078,6.089017,7.3113475,8.099826,8.382772,10.668983,15.652621,17.395575,14.992412,10.782163,10.367173,13.826671,13.5663595,12.234623,11.276376,10.948157,10.416218,9.725827,10.672756,14.109617,19.94964,14.943368,12.027128,11.106608,11.898859,13.951167,14.094527,15.158407,16.950403,18.297232,17.086218,17.859608,19.91946,21.67373,22.028357,20.387266,19.353567,18.580177,20.470263,22.877197,19.104572,15.705438,12.694883,13.864397,18.293459,20.345766,19.840235,17.652113,14.78869,12.381755,11.672502,10.435081,9.978593,17.210714,25.72553,15.803526,17.80679,28.532362,28.819082,18.749947,17.637022,34.583652,26.585688,17.105082,14.169979,10.355856,7.1340337,7.149124,8.167733,9.7220545,13.117417,9.797507,8.756263,7.5490227,5.8626595,5.515578,13.58145,10.989656,7.2170315,5.2854476,1.7655885,1.9994912,2.3692086,2.5125682,2.565385,3.138824,3.0860074,3.2633207,3.029418,2.305074,1.5618668,5.111907,8.627994,9.737145,7.8696957,4.255521,2.0749438,2.686109,2.9501927,2.0108092,1.3204187,2.546522,4.689373,4.817642,3.048281,2.516341,1.6561824,1.750498,2.2899833,2.9916916,3.8141239,3.8405323,3.6066296,3.3727267,3.9612563,6.749226,8.83926,9.178797,11.034928,14.128481,14.64533,14.351066,16.935314,17.08999,13.328684,8.001738,7.0548086,10.665211,14.279386,15.01882,11.68382,8.695901,6.647365,6.5643673,8.111144,9.574923,7.3868,6.304056,6.277648,7.183078,8.82417,9.220296,8.039464,6.7869525,6.1078796,5.7872066,3.6330378,2.6823363,2.4786146,2.3654358,1.4562333,3.7198083,8.722309,12.853333,13.7700815,10.401127,10.227587,11.446144,12.170488,13.008011,17.033401,15.99593,12.528888,10.121953,9.982366,11.053791,11.472552,9.208978,8.786444,11.434827,15.0905,13.826671,12.223305,11.321648,10.902886,9.491924,8.477088,7.798016,8.175279,9.491924,10.7557535,10.03141,8.197914,7.062354,6.8963585,6.417235,5.089271,5.4703064,6.356873,6.8133607,6.1908774,4.8063245,4.647874,5.172269,5.9305663,6.537959,6.3153744,4.4630156,3.1124156,3.5877664,6.387054,5.6778007,4.2819295,3.772625,3.92353,2.6936543,1.8221779,1.3166461,1.177059,1.2487389,1.2298758,1.177059,1.7278622,2.033445,1.8485862,1.5241405,1.6184561,1.8976303,1.569412,0.8865669,1.1393328,1.1506506,1.1129243,1.0450171,0.95824677,0.84884065,1.1846043,1.0035182,0.63002837,0.3055826,0.17731337,0.1659955,0.15845025,0.13958712,0.1056335,0.10186087,0.124496624,0.10186087,0.120724,0.16222288,0.094315626,0.23390275,0.26031113,0.26408374,0.35462674,0.66020936,0.7884786,0.7469798,0.7205714,0.784706,0.9016574,0.8526133,0.7507524,0.60362,0.6111652,1.1431054,1.6146835,1.871222,3.4934506,5.1534057,2.595566,2.9464202,1.659955,0.482896,0.124496624,0.2678564,0.5093044,0.331991,0.3055826,0.543258,0.7092535,0.66020936,0.9695646,1.0902886,1.0186088,1.2713746,1.2713746,0.97710985,0.633801,0.39989826,0.35839936,0.40367088,0.45648763,0.51684964,0.59230214,0.6828451,0.70170826,0.8978847,0.9695646,0.8639311,0.77338815,0.754525,0.724344,0.7130261,0.70170826,0.59230214,0.59607476,0.633801,0.68661773,0.7394345,0.77716076,0.7582976,0.8224323,0.8903395,0.875249,0.69793564,0.7130261,0.7092535,0.6451189,0.5281675,0.422534,0.36971724,0.35085413,0.3470815,0.32821837,0.27917424,0.15845025,0.09808825,0.090543,0.116951376,0.150905,0.17731337,0.4376245,0.694163,0.83752275,0.87147635,1.0487897,1.0978339,1.0374719,0.94692886,0.9507015,1.0676528,0.9695646,0.7394345,0.5319401,0.5696664,0.49421388,0.63002837,0.7884786,0.84129536,0.7432071,0.7507524,0.65643674,0.59230214,0.5696664,0.482896,0.52062225,0.633801,0.66775465,0.573439,0.422534,0.47157812,0.52062225,0.56589377,0.59607476,0.6111652,0.6828451,0.77716076,0.7997965,0.7582976,0.7582976,0.9808825,1.0827434,0.9242931,0.67152727,0.8111144,0.784706,0.8111144,0.77338815,0.6752999,0.663982,0.7092535,0.83752275,1.0336993,1.2562841,1.4109617,1.3355093,1.2789198,1.388326,1.6637276,1.9391292,1.8448136,1.690136,1.5354583,1.3770081,1.1657411,1.1619685,1.0676528,0.9318384,0.814887,0.784706,0.8299775,0.87147635,0.9016574,0.935611,1.0072908,1.0412445,1.0902886,1.2223305,1.4373702,1.6863633,1.7127718,1.6939086,1.6561824,1.6637276,1.8184053,1.7957695,1.7919968,1.7618159,1.8334957,2.3088465,2.8634224,3.1124156,3.308592,3.5538127,3.783943,3.8593953,3.863168,3.7877154,3.6066296,3.2670932,3.1124156,3.097325,3.2029586,3.3727267,3.5047686,3.6292653,3.640583,3.572676,3.4896781,3.4934506,3.440634,3.591539,3.8065786,3.9612563,3.9348478,4.315883,4.6516466,4.7120085,4.606375,4.8025517,4.29702,3.92353,3.7047176,3.7084904,4.032936,4.0291634,4.0593443,3.9386206,3.7160356,3.6481283,0.21503963,0.20372175,0.28294688,0.20372175,0.0,0.0,0.0452715,0.0452715,0.03772625,0.06413463,0.18485862,0.18863125,0.24899325,0.26408374,0.23767537,0.271629,0.3470815,0.55457586,0.6790725,0.7130261,0.8526133,0.77716076,0.7922512,1.086516,1.5203679,1.6260014,1.478869,1.4034165,1.297783,1.1204696,0.8903395,0.97710985,1.5845025,1.8787673,1.6260014,1.2185578,0.5772116,0.2263575,0.090543,0.071679875,0.056589376,0.23013012,0.33953625,0.38858038,0.3961256,0.4074435,0.331991,0.29049212,0.21503963,0.27540162,0.8941121,1.1431054,1.3015556,1.7919968,2.9652832,5.1232247,6.7567716,7.6320205,8.68081,10.110635,11.427281,11.664956,11.898859,11.208468,9.556059,7.748972,8.643084,8.375228,8.816625,11.197151,16.124199,17.169216,16.516552,16.697638,17.746428,17.225805,17.165443,17.199398,14.456699,9.820143,7.8923316,7.5075235,6.1305156,4.7006907,3.7009451,3.1614597,3.4066803,4.6818275,6.085244,6.9265394,6.7454534,6.6360474,6.149379,5.666483,5.50426,5.9192486,6.7831798,7.062354,6.858632,6.40969,6.1116524,6.809588,6.6662283,6.304056,6.1116524,6.217286,5.1345425,5.1269975,6.039973,7.194396,7.3717093,5.6891184,4.6742826,4.074435,3.8971217,4.398881,4.0291634,3.7499893,3.6971724,3.783943,3.6934,2.6785638,2.9313297,3.240685,3.0256453,2.323937,1.7957695,2.6936543,3.6443558,4.285702,5.2552667,3.338773,4.991183,7.7904706,9.5183325,8.167733,8.284684,7.748972,7.1868505,6.8397694,6.5568223,4.447925,3.2255943,3.1727777,4.0782075,5.2364035,7.122716,9.673011,12.079946,13.807808,14.603831,15.396083,15.928022,15.931795,15.486626,15.026365,15.860115,15.614895,15.022593,14.758509,15.411173,14.988639,15.607349,16.746683,17.693611,17.538933,19.429018,20.764528,19.94964,17.833199,17.73511,19.33093,17.327667,14.830189,13.230596,12.238396,9.235386,7.5075235,6.5228686,6.4134626,7.960239,8.024373,8.741172,9.416472,9.865415,10.431308,12.770335,14.769827,16.991903,18.885761,18.79899,17.176762,17.255987,17.13149,16.863634,18.500954,18.414183,18.648085,17.60684,14.803781,10.831206,11.940358,14.354838,15.373446,14.237886,12.14408,11.129244,10.623712,10.401127,9.933322,8.386545,7.9753294,9.186342,10.7557535,10.751981,6.6020937,5.323174,4.8968673,4.236658,3.3538637,3.350091,3.640583,4.146115,4.881777,5.775889,6.651138,7.6848373,8.59404,8.446907,7.303802,6.224831,3.229367,2.9200118,3.0143273,2.5540671,1.9240388,1.9806281,3.3123648,5.9192486,11.691365,24.435291,30.362085,30.871391,27.60807,22.50748,17.7917,16.448645,15.331948,18.055782,20.251451,9.582467,7.032173,8.941121,10.080454,9.303293,9.574923,12.604341,13.807808,12.494934,9.944639,9.4127,12.234623,14.1926155,14.434063,13.588995,13.788944,12.777881,11.102836,10.687846,12.657157,17.33144,14.426518,12.012038,10.26154,10.552032,15.448899,16.852316,19.25925,20.519308,20.88148,22.975286,24.92196,26.359331,26.393284,25.665169,26.336695,26.823364,25.276588,22.401848,19.281887,17.372938,16.301512,14.437836,15.660167,18.87067,18.018057,16.116653,14.735873,13.815352,12.89106,11.106608,7.8998766,7.194396,10.235131,14.5283785,13.864397,14.407655,23.511,27.39303,25.167181,28.834173,30.675215,24.340977,18.765038,17.248442,17.463482,6.7944975,5.010046,7.5112963,11.498961,15.961976,14.781145,9.280658,5.613666,6.145606,9.446653,11.314102,8.428044,6.3417826,6.6020937,6.730363,4.52715,3.9574835,3.6934,3.218049,2.8294687,2.8521044,2.7804246,4.1008434,5.8702044,4.727099,5.4438977,8.892077,11.287694,10.567122,6.428553,3.3123648,2.938875,2.7615614,1.9730829,1.5203679,2.886058,5.7192993,7.1566696,6.6058664,5.745708,3.5839937,3.4179983,3.8707132,4.1008434,3.8103511,4.2630663,4.9987283,6.0362,7.8244243,11.261286,12.113899,10.906659,10.895341,12.67602,14.1926155,16.90136,19.1423,18.719765,15.181043,9.835234,7.7225633,8.371455,9.839006,10.472807,8.907167,6.688864,5.4174895,5.6815734,6.964266,7.6395655,5.9305663,5.1156793,5.3344917,6.432326,7.9300575,7.756517,6.511551,5.43258,5.1043615,5.43258,4.2102494,2.9954643,2.7011995,2.7992878,1.3430545,3.2067313,5.6853456,8.495952,10.367173,9.016574,10.529396,11.7894535,12.019584,12.053536,14.366156,14.909414,11.408418,8.228095,7.2698483,7.99042,7.9715567,7.424526,7.9715567,9.978593,12.562841,12.702429,12.755245,12.543978,11.559323,8.971302,8.959985,8.390318,8.884532,10.393582,11.219787,10.604849,9.242931,8.009283,7.435844,7.6923823,6.730363,5.7192993,6.760544,8.858124,7.9451485,4.9987283,4.5120597,4.961002,5.5382137,6.175787,7.039718,5.3910813,3.9197574,4.4139714,7.7942433,7.9225125,5.149633,3.1048703,2.8898308,3.097325,2.1051247,1.4675511,1.2902378,1.3619176,1.146878,1.0638802,1.4713237,1.8334957,1.7995421,1.2147852,1.2185578,1.5731846,1.3392819,0.67152727,0.8224323,0.86770374,0.8903395,0.86770374,0.80356914,0.72811663,1.0186088,1.0336993,0.8526133,0.56589377,0.241448,0.14713238,0.10940613,0.090543,0.071679875,0.071679875,0.10186087,0.08299775,0.090543,0.120724,0.10940613,0.1659955,0.2263575,0.2678564,0.33576363,0.55080324,0.7167987,0.663982,0.59230214,0.6111652,0.72811663,0.69039035,0.56212115,0.4376245,0.40367088,0.5470306,1.237421,1.6109109,3.429316,5.342037,2.916239,3.0256453,1.9240388,0.7922512,0.18863125,0.030181,0.15467763,0.1659955,0.15845025,0.26408374,0.694163,0.6828451,0.9620194,1.1016065,1.0223814,0.995973,0.90920264,0.784706,0.5998474,0.422534,0.4074435,0.3772625,0.38480774,0.38858038,0.38480774,0.4074435,0.51684964,0.84129536,1.1393328,1.1732863,0.724344,0.7205714,0.66775465,0.66020936,0.68661773,0.6451189,0.6187105,0.6451189,0.6413463,0.60362,0.5998474,0.694163,0.73188925,0.77716076,0.80356914,0.724344,0.66775465,0.58475685,0.47912338,0.38103512,0.34330887,0.271629,0.2565385,0.24899325,0.22258487,0.18863125,0.10940613,0.08299775,0.08677038,0.12826926,0.20749438,0.3169005,0.5281675,0.8111144,1.0299267,0.95447415,0.95447415,0.9997456,1.0487897,1.0148361,0.76584285,0.76207024,0.7809334,0.7167987,0.5885295,0.52062225,0.5357128,0.68661773,0.8639311,0.9620194,0.8903395,0.79602385,0.66775465,0.56589377,0.52062225,0.5357128,0.46026024,0.5583485,0.6752999,0.7054809,0.573439,0.6187105,0.663982,0.663982,0.6375736,0.6790725,0.76584285,0.7432071,0.72811663,0.76584285,0.8337501,0.87147635,0.8262049,0.66020936,0.47535074,0.5357128,0.6752999,0.724344,0.69039035,0.63002837,0.63002837,0.66020936,0.77716076,0.95824677,1.1695137,1.3694628,1.2525115,1.327964,1.4826416,1.6637276,1.8561316,1.7165444,1.6373192,1.6373192,1.6788181,1.6863633,1.3317367,1.1431054,0.995973,0.84884065,0.7205714,0.7469798,0.8639311,0.94692886,0.9695646,1.0148361,1.0676528,1.1506506,1.2600567,1.4109617,1.6410918,1.8184053,1.7844516,1.7052265,1.6825907,1.7391801,1.7316349,1.7089992,1.6637276,1.7052265,2.0636258,2.4861598,2.6974268,2.8785129,3.1199608,3.4142256,3.572676,3.6669915,3.5839937,3.350091,3.1048703,2.9954643,3.0369632,3.097325,3.187868,3.429316,3.410453,3.3764994,3.3538637,3.3350005,3.240685,3.308592,3.519859,3.682082,3.7273536,3.7160356,3.7650797,3.7952607,3.8782585,4.055572,4.3611546,4.093298,3.874486,3.7952607,3.904667,4.1989317,4.085753,4.0517993,3.893349,3.6254926,3.4745877,0.120724,0.16222288,0.29803738,0.2867195,0.14713238,0.13958712,0.08677038,0.0754525,0.0754525,0.071679875,0.090543,0.124496624,0.17354076,0.19240387,0.18863125,0.21503963,0.20749438,0.41876137,0.6111652,0.7054809,0.77716076,0.76207024,0.88279426,1.1204696,1.3845534,1.4864142,1.4222796,1.3732355,1.3505998,1.2902378,1.056335,0.9507015,1.1996948,1.3053282,1.1091517,0.80356914,0.27540162,0.06790725,0.0150905,0.00754525,0.00754525,0.090543,0.15467763,0.19240387,0.24899325,0.40367088,0.32444575,0.29426476,0.25276586,0.32444575,0.814887,1.1129243,1.991946,3.1954134,4.647874,6.462507,8.296002,8.82417,7.91874,7.2283497,10.193633,11.434827,11.295239,9.2995205,6.4247804,5.119452,7.4471617,8.952439,11.231105,14.543469,17.810562,17.150352,17.23335,18.546225,19.934551,18.629223,18.319866,16.24115,12.272349,8.099826,7.1906233,6.270103,4.504514,3.1727777,2.7351532,2.8332415,2.8143783,3.4179983,4.6818275,5.8664317,5.492942,5.956975,5.2326307,4.564876,4.5196047,4.9949555,5.372218,5.3986263,5.6287565,5.9230213,5.455216,5.8400235,5.7872066,5.975838,6.439871,6.5643673,5.926794,6.436098,7.3905725,8.152642,8.137552,6.387054,5.7570257,5.4476705,4.983638,4.191386,3.3048196,2.9426475,3.0143273,3.2935016,3.429316,3.229367,3.5802212,3.3312278,2.323937,1.4071891,1.3732355,2.5993385,3.9197574,4.8629136,5.6476197,3.772625,5.304311,7.3377557,7.835742,5.624984,8.001738,9.1825695,8.907167,7.699928,6.8661776,5.100589,3.7198083,3.2331395,3.8669407,5.564622,7.677292,10.480352,12.751472,13.936077,14.169979,15.9695215,16.36942,15.124454,13.109872,12.31762,13.174006,13.019329,14.509516,17.372938,18.414183,18.557543,18.240643,18.591496,19.595015,20.089228,19.953413,19.76101,19.527107,19.866644,22.020813,21.266287,17.112627,13.106099,10.906659,10.253995,7.122716,5.0251365,4.5761943,5.379763,6.013564,6.730363,7.9225125,8.884532,9.623966,10.853842,12.604341,15.196134,18.444365,20.734346,19.025349,16.81459,16.358103,16.18456,16.569368,19.515789,19.968504,20.138271,18.68204,15.471535,11.593277,12.2119875,14.796235,16.078928,14.958458,12.491161,10.944386,9.733373,9.156161,8.933576,8.201687,8.235641,9.205205,10.106862,9.650374,6.2889657,5.8890676,5.330719,4.4705606,3.591539,3.399135,3.6066296,4.5196047,5.402399,5.6287565,4.6629643,5.240176,7.2358947,9.246704,9.993684,8.348819,6.7756343,6.1418333,4.7836885,2.8558772,2.335255,2.3013012,3.2255943,4.8063245,8.307321,16.55428,23.714722,28.430502,28.58518,25.491627,23.869398,19.01403,16.203424,16.897587,18.214233,12.96274,7.8923316,9.235386,10.880251,10.450171,9.318384,10.982111,13.517315,14.252977,12.600568,10.035183,10.748209,13.977575,16.105335,16.414692,17.071129,15.588487,13.513543,12.642066,13.151371,13.607859,12.453435,12.064855,11.155652,10.948157,15.184815,17.923742,21.83218,23.322369,23.32614,27.279852,31.188292,32.844475,33.048195,33.38773,36.243607,36.632187,33.949852,29.456656,24.793692,21.998177,19.56106,17.572887,17.689838,18.629223,16.173243,13.45318,12.66093,13.2607765,13.970031,12.713746,8.443134,6.8850408,9.291975,14.030393,16.550507,12.034674,16.991903,25.05023,30.750666,29.550972,28.781357,22.97906,19.994913,20.69662,19.002712,7.854605,5.3156285,9.291975,15.656394,18.240643,13.098554,9.556059,7.2660756,6.952948,10.416218,10.86516,9.024119,7.375482,7.122716,8.216777,6.417235,5.945657,6.058836,5.617439,3.078462,2.9237845,2.3013012,3.5085413,5.956975,6.149379,6.952948,10.623712,12.721292,11.480098,7.8017883,4.304565,3.9801195,3.4745877,2.0787163,1.7391801,4.538468,7.888559,9.544742,9.484379,9.903141,6.6850915,6.156924,5.7192993,4.617693,3.942393,4.485651,5.6287565,7.914967,11.038701,13.841762,13.143826,11.800771,11.140562,11.721546,13.313594,17.844517,19.942095,18.576405,14.2077055,8.797762,7.1340337,6.149379,6.0286546,6.4474163,6.5530496,5.745708,5.036454,5.119452,5.975838,6.8699503,4.561104,3.893349,4.4403796,5.5193505,6.2021956,6.270103,5.715527,5.1571784,5.149633,6.1833324,5.032682,3.9612563,3.5500402,3.4330888,2.2711203,3.2784111,3.7914882,5.194905,6.8699503,6.2323766,9.1825695,10.344538,10.197406,9.661693,10.087999,13.170234,10.842525,7.2924843,5.0251365,4.847823,4.447925,4.957229,6.126743,7.5603404,8.722309,9.024119,9.937095,10.216269,9.424017,7.9036493,9.167479,9.035437,9.386291,10.506761,11.102836,11.925267,12.08749,11.604594,10.816116,10.370946,8.314865,6.273875,7.1340337,10.250222,11.461235,7.020855,5.5306683,5.1534057,5.142088,5.8211603,7.333983,6.5040054,4.9949555,4.798779,8.239413,10.193633,6.9454026,3.5123138,2.3163917,3.1840954,2.2371666,1.7580433,1.6373192,1.5920477,1.1657411,1.0714256,1.1959221,1.4260522,1.50905,1.056335,0.95824677,1.3656902,1.3015556,0.76207024,0.68661773,0.76584285,0.7205714,0.6790725,0.69039035,0.7432071,0.7884786,0.8601585,0.8865669,0.77338815,0.39989826,0.15467763,0.07922512,0.06790725,0.06413463,0.060362,0.07922512,0.0754525,0.0754525,0.094315626,0.120724,0.1056335,0.16976812,0.25276586,0.32444575,0.38103512,0.543258,0.5281675,0.5017591,0.52062225,0.52062225,0.482896,0.3772625,0.3169005,0.3169005,0.28294688,0.97333723,1.7429527,3.240685,4.8855495,4.8666863,3.6858547,1.9693103,0.7809334,0.34330887,0.02263575,0.03772625,0.06790725,0.071679875,0.12826926,0.47912338,0.6752999,0.8299775,0.94315624,0.9808825,0.8865669,0.68661773,0.6451189,0.5696664,0.45648763,0.48666862,0.36971724,0.32444575,0.3169005,0.30935526,0.26031113,0.3961256,0.7696155,1.1129243,1.1657411,0.65643674,0.90920264,0.84884065,0.7205714,0.66020936,0.6828451,0.6413463,0.663982,0.6451189,0.5772116,0.56589377,0.66775465,0.6526641,0.67152727,0.7432071,0.76584285,0.724344,0.58098423,0.45648763,0.392353,0.34330887,0.24899325,0.21881226,0.19240387,0.15467763,0.14713238,0.094315626,0.08299775,0.09808825,0.16222288,0.31312788,0.43007925,0.55457586,0.814887,1.0978339,1.0638802,0.95824677,0.8865669,0.91674787,0.9507015,0.7167987,0.5696664,0.5885295,0.5772116,0.4979865,0.4376245,0.5696664,0.7507524,0.8941121,0.935611,0.83752275,0.7507524,0.65643674,0.543258,0.4640329,0.5093044,0.43007925,0.46026024,0.573439,0.70170826,0.7507524,0.663982,0.66020936,0.6526641,0.62625575,0.6375736,0.7167987,0.663982,0.7130261,0.88279426,1.0035182,0.7922512,0.69793564,0.60362,0.49421388,0.45648763,0.56212115,0.56212115,0.55457586,0.58475685,0.65643674,0.73188925,0.814887,0.97710985,1.2110126,1.4373702,1.3204187,1.4449154,1.6222287,1.7429527,1.7995421,1.81086,1.7391801,1.6410918,1.5731846,1.5958204,1.2525115,1.1129243,1.0148361,0.9242931,0.9393836,0.9997456,1.1016065,1.1732863,1.2034674,1.20724,1.2525115,1.2298758,1.2449663,1.3543724,1.5807298,1.7882242,1.7882242,1.7391801,1.6939086,1.6033657,1.6071383,1.5807298,1.5543215,1.5958204,1.780679,2.0447628,2.1994405,2.354118,2.5767028,2.867195,3.127506,3.361409,3.3350005,3.1237335,3.1048703,3.1048703,3.0935526,3.0030096,2.9464202,3.2029586,3.2444575,3.2369123,3.2482302,3.2784111,3.259548,3.3048196,3.519859,3.572676,3.4481792,3.440634,3.429316,3.2369123,3.2218218,3.429316,3.62172,3.591539,3.5575855,3.7914882,4.3385186,4.98741,4.979865,4.5837393,4.08198,3.6254926,3.2331395,0.12826926,0.21881226,0.2867195,0.31312788,0.3055826,0.29803738,0.120724,0.09808825,0.090543,0.049044125,0.0,0.06790725,0.150905,0.20749438,0.23767537,0.29049212,0.24522063,0.31312788,0.3734899,0.4074435,0.47535074,0.8224323,1.116697,1.1204696,1.026154,1.4411428,1.6448646,1.5467763,1.4222796,1.3543724,1.2411937,1.1431054,1.2940104,1.2600567,0.8903395,0.32444575,0.1358145,0.033953626,0.0,0.0,0.0,0.0,0.0,0.018863125,0.08677038,0.26408374,0.35085413,0.36971724,0.35462674,0.3470815,0.3734899,1.0714256,2.8521044,4.636556,5.455216,4.447925,4.0517993,3.802806,3.4179983,4.221567,9.171251,11.593277,11.672502,9.329701,6.2021956,5.643847,8.597813,11.272603,14.7321005,17.810562,17.1164,14.93205,15.264041,17.127718,18.8254,17.935059,18.206688,13.837989,9.646602,7.8432875,8.069645,6.2663302,4.561104,3.2859564,2.6634734,2.806833,2.1202152,1.6184561,2.3163917,3.9725742,5.093044,5.534441,5.0213637,4.5912848,4.4743333,4.115934,3.8367596,3.663219,4.134797,4.8855495,4.6214657,4.06689,3.8480775,4.447925,5.572167,6.1644692,6.749226,7.960239,8.3525915,7.7640624,7.322665,6.2097406,6.0324273,6.047518,5.4665337,3.4594972,1.9051756,1.4562333,1.7655885,2.4786146,3.218049,4.13857,4.508287,3.9310753,2.6597006,1.6109109,1.7769064,1.9278114,2.2371666,2.655928,2.9237845,2.2899833,3.6254926,4.738417,4.4101987,2.4031622,5.8211603,8.371455,8.405409,6.375736,4.847823,4.617693,3.8141239,3.6292653,4.564876,6.4549613,8.22055,10.676529,13.147598,15.184815,16.561823,18.599041,17.297485,13.800262,9.831461,7.7037,8.544995,9.533423,13.185325,18.074646,18.806536,19.681786,18.206688,17.80679,18.919714,18.953669,18.99894,17.89356,17.40689,18.542452,21.541689,19.266796,13.615403,8.75249,6.6322746,6.9869013,5.987156,5.2590394,5.855114,7.0585814,6.356873,6.5756855,7.4999785,8.443134,9.548513,11.774363,12.513797,15.414946,19.836462,22.960196,19.810055,15.562078,13.59654,13.762536,15.98084,20.217497,22.266033,21.78691,19.61765,16.237377,11.751727,12.842015,15.082954,15.633758,14.022847,12.1101265,10.668983,8.899622,7.888559,8.028146,9.039209,10.076681,10.148361,9.684328,8.5563135,6.092789,6.145606,5.643847,4.908185,4.2404304,3.92353,3.5500402,5.111907,6.19465,5.511805,2.897376,3.7273536,5.9720654,8.4544525,10.329447,11.076427,11.00852,9.529651,6.488915,3.4557245,3.7462165,3.5575855,3.187868,4.055572,6.700182,10.767072,17.591751,24.442837,28.928488,30.471493,30.32436,20.832436,18.097282,16.976812,15.667711,15.724301,8.737399,7.8131065,9.239159,10.284176,9.1825695,10.623712,15.4074,18.263277,17.014538,12.608112,10.989656,13.936077,17.191853,19.112118,20.673985,18.259504,16.003475,15.448899,15.663939,13.264549,11.793225,13.109872,13.328684,12.325166,13.728582,17.980331,22.269806,24.401339,25.231316,28.649315,33.45564,36.21343,38.42796,40.94807,43.99258,43.23051,40.48404,37.198082,33.949852,30.456402,24.669195,21.662413,20.270313,19.138527,16.74291,14.079436,13.030646,13.328684,13.807808,12.415709,9.80128,7.111398,9.669238,16.452417,20.085455,11.981857,17.784155,28.219234,32.735065,19.527107,25.5369,21.375692,20.568352,22.499935,12.423254,8.039464,7.8696957,12.261031,17.840744,17.497435,6.5002327,9.273112,10.453944,7.032173,8.382772,14.596286,12.385528,8.495952,6.258785,5.583485,7.3113475,7.8319697,8.431817,8.201687,4.0103,3.3840446,2.4220252,1.7278622,2.0787163,4.395108,7.201941,13.585222,16.77309,14.849052,10.729345,4.9421387,5.5193505,5.2628117,2.6634734,1.8938577,6.198423,9.473062,10.510533,10.578441,13.422999,10.657665,9.374973,7.1868505,4.4894238,4.4630156,4.2064767,4.9534564,7.809334,11.747954,13.592768,11.989402,11.732863,11.819634,11.721546,11.355601,14.928277,17.471025,16.131744,11.242422,6.3342376,6.643593,5.9682927,5.070408,4.6629643,5.372218,6.5643673,6.0550632,5.534441,5.994701,7.745199,5.3458095,3.7914882,3.5764484,4.2328854,4.327201,5.3609,5.6061206,5.617439,6.1041074,7.9225125,6.0248823,5.3458095,4.8138695,4.164978,3.9273026,3.6292653,3.7198083,4.0593443,4.1989317,3.3425457,6.1078796,7.0057645,7.0887623,7.118943,7.5603404,12.792972,10.993429,7.4471617,5.247721,5.27413,4.217795,3.9725742,4.715781,5.8890676,6.187105,5.3156285,5.3269467,5.3156285,5.3458095,6.458734,8.099826,8.733627,9.635284,10.899114,11.457462,13.4644985,14.388792,14.109617,12.826925,11.09529,8.265821,6.560595,6.820906,9.208978,13.241914,9.133525,6.9944468,5.670255,4.881777,5.2062225,6.2927384,6.590776,5.2892203,3.983892,6.7039547,11.042474,8.718536,4.82896,2.5804756,3.2972744,2.3918443,2.1202152,2.0372176,1.8372684,1.358145,1.2902378,1.086516,1.0186088,1.0940613,1.0638802,0.845068,1.388326,1.5015048,0.9808825,0.5998474,0.633801,0.5357128,0.5055317,0.6413463,0.9205205,0.76584285,0.694163,0.73566186,0.7884786,0.6149379,0.2678564,0.116951376,0.0754525,0.071679875,0.056589376,0.06413463,0.06790725,0.06790725,0.0754525,0.1056335,0.090543,0.12826926,0.22258487,0.30935526,0.23013012,0.3772625,0.41876137,0.452715,0.47912338,0.3734899,0.24522063,0.2263575,0.23013012,0.19994913,0.10186087,0.6073926,1.9655377,3.3350005,4.7874613,7.322665,4.504514,1.9806281,0.7205714,0.56589377,0.23390275,0.23390275,0.10940613,0.02263575,0.041498873,0.14335975,0.58475685,0.6752999,0.79602385,0.98465514,0.9205205,0.5885295,0.56212115,0.543258,0.4678055,0.5017591,0.36594462,0.30181,0.31312788,0.35085413,0.30935526,0.34330887,0.58475685,0.73188925,0.6752999,0.5017591,1.0299267,1.0072908,0.784706,0.6187105,0.6488915,0.6111652,0.633801,0.62625575,0.5772116,0.5583485,0.66020936,0.62625575,0.6149379,0.6752999,0.73566186,0.784706,0.6451189,0.51684964,0.44894236,0.36594462,0.27917424,0.22258487,0.17731337,0.14335975,0.14335975,0.116951376,0.11317875,0.150905,0.24522063,0.39989826,0.4640329,0.5696664,0.76207024,0.9922004,1.1091517,0.995973,0.8563859,0.7884786,0.7922512,0.754525,0.60362,0.5017591,0.3961256,0.31312788,0.3772625,0.5772116,0.8111144,0.91674787,0.845068,0.6526641,0.663982,0.62248313,0.513077,0.4074435,0.4376245,0.48666862,0.49044126,0.51684964,0.62625575,0.87147635,0.63002837,0.56589377,0.5696664,0.55457586,0.49044126,0.573439,0.59230214,0.7167987,0.9393836,1.0751982,0.77338815,0.73566186,0.69039035,0.55080324,0.39989826,0.331991,0.32444575,0.41498876,0.5583485,0.60362,0.79602385,0.8941121,1.0638802,1.327964,1.5543215,1.4147344,1.4298248,1.5052774,1.5958204,1.6788181,1.8485862,1.7618159,1.4750963,1.1317875,0.935611,0.9997456,1.0450171,1.0487897,1.0789708,1.2864652,1.3392819,1.3505998,1.358145,1.3770081,1.388326,1.3996439,1.2751472,1.2298758,1.3392819,1.5165952,1.7052265,1.7957695,1.780679,1.6788181,1.5316857,1.5580941,1.5430037,1.5052774,1.4901869,1.5580941,1.750498,1.9089483,2.0485353,2.2069857,2.4371157,2.6936543,2.987919,3.048281,2.9464202,3.1048703,3.187868,3.1124156,2.987919,2.9351022,3.0445085,3.2784111,3.3048196,3.229367,3.199186,3.3878171,3.240685,3.4330888,3.3878171,3.0822346,3.0218725,3.2218218,3.0709167,2.8936033,2.8256962,2.8256962,2.9803739,3.1425967,3.663219,4.557331,5.5004873,5.828706,5.3873086,4.6931453,3.9914372,3.2142766,0.090543,0.056589376,0.056589376,0.060362,0.06790725,0.090543,0.17731337,0.150905,0.071679875,0.0,0.0,0.0,0.03772625,0.09808825,0.181086,0.29049212,0.21503963,0.181086,0.29426476,0.5357128,0.73188925,0.9507015,0.68661773,0.4678055,0.5357128,0.8563859,1.478869,1.8900851,1.6825907,1.0110635,0.59607476,0.935611,1.0487897,0.77338815,0.2867195,0.090543,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.0452715,0.08299775,0.18485862,0.24522063,0.3470815,0.76207024,1.8749946,4.274384,6.5756855,7.496206,5.873977,1.4562333,0.633801,1.6524098,3.482133,5.8136153,9.9257765,8.492179,6.7341356,6.790725,7.7037,8.571404,10.884023,11.796998,10.819888,9.842778,12.344029,13.034419,11.155652,8.36391,8.744945,9.024119,8.269594,8.099826,8.458225,7.6282477,5.1043615,4.425289,3.6669915,2.3201644,1.2826926,1.6976813,1.4071891,2.505023,4.2630663,3.127506,2.6031113,5.1081343,7.145352,7.009537,4.776143,2.9954643,2.897376,4.2328854,6.2436943,7.6584287,5.4250345,3.7047176,2.7238352,2.3805263,2.2598023,3.270866,3.663219,4.5950575,6.2851934,7.9941926,6.8737226,6.0626082,5.3269467,4.22534,2.0900342,1.1619685,1.4600059,1.5052774,1.327964,2.4861598,4.244203,4.08198,2.9200118,1.7467253,1.5882751,1.4901869,1.6033657,1.4864142,1.0676528,0.6413463,1.0299267,1.569412,2.4484336,3.3161373,3.2821836,6.5530496,8.311093,7.752744,5.553304,3.904667,5.247721,5.27413,4.7044635,5.247721,9.567377,11.521597,13.573905,17.139036,21.420965,23.420456,23.752447,20.813572,16.795727,14.2077055,15.8676605,16.724047,16.26756,15.494171,14.449154,12.253486,15.109364,15.660167,16.531643,17.512526,15.55076,16.98813,15.656394,12.683565,9.64283,8.529905,11.057564,8.986393,6.779407,6.2399216,6.5455046,5.753253,6.779407,7.77538,7.5037513,5.3571277,5.772116,6.3342376,7.7301087,9.7220545,11.140562,11.076427,14.320885,18.010511,20.357084,20.673985,15.120681,12.019584,12.96274,16.116653,16.252468,14.7736,15.230087,15.033911,13.521088,11.947904,12.815607,13.517315,12.479843,10.438853,10.438853,9.386291,8.235641,7.6622014,8.416726,11.321648,13.970031,12.162943,9.348565,7.2283497,5.753253,5.3269467,4.3686996,3.9876647,4.315883,4.485651,3.5462675,4.8025517,6.221059,6.228604,3.7386713,4.9723196,6.221059,8.035691,11.676274,19.134754,9.307066,3.9499383,2.4371157,3.6745367,6.1041074,5.2628117,4.776143,5.2137675,5.994701,5.372218,10.155907,20.598532,26.73282,26.091475,23.695858,24.220253,21.900087,18.534906,15.663939,14.543469,10.023865,6.3417826,5.7607985,7.4018903,7.2170315,9.488152,12.593022,15.380992,17.18808,17.82188,12.596795,14.652876,18.28214,21.28515,24.94837,21.322876,18.372684,16.957949,16.780636,16.403374,15.241405,14.916959,14.305794,13.249459,12.543978,18.244415,21.73032,24.280615,26.219744,26.917679,30.237589,35.74562,39.68047,40.52554,39.001396,39.72197,40.680214,37.55648,31.663641,29.969732,27.110083,26.068838,25.687803,25.042685,23.405365,19.56106,15.818617,13.615403,12.257258,8.91094,11.072655,7.5112963,5.66271,7.533932,9.7220545,11.502733,37.873383,43.543636,23.273323,11.872451,11.751727,17.799244,23.963715,23.643042,9.688101,10.140816,11.1782875,10.970794,9.548513,8.805306,4.214022,6.7379084,8.503497,7.5037513,7.6131573,16.014793,13.324911,8.118689,5.240176,5.8136153,9.378746,9.390063,8.45068,7.3188925,4.9119577,3.2520027,3.1237335,2.516341,1.4901869,2.1353056,2.2107582,16.52787,29.796192,32.42194,20.50799,6.4549613,6.488915,6.8661776,3.3953626,1.418507,3.2142766,4.8063245,7.4999785,10.997202,13.411682,14.475562,12.030901,7.6584287,3.802806,3.7537618,2.4823873,3.0633714,5.5797124,8.744945,9.918231,8.744945,9.26934,10.152134,10.231359,8.499724,10.438853,11.457462,10.393582,8.043237,7.141579,9.276885,9.654147,8.062099,5.8098426,5.7381625,9.314611,8.552541,7.0359454,6.8925858,8.7600355,10.638803,6.651138,3.6179473,3.6066296,3.9386206,5.7796617,5.847569,6.1833324,7.4811153,9.0957985,6.7869525,5.836251,5.1873593,4.67051,4.991183,4.183841,6.300284,5.692891,2.1956677,1.0827434,2.2673476,2.425798,4.036709,7.7338815,12.298758,14.569878,10.804798,8.469543,10.269085,14.173752,10.291721,7.77538,7.032173,7.3113475,6.7152724,3.4179983,2.4220252,2.2183034,3.0520537,6.8963585,6.360646,7.250985,10.265312,13.664448,13.275867,12.664702,11.706455,9.367428,6.470052,5.6778007,5.43258,5.0138187,4.738417,5.3458095,7.9791017,8.480861,7.84706,6.3153744,4.4139714,2.9615107,3.9008942,4.859141,4.395108,3.078462,3.4934506,9.597558,9.329701,6.1116524,3.2972744,4.164978,3.0897799,2.384299,2.04099,1.991946,2.0900342,1.7467253,1.20724,0.935611,0.98842776,0.97710985,0.86770374,1.3430545,1.4939595,1.0299267,0.26031113,0.43007925,0.47157812,0.47157812,0.60362,1.1280149,0.83752275,0.5998474,0.543258,0.663982,0.80734175,0.6375736,0.31312788,0.1056335,0.071679875,0.0452715,0.033953626,0.030181,0.030181,0.033953626,0.0452715,0.056589376,0.08677038,0.181086,0.2678564,0.18485862,0.3169005,0.48666862,0.55080324,0.482896,0.3961256,0.29803738,0.26408374,0.28294688,0.28294688,0.1358145,0.36971724,1.7278622,3.5651307,5.613666,7.9791017,5.270357,2.897376,1.4034165,0.87147635,0.9318384,0.88279426,0.392353,0.05281675,0.02263575,0.0452715,0.4376245,0.73566186,1.0336993,1.2034674,0.8865669,0.543258,0.4376245,0.44516975,0.45648763,0.38103512,0.38103512,0.3734899,0.35839936,0.38103512,0.5017591,0.331991,0.20749438,0.1659955,0.19994913,0.26031113,0.44139713,0.56212115,0.6111652,0.6149379,0.62625575,0.5772116,0.58475685,0.5885295,0.5696664,0.5357128,0.754525,0.83752275,0.7884786,0.6488915,0.5017591,0.6488915,0.7054809,0.6375736,0.5017591,0.42630664,0.34330887,0.24899325,0.18485862,0.1659955,0.1659955,0.181086,0.19240387,0.29049212,0.41121614,0.35085413,0.4376245,0.66775465,0.80356914,0.84129536,1.0374719,0.9507015,0.9205205,0.8601585,0.72811663,0.5357128,0.65643674,0.55080324,0.43385187,0.42630664,0.55080324,0.573439,0.7167987,0.80356914,0.7507524,0.58098423,0.543258,0.47912338,0.43007925,0.42630664,0.48666862,0.58475685,0.70170826,0.73188925,0.72811663,0.8865669,0.69039035,0.60362,0.5357128,0.45648763,0.38103512,0.5017591,0.48666862,0.49421388,0.58475685,0.73188925,0.5998474,0.5281675,0.45648763,0.3772625,0.35085413,0.31312788,0.3772625,0.543258,0.69039035,0.58098423,0.8601585,1.0299267,1.1732863,1.3317367,1.5430037,1.4298248,1.4675511,1.4939595,1.5203679,1.7391801,1.5203679,1.4637785,1.3619176,1.1053791,0.70170826,0.935611,1.0940613,1.2562841,1.3694628,1.237421,1.1242423,1.1091517,1.1016065,1.1091517,1.20724,1.3166461,1.4600059,1.539231,1.4939595,1.297783,1.7014539,1.8749946,1.8259505,1.6788181,1.6788181,1.7165444,1.6788181,1.5920477,1.50905,1.4939595,1.5920477,1.7165444,1.8033148,1.9240388,2.305074,2.41448,2.4974778,2.4974778,2.493705,2.7011995,2.8332415,3.0331905,3.4255435,3.8141239,3.6934,3.742444,3.5802212,3.3048196,3.169005,3.5689032,3.180323,3.229367,3.187868,2.9841464,3.0218725,3.1425967,3.1539145,2.8747404,2.4484336,2.3503454,2.546522,2.9426475,3.3953626,3.7047176,3.6330378,4.1083884,5.372218,5.945657,5.300538,3.8593953,0.12826926,0.13204187,0.16976812,0.16976812,0.14713238,0.19994913,0.18863125,0.090543,0.060362,0.116951376,0.14713238,0.030181,0.00754525,0.08299775,0.21503963,0.32821837,0.331991,0.2867195,0.29049212,0.35085413,0.3772625,0.34330887,0.5055317,0.7507524,0.8978847,0.7092535,1.2902378,1.4901869,1.056335,0.331991,0.23013012,0.49421388,0.5772116,0.44894236,0.19994913,0.056589376,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.033953626,0.049044125,0.060362,0.094315626,0.23013012,0.56589377,0.995973,3.5424948,7.54525,9.876732,4.9345937,1.7354075,2.9351022,5.198677,6.571913,6.458734,4.979865,3.9688015,3.5689032,3.7084904,4.104616,3.8178966,3.9989824,4.0404816,3.9461658,4.3385186,7.2396674,8.571404,7.696155,5.9984736,6.862405,10.114408,10.121953,7.914967,5.1043615,3.893349,2.7728794,2.3163917,2.384299,2.8294687,3.4896781,4.9987283,4.696918,3.3878171,2.3390274,3.2746384,2.886058,3.1124156,3.3010468,3.229367,3.1048703,2.474842,2.252257,2.637065,3.2784111,3.2784111,2.8596497,3.0218725,3.199186,3.1124156,2.746471,2.7238352,2.3163917,2.0975795,2.4182527,3.3953626,3.5689032,4.1800685,4.5309224,4.3875628,3.9688015,3.5877664,3.6443558,3.2633207,2.4522061,2.1088974,2.7728794,2.4069347,1.9579924,1.8184053,1.8561316,2.022127,2.3918443,2.6068838,2.4899325,2.0447628,2.173032,2.071171,1.9051756,1.9730829,2.7200627,4.7120085,7.0548086,8.13378,7.7112455,6.9227667,8.99771,9.548513,10.235131,11.604594,13.083464,15.912932,19.066847,23.065828,26.385738,25.450129,26.695095,25.370903,23.80149,22.469755,20.017548,18.51227,18.014284,16.248695,13.88326,14.547242,16.720274,18.776354,18.02183,15.55076,16.218515,15.422491,12.917468,9.81637,7.4207535,7.1981683,8.22055,6.115425,4.5497856,4.776143,5.617439,6.2097406,7.1340337,7.322665,6.8133607,6.7341356,5.4703064,5.1798143,5.5268955,6.643593,9.110889,9.265567,11.16697,13.70972,15.577168,15.230087,14.803781,12.200669,11.902632,14.053028,14.479335,14.166207,15.350811,16.086473,15.856343,15.562078,14.396337,12.619431,11.457462,11.476325,12.596795,10.257768,9.205205,10.680302,14.124708,17.157898,16.652367,13.072145,9.491924,7.594294,7.6697464,9.175024,7.284939,6.4964604,7.4584794,6.964266,6.530414,10.442626,13.226823,11.834724,5.643847,5.832478,6.7680893,8.224322,9.590013,9.869187,4.7610526,6.8359966,6.858632,3.7613072,4.640329,6.7944975,7.2698483,7.122716,7.141579,7.84706,8.952439,14.241659,19.90437,22.960196,21.281378,22.167944,19.493153,15.814844,13.20796,13.298503,10.303039,7.043491,5.7192993,6.3644185,6.8774953,8.52236,10.518079,11.800771,13.607859,19.444109,16.105335,15.252723,16.542961,20.006231,26.057522,23.8279,20.617395,17.999193,16.59955,16.086473,18.980076,18.670721,17.199398,15.743164,14.603831,18.293459,20.50799,22.711203,25.125683,26.710184,29.34725,34.843964,39.661606,41.072567,37.18299,38.880672,38.941036,35.855026,31.429739,30.799711,30.294178,28.000423,26.034885,24.307022,20.515535,19.01403,17.025856,14.758509,12.264804,9.446653,12.47607,8.83926,7.273621,10.054046,12.989148,10.487898,18.02183,18.304777,10.242677,8.929804,7.3415284,12.593022,15.00373,12.200669,9.125979,6.228604,6.300284,6.515323,7.009537,10.842525,8.431817,6.56814,6.405917,6.9189944,4.927048,6.7756343,7.1340337,8.650629,11.174516,11.759273,12.577931,8.171506,7.575431,10.461489,7.111398,3.7009451,3.3915899,2.8747404,1.8221779,2.8822856,3.6481283,6.5756855,11.619685,17.87847,23.620405,11.121698,6.156924,5.05909,4.927048,3.651901,4.236658,6.156924,8.341274,9.9257765,10.26154,9.420244,7.2924843,4.5120597,2.173032,1.7995421,1.116697,1.1619685,2.493705,4.9534564,7.647111,7.677292,6.9189944,6.56814,7.069899,8.107371,10.001229,10.895341,10.729345,10.020092,9.839006,10.921749,10.521852,8.929804,7.2887115,7.61693,9.435335,8.612903,8.254503,9.703192,12.566614,12.151625,10.11818,8.929804,9.469289,11.042474,10.287949,9.046755,8.088508,8.043237,9.4127,7.122716,6.9755836,6.360646,5.191132,5.8702044,4.9647746,5.8098426,5.873977,4.738417,4.085753,5.349582,3.9008942,4.436607,8.477088,14.347293,14.958458,12.494934,9.74469,8.439363,9.280658,8.258276,7.643338,8.68081,10.559577,10.412445,6.1795597,4.4177437,3.6330378,3.5953116,5.3609,6.1795597,6.911449,8.416726,10.012547,9.454198,7.4471617,6.617184,5.300538,3.4934506,2.8558772,4.447925,4.5120597,3.8065786,3.6368105,5.8437963,6.900131,6.515323,5.3948536,3.9574835,2.3390274,2.4182527,3.4896781,3.3689542,2.3088465,3.006782,6.8925858,8.428044,7.3000293,4.678055,3.2029586,2.6446102,2.1466236,1.8372684,1.8184053,2.1503963,2.003264,1.569412,1.4335974,1.6146835,1.5618668,1.1506506,1.3015556,1.3656902,1.0789708,0.56589377,0.69793564,0.79602385,0.76584285,0.7432071,1.0940613,0.965792,0.8111144,0.7469798,0.80734175,0.94315624,0.76207024,0.43385187,0.19994913,0.14335975,0.1659955,0.06790725,0.033953626,0.02263575,0.00754525,0.02263575,0.05281675,0.05281675,0.0754525,0.11317875,0.08677038,0.150905,0.33576363,0.3961256,0.35839936,0.5055317,0.44894236,0.32821837,0.27540162,0.26408374,0.1358145,0.1358145,0.56212115,1.5015048,3.308592,6.6247296,9.627739,7.250985,3.6896272,1.7052265,2.6144292,3.6783094,2.1503963,0.58098423,0.0150905,0.02263575,0.35462674,0.6149379,0.7696155,0.8337501,0.8978847,0.83752275,0.7469798,0.7394345,0.7167987,0.38103512,0.41121614,0.39989826,0.41498876,0.452715,0.4678055,0.36594462,0.33576363,0.29049212,0.241448,0.32067314,0.38480774,0.482896,0.5357128,0.543258,0.56589377,0.58475685,0.5998474,0.59230214,0.5583485,0.52062225,0.6451189,0.7394345,0.77338815,0.724344,0.5772116,0.73188925,0.80356914,0.724344,0.55080324,0.48666862,0.38480774,0.24899325,0.15845025,0.12826926,0.120724,0.150905,0.21881226,0.35462674,0.49421388,0.47157812,0.5093044,0.56212115,0.6451189,0.7507524,0.8186596,0.76207024,0.80356914,0.7696155,0.6111652,0.422534,0.4678055,0.4678055,0.482896,0.543258,0.633801,0.6488915,0.7394345,0.7130261,0.573439,0.52062225,0.65643674,0.6828451,0.663982,0.66020936,0.7205714,0.72811663,0.7432071,0.7054809,0.68661773,0.8865669,0.77716076,0.68661773,0.65643674,0.6413463,0.49044126,0.48666862,0.47535074,0.43385187,0.39989826,0.48666862,0.5093044,0.60362,0.6375736,0.5772116,0.48666862,0.4979865,0.56589377,0.70170826,0.8262049,0.77338815,0.8299775,0.87147635,0.90543,1.0110635,1.3468271,1.4109617,1.478869,1.4147344,1.2600567,1.2147852,1.3958713,1.3807807,1.2298758,1.056335,1.0450171,0.935611,0.8299775,0.8111144,0.875249,0.95447415,1.177059,1.0827434,1.0751982,1.2298758,1.2789198,1.3091009,1.3732355,1.4600059,1.5618668,1.6524098,1.7429527,1.8070874,1.8674494,1.9655377,2.1805773,1.9429018,1.961765,2.033445,2.0485353,2.0070364,2.173032,2.2371666,2.1013522,1.9127209,2.0372176,2.2220762,2.3616633,2.4974778,2.6144292,2.6144292,2.7691069,3.0369632,3.4670424,3.8367596,3.6556737,3.7348988,3.9159849,3.92353,3.7990334,3.8895764,3.4179983,3.270866,3.1916409,3.0709167,2.9615107,2.8106055,2.5201135,2.252257,2.1013522,2.082489,2.2484846,2.5767028,3.1312788,3.6669915,3.6443558,3.874486,5.028909,5.5268955,4.9760923,4.142342,0.12826926,0.14713238,0.14335975,0.120724,0.1056335,0.12826926,0.11317875,0.08299775,0.090543,0.12826926,0.1358145,0.06413463,0.06790725,0.116951376,0.17354076,0.181086,0.26408374,0.27917424,0.26408374,0.2678564,0.33576363,0.392353,0.5357128,0.6828451,0.70170826,0.41498876,0.7394345,0.7167987,0.43007925,0.09808825,0.08299775,0.20372175,0.23767537,0.19240387,0.094315626,0.018863125,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.02263575,0.018863125,0.02263575,0.049044125,0.14713238,0.39989826,0.694163,2.6898816,6.7039547,9.582467,4.719554,1.3920987,2.7841973,5.8136153,7.6207023,5.5495315,2.7653341,2.5389767,2.7804246,2.5389767,2.022127,1.7882242,1.5505489,1.6146835,1.9391292,2.1353056,3.361409,4.1498876,4.172523,3.9008942,4.6252384,6.4926877,8.088508,7.809334,6.047518,5.1571784,3.3425457,2.5276587,2.2409391,2.493705,3.7688525,4.459243,4.7535076,4.3686996,4.063117,5.6551647,4.7648253,3.150142,2.1994405,2.4333432,3.5085413,2.9766011,2.444661,2.2371666,2.233394,1.8448136,1.8297231,2.3805263,2.8407867,3.0030096,3.1237335,2.4484336,2.0145817,2.0598533,2.5729303,3.2784111,4.3875628,4.927048,4.930821,4.640329,4.504514,2.9426475,2.7011995,2.6974268,2.3654358,1.6373192,1.8749946,1.7844516,1.5958204,1.5769572,2.04099,2.5502944,2.8181508,2.7426984,2.795515,4.006528,5.7079816,5.9192486,4.8629136,3.712263,4.5912848,6.6322746,9.529651,11.819634,12.649611,11.778135,11.114153,10.751981,12.23085,14.713238,15.015047,15.965749,18.72731,22.782883,26.461191,26.962952,31.410875,34.874146,35.88521,33.376415,26.706413,23.280869,21.337967,18.874443,16.573141,17.82188,18.270823,18.161417,16.848543,15.033911,14.777372,14.045483,11.197151,8.080963,6.405917,7.7187905,7.8810134,6.5002327,4.727099,3.5877664,3.99521,5.168496,6.4964604,7.677292,8.348819,8.07719,6.590776,5.6589375,5.379763,5.772116,6.7944975,7.0359454,8.3525915,9.997457,11.555551,12.917468,13.230596,12.73261,12.694883,13.249459,13.358865,15.641303,16.720274,16.822134,16.675003,17.48989,14.864142,12.1101265,10.910432,11.434827,12.332711,12.298758,13.43809,16.403374,20.96825,26.004704,21.632233,14.600059,9.786189,8.835487,10.170997,11.25374,9.009028,7.4509344,8.043237,9.688101,11.910177,17.08999,18.602814,14.151116,5.753253,5.692891,6.4926877,8.024373,9.2844305,8.375228,5.5306683,7.281166,6.820906,4.0178456,5.406172,8.488406,9.224068,9.476834,9.906913,9.933322,8.7600355,11.18206,17.463482,24.838963,27.506208,26.049976,20.88148,15.878979,13.038192,12.453435,10.295494,7.1868505,5.7909794,6.4964604,7.413208,9.590013,12.649611,13.29473,12.442118,15.218769,16.373192,15.660167,15.705438,17.91997,22.537663,22.488617,21.202152,19.180025,17.444618,17.56157,22.349031,21.337967,19.794964,19.300749,17.784155,19.821371,22.99415,25.227543,26.185791,27.287397,28.562544,31.765503,33.78763,33.953625,34.03662,36.224747,36.82082,35.221226,33.02933,34.06303,30.94307,27.2044,25.921707,25.359585,18.976303,17.512526,16.101564,14.18507,11.966766,10.416218,10.412445,10.084227,12.408164,15.618668,13.215506,10.759526,11.5857315,10.212496,6.7756343,7.032173,13.12119,14.128481,12.951422,11.136789,8.8769865,5.0779533,3.99521,3.6858547,4.2404304,7.8017883,8.45068,8.0206,7.432071,6.6549106,4.7044635,5.1835866,6.983129,10.306811,13.117417,11.140562,10.789707,7.1604424,5.9682927,7.6093845,7.1566696,3.3764994,2.5201135,2.3767538,2.1353056,2.3805263,3.7537618,5.481624,10.457717,17.244669,20.104319,13.788944,9.7220545,7.3679366,5.9494295,4.4403796,4.2517486,5.2590394,7.3490734,8.726082,5.915476,6.156924,6.802043,6.6247296,5.0779533,2.282438,0.8224323,0.543258,1.4939595,3.682082,7.043491,9.797507,8.465771,6.0776987,4.9647746,6.7567716,10.446399,14.143571,14.57365,12.3893,12.196897,13.045737,12.751472,11.921495,11.072655,10.661438,10.589758,8.75249,8.692128,11.11038,13.8870325,13.841762,12.691111,11.796998,11.9064045,13.128735,12.185578,10.589758,9.250477,8.60913,8.650629,7.6093845,7.624475,6.851087,5.7570257,7.1038527,4.930821,5.383536,6.3153744,6.5228686,5.7419353,7.069899,5.3948536,4.7648253,6.8925858,11.18206,14.109617,12.808062,9.258021,5.907931,5.666483,5.7872066,6.515323,8.156415,9.948412,10.072908,8.243186,6.387054,4.515832,3.2972744,4.06689,6.255012,6.9454026,7.99042,9.1825695,8.262049,5.240176,5.0515447,4.961002,3.8292143,2.123988,3.802806,4.142342,3.7575345,3.429316,4.13857,4.425289,4.29702,4.0103,3.5689032,2.7125173,2.2711203,3.0105548,3.2255943,2.6597006,2.4899325,4.930821,6.8737226,6.8850408,4.991183,2.686109,2.2447119,1.931584,1.720317,1.6675003,1.9089483,1.8787673,1.5241405,1.3920987,1.5430037,1.5731846,1.0978339,1.1280149,1.20724,1.0450171,0.513077,0.52439487,0.754525,0.875249,0.88279426,1.1016065,0.9808825,0.88279426,0.875249,0.95447415,1.0676528,0.9507015,0.6526641,0.3470815,0.16222288,0.20749438,0.17354076,0.094315626,0.033953626,0.00754525,0.00754525,0.026408374,0.02263575,0.02263575,0.041498873,0.05281675,0.056589376,0.17731337,0.23013012,0.22258487,0.34330887,0.5055317,0.392353,0.26408374,0.23013012,0.23767537,0.1056335,0.13958712,0.5696664,1.6750455,3.7688525,6.647365,6.85486,5.349582,3.3915899,2.5502944,3.0822346,1.8900851,0.6375736,0.06790725,0.02263575,0.2263575,0.4979865,0.663982,0.724344,0.8526133,0.9016574,0.8941121,0.8186596,0.6526641,0.392353,0.41876137,0.48666862,0.5394854,0.51684964,0.32067314,0.2565385,0.26408374,0.271629,0.28294688,0.392353,0.392353,0.47912338,0.58098423,0.6375736,0.59607476,0.543258,0.5470306,0.58475685,0.63002837,0.63002837,0.59607476,0.6828451,0.8865669,1.026154,0.7432071,0.84129536,0.91297525,0.8186596,0.59230214,0.45648763,0.35462674,0.24899325,0.18485862,0.1659955,0.16222288,0.19240387,0.29426476,0.3961256,0.46026024,0.47535074,0.5583485,0.59230214,0.6187105,0.67152727,0.7432071,0.66020936,0.6488915,0.6488915,0.62625575,0.5998474,0.58475685,0.47912338,0.46026024,0.55080324,0.63002837,0.68661773,0.7507524,0.69039035,0.5394854,0.49421388,0.6111652,0.663982,0.66775465,0.6752999,0.7582976,0.9318384,0.95824677,0.875249,0.7696155,0.80356914,0.7394345,0.7092535,0.66775465,0.5772116,0.4376245,0.43007925,0.44894236,0.43385187,0.3961256,0.4074435,0.45648763,0.59230214,0.633801,0.5470306,0.44516975,0.543258,0.58098423,0.70170826,0.9016574,1.026154,0.9507015,0.935611,0.9620194,1.0336993,1.1959221,1.2751472,1.2562841,1.1053791,0.9393836,0.9922004,1.3015556,1.2713746,1.0487897,0.814887,0.7922512,0.76207024,0.7696155,0.724344,0.633801,0.5998474,0.7884786,0.8299775,0.8941121,1.0072908,1.0487897,1.1053791,1.20724,1.3543724,1.5241405,1.6863633,1.901403,1.8561316,1.7731338,1.8146327,2.082489,1.9542197,1.9881734,2.082489,2.1277604,1.9994912,1.9466745,1.8749946,1.780679,1.6939086,1.6750455,1.81086,1.9504471,2.0598533,2.1503963,2.3013012,2.6634734,3.029418,3.3689542,3.5689032,3.4557245,3.6443558,3.9876647,4.13857,4.085753,4.142342,3.7613072,3.4179983,3.127506,2.8709676,2.6068838,2.505023,2.233394,1.9730829,1.8372684,1.8599042,2.0183544,2.2748928,2.71629,3.2784111,3.7575345,4.244203,5.032682,5.2628117,4.8063245,4.274384,0.32444575,0.19240387,0.124496624,0.09808825,0.090543,0.060362,0.07922512,0.08677038,0.08299775,0.08299775,0.11317875,0.116951376,0.1358145,0.15467763,0.14335975,0.08677038,0.181086,0.2565385,0.2867195,0.29803738,0.3734899,0.45648763,0.44894236,0.43007925,0.39989826,0.2678564,0.35085413,0.2263575,0.10940613,0.07922512,0.071679875,0.06413463,0.06413463,0.05281675,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.00754525,0.0150905,0.00754525,0.0150905,0.026408374,0.11317875,0.38858038,0.694163,2.4031622,5.5570765,7.6886096,3.832987,1.0638802,2.7389257,5.9003854,7.5112963,4.429062,2.233394,2.2673476,2.5691576,2.1994405,1.2525115,1.5543215,1.2600567,1.2525115,1.5618668,1.3958713,1.5015048,1.8485862,2.3993895,3.2746384,4.7421894,5.481624,6.436098,6.8473144,6.8963585,7.7225633,5.383536,3.5274043,2.5125682,2.637065,4.1272516,3.3651814,3.5387223,4.1574326,4.9949555,6.0814714,5.402399,3.2670932,1.8184053,1.8448136,2.757789,2.3277097,1.9127209,1.6675003,1.5316857,1.2336484,1.20724,1.6788181,2.2748928,2.8747404,3.5839937,3.0369632,2.474842,2.4182527,2.8596497,3.2520027,4.395108,4.8063245,4.908185,4.5799665,3.169005,1.4977322,1.7731338,2.0447628,1.6561824,1.237421,1.4449154,1.7354075,1.9466745,2.305074,3.451952,4.3611546,4.908185,5.0025005,5.194905,6.6813188,8.948667,10.295494,9.7220545,8.073418,8.035691,10.570895,12.559069,14.354838,15.682802,15.633758,13.392818,12.6345215,14.347293,17.169216,17.37671,18.085964,21.24365,24.857826,27.596752,28.788902,33.893265,37.099995,38.910854,38.390232,33.1576,29.63397,25.914162,21.511507,17.731337,17.663431,16.87118,14.403882,12.879742,13.166461,14.366156,12.272349,9.650374,7.3151197,6.319147,7.9300575,7.4169807,6.519096,5.0553174,3.682082,3.904667,4.1498876,6.115425,8.424272,9.639057,8.254503,6.63982,5.515578,5.2364035,5.353355,4.5912848,5.462761,6.802043,8.126234,9.544742,11.759273,11.793225,12.917468,13.758763,13.849306,13.630494,15.365902,15.9695215,16.03743,16.014793,16.22606,13.343775,11.676274,11.623458,12.577931,12.917468,15.098045,18.489635,23.356321,28.739857,32.459667,23.7864,16.16947,12.740154,13.2607765,14.162435,13.008011,11.710228,11.653639,13.4644985,17.037174,18.863125,20.534397,18.746174,12.925014,5.240176,6.0512905,6.5341864,7.914967,9.65792,9.469289,8.062099,8.993938,7.752744,4.745962,5.292993,7.4584794,9.314611,10.9594755,12.095036,11.98563,9.231613,9.835234,15.30554,23.593996,29.105803,27.804247,23.809036,18.097282,12.921241,11.808316,11.812089,9.110889,7.3905725,7.779153,8.854351,11.227332,14.943368,15.690348,13.219278,11.363147,13.822898,14.083209,14.154889,15.531898,19.191343,20.568352,20.33822,19.127209,18.006739,18.459454,21.349285,20.485353,20.036411,20.768301,20.006231,20.764528,25.736847,28.822855,28.554998,28.12492,27.687294,28.44182,28.215462,27.966469,31.784365,34.75342,35.65508,35.47022,35.32309,36.46242,31.448603,27.253443,27.196854,28.01174,19.836462,17.931286,16.735365,15.049001,12.740154,10.7218,9.005256,10.544487,13.2607765,14.566105,11.332966,10.0465,9.688101,8.194141,5.7683434,4.847823,13.973803,13.804035,11.77059,10.502988,7.828197,4.8968673,3.7763977,2.9124665,2.546522,4.7233267,7.0887623,7.54525,6.9152217,6.0512905,5.80607,6.19465,8.6732645,11.027383,11.631002,9.424017,9.7296,7.779153,5.8513412,5.0439997,5.2628117,2.7691069,2.0296721,2.071171,2.1881225,1.9278114,3.2633207,6.802043,12.694883,17.82188,15.79598,14.713238,12.989148,10.79348,8.718536,7.7602897,5.8966126,9.046755,10.612394,8.741172,6.3455553,8.703445,9.382519,8.552541,6.4210076,3.229367,1.1091517,0.5394854,1.2789198,3.0633714,5.613666,8.926031,8.812852,6.579458,4.447925,5.572167,9.061845,14.667966,15.83748,12.913695,13.106099,14.083209,14.5283785,14.769827,14.724555,13.951167,12.743927,9.710737,9.0543,11.457462,14.086982,15.403628,14.811326,13.011784,11.529142,12.702429,12.2119875,10.419991,9.1976595,8.922258,8.458225,8.29223,8.420499,7.567886,6.168242,6.3832817,4.4743333,5.028909,6.092789,6.6058664,6.3945994,8.405409,7.6320205,6.360646,6.2625575,8.367682,11.114153,9.937095,6.7379084,3.7198083,3.3651814,3.7537618,4.9459114,6.3531003,7.54525,8.2507305,7.9791017,7.092535,5.160951,3.0709167,3.029418,5.0439997,5.753253,6.609639,7.432071,6.368191,4.353609,4.949684,5.7079816,5.040227,2.2107582,3.2821836,3.682082,3.500996,3.059599,2.897376,2.674791,2.9803739,3.5802212,3.9914372,3.4632697,3.0181,3.2369123,3.561358,3.5877664,3.0746894,4.0178456,5.304311,5.904158,5.142088,2.71629,2.0183544,1.7693611,1.6712729,1.5920477,1.539231,1.6071383,1.3619176,1.1657411,1.1996948,1.448688,1.0450171,1.0148361,1.0827434,0.97333723,0.41498876,0.35462674,0.663982,0.8337501,0.8224323,1.0412445,0.90543,0.76584285,0.72811663,0.77716076,0.8186596,0.7997965,0.60362,0.33576363,0.14713238,0.23013012,0.27540162,0.19240387,0.1056335,0.06413463,0.00754525,0.00754525,0.003772625,0.00754525,0.018863125,0.033953626,0.0150905,0.071679875,0.10940613,0.11317875,0.15845025,0.43385187,0.4074435,0.2867195,0.21503963,0.24899325,0.120724,0.056589376,0.23767537,0.87147635,2.1956677,3.289729,4.6026025,5.111907,4.3649273,2.4974778,2.0900342,1.448688,0.7696155,0.241448,0.030181,0.150905,0.43385187,0.62248313,0.69793564,0.84129536,0.91674787,0.8865669,0.79602385,0.6790725,0.56212115,0.43007925,0.5319401,0.66775465,0.6526641,0.31312788,0.20749438,0.19240387,0.2263575,0.29803738,0.44516975,0.47157812,0.52062225,0.62248313,0.7092535,0.62625575,0.52439487,0.5319401,0.5998474,0.67152727,0.69039035,0.6375736,0.67152727,0.8299775,0.97333723,0.77338815,0.8224323,0.9393836,0.87147635,0.6149379,0.4074435,0.32067314,0.26031113,0.22258487,0.20749438,0.19994913,0.22258487,0.30935526,0.38858038,0.4376245,0.47157812,0.5772116,0.68661773,0.7130261,0.67152727,0.6790725,0.6111652,0.5583485,0.5470306,0.58475685,0.633801,0.62625575,0.5055317,0.47912338,0.6073926,0.7922512,0.76207024,0.7167987,0.67152727,0.633801,0.6149379,0.69039035,0.73188925,0.7809334,0.8262049,0.814887,0.98465514,0.9808825,0.87147635,0.7507524,0.72811663,0.67152727,0.6488915,0.60362,0.51684964,0.41876137,0.41121614,0.4678055,0.482896,0.44516975,0.4376245,0.55457586,0.6488915,0.62625575,0.513077,0.45648763,0.5885295,0.6375736,0.77338815,0.97710985,1.0186088,0.9016574,0.8563859,0.9205205,1.0450171,1.1280149,1.1619685,1.1053791,1.0110635,0.94692886,1.0035182,1.20724,1.1732863,1.0035182,0.814887,0.7432071,0.72811663,0.79602385,0.814887,0.73566186,0.58098423,0.5885295,0.6375736,0.694163,0.7582976,0.8601585,0.935611,0.9997456,1.116697,1.2713746,1.3920987,1.7316349,1.720317,1.6146835,1.6146835,1.8599042,1.8787673,1.9127209,1.9881734,2.0598533,2.003264,1.8448136,1.6675003,1.5882751,1.6184561,1.6260014,1.6146835,1.6184561,1.6146835,1.6712729,1.9391292,2.4333432,2.8445592,3.1350515,3.2935016,3.31991,3.4632697,3.7763977,4.036709,4.1800685,4.2819295,3.953711,3.5160866,3.029418,2.5691576,2.233394,2.1805773,2.0108092,1.8485862,1.7844516,1.8636768,1.931584,2.0749438,2.474842,3.1652324,4.0480266,4.478106,4.983638,5.0854983,4.745962,4.3724723,0.5583485,0.271629,0.17354076,0.15845025,0.1358145,0.06413463,0.10186087,0.0754525,0.03772625,0.033953626,0.11317875,0.15845025,0.14713238,0.150905,0.1659955,0.13204187,0.14713238,0.23390275,0.32444575,0.3772625,0.34330887,0.29426476,0.211267,0.181086,0.20749438,0.24899325,0.21503963,0.13204187,0.094315626,0.11317875,0.094315626,0.030181,0.02263575,0.02263575,0.011317875,0.0,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.018863125,0.02263575,0.0150905,0.011317875,0.011317875,0.00754525,0.011317875,0.10186087,0.45648763,0.94315624,2.6710186,4.689373,5.413717,2.6446102,1.2638294,3.289729,5.802297,6.4474163,3.399135,2.0598533,1.7957695,1.9655377,1.9806281,1.3392819,2.033445,1.7467253,1.4147344,1.3468271,1.20724,1.4373702,1.8561316,2.9803739,5.2628117,9.0957985,9.710737,7.9225125,6.485142,6.8699503,9.231613,7.3453007,4.4743333,2.9916916,3.5236318,4.9421387,3.3651814,2.9992368,3.4632697,4.1612053,4.293247,4.346064,2.7728794,1.3543724,0.80356914,0.79602385,0.7167987,0.7922512,0.9695646,1.1921495,1.4147344,1.6373192,2.252257,3.150142,4.1762958,5.1534057,4.708236,3.4896781,2.5729303,2.2296214,1.9164935,2.4069347,2.867195,3.5160866,3.5575855,1.1581959,0.76207024,1.7052265,1.8184053,0.98842776,1.1581959,1.7580433,2.2975287,2.8596497,3.7160356,5.3571277,6.48137,7.726336,8.880759,9.639057,9.6051035,10.397354,13.094781,14.264296,13.211733,12.00072,14.875461,15.041456,14.84528,15.46399,16.890041,15.886524,16.094019,17.991648,20.628714,21.617142,24.529608,28.317324,30.603535,30.969479,30.94307,32.776566,30.705395,31.520283,35.13823,34.591198,32.316307,28.377686,22.756474,17.1164,14.811326,13.441863,10.340765,9.258021,11.231105,14.596286,10.054046,8.548768,8.22055,8.239413,8.76758,7.4094353,5.987156,5.0741806,4.9232755,5.4665337,4.115934,6.4549613,9.175024,10.057818,7.9753294,6.356873,5.292993,5.172269,5.251494,3.6556737,5.5004873,6.888813,8.096053,9.363655,10.887795,10.850069,12.385528,13.936077,14.720782,14.750964,13.577678,13.671993,14.596286,15.064092,12.936331,11.091517,12.1101265,14.18507,15.762027,15.539442,18.715992,23.537407,30.181,35.598488,33.51977,22.29244,17.833199,18.327412,20.617395,20.202406,17.45971,18.448135,22.269806,27.2044,30.686531,26.302742,20.274086,14.452927,9.529651,5.036454,7.3113475,7.413208,8.009283,9.578695,10.397354,9.880505,11.657412,10.680302,6.7756343,4.6252384,4.5497856,8.047009,11.589504,13.555041,14.2077055,9.865415,9.26934,12.438345,18.112373,23.763765,26.08393,27.60807,22.665932,13.788944,11.714001,14.290704,12.672247,10.846297,10.453944,10.789707,12.166716,15.256495,16.418465,14.335975,10.023865,10.49167,11.378237,12.155397,13.600313,17.818108,19.768555,19.074392,18.025602,17.738882,18.157644,17.395575,17.399347,18.38023,19.798737,20.33822,20.357084,26.366877,30.76953,30.795938,28.475773,26.755457,26.1292,25.585943,26.151836,30.92798,35.994614,36.413376,36.556736,37.503666,37.062267,32.376667,28.683268,28.868126,29.769783,22.179262,20.010002,18.900852,17.172989,14.249205,10.665211,9.507015,10.269085,9.680555,7.835742,8.194141,7.4018903,7.6886096,7.7640624,6.5266414,3.0860074,7.515069,9.21275,8.918486,7.492433,5.9192486,4.5799665,4.4215164,3.6254926,2.493705,3.4594972,6.587003,6.5945487,5.753253,5.704209,7.4471617,7.092535,9.22784,10.47658,10.144588,10.212496,12.404391,9.978593,7.111398,5.2892203,3.2746384,2.5502944,2.3805263,2.2371666,2.0673985,2.293756,3.3727267,9.076936,14.339747,16.075155,13.181552,13.804035,13.355092,12.479843,12.015811,12.97783,8.963757,14.837734,15.226315,9.314611,10.850069,14.554788,12.038446,7.7829256,4.5120597,3.1652324,1.3656902,0.7130261,1.3468271,2.6710186,3.3727267,4.6252384,6.3531003,6.175787,4.5422406,4.708236,6.5756855,12.325166,14.102073,11.6875925,12.510024,13.377728,14.939595,16.25624,16.825907,16.561823,14.841507,11.234878,9.80128,11.3669195,13.521088,16.28265,16.780636,14.656648,12.200669,14.34352,13.630494,10.533169,8.488406,8.397863,8.612903,8.36391,8.741172,8.246958,6.470052,4.093298,4.3196554,5.4703064,5.764571,5.349582,6.3153744,9.439108,10.163452,8.790216,6.8661776,7.164215,6.934085,5.1571784,3.3878171,2.4484336,2.4182527,3.0633714,3.9310753,4.606375,5.281675,6.771862,6.1644692,7.1868505,6.677546,4.323428,2.6408374,2.8445592,3.270866,3.7650797,3.9499383,3.229367,3.5839937,4.678055,5.7494807,5.572167,2.4672968,2.9124665,3.3463185,3.2520027,2.7540162,2.6106565,2.4484336,3.2105038,4.2630663,4.8365054,4.0480266,3.7047176,3.6934,4.168751,4.7233267,4.432834,3.6971724,4.0706625,4.979865,5.247721,3.0935526,2.0749438,1.7014539,1.6524098,1.6184561,1.2902378,1.4034165,1.3317367,1.0902886,0.935611,1.3543724,1.1053791,0.9997456,0.94692886,0.80734175,0.3734899,0.32444575,0.62248313,0.69793564,0.5696664,0.8262049,0.7167987,0.52439487,0.38480774,0.331991,0.28294688,0.33576363,0.27917424,0.1659955,0.1056335,0.23013012,0.32821837,0.29426476,0.2263575,0.150905,0.02263575,0.00754525,0.003772625,0.00754525,0.011317875,0.0150905,0.003772625,0.033953626,0.05281675,0.056589376,0.0754525,0.26031113,0.34330887,0.32067314,0.23390275,0.1659955,0.124496624,0.08299775,0.14335975,0.59230214,1.9089483,2.263575,2.655928,3.3463185,3.8367596,2.8747404,1.8485862,1.4600059,1.086516,0.5319401,0.033953626,0.16222288,0.41876137,0.58098423,0.6451189,0.8224323,0.9205205,0.80734175,0.76584285,0.8299775,0.7922512,0.44894236,0.5093044,0.7054809,0.784706,0.47912338,0.29426476,0.21881226,0.21881226,0.28294688,0.43007925,0.55457586,0.56589377,0.62248313,0.7130261,0.6526641,0.5470306,0.59230214,0.67152727,0.7130261,0.6790725,0.694163,0.6413463,0.58475685,0.5772116,0.66775465,0.724344,0.8526133,0.80356914,0.56212115,0.35839936,0.29426476,0.26408374,0.24522063,0.23013012,0.20749438,0.23767537,0.27540162,0.362172,0.47157812,0.482896,0.55457586,0.7205714,0.7809334,0.70170826,0.58475685,0.5998474,0.56212115,0.5394854,0.543258,0.55080324,0.56589377,0.573439,0.5998474,0.7167987,1.0148361,0.814887,0.6413463,0.62625575,0.72811663,0.7582976,0.80356914,0.83752275,0.9393836,1.0412445,0.95447415,0.8903395,0.77716076,0.66775465,0.6187105,0.6828451,0.6375736,0.5583485,0.51684964,0.5017591,0.42630664,0.3961256,0.482896,0.52439487,0.5017591,0.56589377,0.76207024,0.76207024,0.66020936,0.5470306,0.51684964,0.6149379,0.73188925,0.91674787,1.0450171,0.8224323,0.7582976,0.6752999,0.7394345,0.95824677,1.1921495,1.177059,1.1431054,1.1581959,1.1846043,1.0751982,1.116697,1.0714256,1.0299267,1.0110635,0.9695646,0.814887,0.79602385,0.8563859,0.90543,0.7922512,0.7054809,0.63002837,0.59607476,0.6413463,0.80734175,0.8639311,0.8111144,0.8111144,0.8865669,0.94692886,1.2147852,1.3392819,1.3958713,1.4675511,1.629774,1.7014539,1.750498,1.841041,1.9806281,2.1013522,2.0258996,1.8372684,1.7316349,1.7655885,1.8485862,1.6939086,1.4977322,1.3770081,1.418507,1.6524098,2.1164427,2.4861598,2.7728794,2.9841464,3.1237335,3.1237335,3.3274553,3.6443558,3.9386206,4.0517993,3.7613072,3.4029078,2.8709676,2.2862108,1.9806281,1.8599042,1.7655885,1.7618159,1.8523588,1.9768555,1.9391292,1.9693103,2.3692086,3.169005,4.142342,4.3007927,4.749735,4.9760923,4.8440504,4.587512,0.29049212,0.31312788,0.27540162,0.21503963,0.150905,0.0754525,0.06413463,0.033953626,0.041498873,0.0754525,0.0754525,0.10186087,0.041498873,0.08677038,0.21503963,0.23013012,0.120724,0.12826926,0.24899325,0.35462674,0.18485862,0.03772625,0.06413463,0.120724,0.116951376,0.030181,0.00754525,0.018863125,0.07922512,0.13204187,0.0452715,0.02263575,0.0150905,0.00754525,0.0,0.0,0.011317875,0.00754525,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.0150905,0.011317875,0.0,0.0,0.018863125,0.02263575,0.0754525,0.32067314,1.5882751,2.8030603,3.7763977,4.123479,3.2821836,2.3767538,2.867195,3.7990334,3.9386206,1.7391801,0.6526641,0.34330887,0.814887,1.5580941,1.5731846,1.961765,2.5087957,2.3201644,1.5882751,1.5882751,1.9051756,2.4786146,5.2854476,10.95193,18.75372,17.142809,13.754991,10.578441,8.778898,8.68081,7.5603404,5.2288585,3.99521,4.346064,4.9421387,4.466788,5.089271,4.991183,4.074435,3.953711,3.5236318,2.2748928,1.2223305,0.784706,0.7469798,0.68661773,0.9016574,1.6071383,2.8445592,4.45547,5.515578,6.900131,8.103599,8.975075,9.718282,7.2887115,4.9157305,3.3915899,2.4672968,0.8563859,0.965792,0.69793564,0.48666862,0.6488915,1.4034165,1.4637785,1.0223814,0.80734175,1.1091517,1.7542707,3.4896781,4.014073,3.9084394,3.9273026,4.991183,5.6853456,7.3792543,10.265312,12.800517,11.7026825,9.763554,12.913695,15.626213,15.90916,15.275358,17.972786,17.969013,15.992157,13.996439,15.165953,16.90136,19.183798,22.296213,25.816072,28.626678,33.372643,34.66288,34.055485,32.96897,32.63698,29.354795,25.26527,25.148317,27.438301,24.21648,22.213217,22.337713,21.669958,19.07062,15.150862,12.698656,11.087745,12.404391,14.607604,11.521597,7.858378,9.258021,12.366665,14.6151495,14.237886,11.649866,8.152642,6.1041074,6.039973,6.700182,5.4665337,7.1906233,9.563604,10.831206,9.782416,9.7069645,8.333729,7.364164,6.9869013,5.8890676,7.99042,8.412953,8.639311,9.374973,10.559577,9.7296,11.106608,12.528888,13.441863,14.909414,14.6151495,14.313339,15.418718,16.135517,11.461235,11.521597,15.297995,18.983849,20.458946,19.28566,23.692085,29.37366,35.636215,38.07333,28.566317,20.66644,20.285404,24.00144,28.087193,28.502182,29.185026,33.1576,40.853756,48.802677,49.621338,32.859562,19.508244,10.93684,6.964266,5.828706,8.820397,9.009028,8.031919,7.8696957,10.850069,9.590013,10.925522,12.2270775,11.461235,7.201941,4.3347464,7.745199,12.721292,16.173243,16.663685,10.035183,9.208978,11.012292,14.32843,20.126955,26.265015,33.21042,30.64126,19.723284,13.106099,14.803781,15.226315,15.403628,15.011275,12.37421,11.348056,13.373956,14.543469,13.072145,9.276885,10.023865,11.050018,11.819634,13.143826,17.195625,20.209951,19.334703,17.603067,16.863634,17.7917,17.30503,17.1164,17.784155,18.874443,18.99894,19.130981,23.58645,28.622906,30.878935,27.389257,26.008476,25.389767,25.00496,25.8123,30.241362,40.00869,39.71065,38.563774,39.125893,37.307487,32.425713,28.969988,27.083675,25.819845,23.133736,20.33822,18.859352,17.029629,14.437836,11.947904,10.26154,10.042727,9.152389,6.9982195,4.5309224,3.2029586,5.2326307,11.02361,14.777372,4.5007415,4.0970707,4.115934,5.3269467,6.4436436,4.134797,3.6971724,3.9989824,4.2592936,3.92353,2.655928,8.624221,11.627231,10.401127,7.4811153,9.216523,7.496206,6.900131,10.023865,14.947141,15.226315,19.123436,12.242168,7.2924843,7.1076255,4.6554193,3.5689032,2.9954643,2.4031622,2.1956677,3.7235808,5.7494807,15.848798,21.013521,17.610613,11.3971,10.616167,9.808825,9.7296,11.148107,14.84528,10.38981,10.310584,9.2995205,7.798016,12.0082655,14.671739,9.944639,4.7421894,2.0900342,1.1129243,0.8563859,0.84884065,2.0070364,3.519859,2.8219235,2.1994405,2.9615107,3.187868,2.7540162,3.3425457,7.149124,13.392818,14.588741,11.155652,11.3971,11.204697,13.95494,16.22606,16.976812,17.56157,14.781145,12.068627,11.148107,11.725319,11.506506,15.656394,18.772581,20.145817,21.043703,24.718239,22.239624,14.992412,8.699674,6.1116524,6.9869013,6.1833324,6.677546,7.4282985,6.9491754,3.3123648,5.5193505,8.141325,7.360391,4.436607,5.7079816,9.35611,11.3669195,9.805053,5.9909286,4.5007415,4.3800178,2.8294687,1.8938577,2.1881225,2.8822856,4.6290107,4.9119577,4.696918,4.9760923,6.760544,5.96452,9.1825695,10.993429,8.975075,3.6783094,1.7731338,0.965792,0.77716076,0.87147635,1.0676528,2.203213,3.0558262,4.134797,4.727099,2.8822856,2.957738,3.8103511,4.5120597,4.6214657,4.195159,3.731126,4.5233774,4.9685473,4.587512,4.014073,2.867195,3.5953116,5.028909,5.885295,4.7610526,2.757789,3.2482302,4.3196554,4.6214657,3.3274553,2.4710693,1.780679,1.5920477,1.7316349,1.50905,1.4373702,1.6486372,1.4939595,1.0638802,1.1581959,1.1732863,0.965792,0.663982,0.39989826,0.29049212,0.27917424,0.513077,0.5319401,0.33953625,0.41121614,0.35085413,0.30935526,0.19994913,0.05281675,0.0150905,0.041498873,0.0452715,0.033953626,0.033953626,0.1056335,0.31312788,0.35839936,0.30935526,0.20372175,0.0452715,0.02263575,0.0150905,0.00754525,0.003772625,0.0150905,0.0150905,0.0150905,0.041498873,0.0754525,0.0754525,0.06413463,0.16976812,0.2565385,0.24899325,0.150905,0.150905,0.14335975,0.10186087,0.06413463,0.1358145,2.0183544,2.4597516,2.0749438,1.7769064,2.776652,1.6410918,1.3770081,1.267602,0.875249,0.0452715,0.20372175,0.4074435,0.513077,0.5319401,0.6413463,0.8224323,0.80734175,0.7696155,0.7696155,0.73188925,0.47535074,0.4376245,0.55457586,0.68661773,0.62625575,0.47912338,0.34330887,0.26408374,0.24899325,0.26031113,0.49044126,0.5583485,0.62625575,0.72811663,0.76207024,0.58098423,0.663982,0.83752275,0.9242931,0.7167987,0.59607476,0.45648763,0.38858038,0.44894236,0.65643674,0.7922512,0.7054809,0.5017591,0.30935526,0.26031113,0.24899325,0.23390275,0.241448,0.2565385,0.24522063,0.3055826,0.31312788,0.38480774,0.49421388,0.45648763,0.482896,0.52439487,0.56589377,0.58475685,0.55080324,0.62248313,0.66020936,0.72811663,0.80734175,0.7922512,0.73188925,0.83752275,0.8299775,0.724344,0.80734175,0.62625575,0.55080324,0.5696664,0.6111652,0.55080324,0.48666862,0.55457586,0.6828451,0.8563859,1.1129243,0.845068,0.6488915,0.5696664,0.58475685,0.6111652,0.67152727,0.5772116,0.46026024,0.36594462,0.24522063,0.23013012,0.3470815,0.47157812,0.59230214,0.8224323,0.87147635,0.7469798,0.6488915,0.5885295,0.38103512,0.43007925,0.663982,0.90543,1.0148361,0.87147635,0.9922004,0.83752275,0.76584285,0.9620194,1.448688,1.4147344,1.2940104,1.177059,1.0751982,0.91674787,1.086516,0.91674787,0.8224323,0.87147635,0.8224323,0.69039035,0.63002837,0.573439,0.5357128,0.59607476,0.754525,0.77338815,0.70170826,0.6375736,0.7469798,0.77338815,0.7130261,0.66020936,0.6526641,0.70170826,0.77338815,0.8941121,1.0601076,1.2034674,1.1883769,1.2638294,1.3807807,1.5958204,1.8334957,1.9089483,1.8599042,1.81086,1.8749946,1.9844007,1.8599042,1.7165444,1.478869,1.3241913,1.3355093,1.4939595,1.8976303,2.1466236,2.2598023,2.305074,2.3654358,2.463524,2.7540162,2.9124665,2.9049213,2.9916916,3.0030096,2.9237845,2.5616124,2.052308,1.8448136,1.6373192,1.6222287,1.6712729,1.720317,1.7693611,1.8787673,1.9164935,2.003264,2.335255,3.187868,3.8858037,4.4516973,4.9345937,5.2326307,5.111907,0.120724,0.32067314,0.17731337,0.06413463,0.094315626,0.150905,0.17731337,0.13204187,0.08677038,0.05281675,0.0150905,0.08677038,0.1659955,0.1961765,0.181086,0.20372175,0.056589376,0.08299775,0.16222288,0.2263575,0.27917424,0.27917424,0.211267,0.11317875,0.033953626,0.06790725,0.120724,0.08677038,0.06790725,0.090543,0.08299775,0.03772625,0.011317875,0.0,0.0,0.0,0.041498873,0.049044125,0.030181,0.003772625,0.0150905,0.003772625,0.003772625,0.00754525,0.011317875,0.0,0.0,0.003772625,0.011317875,0.06790725,0.271629,1.7467253,3.0633714,3.0897799,2.1843498,2.1805773,2.04099,1.7165444,1.418507,1.1204696,0.55457586,0.56212115,0.7167987,1.1053791,1.7919968,2.8407867,2.987919,2.637065,2.2258487,2.022127,2.1466236,2.1541688,3.3576362,5.4401255,8.511042,13.124963,12.2270775,10.265312,8.130007,6.3417826,5.0439997,3.8141239,4.1800685,4.7006907,4.636556,3.953711,4.3875628,4.2781568,4.112161,3.8971217,3.169005,1.8259505,1.2034674,0.97710985,1.0223814,1.3958713,2.3088465,2.848332,3.4594972,4.195159,4.7120085,3.8707132,4.8402777,6.356873,7.352846,6.9869013,5.3269467,4.244203,3.6254926,3.3312278,3.1840954,3.7160356,4.0103,3.9386206,3.6141748,3.3915899,3.4330888,3.7990334,4.002755,4.044254,4.429062,6.6586833,7.141579,6.7341356,6.5341864,7.8696957,7.997965,9.061845,10.638803,12.117672,12.668475,9.827688,9.884277,11.41219,13.592768,16.188334,20.545715,23.133736,22.281124,18.938578,16.693865,19.31584,24.35984,27.626932,27.970242,27.317577,30.282862,32.96897,35.73053,37.047176,33.504684,27.027086,21.153109,17.904879,17.297485,17.308804,17.825653,20.590988,22.039675,21.34174,20.402355,18.270823,14.25675,12.132762,12.2270775,11.434827,13.924759,15.169725,15.569623,15.875206,17.225805,17.120173,12.698656,7.635793,4.5761943,5.1345425,6.3832817,8.397863,10.661438,12.96274,15.4074,14.377474,12.427027,10.9594755,10.080454,8.612903,8.428044,6.7643166,6.6813188,8.699674,10.804798,10.49167,14.1926155,16.271332,15.573396,15.456445,15.973294,15.041456,13.641812,12.1252165,10.212496,13.272095,18.97253,22.50748,22.571615,21.360603,25.163408,30.99966,35.36836,36.1757,32.73884,31.50142,33.998898,36.598236,37.55648,37.03586,42.162857,50.481495,57.17036,58.547367,52.050907,31.96168,17.444618,9.537196,7.492433,8.7600355,11.219787,10.691619,8.5563135,6.5228686,6.651138,7.149124,6.9152217,6.541732,5.9607477,4.45547,2.916239,6.477597,12.37421,17.350302,17.663431,9.578695,7.673519,8.488406,10.7218,15.230087,20.862616,28.796446,34.915646,34.900555,24.20139,15.558306,14.211478,14.675511,14.275613,13.132507,11.2650585,12.355347,15.679029,18.28214,14.954685,14.867915,15.124454,14.622695,13.928532,15.267814,19.47429,19.440336,17.708702,17.014538,20.258997,18.101055,17.429527,18.270823,19.406384,18.376457,18.146326,19.972277,23.89958,27.823109,27.476028,28.977533,32.59925,34.474247,34.41766,35.93048,41.283836,41.129158,42.906063,45.467678,39.07685,33.580135,31.33165,31.50142,32.003178,29.49061,25.484081,21.349285,17.901106,15.531898,14.1926155,13.641812,12.351574,10.020092,7.115171,4.8742313,3.1425967,3.3274553,7.0472636,10.872705,6.356873,5.0251365,6.571913,8.465771,9.114662,7.8206515,4.7836885,5.1760416,8.714764,10.9594755,3.3123648,5.6589375,12.611885,14.286931,9.431562,5.4438977,5.6287565,11.936585,15.977067,15.562078,14.739646,21.534143,16.086473,9.25425,6.175787,6.2889657,5.379763,5.311856,4.4403796,2.8181508,2.1956677,4.534695,18.033148,25.646305,21.994404,13.35132,12.453435,9.842778,7.443389,7.326438,11.69891,12.593022,13.721037,11.072655,6.2436943,6.4436436,7.1038527,5.3759904,3.821669,3.3953626,3.4444065,3.9688015,3.7763977,3.4217708,3.6594462,5.4212623,3.199186,2.5125682,2.214531,2.5012503,4.8930945,8.933576,12.826925,13.702174,12.283667,12.887287,9.929549,10.804798,12.97783,15.354584,18.293459,16.576914,14.219024,12.83447,11.774363,8.137552,9.884277,13.030646,15.380992,17.05981,20.50799,24.718239,19.613878,11.853588,6.205968,5.523123,4.696918,4.7836885,5.855114,6.670001,4.7044635,6.1795597,6.609639,5.2288585,3.2746384,3.983892,6.63982,7.61693,6.983129,5.704209,5.6476197,7.5075235,5.172269,2.4974778,1.4222796,1.991946,3.270866,4.164978,5.1760416,6.33801,7.224577,7.1906233,9.4127,11.502733,11.32542,6.9869013,2.425798,1.0374719,0.9922004,1.2449663,1.50905,1.9089483,3.1954134,5.9682927,7.9413757,3.9197574,4.5497856,5.160951,5.9418845,6.8699503,7.7112455,5.1760416,4.2781568,4.191386,4.112161,3.2557755,3.1652324,2.9841464,3.1350515,3.3878171,2.8822856,1.9730829,2.323937,2.7238352,2.6974268,2.5087957,2.0636258,1.4977322,1.3015556,1.50905,1.7316349,1.6071383,1.6976813,1.5769572,1.2940104,1.3430545,1.0412445,0.7922512,0.60362,0.45648763,0.32821837,0.20749438,0.25276586,0.35839936,0.41498876,0.30181,0.20372175,0.150905,0.08677038,0.026408374,0.026408374,0.033953626,0.08299775,0.1056335,0.08299775,0.056589376,0.14713238,0.2565385,0.2565385,0.14713238,0.056589376,0.02263575,0.02263575,0.02263575,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.033953626,0.10186087,0.049044125,0.094315626,0.14335975,0.14713238,0.116951376,0.124496624,0.16222288,0.16976812,0.12826926,0.0754525,0.5696664,0.97333723,1.720317,2.6634734,3.0709167,2.052308,1.4071891,0.8337501,0.30181,0.056589376,0.090543,0.21881226,0.34330887,0.4376245,0.55457586,0.63002837,0.6752999,0.7167987,0.77716076,0.86770374,0.58098423,0.42630664,0.422534,0.513077,0.5885295,0.41498876,0.31312788,0.32067314,0.36594462,0.26031113,0.34330887,0.43385187,0.5093044,0.6073926,0.8111144,0.6790725,0.62625575,0.67152727,0.76207024,0.7922512,0.6375736,0.482896,0.45648763,0.5696664,0.72811663,0.845068,0.70170826,0.48666862,0.3169005,0.26031113,0.20749438,0.18485862,0.20372175,0.24522063,0.27917424,0.31312788,0.3055826,0.32821837,0.392353,0.43385187,0.45648763,0.5017591,0.573439,0.6526641,0.6828451,0.59230214,0.5357128,0.59607476,0.7054809,0.633801,0.66020936,0.7507524,0.7507524,0.6752999,0.7092535,0.58475685,0.58475685,0.60362,0.5998474,0.5998474,0.7130261,0.69039035,0.66775465,0.724344,0.8941121,0.7507524,0.69039035,0.62248313,0.543258,0.5357128,0.52062225,0.39989826,0.32821837,0.32444575,0.27917424,0.3470815,0.482896,0.56212115,0.56212115,0.58098423,0.7167987,0.76584285,0.7582976,0.7167987,0.68661773,0.6752999,0.69039035,0.8262049,1.0148361,1.0148361,0.8563859,0.7997965,0.7922512,0.8639311,1.1581959,1.3920987,1.1732863,0.8941121,0.80356914,1.026154,1.0902886,0.995973,0.8639311,0.754525,0.6790725,0.62248313,0.6073926,0.6187105,0.60362,0.4979865,0.452715,0.45648763,0.4979865,0.55080324,0.5998474,0.5772116,0.513077,0.51684964,0.6073926,0.72811663,0.7696155,0.7432071,0.7507524,0.8299775,0.935611,0.8903395,0.8978847,1.0186088,1.237421,1.4675511,1.6712729,1.81086,1.9429018,2.0749438,2.1805773,2.04099,1.8561316,1.6561824,1.478869,1.3845534,1.6033657,1.8259505,1.9202662,1.901403,1.9127209,1.9240388,2.1994405,2.444661,2.5578396,2.625747,2.5012503,2.3880715,2.191895,1.9429018,1.7731338,1.5354583,1.5580941,1.6373192,1.690136,1.7580433,1.9768555,2.0296721,2.0862615,2.3390274,3.0181,3.6934,4.353609,4.878004,5.1835866,5.2099953,0.094315626,0.24899325,0.18863125,0.10940613,0.1056335,0.13958712,0.13958712,0.116951376,0.11317875,0.116951376,0.090543,0.10940613,0.15845025,0.15845025,0.116951376,0.124496624,0.090543,0.15467763,0.18485862,0.16976812,0.21503963,0.26408374,0.15467763,0.0452715,0.00754525,0.030181,0.060362,0.056589376,0.049044125,0.049044125,0.056589376,0.041498873,0.02263575,0.003772625,0.0,0.0,0.15845025,0.7054809,0.77716076,0.30935526,0.0150905,0.026408374,0.06413463,0.06790725,0.041498873,0.071679875,0.211267,0.116951376,0.071679875,0.23767537,0.6526641,1.5354583,2.3465726,2.3767538,1.8674494,2.0070364,1.6260014,1.0978339,0.7167987,0.56589377,0.52439487,1.1808317,1.8749946,2.7351532,3.561358,3.8367596,3.31991,2.7728794,2.3578906,2.203213,2.3880715,2.1768045,3.3953626,4.878004,6.5266414,9.337247,10.608622,10.020092,8.013056,5.4212623,3.4859054,2.2220762,3.561358,4.274384,3.4632697,2.5729303,3.3915899,3.4594972,2.9049213,2.1353056,1.8146327,1.4034165,1.6335466,2.161714,2.6898816,2.9766011,5.0741806,7.0963078,8.563859,9.291975,9.390063,9.0957985,8.91094,9.06939,8.816625,6.4210076,4.8968673,3.2331395,2.795515,3.7235808,4.930821,6.900131,7.9451485,8.156415,7.6508837,6.609639,6.530414,6.903904,6.858632,6.2927384,5.847569,7.4282985,7.333983,7.24344,7.967784,9.461743,10.27663,11.529142,12.294985,12.581704,13.313594,12.83447,10.782163,11.091517,14.784918,19.960958,23.246916,25.985842,25.661396,22.537663,19.655376,21.813318,24.755966,26.07261,25.789665,26.37065,30.546946,36.115337,39.118347,37.216946,29.694332,24.827644,21.639776,18.531134,15.656394,14.928277,15.015047,15.69412,17.022083,20.285404,27.985332,31.30147,24.861599,15.946886,9.740918,9.318384,15.082954,17.4333,17.935059,18.221779,19.998686,19.112118,13.189097,7.654656,5.149633,5.534441,6.881268,9.363655,11.5857315,13.117417,14.517061,14.977322,13.287186,11.69891,10.589758,8.488406,7.8621507,7.273621,7.8395147,9.273112,9.922004,11.751727,14.667966,15.648849,14.864142,15.675257,17.033401,16.29774,15.041456,14.019074,13.170234,16.131744,20.82489,25.363358,28.78513,31.044931,29.977278,30.690304,31.493874,32.055996,33.399048,34.20639,35.817303,40.020004,46.312744,51.922638,59.67538,71.838326,76.3353,68.60519,51.59442,33.538635,20.70794,12.89106,9.1825695,7.99042,7.8244243,6.5530496,4.870459,3.4783602,3.0897799,4.032936,3.6028569,3.229367,3.218049,2.7879698,1.9994912,5.915476,13.834216,22.028357,23.744902,10.668983,7.145352,7.8734684,10.121953,13.713491,16.58446,25.238861,34.40257,37.398033,26.163155,17.172989,14.992412,15.124454,15.030138,14.0983,12.472299,13.588995,17.286167,20.583443,17.72002,17.557796,17.271078,16.595778,15.739391,15.380992,19.247932,20.372175,19.889278,19.67424,22.330168,19.681786,18.519815,19.319613,20.48158,18.327412,18.21046,19.538425,23.624178,28.31355,27.989105,28.358822,30.761984,31.376923,30.373404,31.923952,37.390488,37.95638,43.351234,51.183205,46.961636,42.585392,39.065533,37.76775,37.72625,35.651306,32.206898,27.117628,22.643295,19.662922,17.674747,16.199652,13.128735,9.612649,6.560595,4.647874,3.2105038,2.6672459,3.9763467,6.0701537,5.8400235,5.6551647,7.5301595,8.560086,7.696155,5.7607985,5.081726,6.4134626,9.408927,12.404391,12.404391,7.7150183,10.895341,14.060574,13.072145,7.5037513,6.1644692,10.770844,12.113899,9.699419,11.744182,26.996904,19.470518,9.582467,6.549277,8.375228,7.5792036,5.5457587,4.3083377,4.0216184,2.987919,4.349837,14.022847,20.209951,18.116146,9.940866,9.5183325,9.80128,10.767072,11.955449,12.483616,12.559069,11.321648,7.9225125,4.036709,3.8593953,5.1043615,4.496969,3.9159849,4.115934,4.715781,5.7004366,6.0512905,5.3759904,4.7233267,6.56814,5.3986263,3.610402,2.2598023,2.1390784,3.7613072,7.277394,9.295748,10.536942,11.551778,12.736382,9.367428,9.567377,11.751727,15.135772,19.742147,18.202915,14.743419,12.577931,11.631002,8.529905,9.224068,11.895086,14.260523,16.014793,18.814081,25.348267,24.484337,18.010511,9.650374,5.0477724,4.2706113,3.8820312,5.1760416,7.333983,7.4396167,7.424526,7.122716,5.7079816,3.874486,3.8480775,4.949684,5.7570257,5.798525,5.534441,6.33801,7.492433,5.8626595,3.6556737,2.0749438,1.3204187,2.6332922,3.1350515,3.500996,3.9801195,4.38379,4.5988297,5.8928404,6.9982195,6.8435416,4.534695,1.9466745,1.0940613,1.1846043,1.539231,1.5618668,2.0108092,3.4255435,5.670255,7.61693,7.1378064,6.700182,6.1606965,5.692891,5.6061206,6.349328,4.063117,3.1765501,3.4670424,4.285702,4.5497856,4.2291126,3.4255435,3.1916409,3.4368613,2.9426475,2.3880715,1.9504471,1.690136,1.6637276,1.901403,1.6109109,1.2147852,1.1016065,1.3355093,1.6675003,1.4524606,1.3996439,1.388326,1.3053282,1.0789708,0.90543,0.66775465,0.482896,0.362172,0.24522063,0.12826926,0.1056335,0.20372175,0.30935526,0.211267,0.094315626,0.060362,0.0452715,0.033953626,0.041498873,0.06790725,0.090543,0.094315626,0.07922512,0.03772625,0.05281675,0.1659955,0.21503963,0.15845025,0.071679875,0.026408374,0.0150905,0.011317875,0.00754525,0.00754525,0.0150905,0.0150905,0.011317875,0.018863125,0.05281675,0.041498873,0.05281675,0.060362,0.060362,0.071679875,0.0754525,0.10940613,0.14335975,0.150905,0.116951376,0.1659955,0.3772625,0.9922004,1.7655885,1.9730829,1.2902378,0.79602385,0.38858038,0.090543,0.041498873,0.056589376,0.14713238,0.271629,0.38858038,0.48666862,0.543258,0.59230214,0.70170826,0.84129536,0.88279426,0.5885295,0.3961256,0.3169005,0.33953625,0.3961256,0.33953625,0.28294688,0.2867195,0.3169005,0.24899325,0.29049212,0.3734899,0.4376245,0.5055317,0.66775465,0.6413463,0.6413463,0.68661773,0.7507524,0.76207024,0.62625575,0.52062225,0.5319401,0.6488915,0.77338815,0.663982,0.5470306,0.44139713,0.34330887,0.23013012,0.18485862,0.16976812,0.18485862,0.21503963,0.23390275,0.25276586,0.26408374,0.29049212,0.32821837,0.392353,0.47912338,0.65643674,0.70170826,0.62248313,0.633801,0.58098423,0.5055317,0.52439487,0.6073926,0.56589377,0.5357128,0.5885295,0.6451189,0.66775465,0.6790725,0.5394854,0.55457586,0.5583485,0.5319401,0.5998474,0.7092535,0.663982,0.62625575,0.663982,0.77338815,0.6451189,0.5772116,0.5394854,0.5093044,0.482896,0.47535074,0.36971724,0.32821837,0.38103512,0.4376245,0.44139713,0.49044126,0.51684964,0.51684964,0.5470306,0.66775465,0.7167987,0.724344,0.7394345,0.80734175,0.7054809,0.663982,0.7167987,0.8224323,0.8601585,0.8941121,0.9205205,0.90920264,0.87902164,0.90920264,1.0299267,0.9016574,0.7394345,0.69039035,0.8337501,0.7507524,0.6488915,0.573439,0.543258,0.5772116,0.52439487,0.5055317,0.5017591,0.49421388,0.47157812,0.45648763,0.45648763,0.47535074,0.5093044,0.5470306,0.5885295,0.6073926,0.5772116,0.55080324,0.6488915,0.694163,0.6828451,0.66020936,0.663982,0.694163,0.7092535,0.73566186,0.814887,0.95824677,1.146878,1.327964,1.50905,1.7127718,1.9542197,2.2296214,2.11267,1.9542197,1.8070874,1.659955,1.4600059,1.4109617,1.5052774,1.5430037,1.5128226,1.6071383,1.6750455,1.81086,1.9655377,2.1164427,2.2484846,2.1843498,2.0108092,1.8485862,1.7240896,1.5731846,1.4750963,1.5430037,1.6033657,1.629774,1.7089992,1.7995421,1.81086,1.8259505,1.9466745,2.2786655,2.8785129,3.4896781,3.9386206,4.191386,4.3649273,0.08677038,0.12826926,0.124496624,0.10186087,0.08299775,0.116951376,0.10940613,0.124496624,0.16222288,0.18863125,0.120724,0.11317875,0.124496624,0.11317875,0.094315626,0.14335975,0.14335975,0.150905,0.14713238,0.1358145,0.14713238,0.18863125,0.17731337,0.14713238,0.09808825,0.0,0.003772625,0.0452715,0.049044125,0.018863125,0.018863125,0.026408374,0.0150905,0.003772625,0.0,0.0,0.14335975,1.1581959,1.9127209,1.8372684,0.91674787,0.43385187,0.35085413,0.3470815,0.271629,0.12826926,0.41498876,0.29803738,0.22258487,0.42630664,0.9393836,1.146878,1.3430545,1.4864142,1.5731846,1.6184561,1.1016065,0.8639311,0.8262049,0.91674787,1.0789708,1.9429018,2.7804246,3.9725742,4.8855495,3.8669407,3.0407357,2.6068838,2.3428001,2.233394,2.4672968,1.9353566,3.0671442,4.798779,6.647365,8.722309,12.551523,12.264804,9.450426,5.8437963,3.308592,1.6222287,2.7011995,3.2255943,2.4597516,2.2560298,3.0897799,2.837014,2.1805773,1.841041,2.595566,3.410453,4.6252384,5.9230213,6.8699503,6.907676,8.778898,10.967021,12.2270775,12.385528,12.336484,12.1101265,10.487898,8.944894,7.605612,5.2326307,3.8782585,2.4220252,2.3314822,3.6330378,4.90064,6.903904,8.771353,9.87296,9.899368,8.854351,8.4544525,8.571404,8.216777,7.2472124,6.3719635,6.9491754,6.1305156,6.258785,7.8961043,9.827688,10.510533,11.136789,11.1631975,11.197151,13.008011,14.373701,11.830952,11.898859,16.18456,21.383238,23.103556,25.989614,26.891272,25.468992,24.186298,25.578398,25.79721,24.465473,22.609343,22.63575,26.495146,31.901318,34.00267,30.954388,23.903353,21.013521,20.006231,18.58395,16.25624,14.332202,12.291212,11.92904,14.079436,21.809546,40.385952,52.073544,40.310497,21.67373,8.028146,6.5341864,11.619685,14.396337,16.316603,17.972786,19.119663,16.0412,10.397354,8.246958,10.212496,11.4838705,9.846551,11.080199,12.781653,13.400364,12.253486,12.604341,11.77059,10.9594755,10.287949,8.76758,8.922258,8.850578,9.0807085,9.854096,11.140562,15.282904,15.924251,15.147089,14.890551,16.965494,17.53139,16.74291,16.350557,16.65614,16.520325,18.029375,21.519053,27.792929,35.315544,40.193546,34.108303,29.596243,26.989359,26.623415,28.837946,30.39604,31.641006,39.69556,53.797634,65.28905,69.269165,77.13509,76.591835,63.76868,43.192783,29.80751,20.545715,13.79649,8.744945,5.383536,3.7613072,2.8219235,2.0598533,1.3694628,1.0412445,1.901403,1.5920477,1.3920987,1.6939086,1.9768555,1.8033148,6.221059,15.829934,26.551735,29.652832,11.891314,7.3717093,8.499724,11.393328,15.897841,19.391293,25.02382,30.237589,31.882454,26.20088,20.349539,16.667458,16.033657,16.950403,15.546988,13.913441,15.120681,18.26705,20.673985,17.87847,18.651857,18.350048,18.218006,18.199142,16.935314,19.300749,21.654867,22.801746,23.337458,25.687803,23.578907,21.918951,21.967995,22.39053,19.255478,18.915941,19.87796,22.945105,27.098766,29.49061,30.652578,30.335678,28.007969,25.472763,26.90636,31.452375,31.750412,37.941288,48.165104,48.538593,46.92768,45.9053,44.80747,43.309734,41.442287,39.095715,33.795174,28.573862,24.740875,21.892544,19.029121,14.641558,10.529396,7.4471617,5.119452,3.5802212,2.686109,2.425798,2.8030603,3.8141239,4.90064,7.24344,8.771353,8.514814,6.6247296,6.530414,6.417235,8.043237,11.41219,14.792462,8.858124,8.190369,10.695392,12.917468,10.038955,7.6810646,9.748463,10.744436,9.955957,11.438599,27.396803,19.57615,9.435335,6.6322746,9.046755,7.54525,4.398881,3.5387223,4.979865,4.8440504,4.6629643,9.371201,13.407909,12.928786,5.802297,5.873977,9.465516,13.113645,14.464244,12.291212,10.178542,7.605612,4.949684,3.240685,4.1612053,7.7414265,6.881268,4.8553686,3.8065786,4.727099,5.281675,6.119198,5.9607477,5.3910813,6.85486,7.5716586,5.4212623,3.1425967,2.3126192,3.3312278,5.564622,6.2851934,7.5301595,9.469289,10.431308,8.684583,9.046755,10.484125,12.951422,17.399347,16.682549,14.422746,13.019329,12.268577,9.348565,9.884277,12.245941,14.517061,16.233604,18.38023,24.457928,25.359585,20.877707,13.204187,6.937857,4.930821,4.244203,6.1644692,9.559832,10.876478,9.325929,8.677037,7.726336,6.1078796,4.293247,4.134797,4.4630156,4.8855495,5.3344917,6.0512905,6.6850915,6.7152724,5.458988,3.187868,1.1317875,1.9730829,1.8297231,1.5769572,1.6109109,1.8599042,1.8749946,2.3503454,2.6068838,2.4107075,1.9881734,1.7127718,1.6750455,1.9240388,2.2409391,2.1541688,2.5389767,3.0671442,3.983892,5.455216,7.5603404,6.9944468,6.7114997,5.7872066,4.5950575,4.8402777,3.5764484,2.8256962,3.078462,4.08198,4.825187,4.2706113,3.410453,3.2520027,3.651901,3.3123648,3.1350515,2.2220762,1.4411428,1.1996948,1.4449154,1.3619176,0.98465514,0.8186596,1.0374719,1.4637785,1.1619685,0.98465514,0.98842776,1.026154,0.7432071,0.694163,0.52439487,0.35839936,0.24522063,0.1358145,0.06413463,0.06790725,0.15845025,0.24899325,0.181086,0.05281675,0.03772625,0.060362,0.08299775,0.10186087,0.094315626,0.071679875,0.056589376,0.05281675,0.02263575,0.018863125,0.09808825,0.19240387,0.23013012,0.16222288,0.07922512,0.026408374,0.00754525,0.00754525,0.018863125,0.0150905,0.018863125,0.018863125,0.0150905,0.0150905,0.030181,0.03772625,0.030181,0.018863125,0.033953626,0.049044125,0.06413463,0.094315626,0.12826926,0.12826926,0.124496624,0.2565385,0.5055317,0.7582976,0.7884786,0.49044126,0.271629,0.12826926,0.06790725,0.08677038,0.05281675,0.1056335,0.211267,0.32821837,0.41498876,0.49421388,0.5470306,0.66020936,0.7997965,0.80734175,0.65643674,0.46026024,0.30935526,0.23767537,0.23767537,0.2678564,0.24899325,0.23767537,0.24899325,0.24522063,0.27540162,0.33953625,0.422534,0.52439487,0.66775465,0.66020936,0.67152727,0.73566186,0.80734175,0.7582976,0.6828451,0.60362,0.5696664,0.6111652,0.72811663,0.65643674,0.58098423,0.45648763,0.3055826,0.19994913,0.15845025,0.14713238,0.15845025,0.181086,0.18485862,0.20372175,0.21503963,0.241448,0.29803738,0.3961256,0.452715,0.63002837,0.6828451,0.59230214,0.56212115,0.5696664,0.47535074,0.43385187,0.4640329,0.45648763,0.42630664,0.5017591,0.6413463,0.76207024,0.7507524,0.6073926,0.5885295,0.5696664,0.5394854,0.6149379,0.65643674,0.5885295,0.543258,0.573439,0.66020936,0.513077,0.4376245,0.44139713,0.47912338,0.452715,0.452715,0.4074435,0.38480774,0.422534,0.4979865,0.4678055,0.47535074,0.4979865,0.5281675,0.5696664,0.59607476,0.62248313,0.63002837,0.6413463,0.7167987,0.6451189,0.5885295,0.60362,0.68661773,0.7809334,0.91674787,0.95447415,0.9205205,0.84129536,0.73188925,0.724344,0.69039035,0.6375736,0.5772116,0.5583485,0.44894236,0.38858038,0.38103512,0.41876137,0.48666862,0.5017591,0.52062225,0.5017591,0.46026024,0.47912338,0.49044126,0.47912338,0.47157812,0.482896,0.51684964,0.5583485,0.60362,0.56212115,0.47912338,0.5017591,0.56212115,0.58098423,0.58098423,0.5772116,0.58475685,0.633801,0.6752999,0.7205714,0.784706,0.87902164,0.95824677,1.116697,1.3166461,1.5316857,1.7429527,1.7882242,1.8523588,1.871222,1.7882242,1.5882751,1.3732355,1.3694628,1.3543724,1.3204187,1.4750963,1.5807298,1.6524098,1.7957695,1.9844007,2.0598533,1.9994912,1.8259505,1.6750455,1.5807298,1.4939595,1.5128226,1.5543215,1.5618668,1.5618668,1.6486372,1.6222287,1.6184561,1.6109109,1.6222287,1.7429527,2.1164427,2.5427492,2.8822856,3.0822346,3.1539145,0.056589376,0.011317875,0.0,0.00754525,0.030181,0.08677038,0.12826926,0.17354076,0.211267,0.211267,0.1056335,0.09808825,0.09808825,0.09808825,0.124496624,0.22258487,0.15845025,0.071679875,0.05281675,0.10940613,0.13958712,0.14335975,0.271629,0.31312788,0.20372175,0.0,0.0150905,0.060362,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,1.0638802,2.9803739,4.5233774,3.3878171,1.8070874,1.0412445,0.76207024,0.6111652,0.20372175,0.4640329,0.45648763,0.41498876,0.5319401,0.94315624,0.9808825,0.73566186,0.6790725,0.83752275,0.7997965,0.6488915,0.9922004,1.3053282,1.5015048,1.9051756,2.7313805,3.3123648,4.183841,4.6629643,2.867195,2.3993895,2.233394,2.1202152,2.052308,2.2711203,1.7316349,3.0407357,5.372218,7.809334,9.333474,14.849052,13.860624,10.110635,6.115425,3.150142,1.3468271,1.7354075,2.2975287,2.4861598,3.2331395,3.5689032,2.595566,2.3993895,3.663219,5.6778007,6.8737226,8.473316,10.140816,11.329193,11.291467,11.815862,12.551523,12.385528,11.502733,11.389555,10.133271,7.7187905,5.643847,4.5761943,4.3649273,2.8936033,2.4861598,2.8709676,3.5651307,3.8820312,4.436607,6.398372,8.13378,8.865668,8.661947,8.345046,8.303548,7.835742,6.888813,6.043745,5.8664317,4.715781,4.908185,6.983129,9.699419,9.314611,8.386545,7.5905213,8.058327,11.3820095,13.181552,11.32542,11.664956,15.316857,18.685812,20.515535,24.378702,26.834682,27.287397,27.974014,28.373913,26.812046,23.09601,18.599041,16.244923,18.006739,20.300495,21.187061,19.953413,17.139036,15.445127,14.905642,15.30554,15.471535,13.264549,9.322156,10.299266,14.053028,23.386503,46.044888,61.131615,46.16561,23.322369,7.2170315,4.8666863,7.1981683,9.574923,12.642066,15.339493,14.905642,10.340765,6.9454026,10.419991,18.71222,22.013268,15.347038,13.479589,13.9888935,14.120935,10.804798,9.654147,9.8239155,10.246449,10.450171,10.567122,11.623458,10.668983,9.88805,10.79348,14.222796,19.1008,17.89356,16.048746,16.248695,18.376457,17.448391,16.72782,16.965494,17.91997,18.365139,18.448135,20.82489,27.559025,36.583145,41.672417,34.11585,27.698612,23.288414,21.258741,21.45869,23.145054,26.419693,39.978508,60.746807,73.868,67.133865,63.14997,56.219658,44.203846,28.487091,20.187317,14.452927,9.820143,5.745708,2.6106565,1.4637785,1.6486372,1.5505489,0.8337501,0.42630664,1.1280149,0.8941121,0.90920264,1.5920477,2.5691576,2.6182017,7.462252,17.836971,29.354795,32.53889,12.694883,7.805561,9.133525,12.7477,19.523335,27.630705,28.275824,26.431011,25.627441,27.940062,25.12191,19.247932,17.372938,19.372429,17.946377,15.803526,16.765545,19.11589,20.296722,16.931541,18.663176,18.87067,19.727057,20.8513,19.31584,19.583696,22.828154,25.616123,27.66466,31.825865,29.860327,27.366621,26.24238,25.604805,21.798227,20.179771,20.138271,20.756983,23.062057,30.033867,35.157093,33.47073,28.8304,24.85028,24.888006,26.246153,25.75571,30.086685,38.27328,41.717686,42.992836,46.644737,47.829338,45.833622,44.06803,43.479504,39.016487,33.836674,29.581152,26.385738,22.401848,17.482344,13.328684,10.137043,6.6058664,4.2517486,3.0407357,2.4333432,2.0787163,1.8146327,3.0445085,5.7381625,9.009028,11.359374,10.687846,8.597813,5.3684454,5.855114,9.246704,9.061845,7.809334,5.7909794,6.296511,9.175024,10.834979,8.695901,10.63503,13.837989,15.577168,13.192869,21.522825,16.28265,9.114662,6.1418333,7.9791017,5.587258,3.2746384,3.399135,5.5004873,6.2851934,4.6931453,6.156924,9.208978,10.412445,4.3724723,5.945657,10.0465,12.596795,12.083718,9.57115,6.4247804,4.930821,4.032936,3.8593953,5.726845,11.98563,10.808571,6.9567204,4.002755,4.323428,3.4745877,4.3007927,5.2326307,6.066381,7.9489207,10.03141,8.612903,6.304056,5.05909,6.198423,6.085244,5.523123,5.9003854,7.039718,7.201941,7.5829763,8.382772,8.6732645,9.073163,11.732863,12.559069,13.754991,14.543469,13.649357,9.295748,9.484379,11.378237,13.415455,15.007503,16.524097,20.68153,20.949387,18.402864,14.351066,10.310584,6.7039547,5.745708,7.986647,11.6875925,12.777881,11.578186,10.782163,10.016319,8.446907,4.779916,4.146115,3.742444,4.1008434,4.825187,4.5912848,5.4438977,6.9491754,6.3832817,3.6254926,1.1431054,1.0751982,0.6413463,0.49044126,0.784706,1.1883769,0.8299775,0.69039035,0.70170826,0.8978847,1.4222796,1.9579924,2.3805263,2.7351532,3.059599,3.3651814,3.3123648,2.3126192,2.003264,2.897376,4.402653,4.979865,6.149379,5.956975,4.5988297,4.4215164,4.1989317,3.3425457,2.9426475,3.2105038,3.4745877,3.0860074,2.6785638,2.746471,3.1539145,3.1199608,3.6330378,2.9351022,1.8938577,1.1695137,1.2185578,1.3694628,0.87147635,0.52439487,0.69793564,1.3015556,0.9695646,0.67152727,0.573439,0.62248313,0.5319401,0.452715,0.35085413,0.24899325,0.15845025,0.056589376,0.041498873,0.094315626,0.18863125,0.2565385,0.18485862,0.060362,0.049044125,0.08299775,0.116951376,0.150905,0.09808825,0.06413463,0.049044125,0.03772625,0.02263575,0.018863125,0.05281675,0.15467763,0.2678564,0.27917424,0.15845025,0.06413463,0.018863125,0.02263575,0.03772625,0.018863125,0.02263575,0.02263575,0.011317875,0.0150905,0.0150905,0.03772625,0.03772625,0.0150905,0.011317875,0.041498873,0.0452715,0.060362,0.08677038,0.08677038,0.094315626,0.24899325,0.35462674,0.32444575,0.18863125,0.15845025,0.094315626,0.06790725,0.09808825,0.13958712,0.03772625,0.056589376,0.13958712,0.24522063,0.33953625,0.44139713,0.5017591,0.5772116,0.66775465,0.7092535,0.77338815,0.60362,0.38103512,0.2263575,0.19240387,0.21503963,0.211267,0.20749438,0.21881226,0.24522063,0.2678564,0.3169005,0.43007925,0.60362,0.7922512,0.7394345,0.69039035,0.72811663,0.80356914,0.754525,0.76584285,0.6790725,0.5696664,0.51684964,0.5998474,0.7884786,0.7884786,0.55080324,0.23390275,0.18863125,0.14335975,0.120724,0.12826926,0.150905,0.16222288,0.18485862,0.181086,0.19240387,0.2678564,0.422534,0.3772625,0.422534,0.51684964,0.5885295,0.52062225,0.52062225,0.40367088,0.32067314,0.30935526,0.30935526,0.38480774,0.55457586,0.76584285,0.935611,0.935611,0.8262049,0.7394345,0.67152727,0.63002837,0.63002837,0.66020936,0.56589377,0.47157812,0.452715,0.5319401,0.41121614,0.3772625,0.4074435,0.452715,0.44139713,0.43007925,0.452715,0.45648763,0.44139713,0.44516975,0.44516975,0.47157812,0.513077,0.5583485,0.58475685,0.49044126,0.5281675,0.55080324,0.5281675,0.5394854,0.6413463,0.56589377,0.543258,0.6451189,0.7922512,0.845068,0.8224323,0.7696155,0.7054809,0.6073926,0.56589377,0.56212115,0.5281675,0.452715,0.39989826,0.331991,0.36971724,0.39989826,0.40367088,0.42630664,0.55080324,0.6488915,0.6375736,0.543258,0.49421388,0.47535074,0.4376245,0.42630664,0.44516975,0.4640329,0.4376245,0.43385187,0.41876137,0.392353,0.362172,0.422534,0.4376245,0.44894236,0.49421388,0.5583485,0.56589377,0.59230214,0.6149379,0.633801,0.68661773,0.7092535,0.80734175,0.91674787,0.9922004,0.995973,1.2713746,1.6448646,1.8372684,1.7995421,1.6788181,1.448688,1.3845534,1.3355093,1.2826926,1.3543724,1.4298248,1.5656394,1.81086,2.052308,2.0296721,1.8636768,1.7655885,1.659955,1.5430037,1.5052774,1.5580941,1.5165952,1.4600059,1.448688,1.50905,1.5165952,1.5618668,1.5430037,1.4939595,1.5845025,1.7278622,1.9579924,2.233394,2.41448,2.2447119,0.030181,0.00754525,0.0,0.030181,0.060362,0.0,0.10940613,0.1659955,0.16976812,0.1659955,0.21503963,0.13958712,0.049044125,0.049044125,0.124496624,0.1358145,0.11317875,0.1056335,0.10186087,0.1056335,0.150905,0.116951376,0.116951376,0.09808825,0.049044125,0.0,0.02263575,0.02263575,0.00754525,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.011317875,0.5281675,3.4029078,7.33021,7.8432875,4.927048,2.372981,0.995973,0.694163,0.47157812,0.30181,0.452715,0.52062225,0.5017591,0.80734175,1.6260014,1.2261031,0.62248313,0.31312788,0.27540162,0.6526641,1.5731846,2.1466236,2.3314822,2.9313297,3.8443048,4.266839,3.8254418,2.6597006,1.388326,1.841041,2.1541688,1.9542197,1.4411428,1.4034165,2.233394,4.191386,5.7419353,6.2436943,5.9494295,10.819888,9.322156,6.1116524,3.4066803,0.97710985,1.1959221,1.599593,2.4786146,3.6594462,4.5007415,3.4029078,2.897376,3.6934,5.824933,8.68081,8.707218,8.729855,9.420244,10.533169,10.925522,11.144334,10.725573,9.623966,8.43559,8.36391,6.7152724,5.515578,5.7570257,7.232122,8.514814,5.3156285,4.2404304,4.236658,4.52715,4.640329,4.5422406,4.398881,4.2894745,4.4516973,5.281675,6.7680893,6.858632,6.428553,5.775889,4.5912848,4.2894745,3.9084394,4.6290107,6.903904,10.469034,9.918231,7.9225125,6.3531003,6.3531003,8.329956,11.125471,9.639057,8.809079,10.506761,13.536179,19.25925,24.133482,26.434784,26.408375,26.276333,24.529608,21.05502,15.731846,10.751981,10.604849,12.521342,13.449409,12.453435,10.155907,8.729855,9.582467,10.344538,11.589504,12.325166,9.993684,6.930312,8.537451,11.16697,14.060574,19.334703,19.28566,16.105335,11.087745,6.6850915,6.515323,8.835487,11.61214,13.913441,14.4152,11.41219,8.473316,7.2962565,14.094527,26.102793,31.569326,20.60985,15.441354,14.245432,13.7851715,9.416472,9.805053,10.480352,11.174516,11.887542,12.864652,13.3626375,12.189351,12.261031,14.030393,15.456445,17.482344,17.010767,16.418465,16.535416,16.633503,17.022083,18.301004,18.94235,18.719765,18.708447,18.391546,17.595524,19.953413,25.231316,29.343477,27.159128,23.809036,20.300495,17.82188,17.761518,17.003222,24.156118,44.13594,69.20503,78.994995,58.12106,43.54741,33.542408,25.487854,15.856343,11.302785,6.1908774,3.3161373,2.6106565,1.1581959,0.6488915,1.0789708,1.1016065,0.513077,0.24522063,0.7696155,0.935611,2.41448,4.851596,5.8890676,4.8138695,9.627739,20.085455,30.939297,31.950361,13.396591,7.586749,7.9791017,11.732863,19.73083,32.010723,32.772793,29.849009,28.502182,31.433512,30.860073,23.646814,19.813826,21.304014,21.986858,19.61765,20.153362,21.911406,22.254715,17.57666,18.029375,18.957441,21.092747,23.163918,21.881226,20.232588,23.435547,28.034376,33.463184,42.068542,37.12263,32.829384,31.180746,30.780848,26.838455,22.213217,21.047476,19.715738,19.217752,25.163408,33.98758,33.98758,30.471493,26.962952,25.19359,24.178753,24.933279,28.566317,33.35755,34.760967,36.054977,37.111313,38.326096,39.14853,38.08465,41.39324,40.42745,37.42444,33.915897,30.731804,25.763256,20.575897,16.546734,13.2607765,8.499724,5.081726,3.6330378,3.4670424,3.4632697,2.0598533,1.7542707,2.8143783,5.907931,9.491924,9.797507,8.280911,4.919503,3.6443558,5.2779026,7.5226145,7.9489207,4.5497856,4.104616,7.7225633,10.834979,7.673519,10.597303,13.015556,12.449662,10.544487,15.071637,12.166716,8.088508,6.085244,6.379509,4.9760923,4.285702,4.8930945,6.039973,5.5985756,3.4029078,2.9728284,6.828451,11.574413,7.888559,14.539697,14.188843,12.034674,9.88805,6.1644692,3.3312278,3.5123138,3.8254418,3.8103511,5.4476705,12.709973,13.272095,11.038701,8.231868,5.3873086,2.5540671,2.7879698,5.2364035,8.888305,12.58925,14.652876,15.358356,14.792462,13.826671,14.143571,10.020092,6.971811,5.66271,5.775889,6.043745,6.2851934,7.043491,7.4018903,7.435844,8.179051,9.876732,12.936331,15.267814,14.728328,9.125979,7.0510364,6.9982195,7.7678347,8.586494,9.125979,10.982111,12.917468,12.789199,11.299012,11.993175,9.601331,7.858378,8.213005,9.774872,9.322156,13.472044,13.430545,11.099063,7.99042,5.2175403,5.036454,4.9345937,4.52715,3.5877664,2.0749438,2.1503963,3.2029586,3.3123648,2.0598533,0.5357128,0.29049212,0.33953625,0.51684964,0.8941121,1.7844516,1.418507,1.0072908,0.90920264,1.1280149,1.3128735,1.7995421,1.8599042,2.0975795,2.9011486,4.4403796,3.9273026,2.2447119,1.1732863,1.1204696,1.0827434,2.1579416,3.2218218,3.6556737,3.3727267,2.8219235,3.712263,3.3689542,2.6182017,2.1164427,2.3503454,2.0673985,2.2447119,2.4974778,2.546522,2.2296214,3.5839937,3.5839937,2.674791,1.6071383,1.448688,1.4750963,0.95824677,0.55457586,0.6526641,1.3732355,1.1431054,0.69039035,0.44516975,0.47157812,0.45648763,0.31312788,0.18485862,0.12826926,0.116951376,0.030181,0.056589376,0.08677038,0.124496624,0.150905,0.1358145,0.041498873,0.0150905,0.026408374,0.041498873,0.030181,0.090543,0.124496624,0.120724,0.08677038,0.060362,0.02263575,0.02263575,0.03772625,0.08299775,0.23013012,0.1659955,0.08677038,0.041498873,0.02263575,0.0,0.011317875,0.0150905,0.00754525,0.003772625,0.0150905,0.0150905,0.02263575,0.02263575,0.011317875,0.0,0.0,0.026408374,0.05281675,0.06413463,0.0754525,0.05281675,0.0452715,0.08299775,0.150905,0.21503963,0.1659955,0.08677038,0.05281675,0.056589376,0.030181,0.00754525,0.03772625,0.090543,0.1659955,0.29049212,0.362172,0.39989826,0.49044126,0.62625575,0.68661773,0.7469798,0.6451189,0.44139713,0.25276586,0.23013012,0.20372175,0.181086,0.181086,0.20749438,0.24522063,0.2565385,0.3055826,0.38480774,0.4979865,0.65643674,0.694163,0.6752999,0.6149379,0.5583485,0.59607476,0.65643674,0.62625575,0.5885295,0.56212115,0.48666862,0.6111652,0.79602385,0.663982,0.2867195,0.21503963,0.17731337,0.15845025,0.13958712,0.124496624,0.1358145,0.16222288,0.17731337,0.17731337,0.20372175,0.35085413,0.362172,0.392353,0.47912338,0.5583485,0.47157812,0.3734899,0.31312788,0.27917424,0.26031113,0.26031113,0.44139713,0.72811663,0.95824677,1.0940613,1.1883769,1.1431054,0.97333723,0.80356914,0.6790725,0.59607476,0.72811663,0.663982,0.51684964,0.4074435,0.45648763,0.44516975,0.46026024,0.46026024,0.44139713,0.44139713,0.43007925,0.47157812,0.52062225,0.5319401,0.45648763,0.45648763,0.44894236,0.4376245,0.4640329,0.6111652,0.47535074,0.48666862,0.55457586,0.5998474,0.56589377,0.8224323,0.7922512,0.6526641,0.5357128,0.5357128,0.7054809,0.6375736,0.55080324,0.52062225,0.47157812,0.362172,0.33576363,0.3772625,0.46026024,0.5357128,0.35085413,0.3772625,0.3961256,0.3772625,0.48666862,0.56212115,0.663982,0.663982,0.56589377,0.52062225,0.52062225,0.47157812,0.41121614,0.36594462,0.36594462,0.392353,0.35839936,0.3169005,0.30181,0.35085413,0.362172,0.3470815,0.3470815,0.3734899,0.41121614,0.39989826,0.452715,0.513077,0.5772116,0.68661773,0.7469798,0.7167987,0.73566186,0.8111144,0.8224323,1.0940613,1.4260522,1.6146835,1.6410918,1.6788181,1.50905,1.327964,1.2223305,1.146878,0.91674787,0.9393836,1.1393328,1.4071891,1.6750455,1.9089483,1.6637276,1.6561824,1.6260014,1.478869,1.297783,1.3694628,1.2864652,1.20724,1.177059,1.1280149,1.3732355,1.50905,1.4600059,1.327964,1.388326,1.6675003,1.9768555,2.2899833,2.4861598,2.3654358,0.00754525,0.0,0.0,0.00754525,0.011317875,0.0,0.02263575,0.15845025,0.22258487,0.181086,0.13958712,0.049044125,0.14335975,0.14335975,0.026408374,0.026408374,0.120724,0.12826926,0.07922512,0.02263575,0.030181,0.02263575,0.13204187,0.14335975,0.041498873,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.116951376,0.9695646,3.1765501,7.232122,6.6586833,3.6254926,1.1695137,0.36971724,0.31312788,0.13204187,0.35462674,0.46026024,0.482896,0.9922004,1.8674494,1.7089992,1.0601076,0.49421388,0.60362,1.5505489,2.6446102,3.429316,3.712263,3.5764484,3.2331395,2.6936543,2.1579416,1.7354075,1.4600059,1.327964,1.297783,1.2336484,1.3543724,2.233394,3.3161373,5.564622,7.2962565,8.190369,9.2844305,11.00852,8.194141,4.5309224,2.0183544,0.965792,1.3317367,2.252257,3.4066803,4.3196554,4.3913355,3.3727267,4.293247,6.8397694,9.978593,11.966766,11.940358,10.152134,8.684583,8.590267,9.88805,9.005256,7.405663,5.926794,5.0553174,4.9459114,3.9688015,4.3686996,5.3571277,6.096562,5.670255,3.7009451,3.0897799,2.9501927,2.8332415,2.6974268,2.9124665,2.746471,2.2107582,1.7429527,2.191895,2.9954643,3.0897799,3.429316,4.0480266,4.044254,3.1237335,3.5575855,4.5761943,5.6363015,6.428553,6.8359966,5.4891696,4.6818275,5.4740787,7.6848373,9.6201935,10.846297,11.559323,12.310076,14.000212,17.222033,18.395319,17.538933,15.754482,15.230087,14.283158,12.393073,10.887795,10.042727,9.0543,10.072908,10.54826,10.559577,10.242677,9.80128,9.680555,10.103089,10.1294985,9.073163,6.515323,5.9720654,8.578949,11.072655,11.827179,10.861387,13.479589,15.988385,17.003222,15.580941,11.23865,11.838497,13.834216,15.286676,14.750964,11.2801485,9.22784,9.291975,11.348056,13.95494,14.347293,12.1252165,12.849561,13.951167,14.437836,14.871688,14.381247,13.505998,13.038192,13.404137,14.634012,15.701665,17.7502,19.074392,18.919714,17.508753,16.029884,16.429781,17.923742,18.55377,15.203679,17.1164,18.75372,19.319613,19.217752,20.074137,19.247932,17.53139,16.731592,16.991903,16.769318,14.320885,13.521088,13.924759,15.328176,17.799244,19.266796,22.356575,34.17621,55.3595,80.07019,61.950275,48.18774,37.23581,28.294687,21.311558,16.316603,8.028146,3.3161373,3.270866,3.1727777,1.8523588,1.8221779,1.5279131,0.6526641,0.120724,0.95824677,1.7316349,2.2975287,3.2935016,6.145606,8.714764,14.618922,21.715229,25.842482,20.832436,8.986393,5.160951,5.2175403,7.413208,12.381755,25.608578,29.596243,27.668432,24.412657,25.68403,33.636726,31.807001,25.182272,21.081429,29.177483,24.348522,24.371157,24.544699,22.877197,20.055275,22.813063,22.198126,22.745155,25.227543,26.676231,23.514772,24.34475,29.407612,38.650543,51.700054,44.49811,39.83892,36.95286,35.160866,33.881947,26.287651,24.620152,23.473272,22.062311,24.24666,33.01424,33.063286,29.95087,28.238098,31.51651,26.457418,24.838963,26.261242,30.003687,35.040142,33.474503,32.55398,32.606796,33.968716,36.998135,39.310753,39.816284,39.00517,37.137722,34.2328,27.400576,21.851044,17.64834,14.305794,10.744436,7.0359454,5.1835866,4.3875628,3.9725742,3.3764994,2.9086938,2.5917933,3.029418,4.6856003,7.8923316,7.394345,4.315883,2.4522061,3.5085413,7.069899,5.20245,5.142088,5.379763,5.915476,8.246958,13.102326,14.4152,13.917213,11.940358,7.4207535,10.970794,10.774617,8.888305,7.8206515,10.514306,7.9489207,5.7381625,4.398881,4.0178456,4.2819295,2.8558772,3.187868,7.0963078,12.042219,11.148107,9.265567,8.224322,8.190369,8.00551,5.198677,3.2067313,3.180323,2.8634224,2.3126192,3.9084394,11.046246,11.012292,9.774872,9.22784,7.194396,3.9310753,3.6783094,6.5832305,10.514306,11.050018,12.868423,13.970031,14.807553,15.339493,15.011275,9.714509,6.3531003,5.4401255,6.2851934,6.9944468,5.5683947,5.3948536,6.006019,6.7831798,6.983129,6.092789,7.654656,10.042727,10.725573,6.304056,3.5839937,3.0558262,3.1237335,3.1048703,3.240685,5.3609,7.432071,7.8244243,7.0510364,7.745199,7.141579,5.6551647,5.353355,6.609639,8.088508,12.581704,14.84528,13.928532,10.397354,6.330465,4.3875628,3.942393,4.1536603,3.9310753,1.9278114,1.2298758,1.7769064,2.1202152,1.690136,0.7922512,0.47912338,0.68661773,0.7696155,0.68661773,0.9922004,1.3770081,1.0450171,0.7394345,0.7054809,0.6526641,0.60362,0.7394345,1.1016065,1.6486372,2.2673476,3.1916409,3.7688525,3.2557755,2.0560806,1.7165444,2.7615614,2.4823873,2.3918443,2.7238352,2.4182527,3.2520027,2.8709676,2.305074,1.991946,1.7769064,2.1503963,2.071171,2.3428001,2.8709676,2.6898816,3.0407357,2.9501927,2.516341,1.9391292,1.5467763,1.4637785,1.0374719,0.6413463,0.56589377,1.0299267,1.0525624,0.754525,0.5281675,0.5055317,0.543258,0.3961256,0.21881226,0.12826926,0.116951376,0.041498873,0.026408374,0.030181,0.041498873,0.06790725,0.11317875,0.0754525,0.041498873,0.0452715,0.06790725,0.06790725,0.049044125,0.116951376,0.13958712,0.08677038,0.02263575,0.00754525,0.003772625,0.011317875,0.049044125,0.1659955,0.1358145,0.056589376,0.00754525,0.003772625,0.0,0.003772625,0.003772625,0.00754525,0.011317875,0.003772625,0.011317875,0.018863125,0.011317875,0.003772625,0.0,0.011317875,0.033953626,0.041498873,0.041498873,0.05281675,0.056589376,0.041498873,0.03772625,0.049044125,0.07922512,0.090543,0.10940613,0.120724,0.10186087,0.018863125,0.0150905,0.026408374,0.06413463,0.120724,0.19240387,0.3055826,0.35839936,0.41876137,0.543258,0.77338815,0.69793564,0.56589377,0.47535074,0.422534,0.30181,0.23767537,0.18863125,0.17354076,0.1961765,0.23013012,0.271629,0.32821837,0.3961256,0.46026024,0.52062225,0.73566186,0.7167987,0.66020936,0.6413463,0.6187105,0.60362,0.6752999,0.7507524,0.7432071,0.56212115,0.70170826,0.7054809,0.5319401,0.27540162,0.1659955,0.116951376,0.120724,0.13958712,0.16222288,0.17354076,0.15845025,0.18863125,0.21503963,0.24522063,0.30181,0.5093044,0.58098423,0.55457586,0.4979865,0.5093044,0.452715,0.331991,0.26408374,0.27540162,0.34330887,0.5470306,0.7130261,0.8526133,0.94692886,0.95824677,1.0751982,1.0676528,0.90543,0.694163,0.65643674,0.5357128,0.41876137,0.3734899,0.36971724,0.31312788,0.33953625,0.36971724,0.39989826,0.44516975,0.55080324,0.44139713,0.3961256,0.38480774,0.3772625,0.32444575,0.35462674,0.36594462,0.3772625,0.43385187,0.5998474,0.5998474,0.5281675,0.47912338,0.5093044,0.6375736,0.7884786,0.754525,0.663982,0.6149379,0.694163,0.80356914,0.7507524,0.633801,0.5281675,0.4979865,0.3470815,0.3055826,0.39989826,0.5470306,0.5357128,0.28294688,0.1961765,0.1961765,0.23767537,0.32821837,0.34330887,0.38480774,0.41876137,0.4376245,0.44516975,0.543258,0.47912338,0.38858038,0.35462674,0.41498876,0.46026024,0.44139713,0.422534,0.42630664,0.4376245,0.4376245,0.4074435,0.36594462,0.3470815,0.362172,0.38858038,0.422534,0.46026024,0.513077,0.6149379,0.73188925,0.77716076,0.754525,0.7130261,0.72811663,0.91674787,1.0676528,1.1695137,1.2185578,1.2261031,1.1732863,1.116697,1.0789708,1.0827434,1.1732863,1.3619176,1.4260522,1.4222796,1.4411428,1.6146835,1.8787673,1.780679,1.6071383,1.4864142,1.3694628,1.4335974,1.3920987,1.2751472,1.1619685,1.1883769,1.3656902,1.569412,1.6788181,1.6260014,1.4147344,1.4411428,1.8599042,2.4597516,2.9086938,2.7691069,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.18485862,0.2263575,0.1659955,0.1056335,0.10186087,0.1056335,0.08677038,0.056589376,0.06413463,0.060362,0.05281675,0.049044125,0.0452715,0.03772625,0.00754525,0.056589376,0.06413463,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.033953626,0.20372175,1.5354583,5.7607985,7.91874,5.168496,1.9579924,0.392353,0.21881226,0.060362,0.18863125,0.34330887,0.4979865,0.8563859,1.3505998,1.1883769,0.754525,0.44516975,0.66020936,2.3767538,3.1199608,3.229367,3.048281,2.916239,2.4107075,1.9127209,1.4826416,1.1732863,1.0299267,1.116697,1.2261031,1.327964,1.5769572,2.2862108,3.6896272,6.089017,7.99042,9.020347,9.9257765,8.446907,5.413717,3.150142,2.3428001,2.0145817,3.097325,3.942393,4.376245,4.2027044,3.2105038,3.2784111,4.3913355,6.417235,8.537451,9.242931,9.250477,8.20546,7.4094353,7.677292,9.325929,8.028146,5.9796104,4.3686996,3.4594972,2.6068838,2.2409391,2.8181508,3.6292653,4.074435,3.6594462,2.8030603,2.4823873,2.1541688,1.7391801,1.6184561,1.931584,1.9278114,1.8448136,1.901403,2.2975287,2.41448,1.991946,1.8636768,2.335255,3.1916409,3.5990841,4.323428,5.534441,6.7831798,7.0170827,6.647365,5.8513412,5.20245,5.1760416,6.149379,6.9680386,9.110889,10.329447,10.03141,9.273112,10.005001,9.559832,8.145098,6.7869525,7.322665,8.00551,8.080963,8.907167,10.099318,9.5183325,9.703192,9.842778,10.27663,10.627484,9.797507,9.567377,9.771099,9.88805,9.450426,8.062099,8.544995,10.167224,11.8045435,12.00072,9.001483,10.804798,13.04951,15.505488,16.463736,12.740154,10.933067,10.797253,11.204697,10.929295,8.635539,8.899622,10.687846,11.951676,12.162943,12.347801,14.381247,14.32843,13.626721,13.532406,15.147089,15.339493,14.505743,13.856852,14.449154,17.206944,20.37972,21.028612,19.628967,18.029375,19.4592,17.87847,17.580433,18.500954,19.289433,17.327667,18.157644,17.421982,17.074902,17.7502,18.749947,18.23687,19.500698,18.666948,15.335721,12.574159,11.517824,11.314102,11.996947,14.034165,18.327412,24.27307,26.219744,32.15031,44.80747,61.69751,57.151497,49.59493,40.940525,33.474503,29.860327,25.944342,16.856089,10.484125,8.816625,7.9262853,3.7348988,2.1503963,2.3465726,2.806833,1.3091009,1.3694628,2.161714,2.71629,3.0105548,3.9763467,5.383536,10.570895,18.323639,28.004196,39.574837,19.598787,8.228095,5.0213637,6.858632,7.907422,14.735873,19.029121,19.43279,18.644312,23.420456,35.232544,38.846718,33.78763,26.608324,30.875162,29.494383,26.680004,23.775084,22.315077,24.008986,26.61587,25.865116,27.604298,31.67496,31.916407,26.845999,26.268787,30.064049,37.416893,46.829594,40.031322,37.028313,36.156837,36.60201,38.409096,31.886227,28.468227,26.763002,26.012249,26.087702,28.57009,28.287142,26.547962,24.92196,25.22377,21.439827,21.967995,25.253952,28.637997,28.362595,26.981813,26.891272,28.064558,30.211182,32.799202,34.72324,36.368107,38.046925,38.68827,35.832394,29.573606,24.812555,21.134245,18.923487,19.353567,11.812089,9.06939,7.2057137,4.8742313,3.3048196,3.3350005,2.897376,2.6182017,3.289729,5.885295,5.2326307,3.742444,2.474842,3.108643,7.9451485,5.6363015,10.401127,11.604594,8.224322,8.843033,17.395575,17.30503,13.177779,8.345046,4.851596,10.035183,12.736382,10.340765,5.8890676,8.073418,9.21275,7.745199,5.764571,4.293247,3.2746384,2.6144292,4.323428,7.8432875,11.581959,12.932558,7.884786,6.3531003,6.579458,6.779407,5.1345425,3.6669915,2.8256962,2.1202152,2.0673985,4.1762958,11.249968,11.442371,11.389555,12.257258,9.767326,6.63982,5.692891,6.541732,8.122461,8.707218,10.684074,11.981857,13.502225,14.7736,13.947394,10.955703,7.8319697,5.7381625,5.4250345,7.224577,6.273875,4.9421387,4.429062,4.7308717,4.659192,3.6858547,3.6707642,4.425289,4.90064,3.1916409,1.7542707,1.9881734,2.746471,3.1161883,2.4182527,4.4441524,5.881522,6.092789,5.3194013,4.67051,4.4441524,3.5990841,3.4783602,4.5535583,6.40969,9.559832,12.762791,13.875714,11.989402,7.4396167,5.036454,3.5387223,3.399135,3.9197574,3.2821836,1.7127718,1.7769064,2.123988,2.637065,4.432834,1.81086,1.3204187,1.3053282,1.0902886,0.98465514,1.5656394,1.3053282,0.8865669,0.68661773,0.7432071,0.48666862,0.47157812,0.6790725,0.9507015,0.97333723,1.5467763,2.7087448,2.8822856,2.1692593,2.372981,4.1574326,3.4255435,3.1954134,3.7537618,2.674791,2.5578396,2.987919,3.2029586,2.746471,1.4600059,1.9504471,1.7618159,1.841041,2.372981,2.7615614,2.214531,1.9806281,1.7580433,1.4713237,1.2600567,1.2751472,1.0940613,0.76584285,0.48666862,0.633801,1.0072908,0.814887,0.56589377,0.4979865,0.59230214,0.4074435,0.23013012,0.13958712,0.13204187,0.120724,0.056589376,0.02263575,0.011317875,0.033953626,0.08677038,0.07922512,0.041498873,0.033953626,0.049044125,0.056589376,0.056589376,0.1961765,0.19240387,0.041498873,0.00754525,0.09808825,0.120724,0.0754525,0.018863125,0.071679875,0.06790725,0.033953626,0.003772625,0.0,0.00754525,0.0150905,0.00754525,0.003772625,0.003772625,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.011317875,0.018863125,0.0150905,0.018863125,0.03772625,0.056589376,0.060362,0.0452715,0.026408374,0.026408374,0.03772625,0.05281675,0.06790725,0.06413463,0.02263575,0.02263575,0.02263575,0.041498873,0.090543,0.15845025,0.23767537,0.28294688,0.33953625,0.4376245,0.6187105,0.59607476,0.59230214,0.55457586,0.44894236,0.27540162,0.2678564,0.23390275,0.20372175,0.19994913,0.23767537,0.27917424,0.362172,0.43007925,0.45648763,0.43385187,0.573439,0.6073926,0.6413463,0.6828451,0.6526641,0.6073926,0.6526641,0.73566186,0.7809334,0.69039035,0.845068,0.76584285,0.543258,0.30181,0.20749438,0.17354076,0.13958712,0.120724,0.13204187,0.1659955,0.21503963,0.2565385,0.27917424,0.30181,0.38103512,0.573439,0.62625575,0.62625575,0.6187105,0.6187105,0.4979865,0.35462674,0.27917424,0.331991,0.5394854,0.58098423,0.6375736,0.7922512,0.9507015,0.87147635,0.9280658,1.0223814,0.9016574,0.6375736,0.5998474,0.452715,0.35085413,0.32067314,0.32821837,0.2565385,0.29426476,0.31312788,0.31312788,0.3169005,0.3772625,0.35462674,0.33953625,0.32067314,0.30181,0.29049212,0.33953625,0.39989826,0.47535074,0.5772116,0.73188925,0.66020936,0.56589377,0.5017591,0.52439487,0.7092535,0.80356914,0.7582976,0.694163,0.6752999,0.7130261,0.68661773,0.6526641,0.58475685,0.51684964,0.52062225,0.5319401,0.5319401,0.55457586,0.6451189,0.8262049,0.76207024,0.42630664,0.23013012,0.2678564,0.3169005,0.32444575,0.331991,0.3734899,0.44139713,0.47157812,0.5055317,0.44139713,0.4074435,0.44516975,0.52062225,0.52439487,0.47157812,0.41498876,0.38480774,0.392353,0.422534,0.4376245,0.41121614,0.362172,0.35085413,0.38858038,0.4376245,0.49421388,0.5583485,0.6413463,0.7167987,0.7922512,0.814887,0.7997965,0.8111144,0.9393836,1.0072908,1.0450171,1.0676528,1.0601076,1.0940613,1.1317875,1.0978339,1.0299267,1.0902886,1.3128735,1.4411428,1.4562333,1.4335974,1.5316857,1.6448646,1.6109109,1.569412,1.5580941,1.5241405,1.4562333,1.3241913,1.2185578,1.177059,1.1959221,1.2449663,1.3543724,1.4600059,1.4939595,1.3807807,1.2789198,1.50905,2.0296721,2.5993385,2.757789,0.0,0.0,0.0,0.0,0.0,0.0,0.07922512,0.13204187,0.13204187,0.1056335,0.116951376,0.1056335,0.041498873,0.030181,0.0754525,0.06413463,0.011317875,0.0,0.018863125,0.0452715,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.049044125,0.033953626,0.06790725,0.875249,3.821669,7.673519,6.0739264,2.8181508,0.43385187,0.20749438,0.05281675,0.124496624,0.36971724,0.6451189,0.7432071,0.8262049,0.6149379,0.4376245,0.52439487,1.0450171,2.6974268,3.0181,2.686109,2.263575,2.1881225,1.7542707,1.3920987,1.0450171,0.7432071,0.58475685,0.9808825,1.3920987,1.7844516,2.123988,2.354118,3.9725742,6.300284,7.466025,7.3905725,7.7829256,5.6098933,4.2027044,3.9122121,4.164978,3.4745877,5.168496,6.066381,5.6476197,4.055572,2.0749438,2.9501927,4.112161,5.342037,6.1305156,5.6853456,5.6815734,5.7872066,6.1003346,6.6549106,7.4509344,6.304056,4.8365054,3.7235808,2.9426475,1.780679,1.5580941,1.690136,1.9806281,2.1881225,2.0108092,1.8221779,1.901403,1.7580433,1.3996439,1.3430545,1.4071891,1.3505998,1.5543215,2.0560806,2.5427492,2.372981,1.6071383,0.95824677,0.97710985,2.0673985,3.470815,4.0895257,4.776143,5.587258,5.775889,4.9534564,4.776143,4.5233774,4.13857,4.255521,4.4931965,5.847569,6.670001,6.300284,5.0779533,4.606375,3.7386713,2.8521044,2.516341,3.5047686,4.7308717,5.5004873,6.5568223,7.6886096,7.7225633,8.179051,8.7751255,9.7296,10.540714,9.95973,10.299266,10.785934,11.068882,11.09529,11.106608,11.555551,11.815862,12.238396,12.219532,10.212496,13.65313,18.85558,21.432283,19.25925,12.50248,9.42779,7.8395147,7.454707,7.575431,7.0849895,8.586494,10.665211,11.861133,12.166716,13.04951,15.437581,14.237886,13.287186,14.102073,15.897841,15.614895,15.358356,15.403628,16.392056,19.327158,24.159891,23.710949,20.583443,18.45568,22.100037,20.096773,18.361366,18.62545,20.462717,21.288923,20.126955,17.595524,16.305285,16.758,17.357847,16.4826,19.515789,19.527107,15.701665,13.324911,14.196388,14.166207,15.486626,18.836716,23.314823,32.62566,35.013733,37.126404,42.947563,53.797634,56.517696,51.620827,43.023014,35.738075,35.911617,32.444576,22.918697,14.9358225,11.551778,11.283921,9.993684,5.3458095,3.7499893,5.119452,2.8709676,1.871222,2.3880715,3.9008942,5.8966126,7.8696957,11.287694,11.295239,13.562587,21.4436,35.96821,18.006739,7.9828744,5.5495315,7.281166,6.700182,7.432071,9.5032425,11.091517,13.283413,20.036411,34.46293,44.071804,43.01547,34.715694,31.852272,33.206646,29.535881,25.676485,24.69183,27.891016,27.030859,26.008476,29.705648,35.93048,35.38345,28.42673,26.751684,28.536135,32.43703,37.58289,34.79115,33.998898,34.644016,36.956635,41.96668,37.307487,31.901318,29.494383,30.343224,31.180746,27.702385,25.842482,24.567333,22.8357,19.606333,17.025856,19.191343,23.937305,27.400576,24.005213,22.567842,23.201643,24.959686,26.955406,28.389004,29.999914,32.357803,35.587173,37.733795,34.772285,29.498156,26.457418,24.382475,23.714722,26.612097,16.463736,13.981348,12.370438,8.726082,4.063117,4.2291126,4.4743333,5.0439997,5.458988,4.5309224,3.7462165,3.2369123,2.6332922,3.1048703,7.3717093,6.175787,11.185833,13.128735,10.740664,10.729345,16.105335,15.192361,11.796998,8.054554,4.436607,8.4544525,12.664702,11.423509,6.0022464,4.5912848,7.8244243,8.75249,7.598067,5.168496,2.8785129,2.3956168,4.6516466,7.3792543,9.740918,12.321393,9.7069645,8.537451,8.065872,7.533932,6.1833324,4.055572,2.8181508,2.3918443,2.9841464,5.119452,11.902632,12.51757,12.815607,13.656902,10.921749,7.8395147,7.1302614,7.066127,6.9567204,7.1566696,9.152389,10.567122,12.219532,13.411682,11.925267,11.031156,9.020347,6.5832305,5.2099953,7.1679873,7.605612,5.8136153,4.115934,3.361409,2.9200118,2.9954643,2.444661,1.81086,1.418507,1.3732355,1.1846043,2.2183034,3.6066296,4.3422914,3.2859564,4.8327327,5.6098933,5.9494295,5.7909794,4.6931453,3.893349,3.259548,3.0671442,3.5575855,4.9119577,6.0512905,8.3525915,10.220041,10.352083,7.7225633,5.674028,3.5877664,2.5691576,3.0218725,4.6516466,3.742444,2.9351022,2.335255,2.686109,5.3571277,2.161714,1.2449663,1.3053282,1.4449154,1.1506506,1.5618668,1.4222796,1.0525624,0.754525,0.83752275,0.6828451,0.6451189,0.7469798,0.8262049,0.5281675,0.51684964,1.2525115,1.659955,1.6788181,2.2598023,4.821415,4.485651,4.1536603,4.2894745,2.897376,1.9994912,2.7879698,3.712263,3.6330378,1.81086,2.022127,1.7693611,1.6260014,1.8900851,2.5616124,1.6410918,1.3241913,1.2261031,1.1242423,0.9507015,0.95447415,0.98465514,0.8111144,0.5093044,0.44516975,0.80356914,0.77716076,0.6187105,0.513077,0.56589377,0.38103512,0.23013012,0.150905,0.15845025,0.22258487,0.11317875,0.0452715,0.018863125,0.02263575,0.05281675,0.056589376,0.030181,0.0150905,0.030181,0.056589376,0.14713238,0.3772625,0.3470815,0.071679875,0.00754525,0.116951376,0.19994913,0.17731337,0.0754525,0.0150905,0.026408374,0.026408374,0.011317875,0.0,0.00754525,0.0150905,0.00754525,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.00754525,0.003772625,0.003772625,0.011317875,0.02263575,0.03772625,0.05281675,0.0452715,0.02263575,0.0150905,0.018863125,0.018863125,0.018863125,0.02263575,0.02263575,0.02263575,0.018863125,0.030181,0.071679875,0.13958712,0.20749438,0.2565385,0.30181,0.36971724,0.49044126,0.5772116,0.58475685,0.5357128,0.4376245,0.2867195,0.3055826,0.271629,0.2263575,0.20749438,0.24522063,0.27917424,0.3470815,0.392353,0.3961256,0.38480774,0.44894236,0.5093044,0.59230214,0.66020936,0.6111652,0.6111652,0.63002837,0.6752999,0.72811663,0.7507524,0.8978847,0.8111144,0.5696664,0.31312788,0.21503963,0.18863125,0.150905,0.116951376,0.1056335,0.12826926,0.19994913,0.26031113,0.29803738,0.34330887,0.4678055,0.5696664,0.573439,0.6149379,0.70170826,0.7054809,0.5093044,0.41498876,0.4074435,0.4979865,0.724344,0.6111652,0.6111652,0.7809334,0.98842776,0.90920264,0.845068,0.9507015,0.8526133,0.5696664,0.5055317,0.3961256,0.31312788,0.2867195,0.28294688,0.23013012,0.26031113,0.26408374,0.24522063,0.2263575,0.2565385,0.33576363,0.35462674,0.32821837,0.28294688,0.28294688,0.36594462,0.4376245,0.5093044,0.59607476,0.7130261,0.663982,0.62625575,0.55457586,0.5017591,0.6073926,0.67152727,0.633801,0.63002837,0.67152727,0.6790725,0.59230214,0.58098423,0.573439,0.55080324,0.5696664,0.6187105,0.6413463,0.66775465,0.7394345,0.90543,1.0827434,0.66775465,0.31312788,0.24522063,0.2565385,0.28294688,0.30935526,0.3470815,0.38858038,0.422534,0.41498876,0.36594462,0.36594462,0.422534,0.45648763,0.452715,0.43385187,0.41498876,0.40367088,0.4074435,0.43385187,0.44516975,0.42630664,0.3961256,0.39989826,0.43007925,0.47535074,0.5357128,0.5998474,0.66020936,0.69039035,0.76207024,0.8262049,0.8601585,0.84884065,0.91297525,0.95447415,0.9620194,0.9507015,0.94315624,1.0072908,1.0450171,1.026154,0.97333723,0.98465514,1.1280149,1.2562841,1.3619176,1.4411428,1.5015048,1.5354583,1.569412,1.6184561,1.6561824,1.599593,1.4222796,1.2298758,1.1431054,1.1544232,1.1581959,1.1204696,1.1280149,1.1695137,1.2034674,1.1732863,1.1695137,1.2864652,1.5920477,1.9957186,2.2711203,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.0452715,0.033953626,0.060362,0.15845025,0.05281675,0.02263575,0.033953626,0.03772625,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.14335975,0.08299775,0.09808825,0.1056335,0.45648763,1.9278114,5.794752,5.7192993,3.169005,0.35462674,0.19994913,0.06790725,0.17354076,0.51684964,0.8639311,0.7582976,0.5696664,0.38858038,0.43007925,0.84129536,1.7089992,2.4371157,2.4899325,2.2409391,1.9278114,1.6675003,1.237421,0.87147635,0.58098423,0.41876137,0.47535074,0.9242931,1.50905,2.1768045,2.686109,2.6106565,4.032936,5.983383,5.9494295,4.429062,4.9232755,4.6742826,5.7004366,6.541732,6.2399216,4.327201,6.2889657,7.809334,7.2094865,4.6214657,1.991946,3.2670932,4.5761943,5.2665844,5.0025005,3.7914882,3.640583,4.1612053,4.67051,4.7535076,4.274384,3.6292653,3.229367,2.987919,2.686109,1.9730829,1.5580941,1.267602,1.116697,1.0110635,0.7130261,0.754525,1.2411937,1.5279131,1.4750963,1.478869,1.1808317,0.86770374,0.94315624,1.4373702,1.9957186,1.9579924,1.1732863,0.392353,0.18863125,0.94315624,2.123988,2.4408884,2.335255,2.1768045,2.2447119,1.7731338,2.0258996,2.3390274,2.474842,2.6295197,3.0105548,3.0935526,3.270866,3.5764484,3.7009451,3.31991,2.6068838,2.3163917,2.5917933,2.969056,3.4670424,3.5689032,3.5085413,3.5462675,3.953711,5.553304,7.066127,8.367682,9.465516,10.518079,11.910177,12.698656,12.570387,12.196897,13.238141,13.389046,13.12119,12.58925,12.298758,13.124963,23.38273,39.857784,43.20033,29.898052,12.294985,9.276885,7.3000293,6.477597,6.7039547,7.6584287,8.544995,9.582467,10.785934,11.996947,12.872196,12.706201,12.257258,14.339747,18.368912,20.330677,18.519815,17.897333,18.255732,19.417702,21.258741,25.521809,25.717985,23.578907,21.881226,24.41643,21.307787,19.263023,20.006231,22.95265,25.186045,22.484844,20.093,18.48209,17.640795,17.074902,16.395828,19.225298,19.87796,17.738882,17.30503,19.236614,19.43279,22.149082,27.343987,30.660124,40.906574,43.47196,42.22699,43.456867,55.880123,58.155014,52.914837,43.422913,35.39854,37.009453,32.286125,23.028103,15.128226,11.46878,11.917723,16.418465,9.378746,5.251494,6.6322746,4.2592936,2.5917933,2.535204,4.8063245,9.0543,13.864397,21.884998,18.395319,12.762791,9.820143,9.876732,5.8211603,5.6476197,6.6586833,7.2698483,6.990674,5.7683434,5.028909,5.8928404,8.922258,14.0983,29.47552,44.607517,49.708107,43.44555,32.9237,35.579628,34.60629,31.852272,29.39252,29.501928,24.382475,23.09601,27.70993,34.79492,35.417404,28.358822,26.031113,26.02734,27.370394,30.51299,33.49714,34.56479,34.798695,36.52278,43.294643,40.167137,33.949852,30.844982,32.69357,36.97927,31.120384,27.068584,25.07664,23.563816,19.108345,15.611122,16.444872,20.06282,23.533634,22.57916,21.009748,22.066084,23.461954,24.382475,25.476536,26.985586,29.384975,32.327625,34.11585,31.701368,27.03463,25.751938,25.544443,25.910389,28.151327,19.010258,17.91997,18.168962,15.192361,6.549277,6.432326,7.250985,8.903395,9.224068,3.9876647,4.666737,3.640583,2.6483827,2.916239,5.138315,6.19465,7.7640624,9.933322,12.351574,14.252977,12.019584,10.748209,11.514051,12.291212,7.964011,5.7494807,9.774872,11.544232,8.318638,3.1237335,4.7006907,7.8998766,8.571404,6.119198,3.4745877,2.3654358,3.8782585,5.6891184,7.4999785,11.050018,13.309821,12.89106,11.672502,10.227587,7.8206515,4.587512,3.731126,3.8141239,4.45547,6.3116016,12.091263,12.796744,12.427027,12.012038,9.631512,6.6247296,6.971811,8.028146,8.216777,7.0284004,8.262049,9.593785,11.012292,11.695138,10.023865,9.303293,8.944894,7.7301087,6.2323766,6.7869525,8.341274,7.17176,5.160951,3.4557245,2.4786146,3.4217708,3.4330888,2.5427492,1.3996439,1.2336484,1.418507,2.6521554,4.104616,4.851596,3.904667,4.8742313,5.2099953,5.96452,6.937857,6.677546,5.1798143,4.429062,3.8556228,3.5500402,4.2404304,3.8971217,4.2630663,5.251494,6.330465,6.5266414,5.3759904,3.904667,2.3805263,1.9504471,4.640329,5.5570765,4.0706625,2.2183034,1.4411428,2.6219745,1.2261031,0.5319401,0.88279426,1.6939086,1.4298248,1.478869,1.4977322,1.2902378,0.9620194,0.9016574,1.0336993,1.0525624,1.0789708,1.0336993,0.633801,0.452715,0.5885295,0.814887,1.0978339,1.599593,4.395108,4.738417,4.2102494,3.5424948,2.6068838,1.6825907,2.093807,3.2821836,4.0480266,2.5616124,2.2409391,1.9881734,1.7769064,1.7618159,2.282438,1.4675511,1.1657411,1.1544232,1.1506506,0.8186596,0.6752999,0.77338815,0.784706,0.62625575,0.4979865,0.5319401,0.69039035,0.6828451,0.5093044,0.44894236,0.3055826,0.19994913,0.14713238,0.17731337,0.32067314,0.16976812,0.08299775,0.033953626,0.0150905,0.02263575,0.030181,0.0150905,0.003772625,0.02263575,0.06413463,0.21881226,0.5281675,0.58098423,0.33576363,0.10186087,0.060362,0.18485862,0.26408374,0.20749438,0.041498873,0.033953626,0.030181,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.011317875,0.02263575,0.02263575,0.0150905,0.0150905,0.026408374,0.02263575,0.018863125,0.018863125,0.0150905,0.0150905,0.0150905,0.026408374,0.060362,0.116951376,0.20749438,0.271629,0.30181,0.33953625,0.4640329,0.5998474,0.5017591,0.422534,0.4074435,0.32821837,0.32821837,0.27917424,0.23390275,0.21881226,0.24899325,0.2867195,0.3169005,0.3169005,0.30935526,0.35085413,0.422534,0.4640329,0.5470306,0.633801,0.58098423,0.60362,0.62248313,0.63002837,0.6526641,0.7432071,0.86770374,0.79602385,0.59607476,0.35462674,0.19240387,0.150905,0.14335975,0.13204187,0.10940613,0.10186087,0.12826926,0.19240387,0.2678564,0.35085413,0.47157812,0.52062225,0.49421388,0.5357128,0.6488915,0.7092535,0.5017591,0.482896,0.5696664,0.6790725,0.754525,0.633801,0.63002837,0.77338815,0.965792,0.97710985,0.8563859,0.91297525,0.8337501,0.5885295,0.422534,0.331991,0.2678564,0.241448,0.241448,0.211267,0.21503963,0.211267,0.20749438,0.21503963,0.27917424,0.3772625,0.38858038,0.33576363,0.271629,0.271629,0.3734899,0.422534,0.44139713,0.4678055,0.5357128,0.62248313,0.663982,0.58475685,0.44516975,0.4376245,0.47535074,0.46026024,0.52062225,0.6375736,0.6451189,0.5885295,0.5885295,0.59230214,0.58475685,0.6111652,0.56589377,0.58098423,0.6790725,0.784706,0.7167987,0.95824677,0.6828451,0.35085413,0.19994913,0.22258487,0.24522063,0.3169005,0.35839936,0.33576363,0.29426476,0.30181,0.2678564,0.26031113,0.28294688,0.28294688,0.32444575,0.392353,0.46026024,0.4979865,0.4678055,0.4678055,0.44894236,0.42630664,0.422534,0.44894236,0.47912338,0.5017591,0.5357128,0.58475685,0.6149379,0.6451189,0.7054809,0.7884786,0.84884065,0.8262049,0.8337501,0.87902164,0.8865669,0.8563859,0.83752275,0.8865669,0.87147635,0.88279426,0.94315624,0.98465514,1.0336993,1.0940613,1.2411937,1.4298248,1.4901869,1.6524098,1.7014539,1.7391801,1.7542707,1.6146835,1.4260522,1.2487389,1.1393328,1.1053791,1.1204696,1.0676528,1.0487897,1.0336993,0.9997456,0.94315624,1.1129243,1.2487389,1.3543724,1.4524606,1.5769572,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.1358145,0.1659955,0.18485862,0.18485862,0.1358145,0.120724,0.071679875,0.0,0.0,0.049044125,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.1056335,0.30181,0.452715,0.41498876,0.35462674,0.73188925,3.0746894,3.7914882,2.4220252,0.19994913,0.030181,0.041498873,0.15467763,0.5281675,0.9318384,0.7469798,0.38103512,0.3169005,0.6451189,1.2826926,1.9542197,1.8787673,1.8070874,1.629774,1.267602,0.65643674,0.39989826,0.33576363,0.29803738,0.3772625,0.91674787,1.20724,1.5580941,2.11267,2.6597006,2.6106565,2.987919,4.172523,4.2517486,3.7386713,5.5683947,7.496206,8.959985,8.582722,6.270103,3.2029586,5.304311,8.152642,8.7600355,6.643593,3.8593953,6.1795597,7.1076255,6.571913,5.0138187,3.4029078,2.8898308,2.9464202,2.4559789,1.5505489,1.5882751,1.4901869,1.2638294,1.3807807,1.750498,1.7391801,1.4826416,1.2826926,1.026154,0.663982,0.21503963,0.4074435,0.80734175,1.056335,1.1242423,1.2826926,1.1242423,0.7922512,0.8563859,1.3732355,1.8599042,1.9579924,1.1129243,0.32067314,0.06413463,0.32067314,0.55080324,0.6828451,1.0186088,1.5618668,2.0145817,1.5618668,1.358145,1.448688,1.7391801,1.9844007,2.8634224,3.4934506,3.9574835,4.191386,3.983892,3.7386713,3.4029078,3.2670932,3.2972744,3.127506,3.1765501,2.7502437,2.354118,2.3692086,3.0520537,5.1760416,6.749226,6.983129,7.1604424,10.650121,13.422999,13.20796,12.00072,11.506506,13.151371,13.898351,14.762281,14.396337,14.237886,18.5085,40.310497,77.38031,82.80534,50.292866,14.173752,11.099063,8.488406,7.33021,7.707473,8.805306,8.216777,8.986393,12.174261,16.263786,17.180534,12.981603,13.407909,19.583696,27.740112,29.20389,27.713703,23.937305,21.790682,22.541435,24.808783,24.699375,25.212452,25.272816,24.574879,23.575134,21.707684,23.38273,25.597261,26.808273,26.93277,24.17121,23.243143,22.46221,20.749437,17.625704,21.651094,25.944342,27.09122,25.325632,24.522062,24.94837,24.823872,26.521553,29.87919,32.21067,41.683735,41.81955,34.63647,28.279596,37.02077,45.478996,46.92391,43.67568,38.352505,33.85931,26.1707,20.549488,17.836971,16.237377,11.306557,10.868933,6.8774953,5.692891,7.3000293,5.311856,3.893349,2.6785638,3.1237335,4.8327327,5.5382137,11.608367,21.251196,22.899834,16.4411,13.245687,13.536179,12.457208,9.9257765,6.7944975,4.8666863,5.832478,5.221313,4.3724723,4.640329,7.3868,17.761518,35.406086,50.206093,52.077316,30.961933,38.66186,42.766476,39.457886,31.052477,25.985842,21.726547,22.01704,24.903097,28.483318,30.897799,28.626678,27.072357,26.412148,26.849771,28.596497,34.538383,36.74914,35.52681,34.044167,38.31478,37.42444,33.383957,29.256706,29.083166,37.873383,33.18401,28.44182,25.92925,24.442837,19.31584,14.068119,10.733118,10.714255,13.377728,16.03743,17.844517,21.553007,23.661903,23.767538,24.597515,27.027086,28.404093,28.660633,28.358822,28.68704,24.695602,23.624178,23.537407,23.375185,22.948877,18.45568,18.184053,20.73812,21.03993,10.344538,10.442626,10.355856,11.02361,10.469034,3.8292143,9.5183325,6.609639,3.0445085,2.3428001,3.6028569,7.5075235,9.857869,11.638548,14.750964,22.00195,15.192361,13.407909,14.811326,17.082445,17.425755,4.7912335,7.9036493,10.54826,7.432071,4.195159,2.6219745,4.991183,7.4282985,7.7602897,5.5382137,3.108643,3.1425967,4.425289,7.2660756,13.502225,16.542961,15.645076,14.558559,13.422999,8.7751255,6.330465,6.307829,5.9003854,5.3571277,7.9941926,11.41219,11.461235,10.038955,8.179051,6.043745,4.0517993,4.9119577,7.213259,9.042982,7.9791017,6.9189944,7.643338,8.654402,9.22784,9.397609,7.2283497,8.047009,8.650629,7.665974,5.553304,6.8246784,7.232122,6.3116016,4.478106,3.0520537,3.429316,4.074435,3.9348478,2.9313297,1.9542197,1.9051756,2.7087448,4.0970707,5.0515447,3.7688525,4.659192,4.508287,4.9421387,6.0550632,6.40969,5.323174,5.1345425,4.8402777,4.459243,5.0213637,5.119452,4.647874,4.2630663,4.0216184,3.3878171,3.6066296,4.255521,3.9348478,2.674791,1.9542197,3.4670424,3.1124156,1.6976813,0.33953625,0.47157812,0.5357128,0.3470815,1.086516,2.3805263,2.3201644,1.9881734,2.071171,2.0183544,1.7467253,1.6486372,2.0145817,1.7014539,1.3241913,1.0751982,0.73188925,0.513077,0.91674787,1.1883769,1.2336484,1.5882751,3.651901,3.9273026,3.1765501,2.142851,1.5580941,1.4222796,1.4600059,2.3956168,3.5274043,2.746471,1.8184053,1.750498,1.81086,1.8297231,2.1956677,1.4411428,1.20724,1.1695137,1.1091517,0.91674787,0.73188925,0.7507524,0.7922512,0.754525,0.59607476,0.5696664,0.76584285,0.68661773,0.33953625,0.23013012,0.15467763,0.10940613,0.090543,0.150905,0.38103512,0.22258487,0.10186087,0.026408374,0.00754525,0.0452715,0.0452715,0.018863125,0.0,0.003772625,0.0150905,0.05281675,0.35462674,0.7997965,1.0299267,0.44139713,0.08677038,0.1358145,0.26408374,0.2867195,0.150905,0.06790725,0.026408374,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.026408374,0.02263575,0.026408374,0.041498873,0.0150905,0.0150905,0.0150905,0.026408374,0.056589376,0.090543,0.1659955,0.23767537,0.2678564,0.29426476,0.42630664,0.4640329,0.41876137,0.35085413,0.29049212,0.23013012,0.27917424,0.27917424,0.2678564,0.26031113,0.26031113,0.30935526,0.38480774,0.392353,0.32821837,0.29049212,0.35085413,0.3734899,0.52062225,0.7507524,0.8224323,0.6413463,0.59607476,0.59607476,0.63002837,0.77716076,0.8639311,0.8111144,0.7130261,0.5696664,0.29049212,0.181086,0.16976812,0.15845025,0.124496624,0.1358145,0.1358145,0.1659955,0.23767537,0.32444575,0.33576363,0.44516975,0.5017591,0.5055317,0.51684964,0.62625575,0.5017591,0.4640329,0.52439487,0.59607476,0.47157812,0.5583485,0.6073926,0.68661773,0.80734175,0.91674787,0.9016574,0.91674787,0.94315624,0.83752275,0.33576363,0.2867195,0.23767537,0.20749438,0.19994913,0.19994913,0.17354076,0.150905,0.16222288,0.21881226,0.3055826,0.29426476,0.271629,0.23390275,0.211267,0.26031113,0.331991,0.38858038,0.41876137,0.4376245,0.48666862,0.52439487,0.55080324,0.55080324,0.55080324,0.6111652,0.5998474,0.5394854,0.5696664,0.66775465,0.65643674,0.58475685,0.52062225,0.47535074,0.47535074,0.55080324,0.573439,0.5998474,0.6526641,0.7054809,0.65643674,0.5357128,0.40367088,0.34330887,0.392353,0.56589377,0.47912338,0.5394854,0.6375736,0.6111652,0.24522063,0.23013012,0.19994913,0.18485862,0.211267,0.32067314,0.41876137,0.47912338,0.5017591,0.47912338,0.38103512,0.392353,0.47157812,0.482896,0.41121614,0.35085413,0.39989826,0.44894236,0.48666862,0.5055317,0.52062225,0.56589377,0.663982,0.77338815,0.875249,0.9620194,0.9507015,1.0110635,1.0336993,0.9808825,0.8865669,0.94692886,0.9620194,0.97333723,0.9997456,1.0223814,1.1581959,1.327964,1.4600059,1.539231,1.5882751,1.6222287,1.7165444,1.8070874,1.8448136,1.7844516,1.6750455,1.50905,1.297783,1.1204696,1.1431054,1.1204696,1.1242423,1.1242423,1.1129243,1.1129243,1.1393328,1.1355602,1.1544232,1.2110126,1.297783,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.026408374,0.056589376,0.08677038,0.03772625,0.06413463,0.08677038,0.07922512,0.03772625,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.23767537,0.5885295,0.845068,0.8601585,0.58475685,0.995973,1.2638294,0.9695646,0.34330887,0.24899325,0.94692886,1.2525115,1.2562841,1.0487897,0.7092535,0.3734899,0.4640329,0.9922004,1.6863633,1.9768555,1.7882242,1.5467763,1.1544232,0.6828451,0.3772625,0.34330887,0.3734899,0.3169005,0.33953625,0.91674787,1.0902886,1.4600059,2.1202152,2.6031113,1.8900851,2.3654358,4.1310244,4.82896,4.7120085,6.6322746,7.183078,8.058327,8.182823,7.24344,5.692891,9.786189,11.332966,10.005001,7.01331,5.13077,4.617693,4.0593443,3.1539145,2.2409391,2.3277097,2.8596497,2.9124665,2.9992368,3.4142256,4.221567,4.4101987,2.9803739,2.425798,3.1425967,3.4255435,2.9803739,2.5729303,2.2447119,1.8146327,0.8865669,0.3961256,0.32067314,0.33953625,0.35839936,0.52439487,0.6413463,0.55080324,0.68661773,1.1280149,1.6184561,1.5505489,0.875249,0.32067314,0.15845025,0.211267,0.32444575,0.56589377,1.0638802,1.690136,2.0636258,2.1956677,2.233394,2.1994405,2.2484846,2.6672459,2.9124665,3.1048703,3.350091,3.5047686,3.2029586,3.1727777,3.1614597,3.1576872,3.097325,2.848332,3.0218725,2.757789,2.4861598,2.6295197,3.6254926,7.232122,9.465516,9.405154,8.118689,8.661947,8.09228,9.050528,9.820143,9.854096,9.782416,9.016574,8.416726,8.446907,9.665465,12.736382,27.985332,49.34971,51.077568,31.83341,14.724555,12.166716,9.363655,7.8395147,7.6018395,7.1566696,6.3153744,8.873214,14.351066,20.549488,23.563816,18.085964,13.70972,15.845025,22.990377,26.740366,29.037895,25.484081,22.401848,22.737612,26.04243,28.26828,31.399557,33.47073,33.75745,32.765247,29.268024,27.611843,25.872662,24.499426,26.310287,26.529099,26.212198,24.752193,23.967487,28.109829,35.466446,39.963417,40.782078,38.94858,37.31126,36.364334,35.77203,38.9184,44.335888,45.697807,45.037598,36.89627,28.898308,26.547962,33.1991,33.278324,32.27858,32.15031,32.516254,30.648806,26.385738,21.839725,16.573141,11.140562,7.1076255,5.0666356,4.504514,6.6662283,10.33322,11.827179,7.092535,9.205205,11.140562,10.065364,7.3453007,7.2396674,10.846297,12.928786,11.317875,6.8963585,10.284176,10.080454,7.3151197,4.5950575,6.1229706,7.4509344,6.952948,5.2854476,3.9763467,5.4438977,12.344029,24.476791,40.517994,51.749096,42.068542,49.681698,53.427914,46.55042,32.138992,23.118647,25.212452,28.939806,35.160866,41.812004,43.898266,37.98656,34.828873,33.16892,32.5653,33.40282,36.654823,40.385952,41.67619,40.21241,38.31478,40.83112,37.43953,32.101265,29.856554,36.798183,32.961426,30.36963,32.097492,35.28159,31.120384,21.869907,15.120681,11.98563,12.151625,13.913441,14.7321005,17.844517,20.972023,23.216734,25.061548,26.29897,27.19308,27.242125,26.585688,26.02734,23.850534,24.442837,23.661903,21.005976,19.591242,17.882242,17.210714,17.852062,17.244669,9.978593,10.438853,9.337247,7.677292,7.8017883,13.373956,11.310329,8.601585,6.3832817,4.7874613,2.9313297,4.659192,6.1795597,9.548513,14.226569,17.082445,12.321393,10.917976,12.898605,17.56157,23.480818,9.476834,6.089017,6.0512905,5.2779026,2.8521044,1.7467253,2.9916916,4.9723196,6.2851934,5.73439,4.0291634,4.3007927,6.089017,9.020347,12.808062,13.162688,14.347293,14.996184,13.773854,9.397609,9.8239155,8.990166,7.4471617,6.598321,8.66572,10.785934,10.823661,9.020347,6.432326,4.930821,3.519859,4.564876,6.228604,7.541477,8.382772,7.9451485,6.356873,6.009792,7.3679366,8.98262,7.515069,8.028146,8.8769865,8.514814,5.492942,5.5797124,8.60913,10.178542,8.684583,5.3344917,4.353609,5.070408,5.6513925,5.0477724,2.9766011,2.293756,2.8219235,3.904667,4.5196047,3.2670932,2.927557,2.6521554,2.727608,3.0671442,3.187868,2.8219235,3.150142,3.5123138,3.85185,4.727099,5.5759397,4.4894238,3.6179473,3.5424948,3.289729,2.3163917,2.584248,3.1425967,3.0218725,1.20724,1.3656902,1.358145,0.9393836,0.32821837,0.23013012,0.56212115,0.38103512,0.44894236,0.8601585,1.0148361,1.1996948,1.4071891,1.3656902,1.1883769,1.3543724,1.2336484,1.1883769,1.1657411,1.0638802,0.73188925,0.66775465,0.9280658,1.0601076,1.1581959,1.8448136,2.4710693,3.451952,3.5651307,2.8445592,2.5691576,1.7429527,0.9507015,1.0525624,1.8297231,1.9655377,1.3996439,1.4298248,1.3355093,1.0902886,1.3656902,1.177059,1.0525624,1.056335,1.1242423,1.0751982,0.7167987,0.573439,0.5583485,0.55457586,0.422534,0.362172,0.33953625,0.32067314,0.2565385,0.120724,0.06413463,0.0754525,0.071679875,0.0754525,0.19994913,0.17731337,0.124496624,0.056589376,0.0,0.00754525,0.18485862,0.17354076,0.08677038,0.011317875,0.003772625,0.030181,0.116951376,0.3169005,0.7092535,1.3958713,0.59230214,0.19994913,0.13958712,0.28294688,0.422534,0.33576363,0.1659955,0.0452715,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.018863125,0.00754525,0.003772625,0.011317875,0.0150905,0.033953626,0.033953626,0.030181,0.049044125,0.1056335,0.15845025,0.23390275,0.27917424,0.29426476,0.34330887,0.36971724,0.38480774,0.38858038,0.3470815,0.23013012,0.23767537,0.28294688,0.29426476,0.27540162,0.28294688,0.35085413,0.38858038,0.3772625,0.31312788,0.23013012,0.271629,0.28294688,0.3772625,0.56212115,0.7507524,0.65643674,0.62625575,0.5998474,0.5772116,0.6073926,0.7130261,0.694163,0.62248313,0.5357128,0.44894236,0.24899325,0.1961765,0.16976812,0.12826926,0.11317875,0.14335975,0.16222288,0.1961765,0.23767537,0.24899325,0.5357128,0.6488915,0.58098423,0.45648763,0.5281675,0.543258,0.5583485,0.5696664,0.56212115,0.4979865,0.52439487,0.543258,0.6413463,0.8186596,0.98842776,0.8111144,0.6828451,0.6526641,0.63002837,0.3734899,0.29426476,0.23767537,0.1961765,0.18485862,0.22258487,0.21881226,0.18485862,0.1659955,0.18863125,0.24522063,0.241448,0.331991,0.39989826,0.40367088,0.392353,0.52439487,0.513077,0.452715,0.392353,0.35462674,0.41121614,0.48666862,0.5357128,0.55080324,0.573439,0.5319401,0.5093044,0.482896,0.452715,0.46026024,0.55457586,0.573439,0.51684964,0.4376245,0.4640329,0.46026024,0.482896,0.49421388,0.482896,0.47157812,0.4979865,0.38103512,0.27540162,0.2678564,0.36971724,0.47912338,0.5319401,0.48666862,0.36594462,0.24522063,0.23013012,0.23013012,0.2678564,0.33576363,0.4074435,0.43385187,0.4074435,0.44894236,0.5281675,0.43007925,0.38480774,0.36594462,0.36594462,0.3734899,0.35085413,0.35085413,0.40367088,0.44516975,0.47535074,0.55457586,0.573439,0.6187105,0.66020936,0.72811663,0.9016574,0.98465514,1.0110635,0.97333723,0.9205205,0.95824677,0.9016574,0.90920264,0.9620194,1.0336993,1.0940613,1.1129243,1.1506506,1.2110126,1.2751472,1.2940104,1.448688,1.6184561,1.7354075,1.7278622,1.5279131,1.5165952,1.6675003,1.6109109,1.297783,1.0110635,1.1996948,1.2562841,1.1883769,1.0789708,1.0902886,1.2411937,1.2826926,1.1808317,1.0374719,1.1016065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.056589376,0.06790725,0.049044125,0.030181,0.026408374,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.23390275,0.7469798,1.1393328,1.3128735,1.4298248,1.3694628,1.4071891,1.116697,0.66020936,0.7997965,1.3656902,1.5505489,1.3430545,0.9318384,0.72811663,0.41498876,0.6488915,1.3128735,1.9655377,1.8749946,1.5015048,1.1016065,0.694163,0.40367088,0.452715,0.8337501,0.7092535,0.5583485,0.63002837,0.91674787,1.0978339,1.7919968,3.108643,3.9197574,1.8448136,1.7844516,3.6443558,4.919503,5.138315,5.8702044,5.4288073,7.6320205,8.926031,8.52236,8.412953,11.16697,10.510533,8.062099,5.353355,3.8178966,2.6332922,2.384299,2.5276587,2.7841973,3.150142,3.3878171,3.1124156,3.0407357,3.470815,4.29702,4.4215164,3.7348988,3.3915899,3.5349495,3.2859564,2.5201135,1.9957186,1.6939086,1.4411428,0.8865669,0.3734899,0.181086,0.12826926,0.1358145,0.23390275,0.30181,0.23390275,0.33953625,0.6526641,0.94315624,0.995973,0.87902164,0.72811663,0.55080324,0.26408374,0.513077,0.7507524,1.0450171,1.3770081,1.6260014,2.323937,2.5880208,2.4899325,2.3465726,2.6898816,2.5729303,2.463524,2.305074,2.233394,2.584248,2.8445592,2.7841973,2.565385,2.4484336,2.7879698,2.7087448,2.2447119,2.4069347,3.2105038,3.6669915,5.934339,7.8734684,8.507269,8.190369,8.612903,7.9036493,8.065872,8.156415,7.7602897,6.983129,5.987156,6.1908774,8.790216,13.426772,18.16519,20.734346,23.816582,22.782883,17.550251,12.555296,9.307066,7.496206,6.8774953,6.8737226,6.579458,5.413717,5.926794,8.348819,11.623458,13.396591,11.314102,8.805306,9.635284,13.890805,17.984104,22.273579,24.431519,26.238607,28.306005,30.07914,33.236828,38.31478,42.204357,44.76597,48.813995,52.152767,46.275017,36.24738,27.857063,27.600525,30.592216,29.486837,28.483318,33.821583,53.782543,79.76084,88.20775,85.09156,74.19621,57.091133,49.71188,48.83286,53.714634,59.29812,56.204567,39.986053,28.490864,21.824636,20.515535,25.521809,24.495655,23.29596,23.895807,26.076384,27.438301,25.080412,21.34174,16.58446,10.963248,4.402653,3.2331395,3.9084394,6.8699503,11.1631975,14.437836,8.379,6.417235,6.3945994,6.7454534,6.488915,6.8774953,12.468526,16.252468,14.603831,7.2887115,7.8017883,7.7640624,7.3453007,7.6395655,10.631257,11.936585,10.816116,7.7678347,4.7950063,5.379763,10.906659,20.889025,33.85931,44.53961,43.87563,49.462887,61.00712,60.373318,45.39977,29.898052,34.485565,42.01195,51.534058,59.011402,57.328808,50.87762,48.670635,46.508923,43.528545,42.177948,44.00767,51.171886,58.39269,58.917084,44.53961,42.09495,39.642742,35.221226,31.407103,35.349495,36.270016,33.840446,34.61006,38.57132,39.171165,28.90208,22.126446,19.047983,19.225298,21.549234,21.134245,22.00195,24.34475,26.740366,26.174473,24.793692,24.642786,25.012505,25.51049,26.046204,24.729557,27.423212,26.729048,22.01704,19.447882,17.972786,16.610868,16.01102,14.807553,9.612649,18.678267,24.069347,19.391293,9.597558,10.948157,12.683565,13.588995,10.895341,6.009792,4.4931965,4.7308717,5.0779533,8.635539,16.867407,29.603788,21.005976,13.472044,14.464244,25.672712,43.01924,16.486372,6.175787,4.0216184,4.8327327,6.270103,2.5427492,2.505023,4.3309736,6.224831,6.4436436,5.7570257,5.511805,6.6360474,8.624221,9.522105,11.45369,15.833707,17.323895,15.150862,13.151371,13.309821,11.087745,8.714764,7.3415284,7.020855,8.529905,8.473316,7.2472124,5.594803,4.617693,3.4632697,3.7235808,4.5460134,5.462761,6.368191,7.1868505,5.9532022,5.523123,6.7379084,8.424272,7.6207023,8.122461,8.790216,8.409182,5.6891184,5.7079816,8.103599,10.167224,10.378491,8.412953,7.696155,8.035691,8.009283,6.862405,4.4894238,2.7691069,2.5880208,3.410453,4.025391,2.5767028,1.81086,1.780679,2.191895,2.5238862,2.04099,1.8599042,2.123988,2.233394,2.173032,2.5012503,2.8596497,2.2447119,1.8184053,1.9881734,2.3880715,1.4750963,1.237421,1.4675511,1.5920477,0.6828451,0.47157812,0.49044126,0.58475685,0.5772116,0.27917424,0.56212115,0.38858038,0.211267,0.2263575,0.3772625,0.5696664,0.7054809,0.6488915,0.513077,0.6790725,0.5281675,0.6073926,0.7432071,0.7922512,0.63002837,0.6073926,0.7922512,0.8601585,0.90920264,1.4600059,1.6976813,2.3314822,2.9086938,3.240685,3.380272,2.0145817,0.83752275,0.47157812,0.8111144,1.0450171,1.1581959,1.1808317,1.0110635,0.83752275,1.1695137,1.3317367,1.0978339,0.87902164,0.83752275,0.875249,0.7130261,0.5319401,0.5017591,0.56212115,0.41876137,0.27917424,0.211267,0.18863125,0.17731337,0.120724,0.056589376,0.05281675,0.0754525,0.094315626,0.08677038,0.094315626,0.06790725,0.033953626,0.00754525,0.00754525,0.09808825,0.124496624,0.08299775,0.0150905,0.00754525,0.026408374,0.030181,0.116951376,0.44139713,1.2298758,0.84129536,0.36594462,0.13204187,0.18863125,0.27917424,0.24899325,0.15467763,0.06790725,0.02263575,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.00754525,0.0150905,0.011317875,0.003772625,0.0,0.00754525,0.030181,0.033953626,0.030181,0.0452715,0.1056335,0.13204187,0.1659955,0.21881226,0.27917424,0.31312788,0.26408374,0.27917424,0.29049212,0.271629,0.23767537,0.23013012,0.23390275,0.24899325,0.29049212,0.39989826,0.4074435,0.38103512,0.3734899,0.36594462,0.2678564,0.23767537,0.23767537,0.31312788,0.4640329,0.6413463,0.6413463,0.6752999,0.66775465,0.6187105,0.6111652,0.7054809,0.7054809,0.59607476,0.452715,0.422534,0.34330887,0.26408374,0.23767537,0.2565385,0.25276586,0.25276586,0.23013012,0.23390275,0.2678564,0.26408374,0.41876137,0.5319401,0.52439487,0.44516975,0.44894236,0.543258,0.9280658,0.95824677,0.6149379,0.52062225,0.59230214,0.7507524,0.86770374,0.91674787,0.9997456,0.8224323,0.76584285,0.7507524,0.6790725,0.44516975,0.27917424,0.19994913,0.16976812,0.1659955,0.19240387,0.20749438,0.17354076,0.15467763,0.17354076,0.23767537,0.2678564,0.3055826,0.35085413,0.38103512,0.362172,0.43007925,0.4376245,0.41498876,0.3772625,0.33953625,0.4074435,0.44139713,0.43385187,0.4074435,0.41876137,0.45648763,0.49044126,0.482896,0.452715,0.45648763,0.49044126,0.5394854,0.55457586,0.5357128,0.52439487,0.49044126,0.48666862,0.49044126,0.47535074,0.4074435,0.41121614,0.34330887,0.32821837,0.38858038,0.45648763,0.4979865,0.5093044,0.45648763,0.3734899,0.33576363,0.271629,0.22258487,0.22258487,0.271629,0.3169005,0.40367088,0.40367088,0.4376245,0.5093044,0.5055317,0.4376245,0.43385187,0.47157812,0.5093044,0.46026024,0.38858038,0.35462674,0.35462674,0.39989826,0.52062225,0.60362,0.6149379,0.5998474,0.6111652,0.7205714,0.7997965,0.9393836,1.0110635,0.98842776,0.9318384,0.9620194,0.9695646,1.0223814,1.1204696,1.2223305,1.2638294,1.297783,1.3694628,1.4864142,1.6146835,1.659955,1.5354583,1.4298248,1.4411428,1.5845025,1.6561824,1.6373192,1.5128226,1.3091009,1.0940613,1.1506506,1.1657411,1.1581959,1.1280149,1.0751982,1.0676528,1.1129243,1.1619685,1.1921495,1.20724,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.056589376,0.049044125,0.018863125,0.0,0.00754525,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.011317875,0.23767537,0.7432071,1.1695137,1.4826416,1.9730829,2.0560806,2.052308,1.6486372,1.1016065,1.2449663,1.9768555,2.033445,1.4750963,0.76207024,0.7582976,0.5281675,0.8299775,1.4222796,1.8523588,1.4600059,1.0412445,0.694163,0.452715,0.3961256,0.62248313,0.9620194,0.814887,0.79602385,1.0299267,1.1581959,1.3732355,2.3692086,3.640583,4.044254,1.8146327,2.3616633,4.014073,5.111907,5.413717,6.1229706,6.1418333,8.620448,9.473062,8.311093,8.469543,9.431562,7.745199,5.4174895,3.5349495,2.2447119,1.1921495,1.267602,1.8674494,2.4522061,2.5767028,2.6672459,2.5691576,2.5729303,2.837014,3.361409,3.4444065,3.519859,3.4330888,3.1539145,2.7540162,1.8636768,1.2525115,0.95447415,0.87902164,0.8224323,0.43007925,0.25276586,0.1659955,0.10940613,0.10186087,0.094315626,0.060362,0.10186087,0.2263575,0.32067314,0.41498876,0.55457586,0.5998474,0.47912338,0.19240387,0.4678055,0.6526641,0.7582976,0.8639311,1.1242423,1.9164935,2.0560806,1.7882242,1.4977322,1.7089992,1.5845025,1.4864142,1.267602,1.1393328,1.6637276,1.901403,1.8146327,1.8674494,2.2220762,2.7426984,2.4861598,2.8822856,3.5123138,3.8971217,3.519859,4.5120597,5.832478,6.9189944,7.665974,8.446907,8.160188,7.9451485,7.6018395,7.0887623,6.5568223,6.94163,8.428044,11.978085,17.093763,21.82841,17.448391,11.415963,8.7600355,9.529651,8.793989,6.983129,7.394345,7.586749,6.851087,6.2436943,4.561104,3.429316,3.31991,3.9989824,4.5460134,5.2062225,5.4665337,6.2814207,8.09228,10.853842,15.433809,21.38701,27.136492,32.606796,39.23153,45.407314,49.82883,57.023228,69.20126,86.238434,94.070404,81.30007,59.320755,39.703106,34.168663,38.424187,36.628418,38.065784,55.219913,103.76982,133.32457,125.35301,110.34551,99.3219,83.80132,67.48849,64.52698,67.06218,66.73396,54.71061,34.07435,23.424229,19.021576,18.255732,19.644058,18.62545,17.825653,18.51227,20.541943,22.352802,22.684793,20.66644,17.784155,13.200415,3.7537618,4.217795,6.2663302,8.888305,11.45369,13.717264,9.058073,4.508287,2.5238862,3.4745877,5.6476197,7.854605,13.751218,18.504726,19.021576,13.93985,10.133271,7.54525,7.254758,8.929804,10.816116,12.064855,14.120935,12.095036,6.9755836,5.6476197,9.612649,17.508753,27.340214,36.243607,40.52554,43.83413,64.32703,76.68237,70.34059,49.50816,46.814503,57.219402,74.64516,88.751,84.95197,69.9671,63.968628,60.41859,56.513924,53.212875,52.522484,58.400234,68.71836,74.034,57.6193,44.505657,40.106777,36.839684,33.202873,33.749905,38.22801,35.817303,33.62541,34.727013,38.178967,29.120892,25.216225,24.76351,25.921707,26.706413,25.26527,24.631468,25.529354,26.857317,25.687803,23.665676,22.790428,22.843245,23.676994,25.212452,26.05375,31.309015,31.671186,26.09902,21.824636,19.04421,17.23335,16.90136,17.172989,15.799753,20.98334,24.925734,21.715229,13.864397,12.283667,14.803781,14.369928,10.79348,6.326692,5.66271,5.6853456,5.149633,6.8699503,13.264549,26.381968,19.263023,12.7477,12.879742,22.326395,40.389725,17.852062,7.7301087,5.3684454,7.01331,9.786189,3.4179983,2.022127,3.5424948,5.745708,6.217286,5.73439,5.4703064,6.3719635,7.907422,8.062099,12.287439,15.724301,16.15438,14.437836,14.543469,13.788944,11.050018,8.646856,7.3453007,6.33801,7.8961043,7.111398,5.907931,5.062863,4.2102494,3.2821836,2.848332,2.9992368,3.5349495,3.9688015,5.5193505,4.983638,4.678055,5.5306683,7.073672,6.549277,7.383027,8.088508,7.696155,5.7419353,5.6589375,6.8737226,8.235641,8.975075,8.669493,8.66572,9.035437,8.707218,7.3717093,5.4665337,4.014073,3.138824,3.2142766,3.5274043,2.2748928,1.3505998,1.2751472,1.7316349,2.123988,1.5580941,1.4637785,1.5203679,1.3015556,0.8639311,0.7432071,0.7092535,0.55457586,0.4979865,0.7130261,1.3317367,0.8941121,0.482896,0.34330887,0.43385187,0.4074435,0.24522063,0.17354076,0.4074435,0.73566186,0.5470306,0.60362,0.39989826,0.18485862,0.14713238,0.44139713,0.46026024,0.38480774,0.24899325,0.14335975,0.20749438,0.21503963,0.30181,0.3961256,0.46026024,0.47912338,0.5394854,0.6413463,0.6413463,0.65643674,1.0751982,1.7240896,1.7844516,2.3918443,3.5689032,4.247976,3.0897799,1.4562333,0.5357128,0.5017591,0.52062225,0.7205714,0.7696155,0.7130261,0.7507524,1.2487389,1.478869,1.2223305,0.87147635,0.70170826,0.88279426,0.754525,0.6413463,0.6375736,0.663982,0.47912338,0.3772625,0.2867195,0.20749438,0.150905,0.150905,0.071679875,0.05281675,0.0754525,0.09808825,0.041498873,0.030181,0.0150905,0.011317875,0.0150905,0.00754525,0.00754525,0.06413463,0.090543,0.0754525,0.071679875,0.09808825,0.056589376,0.05281675,0.20372175,0.65643674,0.70170826,0.482896,0.29803738,0.2263575,0.10186087,0.09808825,0.08299775,0.06413463,0.03772625,0.02263575,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.0,0.00754525,0.011317875,0.00754525,0.0,0.0,0.018863125,0.026408374,0.026408374,0.03772625,0.08677038,0.120724,0.14713238,0.18863125,0.23767537,0.24899325,0.18863125,0.20749438,0.22258487,0.20749438,0.19994913,0.20749438,0.20749438,0.23390275,0.3169005,0.4678055,0.41498876,0.3470815,0.3470815,0.38858038,0.32444575,0.24522063,0.241448,0.29426476,0.392353,0.543258,0.573439,0.6111652,0.66775465,0.7092535,0.67152727,0.633801,0.6413463,0.5583485,0.41498876,0.38103512,0.40367088,0.31312788,0.271629,0.3169005,0.36971724,0.34330887,0.32444575,0.31312788,0.3055826,0.27917424,0.331991,0.46026024,0.5281675,0.49421388,0.41121614,0.49044126,0.9280658,1.0789708,0.88279426,0.8563859,0.724344,0.80734175,0.90543,0.935611,0.9507015,0.86770374,0.84129536,0.784706,0.66775465,0.513077,0.32067314,0.21881226,0.17731337,0.16976812,0.1659955,0.17354076,0.15467763,0.14713238,0.1659955,0.21503963,0.2678564,0.27917424,0.32067314,0.3961256,0.4376245,0.41876137,0.4074435,0.41121614,0.422534,0.39989826,0.41498876,0.3961256,0.36971724,0.35462674,0.3734899,0.40367088,0.4376245,0.45648763,0.452715,0.43385187,0.4376245,0.5055317,0.5583485,0.55457586,0.5017591,0.46026024,0.45648763,0.49044126,0.51684964,0.44516975,0.39989826,0.392353,0.42630664,0.47535074,0.482896,0.47157812,0.47535074,0.45648763,0.41121614,0.40367088,0.30181,0.21881226,0.20372175,0.23767537,0.24522063,0.32821837,0.39989826,0.46026024,0.52439487,0.58098423,0.5470306,0.5281675,0.52062225,0.4979865,0.45648763,0.41498876,0.362172,0.3470815,0.38858038,0.45648763,0.56589377,0.5998474,0.5885295,0.58475685,0.633801,0.67152727,0.8337501,0.95824677,0.98465514,0.97333723,1.0450171,1.0035182,0.9997456,1.0751982,1.1695137,1.1921495,1.2223305,1.2940104,1.418507,1.5731846,1.5656394,1.3317367,1.1393328,1.1393328,1.3694628,1.4298248,1.3694628,1.2902378,1.2185578,1.0940613,1.0601076,1.116697,1.1619685,1.1393328,1.0072908,0.91674787,0.9507015,1.0789708,1.2223305,1.2449663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.02263575,0.21881226,0.59230214,0.9620194,1.2940104,1.7014539,1.9504471,1.9730829,1.720317,1.3770081,1.3543724,2.595566,2.5917933,1.6939086,0.6828451,0.784706,0.663982,0.95447415,1.3128735,1.4034165,0.87147635,0.58098423,0.47535074,0.48666862,0.56212115,0.66775465,0.7092535,0.76584285,1.0072908,1.3656902,1.5354583,1.7391801,2.7426984,3.2633207,2.8785129,2.0070364,4.5460134,5.9984736,6.417235,6.651138,8.333729,9.329701,10.570895,9.763554,7.3113475,6.3153744,5.9418845,4.5912848,3.2520027,2.263575,1.3392819,0.6488915,0.6073926,0.7130261,0.72811663,0.65643674,0.995973,1.3468271,1.6637276,1.9278114,2.142851,2.2220762,2.3428001,2.2711203,2.052308,2.052308,1.4222796,0.87902164,0.5998474,0.6187105,0.80356914,0.5017591,0.35839936,0.2263575,0.07922512,0.0,0.026408374,0.071679875,0.06413463,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.12826926,0.25276586,0.32067314,0.4074435,0.7432071,1.1544232,0.9695646,0.55457586,0.23767537,0.32067314,0.36971724,0.49421388,0.58475685,0.6451189,0.7922512,0.76584285,0.7922512,1.4600059,2.463524,2.6106565,2.8219235,4.4215164,5.1232247,4.4139714,3.5689032,4.0970707,4.9459114,6.0550632,7.122716,7.643338,7.594294,8.246958,8.703445,8.831716,9.261794,11.200924,12.849561,14.449154,16.18456,18.19537,15.396083,11.917723,9.574923,8.167733,5.458988,6.9454026,9.857869,10.110635,7.4773426,5.6061206,3.5160866,2.4974778,2.2409391,2.4823873,3.0105548,4.255521,5.945657,7.5226145,8.91094,10.521852,14.875461,21.371922,29.886736,41.72146,59.63011,69.19749,68.9749,78.91954,105.16192,140.00212,145.51392,123.708145,90.550545,61.535286,51.6661,55.351955,52.812977,56.75537,83.97863,155.34915,164.3959,128.98605,103.46801,104.490395,110.95667,91.64083,84.57848,77.99902,65.05138,43.81904,31.20338,23.186554,20.02132,19.708193,17.99542,15.788436,14.890551,15.558306,16.90136,16.893814,19.640285,19.723284,18.614132,15.098045,5.2590394,6.609639,9.782416,11.604594,11.487643,11.438599,9.42779,6.3229194,4.0593443,3.8065786,5.96452,9.65792,13.4644985,17.38803,20.398582,20.432537,14.166207,8.692128,6.6586833,7.605612,7.964011,8.677037,14.32843,14.7170105,9.231613,6.85486,8.047009,12.615658,20.255224,28.954897,34.964687,37.348988,62.48976,90.04878,102.74367,86.336525,66.77169,71.70251,93.42906,116.16667,116.05727,91.70874,78.77241,72.14768,67.933655,63.4216,59.08308,58.370052,66.647194,77.48595,72.69471,49.938236,40.838665,37.382942,35.08164,33.006695,37.933743,36.613327,31.980541,27.958923,29.44911,22.839472,21.952906,24.110846,26.004704,23.692085,22.254715,21.764273,21.82841,22.337713,23.4695,22.95265,22.054766,21.375692,21.439827,22.692339,26.317833,33.749905,36.021023,31.505192,25.92548,21.375692,19.059301,19.80251,23.375185,28.475773,17.984104,12.189351,13.298503,18.187824,18.399092,17.923742,12.596795,8.405409,7.5603404,8.514814,8.922258,6.8171334,5.7570257,6.9755836,9.363655,7.99042,9.737145,10.020092,10.465261,18.89708,13.20796,8.918486,7.7338815,9.099571,10.208723,4.636556,2.2447119,3.0558262,5.251494,5.160951,4.221567,4.5799665,5.794752,7.3188925,8.492179,13.343775,13.211733,12.00072,11.638548,12.049765,10.929295,9.005256,7.635793,7.4509344,8.326183,9.97482,8.050782,6.017337,4.9723196,3.640583,2.806833,2.2107582,2.1277604,2.4182527,2.516341,3.863168,3.3048196,2.8407867,3.410453,4.8930945,4.587512,5.7570257,6.688864,6.5266414,5.2628117,4.957229,5.8211603,6.156924,5.7192993,5.7381625,6.013564,6.673774,6.8473144,6.3153744,5.523123,5.2628117,4.217795,3.4066803,3.0445085,2.546522,1.4449154,0.935611,0.9695646,1.2298758,1.1581959,1.1695137,1.086516,0.79602385,0.40367088,0.23013012,0.3961256,0.62625575,0.5017591,0.2263575,0.6149379,0.5055317,0.24899325,0.120724,0.1961765,0.35462674,0.70170826,0.3961256,0.3470815,0.69039035,0.7884786,0.62248313,0.3772625,0.1961765,0.2565385,0.76584285,0.7507524,0.47535074,0.23390275,0.1358145,0.09808825,0.2263575,0.271629,0.24522063,0.21503963,0.31312788,0.49044126,0.52062225,0.47157812,0.5017591,0.8563859,1.9504471,1.7769064,2.1843498,3.6292653,5.149633,4.485651,2.516341,1.0827434,0.694163,0.52439487,0.23013012,0.29049212,0.4074435,0.58475685,1.1280149,1.3128735,1.2751472,1.0789708,0.9393836,1.2034674,0.87902164,0.86770374,0.9280658,0.86770374,0.5470306,0.5470306,0.422534,0.271629,0.1659955,0.15467763,0.0754525,0.060362,0.0754525,0.07922512,0.03772625,0.00754525,0.0,0.00754525,0.011317875,0.0,0.0,0.0452715,0.09808825,0.13958712,0.14335975,0.21503963,0.150905,0.06790725,0.05281675,0.16976812,0.331991,0.49044126,0.5093044,0.35462674,0.08299775,0.06413463,0.06413463,0.071679875,0.06413463,0.030181,0.00754525,0.00754525,0.00754525,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.00754525,0.00754525,0.0,0.003772625,0.011317875,0.026408374,0.030181,0.030181,0.060362,0.12826926,0.1961765,0.22258487,0.20749438,0.16976812,0.15467763,0.18485862,0.21503963,0.211267,0.14713238,0.1659955,0.20372175,0.24899325,0.30935526,0.422534,0.40367088,0.331991,0.32067314,0.35839936,0.3470815,0.2678564,0.2678564,0.2867195,0.32067314,0.44894236,0.482896,0.4678055,0.5696664,0.7394345,0.7205714,0.5281675,0.5319401,0.52062225,0.44139713,0.38480774,0.422534,0.3470815,0.27917424,0.29803738,0.39989826,0.38858038,0.41121614,0.38480774,0.30935526,0.2565385,0.36971724,0.5281675,0.60362,0.55080324,0.4376245,0.4678055,0.5885295,0.88279426,1.2638294,1.4901869,1.026154,0.77716076,0.7432071,0.83752275,0.875249,0.90920264,0.8111144,0.6752999,0.5696664,0.5583485,0.39989826,0.28294688,0.21503963,0.18485862,0.1659955,0.14713238,0.150905,0.16222288,0.17354076,0.18485862,0.2565385,0.32444575,0.3961256,0.47157812,0.56589377,0.5093044,0.44139713,0.43007925,0.45648763,0.43007925,0.3772625,0.33953625,0.35085413,0.40367088,0.44894236,0.3734899,0.36971724,0.392353,0.3961256,0.34330887,0.39989826,0.482896,0.513077,0.4640329,0.3734899,0.362172,0.38103512,0.43385187,0.49421388,0.4979865,0.43007925,0.44894236,0.45648763,0.41498876,0.35839936,0.38103512,0.41876137,0.41876137,0.38858038,0.4074435,0.30181,0.23013012,0.23767537,0.2867195,0.2678564,0.29049212,0.41498876,0.5281675,0.5885295,0.6149379,0.6187105,0.5583485,0.452715,0.35839936,0.35839936,0.39989826,0.39989826,0.41498876,0.44516975,0.43007925,0.49044126,0.543258,0.5696664,0.5772116,0.62625575,0.62248313,0.694163,0.7582976,0.8262049,0.98842776,1.026154,0.95824677,0.91297525,0.9242931,0.9393836,0.8978847,0.8903395,0.9242931,0.995973,1.0789708,1.1581959,1.1242423,1.0487897,0.98465514,0.9507015,0.9318384,1.0186088,1.0940613,1.0940613,1.0035182,1.0223814,1.1393328,1.1808317,1.0902886,0.9280658,0.8978847,0.90543,0.94692886,1.0110635,1.0789708,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1961765,0.5017591,0.7130261,0.7997965,0.8865669,0.995973,0.9016574,0.86770374,0.965792,1.0978339,2.173032,2.0485353,1.388326,0.79602385,0.80734175,0.69793564,0.9808825,1.1544232,0.9922004,0.56589377,0.44139713,0.5394854,0.7092535,0.754525,0.41121614,0.9620194,1.20724,1.3656902,1.50905,1.5731846,1.7165444,2.1956677,2.5314314,2.776652,3.5085413,8.099826,9.812597,10.303039,10.691619,11.581959,11.080199,11.604594,11.012292,8.729855,5.753253,3.410453,2.1013522,1.4449154,1.0827434,0.65643674,0.76584285,1.0035182,0.98465514,0.754525,0.77716076,0.76584285,0.56212115,0.44139713,0.47157812,0.52062225,0.32444575,0.24899325,0.16976812,0.09808825,0.18485862,0.2678564,0.25276586,0.23390275,0.29049212,0.47157812,0.38858038,0.27540162,0.12826926,0.0,0.0,0.1358145,0.13204187,0.094315626,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.15845025,0.25276586,0.41121614,0.422534,0.34330887,0.241448,0.150905,0.0754525,0.026408374,0.20749438,0.48666862,0.80356914,1.1431054,1.1204696,1.2789198,1.780679,2.3692086,2.3805263,4.406426,4.666737,4.4818783,4.4139714,4.2404304,3.7047176,4.561104,6.1342883,7.4471617,7.201941,8.375228,10.38981,11.993175,13.106099,14.815099,15.279131,14.517061,12.521342,10.163452,9.186342,10.235131,14.203933,15.535669,12.147853,5.4476705,8.243186,11.981857,11.619685,7.3151197,4.4101987,2.7502437,2.052308,1.9089483,2.1654868,2.897376,4.889322,7.960239,11.517824,15.30554,19.410156,25.253952,33.814037,50.25514,74.498024,101.19312,107.636765,97.96375,104.31686,137.2066,185.4962,183.75325,153.60997,118.24916,93.54978,88.05684,89.98465,84.82748,86.65343,106.81433,153.94574,130.65732,99.619934,88.02289,101.800514,125.63973,123.5497,111.89606,88.46429,59.113262,37.748886,31.622143,23.92976,18.251959,16.678776,19.791191,16.750456,14.709465,14.524607,15.611122,15.931795,16.380737,16.686321,16.060064,13.645585,8.529905,8.748717,9.684328,10.18986,10.167224,10.559577,8.801534,7.3377557,6.428553,6.2814207,7.0510364,13.909668,21.53037,22.688566,17.697384,14.388792,9.616421,7.6810646,7.5527954,8.929804,12.238396,10.725573,9.027891,8.284684,9.137298,11.747954,9.224068,9.899368,14.0983,21.062565,28.947351,33.255688,54.876602,93.87423,134.65253,145.99304,106.21071,83.75227,85.12551,102.85307,115.44987,106.35407,93.779915,82.243225,73.85668,68.32978,61.52774,54.401253,57.147724,69.24276,79.4213,58.841633,45.77703,39.446568,37.281082,34.911873,38.499638,39.88419,35.175957,26.287651,20.904116,16.754227,13.985121,14.211478,15.69412,13.35132,14.120935,14.871688,16.097792,18.21046,21.53037,21.568098,21.228561,21.032385,20.945614,20.387266,23.767538,31.305243,35.896526,35.043915,30.867619,25.216225,21.194607,21.598278,28.038149,40.936752,25.155863,16.0827,15.912932,19.742147,15.580941,21.41342,18.761265,14.154889,13.041965,19.806282,19.304522,12.313848,10.340765,14.5283785,15.641303,10.95193,14.743419,16.293968,15.086727,20.813572,9.80128,6.519096,5.4740787,4.715781,5.8136153,8.329956,6.119198,5.73439,7.383027,4.927048,4.3422914,4.9459114,5.5759397,5.9192486,6.515323,9.092027,11.0613365,11.295239,9.876732,8.118689,7.069899,6.779407,7.533932,9.58624,13.13628,13.70972,11.208468,8.390318,6.1795597,3.6783094,2.3465726,1.8938577,2.1654868,2.674791,2.6408374,3.1652324,2.0787163,1.2713746,1.50905,2.425798,3.3048196,4.1008434,4.7308717,4.847823,3.8593953,4.1762958,5.594803,5.485397,3.6858547,2.5012503,2.0258996,2.082489,2.9237845,4.195159,4.9119577,4.2894745,4.191386,3.5500402,2.6597006,3.1576872,1.841041,1.0072908,0.72811663,0.8639311,1.0827434,1.0110635,0.83752275,0.58098423,0.3055826,0.120724,0.694163,2.2296214,1.931584,0.18863125,0.58098423,0.3734899,0.1659955,0.056589376,0.120724,0.42630664,2.4031622,1.4524606,0.5055317,0.543258,0.58098423,0.43385187,0.23013012,0.10940613,0.15467763,0.41121614,0.8262049,0.63002837,0.32444575,0.14713238,0.060362,0.10940613,0.1659955,0.181086,0.15467763,0.1659955,0.31312788,0.38858038,0.44139713,0.49044126,0.5017591,0.79602385,1.0072908,1.4637785,2.7691069,5.783434,4.3686996,3.1350515,1.9240388,0.9507015,0.7922512,0.35462674,0.16976812,0.13958712,0.17354076,0.19994913,0.6488915,1.0638802,1.3807807,1.5430037,1.4939595,1.1431054,1.1091517,1.2902378,1.327964,0.59607476,0.5093044,0.4074435,0.28294688,0.1659955,0.1056335,0.0452715,0.056589376,0.10186087,0.120724,0.060362,0.011317875,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.1056335,0.26408374,0.26031113,0.18485862,0.10940613,0.060362,0.18485862,0.43385187,0.45648763,0.26408374,0.23013012,0.23013012,0.23013012,0.18485862,0.1056335,0.030181,0.018863125,0.00754525,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.033953626,0.0452715,0.049044125,0.060362,0.14713238,0.241448,0.29049212,0.2678564,0.18485862,0.14713238,0.12826926,0.15845025,0.20749438,0.18485862,0.1358145,0.13958712,0.1659955,0.20372175,0.29049212,0.47157812,0.41876137,0.35085413,0.3470815,0.33576363,0.27540162,0.26031113,0.26408374,0.27917424,0.29049212,0.46026024,0.4678055,0.46026024,0.5357128,0.73188925,0.6451189,0.62625575,0.5772116,0.482896,0.3961256,0.44516975,0.422534,0.36594462,0.33953625,0.41121614,0.44894236,0.44894236,0.392353,0.3055826,0.24522063,0.4640329,0.59230214,0.59230214,0.52062225,0.5357128,0.6451189,0.6149379,0.8601585,1.4411428,2.0749438,1.7580433,1.1921495,0.7922512,0.7054809,0.83752275,0.9507015,0.8299775,0.7092535,0.65643674,0.59607476,0.38858038,0.27917424,0.20749438,0.150905,0.150905,0.150905,0.16976812,0.20749438,0.24899325,0.26031113,0.36971724,0.5055317,0.5055317,0.3961256,0.3961256,0.3470815,0.33576363,0.32444575,0.29426476,0.26031113,0.28294688,0.27917424,0.29426476,0.33953625,0.41121614,0.32821837,0.35085413,0.38858038,0.38103512,0.32067314,0.35839936,0.422534,0.44516975,0.41121614,0.35085413,0.3734899,0.392353,0.36594462,0.33953625,0.41121614,0.32821837,0.26031113,0.23390275,0.24899325,0.27540162,0.27540162,0.30181,0.32821837,0.34330887,0.38103512,0.30935526,0.24522063,0.24522063,0.3055826,0.36594462,0.42630664,0.56212115,0.6413463,0.63002837,0.58098423,0.49421388,0.4640329,0.452715,0.44516975,0.45648763,0.422534,0.392353,0.41876137,0.47912338,0.5017591,0.51684964,0.45648763,0.39989826,0.392353,0.44139713,0.43007925,0.45648763,0.5093044,0.573439,0.6111652,0.7432071,0.87902164,0.9393836,0.9016574,0.7922512,0.7809334,0.7884786,0.7922512,0.8224323,0.94692886,1.0940613,1.2562841,1.2826926,1.1581959,1.0374719,0.98842776,0.9507015,0.935611,0.9808825,1.1129243,1.1129243,1.0487897,1.0299267,1.0487897,0.97710985,0.9280658,0.87902164,0.8186596,0.77338815,0.8224323,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14713238,0.36594462,0.55080324,0.65643674,0.7130261,0.88279426,0.97333723,1.0412445,1.056335,0.91674787,1.0714256,1.2751472,1.146878,0.9280658,1.4675511,1.327964,1.2298758,1.0223814,0.73566186,0.5998474,0.5281675,0.573439,0.62625575,0.663982,0.7432071,0.9016574,1.0412445,1.3770081,1.9164935,2.4861598,3.1614597,3.1916409,3.169005,3.187868,2.837014,5.1345425,6.990674,8.699674,9.4127,7.1378064,5.621211,5.7607985,6.1644692,5.836251,4.164978,1.9278114,0.875249,0.5281675,0.56212115,0.7922512,0.7432071,0.73188925,0.66775465,0.5696664,0.5357128,0.43385187,0.362172,0.3772625,0.452715,0.482896,0.36594462,0.2565385,0.181086,0.12826926,0.03772625,0.05281675,0.049044125,0.06790725,0.116951376,0.19240387,0.23390275,0.20372175,0.15845025,0.14335975,0.18485862,0.211267,0.21503963,0.1358145,0.011317875,0.0,0.0,0.0,0.0,0.011317875,0.049044125,0.06790725,0.116951376,0.241448,0.43385187,0.63002837,0.60362,0.35462674,0.15467763,0.08677038,0.06413463,0.033953626,0.08677038,0.211267,0.40367088,0.65643674,0.67152727,1.0751982,1.5015048,2.04099,3.2331395,3.289729,3.640583,3.6141748,3.1199608,2.655928,3.3764994,5.036454,6.7114997,7.7037,7.5565677,8.601585,9.88805,10.899114,12.117672,15.0376835,12.970284,11.385782,10.842525,11.415963,12.67602,17.701157,30.316814,34.353523,24.895552,8.29223,6.7114997,6.8246784,6.085244,4.195159,3.0671442,2.1277604,1.6863633,1.6109109,2.1051247,3.6556737,7.069899,13.238141,21.194607,29.57738,36.620872,52.23954,77.55008,108.93077,139.91158,161.18918,141.68848,110.783134,93.051796,98.14484,120.77304,126.330124,120.92017,119.479034,126.79415,137.49332,128.53334,127.95612,139.10046,156.08481,163.79607,123.71947,100.76304,108.719505,147.12483,201.24313,211.5575,173.26535,118.81128,70.74804,41.69128,33.90458,24.397566,16.950403,15.184815,22.575388,17.923742,15.120681,16.01102,19.025349,19.176252,20.655123,19.794964,15.894069,11.246195,11.129244,12.736382,11.876224,10.808571,11.099063,13.645585,12.623203,10.880251,11.54046,13.93985,13.615403,16.444872,21.202152,21.78691,18.176508,16.4411,15.241405,12.325166,8.918486,6.6020937,7.2924843,8.809079,10.650121,10.370946,9.593785,14.030393,13.664448,12.419481,13.185325,17.516298,25.63876,32.142765,48.00288,84.155945,137.76117,192.16997,172.09206,126.379166,100.480095,106.5842,123.61383,120.85604,103.56233,90.81086,87.555084,84.62375,77.97261,62.565212,53.186466,56.04989,68.827774,57.913567,47.169132,41.423424,40.208637,37.779068,41.027298,43.268234,43.313507,39.13344,27.860836,19.610106,14.139798,11.955449,11.887542,11.117926,12.404391,13.555041,14.875461,16.399601,17.89356,18.97253,20.11941,20.65135,20.217497,18.787672,21.036158,27.272306,32.68225,34.108303,30.048958,31.64478,22.782883,17.14658,19.040438,23.39782,26.793182,19.108345,15.313085,17.780382,16.324148,21.51528,16.188334,10.518079,9.540969,13.189097,24.397566,17.89356,12.943876,15.641303,18.900852,11.487643,12.472299,16.143063,19.866644,24.107073,10.676529,6.0701537,4.8629136,4.508287,5.311856,6.7944975,5.934339,6.1908774,7.7037,7.3075747,6.6360474,6.017337,6.1041074,6.6360474,6.4549613,5.836251,7.1340337,8.284684,8.050782,6.0286546,6.7756343,6.6662283,7.0057645,8.118689,9.318384,9.473062,9.039209,7.1679873,4.293247,2.1503963,1.659955,1.418507,1.7655885,2.655928,3.663219,3.7990334,3.0105548,1.9768555,1.3015556,1.5241405,1.931584,2.444661,3.169005,3.7650797,3.4217708,3.2029586,4.357382,4.606375,3.3727267,1.8184053,1.20724,0.95447415,1.2223305,1.9693103,2.9728284,2.2409391,2.3805263,2.2598023,2.0787163,3.3425457,1.9164935,1.2034674,0.98465514,0.9318384,0.59607476,0.513077,0.38858038,0.271629,0.17731337,0.071679875,0.76584285,2.263575,2.022127,0.331991,0.32444575,1.3166461,0.91297525,0.29426476,0.056589376,0.1961765,1.0299267,0.8111144,0.43007925,0.29049212,0.29803738,0.29049212,0.18863125,0.14335975,0.18485862,0.21503963,0.3961256,0.38103512,0.2565385,0.16976812,0.32821837,0.30935526,0.18863125,0.08299775,0.049044125,0.071679875,0.18863125,0.26031113,0.3169005,0.36971724,0.43007925,0.65643674,1.0902886,1.4600059,2.252257,4.708236,3.6745367,2.6031113,1.6146835,0.995973,1.20724,0.58475685,0.271629,0.13958712,0.08677038,0.06413463,0.36971724,0.6073926,0.8865669,1.1355602,1.1053791,0.8563859,0.7922512,0.80356914,0.724344,0.31312788,0.20749438,0.17354076,0.14335975,0.09808825,0.0452715,0.02263575,0.02263575,0.041498873,0.06413463,0.060362,0.02263575,0.00754525,0.00754525,0.011317875,0.0,0.030181,0.0150905,0.0,0.0150905,0.056589376,0.12826926,0.150905,0.12826926,0.071679875,0.02263575,0.049044125,0.120724,0.14713238,0.14335975,0.25276586,0.1961765,0.120724,0.07922512,0.071679875,0.06790725,0.094315626,0.056589376,0.018863125,0.018863125,0.041498873,0.0754525,0.049044125,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.02263575,0.041498873,0.060362,0.071679875,0.13958712,0.20749438,0.271629,0.31312788,0.3055826,0.19994913,0.1659955,0.1659955,0.17731337,0.18485862,0.11317875,0.10186087,0.13204187,0.181086,0.23013012,0.34330887,0.35839936,0.33953625,0.32821837,0.33576363,0.28294688,0.24899325,0.241448,0.25276586,0.26408374,0.32821837,0.42630664,0.49421388,0.52439487,0.573439,0.6149379,0.62625575,0.55080324,0.452715,0.49421388,0.47535074,0.42630664,0.44516975,0.5093044,0.48666862,0.44516975,0.41498876,0.4074435,0.3961256,0.36594462,0.5470306,0.6451189,0.6488915,0.60362,0.6073926,0.66020936,0.5281675,0.56212115,0.9280658,1.6109109,2.0447628,1.9994912,1.5316857,0.9205205,0.6451189,0.7130261,0.70170826,0.66775465,0.6187105,0.5093044,0.38858038,0.362172,0.32067314,0.23767537,0.18863125,0.18863125,0.16976812,0.1961765,0.26031113,0.28294688,0.35462674,0.4678055,0.47157812,0.4074435,0.49421388,0.3961256,0.32821837,0.29803738,0.2867195,0.26031113,0.27540162,0.28294688,0.29049212,0.3055826,0.35085413,0.392353,0.43385187,0.44516975,0.4074435,0.30935526,0.2678564,0.25276586,0.24899325,0.23767537,0.21503963,0.271629,0.32067314,0.29803738,0.23390275,0.27917424,0.33953625,0.35839936,0.3772625,0.3961256,0.35839936,0.36971724,0.38480774,0.36971724,0.33953625,0.35839936,0.35085413,0.29803738,0.2678564,0.29426476,0.35462674,0.41498876,0.44516975,0.5055317,0.56589377,0.5055317,0.41121614,0.4074435,0.44516975,0.47912338,0.482896,0.513077,0.52439487,0.51684964,0.4979865,0.49044126,0.49421388,0.47535074,0.4678055,0.47535074,0.4678055,0.47535074,0.51684964,0.5470306,0.56212115,0.6111652,0.68661773,0.7469798,0.7884786,0.80356914,0.7809334,0.72811663,0.72811663,0.68661773,0.633801,0.6790725,0.754525,0.7997965,0.8299775,0.84129536,0.80734175,0.7167987,0.76207024,0.8262049,0.88279426,1.0148361,1.0638802,1.0638802,0.97333723,0.8337501,0.7809334,0.8111144,0.73566186,0.6526641,0.6073926,0.6149379,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.120724,0.241448,0.35839936,0.45648763,0.543258,0.69793564,0.9205205,1.0601076,1.0336993,0.84129536,1.0412445,1.1053791,1.0374719,1.2223305,2.4182527,1.9579924,1.5241405,1.1280149,0.84129536,0.7582976,0.784706,0.98842776,1.1506506,1.2034674,1.2525115,1.3732355,1.5920477,2.0108092,2.565385,3.0256453,3.218049,3.2670932,3.4934506,3.5424948,2.3880715,2.7540162,3.5387223,4.6214657,5.1156793,3.3915899,2.3692086,2.1202152,2.3088465,2.4559789,1.9579924,0.7884786,0.26408374,0.1358145,0.21503963,0.38480774,0.43007925,0.392353,0.33953625,0.30935526,0.3169005,0.26031113,0.24899325,0.36971724,0.56212115,0.59230214,0.5394854,0.32444575,0.13958712,0.05281675,0.0,0.0,0.0,0.011317875,0.030181,0.049044125,0.07922512,0.0754525,0.06790725,0.071679875,0.090543,0.19240387,0.52062225,0.6526641,0.4376245,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.071679875,0.124496624,0.271629,0.482896,0.66775465,0.573439,0.32444575,0.1358145,0.06790725,0.041498873,0.049044125,0.0754525,0.23767537,0.5583485,0.97333723,0.95447415,1.5052774,2.1768045,2.8106055,3.531177,3.1954134,3.006782,3.0822346,3.2859564,3.2482302,4.3875628,5.8626595,6.9680386,7.3113475,6.802043,7.3113475,8.27714,9.333474,10.552032,12.472299,11.18206,10.284176,9.563604,9.020347,8.892077,12.30253,24.061802,29.135983,22.198126,7.6282477,6.700182,5.6287565,4.402653,3.3236825,3.0143273,1.8485862,1.3807807,1.6146835,2.686109,4.851596,8.778898,14.996184,22.39053,30.343224,38.76372,57.362762,81.79051,109.00246,133.17366,145.73651,124.538124,102.60786,89.30935,88.89813,100.548004,114.45767,124.24009,134.88266,140.5152,124.4174,96.15289,94.06286,113.12971,140.07379,153.37984,128.89174,110.239876,120.90508,164.92407,226.87434,234.47241,196.19914,137.73099,81.50379,46.671143,33.764996,24.080666,17.452164,15.226315,20.22127,17.357847,15.845025,17.157898,19.293203,16.776863,18.09351,20.768301,18.101055,11.41219,10.050273,11.608367,10.646348,10.8576145,12.510024,12.479843,10.79348,10.008774,10.250222,11.638548,14.27184,16.91645,18.229324,18.8254,18.689585,17.172989,13.65313,10.352083,7.462252,5.715527,6.368191,6.749226,10.121953,14.815099,17.237123,11.864905,16.365646,17.48989,16.531643,17.14658,25.359585,37.51121,49.315754,76.85592,125.46619,189.71399,224.64096,200.1453,161.09486,138.09317,147.45305,152.3386,131.72874,124.741844,135.78809,134.58086,105.165695,76.576744,56.823277,50.436222,58.460598,55.63867,47.867065,42.883427,42.924927,44.732014,45.28659,43.03056,42.890972,42.66839,33.051968,23.835445,17.637022,14.543469,13.389046,11.747954,11.898859,12.551523,13.773854,15.339493,16.735365,17.640795,18.89708,20.69662,21.322876,17.176762,18.595268,25.435038,31.550463,34.08944,33.482048,34.75342,25.378448,20.157135,21.734093,20.587215,29.524563,21.85859,18.693357,24.024076,24.729557,21.028612,19.383747,15.490398,11.966766,18.372684,20.907888,17.723793,15.0905,15.418718,17.252214,12.770335,10.627484,16.501461,26.8045,28.694586,13.219278,9.733373,8.722309,6.8774953,7.0812173,5.0968165,6.368191,7.816879,8.6732645,10.495442,9.608876,7.1264887,6.8473144,8.635539,8.424272,6.519096,6.7454534,8.326183,9.088254,5.462761,5.5759397,5.13077,4.6629643,4.436607,4.4630156,4.2894745,4.5460134,3.832987,2.2447119,1.358145,1.2298758,0.95447415,1.0110635,1.6033657,2.6295197,3.2520027,3.338773,2.5729303,1.4637785,1.3430545,1.1581959,1.3430545,2.1088974,3.150142,3.640583,3.7047176,3.7952607,3.5689032,2.8785129,1.8033148,1.8749946,1.2110126,0.8563859,1.0751982,1.3430545,1.026154,1.1280149,1.2185578,1.358145,2.0787163,1.3958713,1.0336993,0.94315624,0.8941121,0.5017591,0.2678564,0.15845025,0.116951376,0.09808825,0.041498873,0.72811663,1.8485862,1.7769064,0.60362,0.150905,1.6033657,1.6184561,0.86770374,0.08677038,0.071679875,0.34330887,0.35839936,0.26408374,0.17354076,0.17354076,0.3734899,0.23767537,0.124496624,0.1358145,0.11317875,0.26408374,0.30181,0.241448,0.17354076,0.27917424,0.31312788,0.19994913,0.11317875,0.10940613,0.12826926,0.17354076,0.24522063,0.35462674,0.4376245,0.35839936,0.6149379,1.478869,1.9579924,2.1277604,3.1124156,2.957738,2.1881225,1.3505998,0.8941121,1.146878,0.80734175,0.41876137,0.18485862,0.11317875,0.041498873,0.241448,0.44894236,0.5583485,0.5696664,0.5583485,0.6451189,0.8601585,0.9318384,0.7582976,0.392353,0.15467763,0.1056335,0.090543,0.049044125,0.02263575,0.00754525,0.011317875,0.0150905,0.018863125,0.02263575,0.018863125,0.00754525,0.003772625,0.003772625,0.0,0.02263575,0.0150905,0.003772625,0.003772625,0.026408374,0.14335975,0.17354076,0.13204187,0.056589376,0.0150905,0.00754525,0.018863125,0.026408374,0.060362,0.17731337,0.16222288,0.08677038,0.041498873,0.08299775,0.21503963,0.18485862,0.120724,0.06413463,0.033953626,0.026408374,0.041498873,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.041498873,0.0754525,0.094315626,0.13958712,0.21881226,0.28294688,0.30935526,0.29803738,0.22258487,0.19240387,0.17354076,0.15467763,0.14713238,0.10186087,0.08677038,0.10940613,0.16222288,0.20372175,0.24899325,0.3169005,0.35839936,0.35462674,0.30935526,0.23767537,0.23767537,0.25276586,0.26408374,0.27917424,0.2867195,0.31312788,0.38858038,0.47157812,0.46026024,0.4678055,0.52439487,0.573439,0.573439,0.49044126,0.44894236,0.36971724,0.3772625,0.49044126,0.63002837,0.5394854,0.43007925,0.3772625,0.39989826,0.43385187,0.5885295,0.68661773,0.663982,0.55457586,0.48666862,0.47912338,0.362172,0.33953625,0.4979865,0.8262049,1.177059,1.5958204,1.5052774,0.97333723,0.694163,0.6752999,0.59607476,0.55080324,0.5470306,0.4979865,0.392353,0.35839936,0.30935526,0.23767537,0.20749438,0.20749438,0.20372175,0.2565385,0.36594462,0.45648763,0.45648763,0.4678055,0.41876137,0.34330887,0.3734899,0.33576363,0.3169005,0.3169005,0.3169005,0.2867195,0.23390275,0.24899325,0.31312788,0.38103512,0.4074435,0.43007925,0.44894236,0.4074435,0.32067314,0.27917424,0.3055826,0.29426476,0.27540162,0.26408374,0.23013012,0.21503963,0.22258487,0.23390275,0.24899325,0.26408374,0.38103512,0.47535074,0.52062225,0.4979865,0.38103512,0.35839936,0.35085413,0.331991,0.3055826,0.2867195,0.28294688,0.30181,0.3169005,0.32444575,0.3055826,0.41876137,0.392353,0.3961256,0.47157812,0.543258,0.46026024,0.4678055,0.48666862,0.482896,0.47157812,0.5394854,0.6111652,0.62248313,0.5772116,0.543258,0.5583485,0.5470306,0.52062225,0.49421388,0.5017591,0.482896,0.44894236,0.41121614,0.3961256,0.44516975,0.5357128,0.5583485,0.5583485,0.5998474,0.7582976,0.77338815,0.724344,0.6187105,0.55080324,0.6828451,0.5998474,0.5319401,0.55080324,0.633801,0.6752999,0.56212115,0.5998474,0.65643674,0.7054809,0.8186596,0.814887,0.8224323,0.8224323,0.7809334,0.6488915,0.6413463,0.5470306,0.4640329,0.44139713,0.4640329,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06413463,0.1659955,0.2263575,0.2565385,0.3470815,0.482896,0.72811663,0.95824677,1.1129243,1.2034674,1.7165444,1.5203679,1.478869,2.022127,3.097325,2.323937,1.9881734,1.8221779,1.6486372,1.4147344,1.3468271,1.5316857,1.6260014,1.5618668,1.5354583,1.7919968,2.0145817,2.4710693,3.0709167,3.3764994,3.1840954,3.127506,3.2255943,3.0746894,1.8561316,1.3996439,1.3845534,1.690136,1.8825399,1.1732863,0.79602385,0.482896,0.3734899,0.4376245,0.44894236,0.16222288,0.03772625,0.0150905,0.0452715,0.08677038,0.18485862,0.17354076,0.14335975,0.14335975,0.17731337,0.1659955,0.1659955,0.25276586,0.38103512,0.40367088,0.38858038,0.21881226,0.06413463,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.033953626,0.026408374,0.0150905,0.0,0.0,0.150905,0.52062225,0.66775465,0.4376245,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.03772625,0.0754525,0.19994913,0.38480774,0.55080324,0.422534,0.23390275,0.09808825,0.0452715,0.02263575,0.05281675,0.17354076,0.5093044,0.94315624,1.1091517,1.1431054,1.901403,2.916239,3.7235808,3.874486,3.4670424,3.451952,3.7386713,4.146115,4.3686996,5.564622,7.624475,8.831716,8.563859,7.2887115,7.2472124,7.907422,8.631766,9.107117,9.348565,9.623966,10.114408,9.955957,8.83926,7.020855,7.1793056,12.559069,15.46399,12.743927,5.7796617,6.255012,5.413717,4.538468,4.7006907,6.7756343,4.478106,4.3385186,4.5535583,4.870459,6.5568223,10.748209,15.015047,20.22127,27.057266,36.054977,49.621338,66.6057,86.2573,104.29044,112.87317,97.2545,88.88682,86.11394,88.045525,94.541985,101.97783,109.919205,116.55525,112.82412,82.45449,53.73727,50.41359,66.137886,91.3013,113.04294,108.39129,100.23865,109.22504,141.90352,190.74014,194.28264,173.26158,132.69453,85.12928,50.6324,32.82561,23.61286,19.58747,18.16519,17.591751,16.720274,16.708956,18.617905,20.7268,18.516043,17.746428,20.013775,18.938578,14.290704,12.00072,13.321139,12.774108,14.264296,16.803272,14.505743,12.679792,11.993175,10.585986,9.35611,11.940358,13.717264,12.989148,13.389046,15.290449,15.83748,10.782163,8.303548,6.7114997,5.987156,7.7602897,7.4471617,8.763808,13.230596,16.878725,10.231359,15.90916,19.055529,18.700903,18.912169,28.78513,42.460896,50.334362,64.97592,96.20571,151.09363,233.76317,243.1155,213.74184,179.9693,175.81564,174.98944,151.93115,150.64468,174.416,185.84705,139.56071,101.09126,73.634094,59.54711,60.339363,54.027763,47.335125,43.479504,44.418888,50.858757,48.723454,42.28358,40.650036,42.67216,36.930225,27.491117,20.877707,17.229578,15.501716,13.45318,14.226569,14.34352,14.977322,16.618414,19.078165,18.802763,19.447882,22.941332,25.370903,16.999449,18.489635,24.393793,29.841463,32.64075,33.267006,33.44432,26.08393,22.07363,23.054512,21.405874,28.702131,23.314823,21.454918,27.072357,31.829638,19.670467,18.48209,16.490145,12.785426,17.323895,16.791954,16.022339,14.939595,13.973803,14.034165,11.744182,8.507269,14.000212,24.657877,23.68454,12.638294,11.378237,11.242422,9.691874,10.280403,5.4665337,6.628502,7.6508837,7.5188417,10.329447,9.759781,6.8925858,6.270103,8.07719,8.114917,6.4210076,6.398372,7.8696957,8.627994,4.436607,3.9008942,3.3689542,2.584248,1.7731338,1.6524098,1.2826926,1.4675511,1.358145,0.9205205,0.9507015,0.9242931,0.69793564,0.59607476,0.8224323,1.4637785,2.191895,2.7200627,2.3201644,1.327964,1.1544232,0.8224323,0.7696155,1.569412,3.1010978,4.538468,4.436607,3.6141748,2.8106055,2.2371666,1.5882751,1.9542197,1.5203679,1.5241405,1.841041,0.9808825,0.5281675,0.46026024,0.5772116,0.77338815,1.0412445,1.1242423,0.88279426,0.73566186,0.7809334,0.7809334,0.47912338,0.29803738,0.20372175,0.17354076,0.1659955,0.6073926,1.2638294,1.3920987,0.8865669,0.25276586,1.1996948,1.6335466,1.1808317,0.26031113,0.090543,0.14335975,0.17354076,0.18863125,0.1961765,0.21503963,0.38103512,0.24899325,0.124496624,0.120724,0.120724,0.23767537,0.2867195,0.2565385,0.20749438,0.271629,0.362172,0.32067314,0.23013012,0.15467763,0.15845025,0.17354076,0.19240387,0.2867195,0.4074435,0.3734899,0.5055317,1.267602,2.082489,2.5314314,2.3616633,2.2748928,1.8485862,1.3505998,1.0336993,1.1431054,1.0638802,0.6451189,0.3055826,0.17731337,0.120724,0.25276586,0.422534,0.45648763,0.362172,0.362172,0.5696664,0.97333723,1.2110126,1.0978339,0.6526641,0.35085413,0.211267,0.124496624,0.05281675,0.0150905,0.003772625,0.003772625,0.003772625,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.011317875,0.018863125,0.018863125,0.011317875,0.00754525,0.12826926,0.18485862,0.15845025,0.071679875,0.0150905,0.011317875,0.02263575,0.018863125,0.0150905,0.071679875,0.116951376,0.116951376,0.14713238,0.2263575,0.33576363,0.20372175,0.13958712,0.10186087,0.071679875,0.056589376,0.06413463,0.049044125,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.00754525,0.011317875,0.03772625,0.071679875,0.08299775,0.124496624,0.19994913,0.2678564,0.3055826,0.27917424,0.2678564,0.24522063,0.21881226,0.181086,0.116951376,0.10940613,0.08299775,0.08299775,0.124496624,0.16222288,0.18485862,0.26408374,0.33953625,0.362172,0.29049212,0.22258487,0.24899325,0.28294688,0.2867195,0.29049212,0.2678564,0.241448,0.2867195,0.38103512,0.4074435,0.43385187,0.5017591,0.6073926,0.6828451,0.5772116,0.47912338,0.38480774,0.36971724,0.46026024,0.63002837,0.59607476,0.44516975,0.3470815,0.36971724,0.47535074,0.6451189,0.72811663,0.70170826,0.5998474,0.49421388,0.41498876,0.33576363,0.29803738,0.29803738,0.32067314,0.43385187,0.845068,0.97333723,0.77338815,0.7394345,0.7092535,0.56589377,0.49421388,0.52062225,0.51684964,0.3772625,0.3169005,0.27917424,0.241448,0.24522063,0.26031113,0.26408374,0.3169005,0.41498876,0.51684964,0.49044126,0.4376245,0.36594462,0.30181,0.2867195,0.271629,0.29049212,0.32821837,0.35462674,0.33576363,0.30181,0.29049212,0.32821837,0.39989826,0.45648763,0.41498876,0.41498876,0.3734899,0.29803738,0.27917424,0.33953625,0.32821837,0.29426476,0.26408374,0.23390275,0.18485862,0.15845025,0.1961765,0.271629,0.3169005,0.392353,0.49044126,0.543258,0.5319401,0.45648763,0.4678055,0.44139713,0.3772625,0.30935526,0.2867195,0.27540162,0.32821837,0.38480774,0.38858038,0.3055826,0.3772625,0.32821837,0.29426476,0.35085413,0.49421388,0.43007925,0.44139713,0.4678055,0.47157812,0.45648763,0.513077,0.6073926,0.6526641,0.6451189,0.6451189,0.66775465,0.6526641,0.6187105,0.5772116,0.543258,0.48666862,0.4376245,0.38480774,0.33953625,0.3470815,0.41876137,0.43007925,0.422534,0.46026024,0.6149379,0.69039035,0.67152727,0.58098423,0.513077,0.6413463,0.58475685,0.49421388,0.452715,0.47535074,0.5093044,0.44516975,0.48666862,0.55080324,0.6111652,0.7092535,0.663982,0.6752999,0.73188925,0.754525,0.5998474,0.52439487,0.482896,0.422534,0.35839936,0.3734899,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10940613,0.14335975,0.09808825,0.14713238,0.29803738,0.47157812,0.7394345,1.1280149,1.599593,2.1315331,1.9240388,2.1579416,2.9501927,3.3312278,2.474842,2.4861598,2.7313805,2.8106055,2.5578396,2.305074,2.2258487,2.0749438,1.8636768,1.8749946,1.9391292,1.9353566,2.4031622,3.169005,3.350091,3.2331395,2.8822856,2.4597516,1.9655377,1.2261031,0.91674787,0.7922512,0.8563859,0.88279426,0.4376245,0.29049212,0.18863125,0.11317875,0.06413463,0.018863125,0.003772625,0.011317875,0.018863125,0.030181,0.060362,0.10186087,0.08677038,0.07922512,0.090543,0.116951376,0.1056335,0.1056335,0.071679875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.08677038,0.06413463,0.05281675,0.030181,0.0,0.0,0.09808825,0.1961765,0.14713238,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0754525,0.22258487,0.3734899,0.2565385,0.12826926,0.0452715,0.018863125,0.0150905,0.05281675,0.3169005,0.7922512,1.1959221,0.9695646,1.1959221,2.161714,3.3878171,4.29702,4.2102494,4.134797,5.142088,5.7872066,5.726845,5.715527,6.8699503,9.578695,10.948157,10.167224,8.507269,8.36391,8.82417,8.971302,8.492179,7.6886096,8.748717,9.906913,10.597303,10.220041,8.130007,6.417235,5.9305663,5.621211,5.342037,5.8211603,7.115171,7.413208,7.4207535,8.348819,11.9064045,9.159933,9.854096,9.910686,8.465771,7.8508325,13.079691,14.875461,18.010511,25.027594,36.220974,40.023777,49.02149,63.12356,78.62905,88.20397,76.80687,72.90221,73.9774,77.53122,81.111435,72.28349,68.37505,65.47768,58.339874,40.34068,30.113092,28.102283,32.154083,41.63469,57.43067,63.43669,68.97113,77.10868,92.18409,119.78839,126.41689,124.873886,108.379974,79.86647,51.983,32.27858,23.099783,21.934042,24.065575,22.571615,22.854563,22.269806,22.982832,24.725784,24.801237,21.50019,18.991394,17.614386,16.886269,15.528125,17.05981,17.139036,18.595268,20.447628,17.931286,16.705183,15.369675,12.808062,9.899368,9.495697,9.4013815,8.865668,9.635284,12.057309,15.098045,11.106608,9.559832,8.058327,6.9152217,9.171251,10.61994,8.367682,7.224577,8.650629,10.7557535,13.837989,16.497688,17.637022,20.111864,30.731804,41.33665,45.267727,48.100967,60.395954,97.69967,191.96625,223.96942,220.0459,202.43529,189.25374,172.20525,148.0793,146.72493,171.1791,197.6516,160.72891,123.56856,93.629005,75.57323,71.249794,52.48476,44.577335,41.940273,43.298416,51.688736,48.632908,40.94807,38.499638,41.098976,38.50341,29.728285,22.816835,18.523588,16.392056,14.724555,18.663176,19.25925,18.489635,18.565088,21.918951,21.224789,21.749184,27.56657,32.248398,18.874443,20.11941,23.360094,27.223263,29.773556,28.509727,28.664404,24.322113,20.68153,19.723284,20.22127,24.325886,24.80501,24.699375,26.551735,32.399303,18.69713,14.498198,13.023102,11.057564,8.959985,14.471789,14.675511,13.479589,12.528888,11.204697,9.473062,7.3981175,9.242931,13.264549,11.7026825,10.325675,10.544487,11.336739,12.113899,12.706201,7.466025,6.511551,5.7117543,4.847823,7.5829763,7.6093845,5.4476705,4.4215164,5.0666356,5.138315,4.3007927,4.7346444,5.753253,5.881522,2.8521044,2.3088465,2.2786655,2.0787163,1.7354075,1.9730829,1.3430545,1.0525624,0.7922512,0.56589377,0.69039035,0.66775465,0.6375736,0.633801,0.7092535,0.935611,1.1355602,1.4637785,1.3241913,0.814887,0.724344,0.6790725,0.56212115,1.3317367,3.0822346,5.0175915,4.5422406,3.5462675,2.4823873,1.6146835,1.0148361,1.1129243,1.3958713,2.3277097,3.1124156,1.6750455,0.543258,0.271629,0.3169005,0.46026024,0.7809334,1.1544232,0.8299775,0.55080324,0.6752999,1.1581959,0.8865669,0.5885295,0.38480774,0.33576363,0.452715,0.5017591,0.77338815,1.0186088,1.0223814,0.573439,0.59230214,1.0789708,1.056335,0.47535074,0.19240387,0.2263575,0.21881226,0.23767537,0.2867195,0.30181,0.24522063,0.19240387,0.15467763,0.150905,0.19994913,0.21503963,0.2565385,0.25276586,0.2565385,0.4376245,0.4979865,0.4979865,0.362172,0.16222288,0.120724,0.14335975,0.08677038,0.10186087,0.26031113,0.573439,0.4678055,0.62248313,1.629774,2.8898308,2.5917933,1.7165444,1.4939595,1.4034165,1.2562841,1.20724,1.1921495,0.814887,0.4376245,0.24522063,0.25276586,0.35462674,0.422534,0.482896,0.5281675,0.52062225,0.55457586,0.87147635,1.1695137,1.2147852,0.83752275,0.56212115,0.34330887,0.18863125,0.08677038,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.02263575,0.030181,0.02263575,0.0,0.05281675,0.1358145,0.150905,0.08299775,0.011317875,0.02263575,0.071679875,0.07922512,0.033953626,0.003772625,0.0754525,0.15845025,0.2867195,0.41876137,0.422534,0.20749438,0.13958712,0.12826926,0.124496624,0.116951376,0.150905,0.19994913,0.16222288,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.00754525,0.026408374,0.05281675,0.049044125,0.094315626,0.1358145,0.20749438,0.29049212,0.28294688,0.32067314,0.29803738,0.26031113,0.211267,0.1056335,0.116951376,0.0754525,0.056589376,0.08299775,0.10940613,0.13958712,0.20372175,0.27540162,0.31312788,0.271629,0.24899325,0.271629,0.29426476,0.29049212,0.27917424,0.24899325,0.23013012,0.23390275,0.27540162,0.36594462,0.47912338,0.52439487,0.58475685,0.67152727,0.70170826,0.55457586,0.46026024,0.44139713,0.482896,0.5319401,0.56589377,0.43007925,0.32067314,0.33953625,0.5055317,0.7130261,0.7582976,0.76207024,0.754525,0.6828451,0.5583485,0.47912338,0.40367088,0.32067314,0.23013012,0.24899325,0.30935526,0.36971724,0.45648763,0.663982,0.7130261,0.59230214,0.5055317,0.5055317,0.4979865,0.33576363,0.27917424,0.2678564,0.27540162,0.29803738,0.331991,0.33576363,0.36594462,0.422534,0.47912338,0.49044126,0.422534,0.3470815,0.30181,0.30181,0.2565385,0.29049212,0.34330887,0.38103512,0.3734899,0.41498876,0.36971724,0.33576363,0.3772625,0.4979865,0.41498876,0.40367088,0.3961256,0.362172,0.29426476,0.3169005,0.29049212,0.241448,0.1961765,0.18863125,0.16222288,0.150905,0.17731337,0.25276586,0.36971724,0.35839936,0.39989826,0.44894236,0.49044126,0.5357128,0.633801,0.60362,0.47535074,0.331991,0.32821837,0.32067314,0.35839936,0.40367088,0.41498876,0.34330887,0.30935526,0.2565385,0.22258487,0.241448,0.35462674,0.32067314,0.33576363,0.38480774,0.44139713,0.45648763,0.46026024,0.5319401,0.6073926,0.66775465,0.7469798,0.7696155,0.7582976,0.7394345,0.7054809,0.60362,0.52062225,0.52062225,0.4979865,0.43007925,0.38480774,0.38858038,0.38858038,0.39989826,0.41876137,0.4074435,0.482896,0.5394854,0.5281675,0.47912338,0.5017591,0.59230214,0.55457586,0.452715,0.35085413,0.34330887,0.38858038,0.44516975,0.5017591,0.56589377,0.6488915,0.6187105,0.6451189,0.6790725,0.68661773,0.62625575,0.52062225,0.5319401,0.47912338,0.35462674,0.331991,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21881226,0.29426476,0.3734899,0.56212115,0.91674787,0.694163,1.1732863,2.033445,2.9049213,3.3576362,2.7691069,2.5880208,2.7879698,3.2520027,3.7537618,3.7047176,3.399135,3.180323,3.169005,3.2821836,1.9730829,1.4449154,1.9051756,2.71629,2.4107075,2.4107075,2.0447628,1.6712729,1.3355093,0.76207024,0.5319401,0.392353,0.35839936,0.362172,0.23013012,0.14335975,0.1056335,0.08677038,0.07922512,0.090543,0.018863125,0.056589376,0.09808825,0.08677038,0.0,0.0,0.0,0.0,0.018863125,0.090543,0.07922512,0.1056335,0.1056335,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.1659955,0.27540162,0.18863125,0.13958712,0.090543,0.041498873,0.0150905,0.05281675,0.392353,0.694163,0.935611,1.3732355,1.8599042,2.7615614,3.8405323,4.5120597,3.8292143,5.904158,7.7414265,8.7751255,8.865668,8.314865,9.4013815,9.646602,8.699674,7.2623034,7.0812173,7.8244243,8.771353,9.352338,9.435335,9.337247,9.740918,8.816625,7.3453007,5.956975,5.1269975,5.0175915,7.2887115,8.582722,8.89585,11.581959,14.694374,17.093763,16.957949,14.3095665,11.000975,11.5857315,13.317367,13.996439,12.1101265,6.8359966,15.211224,15.977067,17.30503,25.404858,44.50943,41.604507,43.011696,48.614044,56.879868,64.851425,56.012165,45.784576,40.891483,42.70989,47.274765,38.337414,34.108303,31.576872,28.192827,21.881226,22.028357,22.035902,21.805773,22.284895,25.484081,34.2743,40.67267,46.769234,57.31372,79.71557,99.77084,99.29172,86.642105,68.45051,49.591156,32.904835,22.115128,21.851044,31.678732,46.093933,47.802933,41.842182,34.77983,29.79242,26.657368,24.069347,20.243906,16.301512,13.04951,10.985884,13.219278,14.7321005,15.041456,13.9888935,11.717773,10.374719,9.940866,9.390063,8.888305,9.767326,10.70671,12.23085,16.31283,21.1267,21.03993,17.64834,14.347293,10.763299,7.816879,7.707473,12.808062,11.189606,8.401636,8.035691,11.732863,14.637785,14.66042,14.667966,16.33924,20.172226,29.732058,31.022295,32.42194,40.461403,59.848923,114.36713,142.01292,156.49603,163.36221,160.00458,136.56903,114.34072,102.815346,105.68632,120.81077,131.3779,114.26149,91.25603,75.75431,72.73998,47.81425,38.12992,36.077614,37.79793,43.166374,42.15531,35.78712,33.527317,36.07384,35.353268,30.788393,24.97855,20.225042,17.082445,14.358611,22.14531,25.46522,22.133991,16.252468,18.218006,21.19838,23.865625,33.150055,40.638718,22.598024,20.228815,22.156626,25.702894,27.860836,25.299223,23.443092,21.835953,20.07791,18.244415,16.874952,21.051247,30.003687,35.24009,33.146282,24.97855,20.915434,19.33093,16.686321,12.464753,9.156161,10.827434,13.2607765,14.535924,13.411682,9.322156,11.117926,10.578441,6.8171334,3.5123138,8.89585,13.875714,12.438345,12.623203,14.618922,10.789707,7.9941926,6.379509,4.9987283,4.666737,7.9489207,7.6923823,4.4441524,2.9237845,3.6745367,3.0520537,2.3805263,2.5238862,3.1954134,3.6066296,2.4710693,1.4713237,2.4823873,3.712263,4.327201,4.485651,3.1539145,2.071171,1.2864652,0.77338815,0.45648763,0.44516975,0.543258,0.67152727,0.7394345,0.6413463,0.482896,0.543258,0.55080324,0.43007925,0.32067314,0.392353,0.422534,0.9393836,1.9429018,2.867195,3.5651307,3.3463185,2.4522061,1.3317367,0.6111652,0.7696155,1.1846043,1.7693611,2.2258487,2.0296721,0.77338815,0.31312788,0.2565385,0.40367088,0.73188925,0.7432071,0.663982,0.6149379,0.7205714,1.0978339,0.7582976,0.44139713,0.27917424,0.36594462,0.7922512,0.56212115,0.6488915,0.76584285,0.7922512,0.7922512,0.7922512,0.84884065,0.7432071,0.47157812,0.23013012,0.39989826,0.35839936,0.3055826,0.27917424,0.1659955,0.13204187,0.13958712,0.150905,0.17354076,0.26031113,0.19994913,0.14713238,0.1358145,0.25276586,0.65643674,0.5696664,0.513077,0.41498876,0.2678564,0.120724,0.071679875,0.060362,0.060362,0.2565385,1.0374719,0.9393836,0.7582976,1.0714256,1.8938577,2.7011995,1.4071891,0.9922004,0.9016574,0.8563859,0.8563859,0.8186596,0.62625575,0.422534,0.31312788,0.35085413,0.46026024,0.38858038,0.41876137,0.5583485,0.5357128,0.39989826,0.33953625,0.32067314,0.3734899,0.58098423,0.32444575,0.22258487,0.15467763,0.0754525,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.0452715,0.00754525,0.018863125,0.02263575,0.011317875,0.0,0.011317875,0.041498873,0.041498873,0.011317875,0.0,0.011317875,0.1358145,0.20749438,0.16222288,0.0150905,0.0754525,0.090543,0.20749438,0.422534,0.58098423,0.38480774,0.26408374,0.18485862,0.12826926,0.090543,0.116951376,0.51684964,0.52062225,0.10940613,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.060362,0.09808825,0.09808825,0.12826926,0.19994913,0.26031113,0.29426476,0.24899325,0.18863125,0.13958712,0.090543,0.06790725,0.05281675,0.056589376,0.08677038,0.120724,0.120724,0.150905,0.18485862,0.211267,0.19994913,0.23390275,0.24522063,0.24899325,0.25276586,0.23013012,0.23013012,0.211267,0.18485862,0.18485862,0.24522063,0.3169005,0.34330887,0.38858038,0.47157812,0.58098423,0.5319401,0.44516975,0.42630664,0.5055317,0.6413463,0.5319401,0.35839936,0.26408374,0.32444575,0.52062225,0.7130261,0.7432071,0.76207024,0.8186596,0.8526133,0.80734175,0.63002837,0.48666862,0.39989826,0.23013012,0.23013012,0.24899325,0.28294688,0.35839936,0.5017591,0.6149379,0.5583485,0.44139713,0.35085413,0.35085413,0.27917424,0.24899325,0.2678564,0.31312788,0.33576363,0.3470815,0.3772625,0.44516975,0.5394854,0.62625575,0.724344,0.58475685,0.39989826,0.29049212,0.29049212,0.31312788,0.38480774,0.43385187,0.422534,0.33576363,0.31312788,0.3055826,0.36594462,0.4979865,0.65643674,0.58098423,0.5357128,0.482896,0.392353,0.26031113,0.271629,0.2565385,0.2263575,0.18863125,0.150905,0.1659955,0.150905,0.1358145,0.17354076,0.32067314,0.32067314,0.31312788,0.33576363,0.38858038,0.41121614,0.47157812,0.47157812,0.3772625,0.25276586,0.23013012,0.25276586,0.26031113,0.26408374,0.28294688,0.32067314,0.28294688,0.24899325,0.22258487,0.23013012,0.3055826,0.34330887,0.34330887,0.3470815,0.38103512,0.44139713,0.41876137,0.47535074,0.56212115,0.6488915,0.7469798,0.80734175,0.814887,0.77338815,0.7130261,0.70170826,0.6149379,0.5583485,0.52062225,0.49421388,0.45648763,0.43385187,0.38103512,0.34330887,0.34330887,0.38103512,0.36971724,0.3772625,0.39989826,0.4376245,0.48666862,0.40367088,0.41876137,0.38858038,0.3169005,0.36594462,0.5017591,0.46026024,0.38103512,0.34330887,0.38103512,0.36971724,0.422534,0.482896,0.55080324,0.68661773,0.6488915,0.5017591,0.38103512,0.331991,0.32067314,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.21881226,0.23390275,0.26031113,0.91674787,1.2411937,1.3807807,1.5279131,1.9127209,2.795515,2.9124665,2.3126192,1.9994912,2.4786146,3.731126,3.7763977,3.6141748,3.5424948,3.4029078,2.584248,1.8561316,1.8297231,2.1956677,2.5389767,2.3503454,2.5540671,2.033445,1.2638294,0.62248313,0.4074435,0.28294688,0.19240387,0.1659955,0.16222288,0.0452715,0.07922512,0.06790725,0.060362,0.071679875,0.1056335,0.07922512,0.0754525,0.07922512,0.06413463,0.0,0.0,0.0,0.02263575,0.06790725,0.1056335,0.071679875,0.09808825,0.09808825,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.13204187,0.19994913,0.1056335,0.06790725,0.056589376,0.05281675,0.08677038,0.15467763,0.36971724,0.7130261,1.3505998,2.6182017,3.078462,3.6254926,4.447925,5.515578,6.6020937,8.635539,10.106862,10.623712,10.216269,9.318384,7.8244243,7.01331,6.9265394,7.7414265,9.763554,10.246449,10.050273,10.355856,11.144334,11.193378,12.064855,13.140053,13.958713,13.389046,9.6201935,11.374464,16.25624,17.89356,15.648849,14.64533,20.568352,18.384,14.124708,11.827179,13.528633,14.11339,17.53516,21.681276,22.598024,14.50197,16.429781,18.018057,30.901571,51.669872,61.878593,41.925182,32.58039,32.55021,36.87364,36.934,33.331142,27.113855,23.314823,23.959942,28.045694,24.608833,22.662159,19.749691,15.611122,12.200669,14.78869,16.361876,16.0412,14.792462,15.411173,19.357338,25.344494,32.66716,43.441776,62.599167,83.63155,82.431854,69.48421,55.570766,51.737778,42.777794,30.84121,29.630198,43.37387,66.82073,73.24929,63.331055,49.361027,37.258446,26.585688,22.394302,24.242887,25.646305,23.94485,20.300495,15.452672,13.845533,15.158407,17.21826,16.003475,19.055529,17.814335,16.59955,15.358356,9.654147,11.046246,13.992666,16.52787,18.070873,19.429018,18.029375,15.328176,12.0724,9.574923,9.7069645,13.932304,11.378237,8.865668,10.072908,15.516807,22.571615,19.772327,15.897841,14.939595,16.109108,18.361366,22.258488,26.936543,32.991604,42.475986,68.46937,86.90619,102.04196,112.07337,109.11563,104.486626,96.76406,83.273155,71.11775,77.18036,88.51333,81.85087,71.24225,63.949768,60.44877,45.539356,40.608536,39.016487,38.34496,40.39727,40.985798,37.62439,35.28159,33.942307,28.592726,26.4876,25.665169,24.669195,21.534143,13.773854,15.878979,22.88097,24.09953,20.349539,23.95617,26.838455,26.683777,29.535881,33.338688,27.932516,25.46522,24.122164,24.857826,25.419947,20.368402,18.621677,18.334957,18.233097,17.82188,17.399347,19.097027,30.863846,36.5756,32.61057,27.872154,28.736084,25.699121,19.270569,12.691111,11.902632,8.009283,8.001738,11.18206,16.086473,20.492899,29.501928,21.896315,10.306811,4.195159,9.87296,11.348056,15.712983,17.463482,14.607604,8.677037,8.028146,7.1264887,5.5268955,4.4403796,6.7152724,10.446399,7.575431,4.1762958,3.029418,3.6368105,3.9348478,3.6292653,3.500996,3.3576362,2.0560806,1.4373702,1.5580941,1.8599042,2.173032,2.6936543,2.6106565,3.0709167,3.6594462,3.6783094,2.1315331,1.0148361,0.7205714,0.67152727,0.58475685,0.45648763,0.27917424,0.2263575,0.20749438,0.17354076,0.11317875,0.23390275,0.27540162,0.41876137,0.784706,1.4411428,2.3993895,2.795515,2.5427492,1.9542197,1.7316349,1.9202662,1.8297231,1.629774,1.5279131,1.7731338,0.995973,0.72811663,0.6073926,0.4979865,0.47535074,0.7696155,1.0638802,1.1204696,1.0148361,1.0978339,0.5319401,0.271629,0.1961765,0.23767537,0.40367088,0.35462674,0.543258,0.83752275,1.1016065,1.1581959,0.7582976,0.60362,0.49044126,0.36971724,0.33953625,0.5583485,0.5017591,0.44516975,0.43007925,0.25276586,0.17731337,0.1056335,0.056589376,0.0452715,0.06413463,0.13958712,0.23013012,0.21881226,0.20372175,0.4979865,0.5885295,0.47912338,0.33576363,0.23013012,0.1358145,0.33953625,0.271629,0.1358145,0.1358145,0.47535074,0.73188925,0.69039035,0.77716076,1.116697,1.5430037,1.1959221,0.88279426,0.7130261,0.6828451,0.6828451,0.52062225,0.362172,0.3772625,0.47912338,0.35085413,0.3734899,0.34330887,0.32444575,0.32067314,0.26408374,0.21881226,0.27540162,0.27540162,0.21503963,0.23767537,0.18863125,0.29049212,0.3169005,0.1961765,0.026408374,0.003772625,0.0,0.0,0.003772625,0.02263575,0.02263575,0.018863125,0.00754525,0.00754525,0.033953626,0.0150905,0.00754525,0.003772625,0.003772625,0.0,0.003772625,0.0150905,0.033953626,0.041498873,0.0,0.003772625,0.033953626,0.1358145,0.24522063,0.18485862,0.08299775,0.056589376,0.13204187,0.3772625,0.8978847,0.56589377,0.27540162,0.12826926,0.10940613,0.1056335,0.06790725,0.271629,0.28294688,0.08677038,0.071679875,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.011317875,0.03772625,0.0452715,0.0452715,0.06790725,0.12826926,0.19994913,0.23390275,0.2263575,0.20749438,0.181086,0.090543,0.049044125,0.041498873,0.049044125,0.060362,0.08677038,0.1056335,0.1358145,0.1659955,0.1659955,0.124496624,0.16222288,0.20749438,0.23767537,0.241448,0.21503963,0.1961765,0.1659955,0.14335975,0.13958712,0.16976812,0.2263575,0.29803738,0.3734899,0.44894236,0.52062225,0.6451189,0.52439487,0.4376245,0.52439487,0.77338815,0.6451189,0.44516975,0.32444575,0.36971724,0.60362,0.8186596,0.8903395,0.8903395,0.8224323,0.633801,0.5772116,0.573439,0.5885295,0.56589377,0.422534,0.29803738,0.25276586,0.3055826,0.46026024,0.73566186,0.7582976,0.68661773,0.58098423,0.47157812,0.362172,0.271629,0.26031113,0.271629,0.29426476,0.3470815,0.38103512,0.35462674,0.36594462,0.44139713,0.56589377,0.67152727,0.6149379,0.49044126,0.38103512,0.362172,0.30935526,0.35839936,0.41498876,0.44139713,0.49421388,0.34330887,0.27540162,0.29803738,0.40367088,0.5696664,0.59607476,0.51684964,0.422534,0.36594462,0.36971724,0.3734899,0.3169005,0.24899325,0.18863125,0.150905,0.14713238,0.13204187,0.120724,0.1358145,0.22258487,0.25276586,0.2565385,0.2678564,0.28294688,0.27917424,0.3772625,0.5017591,0.4979865,0.3734899,0.29049212,0.2867195,0.32821837,0.32821837,0.29049212,0.30935526,0.30181,0.26408374,0.24522063,0.26031113,0.3055826,0.38103512,0.35462674,0.32444575,0.35085413,0.43007925,0.42630664,0.47535074,0.52062225,0.5470306,0.5772116,0.7167987,0.7130261,0.6752999,0.663982,0.70170826,0.65643674,0.56212115,0.51684964,0.52439487,0.5055317,0.513077,0.5017591,0.47535074,0.44139713,0.41876137,0.45648763,0.45648763,0.44516975,0.44139713,0.5017591,0.49421388,0.44894236,0.4074435,0.38480774,0.36594462,0.452715,0.45648763,0.38858038,0.28294688,0.22258487,0.24899325,0.31312788,0.3961256,0.482896,0.5394854,0.7092535,0.7394345,0.6451189,0.4979865,0.41876137,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.0452715,0.0,0.10940613,0.513077,0.8526133,0.98465514,1.0072908,1.1431054,1.2713746,1.3166461,1.5656394,2.674791,3.2369123,2.1541688,1.448688,1.9730829,3.4217708,3.772625,4.0480266,4.1536603,3.9273026,3.1350515,2.8558772,2.2899833,1.9504471,1.9202662,1.8863125,1.7919968,1.2638294,0.7167987,0.36971724,0.24899325,0.11317875,0.056589376,0.049044125,0.0452715,0.0,0.02263575,0.02263575,0.02263575,0.026408374,0.041498873,0.03772625,0.033953626,0.049044125,0.06790725,0.03772625,0.0452715,0.018863125,0.0452715,0.10940613,0.08677038,0.03772625,0.06790725,0.06790725,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.13204187,0.17354076,0.14335975,0.06413463,0.0,0.03772625,0.07922512,0.08677038,0.0754525,0.090543,0.06790725,0.05281675,0.049044125,0.08299775,0.19994913,0.26408374,0.5055317,0.90920264,1.750498,3.6066296,4.0291634,4.6818275,5.4212623,6.507778,8.575176,9.691874,10.34831,10.265312,9.469289,8.27714,7.8017883,7.677292,8.114917,9.420244,11.966766,12.272349,12.811834,14.196388,15.577168,14.652876,17.338985,20.89657,24.020304,24.714466,20.289177,18.116146,23.416683,31.31656,40.68776,54.144714,56.49506,37.315033,21.334194,18.059555,21.741638,20.157135,29.117119,39.827602,45.939255,43.55118,34.511974,25.344494,35.519264,58.33233,60.90526,39.774784,29.47552,29.056757,31.41842,23.29596,19.595015,16.143063,13.6682205,12.925014,14.690601,15.196134,14.286931,11.77059,8.624221,6.9793563,9.978593,12.174261,12.310076,10.79348,9.661693,11.729091,17.84829,25.1785,33.1991,43.71718,55.152004,53.005383,45.85626,42.332626,51.115295,49.45157,36.04366,29.96596,37.514984,52.22445,58.728455,58.419098,53.288326,43.524776,27.498663,18.765038,19.73083,22.673477,24.250433,25.514263,20.455173,16.625957,15.015047,14.966003,14.143571,18.663176,21.209698,21.926497,20.198635,14.671739,18.297232,19.640285,20.26277,19.94964,16.720274,18.931032,17.618158,15.169725,12.755245,10.336992,12.97783,12.340257,10.355856,10.465261,17.637022,27.95515,23.4695,15.99593,11.849815,11.823407,13.196642,16.708956,21.085201,26.20088,33.104786,45.47145,55.61604,64.5383,70.55186,69.2918,76.05989,89.05659,86.23089,71.246025,73.48319,82.09232,76.55033,70.49905,68.31092,65.07024,54.046627,51.36429,49.3233,45.392223,42.204357,42.751385,44.060486,45.19982,42.906063,31.542917,25.982069,23.273323,21.941587,19.794964,13.936077,18.09351,18.334957,17.73511,19.787418,28.411638,32.73884,28.211689,26.744139,30.365858,31.214699,25.027594,22.567842,23.993895,24.884235,16.252468,16.946632,17.96524,17.991648,17.482344,18.678267,23.84299,32.199356,35.809757,33.338688,30.048958,30.090458,30.614851,27.053493,20.36463,17.029629,11.00852,7.183078,8.258276,14.584969,24.156118,23.888262,17.074902,9.061845,4.146115,5.5759397,10.186088,19.960958,19.206434,9.258021,8.477088,8.469543,6.6247296,4.779916,3.9159849,4.1574326,9.7069645,8.246958,4.7421894,2.7125173,4.214022,5.409944,4.859141,4.0291634,3.3953626,2.4107075,2.0108092,1.6184561,1.3053282,1.3204187,2.1051247,2.7841973,2.9992368,3.5085413,3.9273026,2.7238352,1.5354583,1.0223814,0.76207024,0.52439487,0.27540162,0.181086,0.150905,0.13204187,0.094315626,0.060362,0.14335975,0.2565385,0.2867195,0.331991,0.69793564,1.6222287,2.3201644,2.4031622,2.071171,2.1315331,2.4182527,1.9202662,1.3053282,1.0374719,1.3694628,1.3128735,1.2261031,1.0148361,0.69793564,0.41121614,0.77716076,1.1506506,1.2298758,1.0450171,0.9695646,0.5093044,0.241448,0.19240387,0.28294688,0.32444575,0.23390275,0.31312788,0.69793564,1.1619685,1.1317875,1.0940613,0.98465514,0.87147635,0.76584285,0.6149379,0.5885295,0.5357128,0.56589377,0.6488915,0.6149379,0.35085413,0.18485862,0.08299775,0.033953626,0.041498873,0.124496624,0.18485862,0.16222288,0.11317875,0.23013012,0.32821837,0.271629,0.181086,0.116951376,0.090543,0.30181,0.34330887,0.24522063,0.10940613,0.14335975,0.4640329,0.6828451,0.76584285,0.8186596,1.0940613,1.2713746,1.1016065,0.875249,0.7884786,0.935611,0.73188925,0.392353,0.29426476,0.40367088,0.2678564,0.33576363,0.331991,0.30935526,0.2678564,0.16976812,0.124496624,0.14335975,0.15845025,0.15467763,0.181086,0.08299775,0.13958712,0.16976812,0.11317875,0.02263575,0.018863125,0.00754525,0.0,0.00754525,0.030181,0.13204187,0.08299775,0.018863125,0.003772625,0.011317875,0.02263575,0.0150905,0.003772625,0.0,0.00754525,0.0,0.018863125,0.0452715,0.049044125,0.00754525,0.0,0.003772625,0.08299775,0.20749438,0.23013012,0.15467763,0.08299775,0.094315626,0.29426476,0.7922512,0.5281675,0.27917424,0.14335975,0.10940613,0.07922512,0.05281675,0.150905,0.20749438,0.25276586,0.513077,0.271629,0.08299775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.003772625,0.02263575,0.030181,0.041498873,0.06413463,0.09808825,0.12826926,0.19994913,0.24899325,0.26031113,0.22258487,0.120724,0.06413463,0.0452715,0.03772625,0.033953626,0.056589376,0.08299775,0.1056335,0.124496624,0.1358145,0.116951376,0.13958712,0.16222288,0.1961765,0.22258487,0.20372175,0.15845025,0.12826926,0.116951376,0.116951376,0.124496624,0.150905,0.19240387,0.25276586,0.32067314,0.3772625,0.5319401,0.4640329,0.38858038,0.4376245,0.6451189,0.52439487,0.38480774,0.32067314,0.38103512,0.5885295,0.8601585,0.90543,0.84129536,0.7469798,0.67152727,0.5281675,0.5017591,0.5281675,0.5772116,0.6111652,0.362172,0.27917424,0.31312788,0.44139713,0.663982,0.6375736,0.5885295,0.55080324,0.5093044,0.40367088,0.31312788,0.32444575,0.35839936,0.3734899,0.35839936,0.41876137,0.43007925,0.42630664,0.43385187,0.5017591,0.5319401,0.49421388,0.44894236,0.4376245,0.47157812,0.44516975,0.452715,0.44894236,0.43007925,0.43385187,0.30181,0.25276586,0.2565385,0.29049212,0.36594462,0.51684964,0.543258,0.52439487,0.5055317,0.5055317,0.38858038,0.2867195,0.21881226,0.1961765,0.181086,0.1659955,0.13958712,0.116951376,0.116951376,0.16222288,0.18485862,0.2263575,0.26031113,0.26408374,0.25276586,0.29803738,0.40367088,0.4640329,0.44139713,0.35839936,0.29803738,0.30935526,0.32067314,0.30935526,0.31312788,0.32821837,0.33576363,0.35462674,0.38480774,0.4074435,0.40367088,0.35462674,0.331991,0.36971724,0.45648763,0.47535074,0.482896,0.52062225,0.56212115,0.5055317,0.5772116,0.66020936,0.67152727,0.6111652,0.573439,0.6526641,0.7092535,0.69039035,0.5998474,0.5017591,0.5055317,0.58475685,0.58098423,0.52062225,0.6111652,0.5696664,0.5357128,0.49421388,0.46026024,0.48666862,0.47535074,0.41876137,0.3734899,0.3470815,0.31312788,0.36971724,0.41876137,0.39989826,0.31312788,0.18485862,0.18485862,0.22258487,0.27917424,0.34330887,0.40367088,0.55080324,0.6111652,0.62625575,0.63002837,0.6451189,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041498873,0.090543,0.041498873,0.27540162,1.1280149,1.9051756,2.0636258,1.2336484,1.2411937,1.3920987,1.5241405,1.7769064,2.5993385,3.5990841,2.3163917,1.3015556,1.6524098,3.006782,3.62172,4.432834,4.9534564,4.878004,4.074435,3.4444065,2.2107582,1.418507,1.3015556,1.2525115,0.87902164,0.5093044,0.3055826,0.241448,0.120724,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.049044125,0.060362,0.06790725,0.049044125,0.06413463,0.10186087,0.0754525,0.0150905,0.026408374,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14335975,0.2263575,0.20749438,0.1056335,0.0,0.060362,0.116951376,0.13958712,0.11317875,0.03772625,0.0452715,0.0452715,0.1056335,0.24899325,0.46026024,0.79602385,1.6788181,2.493705,3.2029586,4.3649273,5.3269467,7.4094353,8.639311,9.114662,11.012292,11.936585,11.019837,9.971047,9.378746,8.692128,8.99771,9.0957985,9.020347,9.733373,13.094781,15.739391,17.803017,20.50799,24.925734,32.00695,38.405323,37.29617,36.36056,37.2094,35.360813,34.413887,40.88771,50.311726,61.35797,75.87503,75.51286,50.191,33.2406,34.31957,39.386204,37.696068,44.445293,51.775505,56.487514,60.03001,43.479504,28.060785,29.928234,44.528294,46.603237,32.044678,24.510744,23.94485,24.627695,15.173498,11.84227,10.933067,9.808825,8.080963,7.6207023,9.552286,8.801534,6.617184,4.6290107,4.8440504,8.0206,10.431308,10.3634,8.280911,6.8171334,10.438853,16.052519,21.077656,24.914415,28.928488,32.569073,31.342968,29.358568,31.565554,43.739815,45.554447,32.49739,25.427492,30.429993,38.81654,40.71417,46.63342,49.02526,43.14751,27.061039,22.08872,24.427748,24.37493,21.002203,22.156626,23.1526,21.719002,18.689585,15.23386,12.857106,16.229834,20.06282,21.571869,20.285404,18.03692,22.111355,23.480818,24.178753,22.95265,15.279131,17.48989,18.135008,17.969013,16.724047,13.087236,12.306303,12.781653,11.649866,10.457717,15.165953,24.133482,19.640285,12.464753,8.635539,9.424017,10.265312,12.992921,15.799753,18.957441,24.812555,31.154337,36.726505,41.50642,45.663853,49.576065,62.335083,78.68187,79.772156,67.97893,66.91128,78.014114,80.68513,81.44343,81.40193,76.29757,69.32953,66.19825,60.603447,52.035816,45.784576,44.90933,46.339153,48.30469,47.78784,40.52554,30.445084,21.817091,16.595778,14.264296,11.827179,15.912932,13.3626375,12.645839,18.040693,29.66415,32.716206,26.966724,24.340977,27.657114,30.618624,23.431774,20.98334,22.511253,23.401592,15.150862,17.278622,18.402864,18.516043,19.176252,23.473272,30.199863,35.52681,37.2509,35.97198,35.092957,33.855537,37.23581,35.579628,27.891016,21.87368,16.437326,8.892077,6.4926877,11.02361,18.810308,13.660675,10.955703,8.246958,5.4967146,5.0854983,12.095036,18.191597,14.818871,6.156924,9.107117,8.341274,7.1868505,7.0246277,7.0472636,4.247976,8.273367,8.567632,5.987156,3.0030096,3.7386713,6.609639,6.4134626,5.194905,3.8103511,1.9164935,1.8863125,1.569412,1.2034674,1.2600567,2.4371157,2.776652,2.2748928,2.1353056,2.3956168,1.9353566,1.3091009,0.95824677,0.663982,0.35839936,0.12826926,0.1358145,0.20372175,0.27540162,0.30935526,0.27917424,0.29426476,0.4074435,0.44894236,0.43385187,0.5772116,1.3920987,2.3465726,2.535204,2.0183544,1.8221779,2.0108092,1.4939595,0.98465514,0.84129536,1.0450171,1.5656394,1.6448646,1.4449154,1.1280149,0.8526133,0.8563859,0.8941121,0.8526133,0.7469798,0.7130261,0.58475685,0.3169005,0.23767537,0.41121614,0.6451189,0.27540162,0.21881226,0.5470306,1.0299267,1.1016065,1.4109617,1.4147344,1.2600567,1.0789708,0.9808825,0.7922512,0.7394345,0.7469798,0.79602385,0.91674787,0.6752999,0.4376245,0.241448,0.1056335,0.056589376,0.10940613,0.13204187,0.11317875,0.0754525,0.05281675,0.094315626,0.09808825,0.071679875,0.03772625,0.03772625,0.241448,0.30935526,0.25276586,0.12826926,0.0452715,0.24899325,0.6187105,0.8224323,0.8903395,1.2185578,1.3656902,1.4147344,1.2562841,1.1053791,1.5203679,1.0676528,0.5093044,0.24522063,0.2678564,0.18485862,0.26031113,0.32821837,0.35839936,0.33953625,0.2867195,0.181086,0.11317875,0.120724,0.18863125,0.26031113,0.0754525,0.030181,0.030181,0.030181,0.0150905,0.02263575,0.011317875,0.0,0.003772625,0.018863125,0.1659955,0.17731337,0.09808825,0.003772625,0.0,0.018863125,0.02263575,0.018863125,0.011317875,0.0150905,0.00754525,0.049044125,0.06413463,0.03772625,0.00754525,0.0,0.0,0.03772625,0.10186087,0.150905,0.24899325,0.26408374,0.24899325,0.3169005,0.6413463,0.45648763,0.27540162,0.1659955,0.116951376,0.06790725,0.09808825,0.13204187,0.15845025,0.241448,0.49421388,0.27540162,0.1056335,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.033953626,0.049044125,0.06413463,0.0754525,0.07922512,0.15845025,0.23013012,0.2678564,0.25276586,0.1659955,0.10186087,0.060362,0.033953626,0.026408374,0.06413463,0.0754525,0.08299775,0.10186087,0.120724,0.120724,0.124496624,0.116951376,0.14713238,0.1961765,0.19240387,0.120724,0.090543,0.08299775,0.08677038,0.08677038,0.094315626,0.10940613,0.14713238,0.19994913,0.25276586,0.35462674,0.35839936,0.331991,0.3470815,0.47157812,0.47157812,0.39989826,0.331991,0.33953625,0.48666862,0.8111144,0.84129536,0.76207024,0.7054809,0.76207024,0.5772116,0.48666862,0.46026024,0.482896,0.55457586,0.35839936,0.30181,0.3470815,0.44894236,0.58098423,1.2638294,0.8563859,0.5017591,0.5319401,0.482896,0.3734899,0.36594462,0.3961256,0.41121614,0.3772625,0.44139713,0.58098423,0.6187105,0.5583485,0.5885295,0.52439487,0.4640329,0.44516975,0.4640329,0.47912338,0.49421388,0.49044126,0.46026024,0.422534,0.40367088,0.30935526,0.2565385,0.23767537,0.241448,0.26408374,0.422534,0.58098423,0.6526641,0.6413463,0.6149379,0.44894236,0.3055826,0.241448,0.24899325,0.25276586,0.211267,0.15845025,0.120724,0.116951376,0.13204187,0.14335975,0.19994913,0.24522063,0.2565385,0.25276586,0.2678564,0.30181,0.35462674,0.39989826,0.3734899,0.29049212,0.27540162,0.29426476,0.32067314,0.32067314,0.36971724,0.3961256,0.43007925,0.4678055,0.5017591,0.47535074,0.4678055,0.4640329,0.4678055,0.48666862,0.5055317,0.48666862,0.5017591,0.5394854,0.47157812,0.422534,0.513077,0.58098423,0.56212115,0.47535074,0.56589377,0.694163,0.694163,0.5696664,0.5017591,0.5357128,0.62248313,0.663982,0.66775465,0.7582976,0.6828451,0.6073926,0.52062225,0.46026024,0.47157812,0.47157812,0.45648763,0.392353,0.3169005,0.32444575,0.38103512,0.38103512,0.38480774,0.3734899,0.26408374,0.16976812,0.181086,0.2263575,0.271629,0.34330887,0.4678055,0.5281675,0.58475685,0.663982,0.72811663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.094315626,0.08677038,0.42630664,1.6637276,2.7351532,2.9086938,1.7919968,2.2560298,2.1881225,2.1202152,2.3314822,2.8521044,4.0103,2.8596497,1.6109109,1.4675511,2.6332922,3.4972234,4.7572803,5.7796617,6.0550632,5.1835866,3.6783094,2.022127,1.0978339,0.9318384,0.67152727,0.26031113,0.11317875,0.10186087,0.09808825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.049044125,0.049044125,0.0754525,0.0754525,0.056589376,0.08677038,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.1056335,0.12826926,0.07922512,0.00754525,0.06413463,0.090543,0.14713238,0.18863125,0.05281675,0.0452715,0.11317875,0.38480774,0.8601585,1.4147344,2.3201644,3.8367596,5.0666356,5.802297,6.537959,8.126234,11.16697,12.713746,12.823153,14.539697,15.064092,13.174006,13.230596,15.173498,14.498198,11.98563,10.7557535,9.695646,9.948412,14.913187,22.945105,26.540417,29.939552,38.23178,57.336353,65.48145,54.831333,46.188248,47.531303,53.99381,59.426388,63.40651,64.91556,64.855194,66.036026,65.572,48.357506,41.630917,50.477722,57.834343,57.690983,53.454323,49.142212,48.357506,54.261665,37.69984,26.034885,22.043447,24.586197,28.581408,21.398329,17.40689,15.984612,14.588741,8.782671,8.311093,9.997457,9.7296,7.0585814,5.198677,6.900131,6.096562,4.044254,2.8709676,5.5457587,8.254503,9.948412,8.9788475,6.515323,6.530414,12.826925,16.765545,17.886015,17.667202,19.553514,21.900087,23.258234,23.793945,25.382221,31.59196,33.14251,23.235598,20.296722,28.385231,37.17922,32.157856,36.066296,39.144756,35.673943,24.005213,27.498663,33.391502,29.5472,17.946377,14.68683,23.92976,26.763002,24.208935,18.866898,14.928277,13.864397,15.331948,16.51278,17.025856,18.938578,20.790936,24.091984,27.310032,27.24967,19.074392,17.659658,18.776354,20.258997,20.353312,17.73511,12.1101265,11.427281,11.268831,10.167224,9.623966,12.974057,9.918231,6.63982,6.175787,8.409182,7.8696957,10.518079,12.525115,13.505998,16.535416,19.655376,23.820354,28.464457,34.787376,45.739307,63.13488,69.2918,64.957054,54.820015,47.508667,61.158024,76.595604,88.66801,94.90793,95.5455,98.24293,90.01861,75.32046,60.13187,51.983,47.323807,44.50943,43.622864,44.464157,46.531555,34.655334,21.345512,12.238396,8.782671,8.231868,8.718536,9.782416,12.079946,17.006994,26.691322,26.47251,23.114874,21.58696,23.360094,26.408375,22.782883,20.938068,21.307787,21.511507,16.376965,18.546225,19.413929,20.051502,22.711203,30.844982,36.341698,40.8198,41.687508,40.25391,41.740322,41.657326,44.837646,41.744095,31.742867,23.126192,19.538425,10.570895,6.0776987,8.096053,10.808571,9.695646,11.038701,10.9594755,9.035437,8.307321,13.004238,10.925522,9.027891,9.986138,12.219532,8.156415,8.409182,11.498961,13.45318,7.7829256,7.3981175,8.66572,7.2924843,3.62172,2.637065,6.881268,7.586749,6.579458,4.5799665,1.1996948,1.237421,1.3128735,1.237421,1.358145,2.5880208,2.161714,1.4675511,0.8526133,0.5319401,0.55457586,0.5093044,0.513077,0.3772625,0.14335975,0.0754525,0.124496624,0.29426476,0.55457586,0.76207024,0.694163,0.6413463,0.6752999,0.8111144,0.97710985,1.0110635,1.6410918,2.71629,2.886058,2.0145817,1.1921495,1.1242423,0.8903395,0.80734175,0.9242931,1.0450171,1.6637276,1.8033148,1.7240896,1.6335466,1.6675003,1.2223305,0.7884786,0.5319401,0.4640329,0.47157812,0.73188925,0.49044126,0.32067314,0.49421388,0.9808825,0.392353,0.26031113,0.47157812,0.8337501,1.0940613,1.5241405,1.6335466,1.478869,1.2713746,1.3845534,1.0751982,0.97710985,0.86770374,0.754525,0.8941121,0.8639311,0.62248313,0.35462674,0.15845025,0.041498873,0.07922512,0.11317875,0.120724,0.094315626,0.011317875,0.0150905,0.030181,0.049044125,0.05281675,0.0,0.20749438,0.19240387,0.15467763,0.15467763,0.08299775,0.124496624,0.44894236,0.7432071,0.9695646,1.3656902,1.3053282,1.5467763,1.50905,1.358145,1.9730829,1.2940104,0.6187105,0.26031113,0.20749438,0.14713238,0.150905,0.2867195,0.38858038,0.41121614,0.44139713,0.29049212,0.16976812,0.15467763,0.23390275,0.3055826,0.120724,0.030181,0.003772625,0.011317875,0.0150905,0.0150905,0.00754525,0.003772625,0.003772625,0.0,0.10186087,0.2565385,0.22258487,0.03772625,0.00754525,0.011317875,0.02263575,0.026408374,0.02263575,0.011317875,0.011317875,0.06413463,0.06790725,0.0150905,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.26031113,0.4640329,0.5055317,0.45648763,0.5885295,0.39989826,0.24899325,0.15845025,0.11317875,0.07922512,0.16976812,0.150905,0.09808825,0.05281675,0.041498873,0.030181,0.041498873,0.030181,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.033953626,0.041498873,0.0452715,0.0452715,0.056589376,0.1056335,0.150905,0.20749438,0.24899325,0.21503963,0.14335975,0.07922512,0.03772625,0.030181,0.07922512,0.06790725,0.06790725,0.08677038,0.11317875,0.116951376,0.1056335,0.08299775,0.1056335,0.15845025,0.17354076,0.094315626,0.056589376,0.0452715,0.05281675,0.056589376,0.056589376,0.071679875,0.09808825,0.124496624,0.17731337,0.21503963,0.26031113,0.27917424,0.28294688,0.34330887,0.48666862,0.4640329,0.3734899,0.31312788,0.39989826,0.694163,0.72811663,0.7205714,0.754525,0.7884786,0.67152727,0.5470306,0.43385187,0.35085413,0.32444575,0.30181,0.32067314,0.392353,0.49044126,0.55080324,1.9693103,1.1883769,0.47535074,0.55457586,0.60362,0.44894236,0.3961256,0.4074435,0.44516975,0.44894236,0.47912338,0.70170826,0.77716076,0.68661773,0.72811663,0.6187105,0.5470306,0.52439487,0.51684964,0.49044126,0.49044126,0.47912338,0.46026024,0.452715,0.4640329,0.392353,0.29803738,0.2565385,0.27540162,0.30935526,0.392353,0.6187105,0.7432071,0.7130261,0.68661773,0.55457586,0.392353,0.3169005,0.32821837,0.31312788,0.23767537,0.17731337,0.150905,0.14713238,0.1358145,0.13204187,0.1659955,0.211267,0.23767537,0.24522063,0.27917424,0.2565385,0.25276586,0.29426476,0.34330887,0.2867195,0.271629,0.29426476,0.32067314,0.32821837,0.40367088,0.422534,0.4376245,0.47912338,0.5583485,0.58098423,0.633801,0.6413463,0.5885295,0.513077,0.5093044,0.49421388,0.48666862,0.47912338,0.45648763,0.33953625,0.3470815,0.42630664,0.4979865,0.4376245,0.44139713,0.5319401,0.5357128,0.4678055,0.5357128,0.6375736,0.6790725,0.7507524,0.8337501,0.784706,0.7922512,0.70170826,0.573439,0.49421388,0.56212115,0.5470306,0.543258,0.45648763,0.3470815,0.392353,0.45648763,0.36594462,0.33576363,0.3961256,0.3734899,0.20749438,0.20749438,0.24522063,0.27917424,0.33953625,0.5017591,0.573439,0.60362,0.633801,0.66020936,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.47535074,1.3807807,2.3465726,3.0105548,3.0369632,4.768598,3.99521,2.927557,2.897376,4.3649273,4.644101,3.7084904,2.2975287,1.4373702,2.425798,3.8178966,5.27413,6.3832817,6.9265394,6.8661776,5.2062225,3.218049,1.7089992,0.8903395,0.36594462,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.056589376,0.02263575,0.120724,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.071679875,0.06790725,0.06790725,0.0754525,0.0754525,0.08677038,0.40367088,1.1732863,2.4182527,4.0291634,5.564622,6.006019,6.609639,8.650629,13.411682,14.120935,13.151371,13.011784,14.988639,19.164934,15.599804,16.376965,24.774828,34.576107,30.075367,18.233097,14.18507,13.502225,15.158407,21.53037,36.639732,41.280064,44.14726,51.36806,66.46611,66.137886,53.2921,45.090412,51.700054,76.30888,82.33754,68.31092,53.756134,48.214146,51.23979,49.5572,38.212917,35.436268,44.96969,56.076298,54.088123,39.646515,31.844728,35.45136,40.895256,31.859818,28.898308,28.977533,28.041922,21.013521,16.301512,16.825907,16.927769,13.373956,5.342037,8.439363,12.310076,11.5857315,6.6624556,3.7084904,6.221059,6.1078796,4.6026025,4.459243,9.963503,8.963757,7.375482,5.9532022,6.0286546,9.522105,14.539697,15.754482,13.853079,11.302785,12.37421,16.939087,20.070366,23.163918,25.170954,22.582933,23.695858,19.549744,20.557034,27.574116,31.90509,22.469755,23.378958,26.32915,25.616123,18.157644,16.32792,19.002712,18.776354,15.543215,16.493916,28.626678,28.373913,23.552498,19.53088,19.225298,8.729855,9.016574,12.498707,16.361876,22.552752,21.319103,24.325886,31.052477,36.99436,33.65936,30.203636,26.438557,23.688313,22.03213,20.30804,10.397354,7.039718,7.462252,8.571404,6.971811,4.8742313,3.6707642,3.6896272,4.6516466,5.6778007,6.579458,9.488152,13.200415,15.482853,13.091009,13.456953,15.490398,18.938578,25.793438,40.28409,67.050865,80.7304,75.85995,56.89496,38.209145,35.390995,46.6221,68.95227,99.601074,135.99936,158.51816,136.83311,104.78843,80.289,65.27773,52.277264,47.406807,44.20762,39.86533,35.202362,27.000677,17.953922,11.506506,8.624221,7.7829256,8.160188,9.673011,12.932558,16.999449,19.379974,19.598787,18.444365,17.40312,17.829426,20.964478,22.760246,22.100037,22.767792,23.163918,16.32792,19.757236,22.865881,23.89958,25.78212,36.1342,43.736042,46.508923,46.373108,45.022507,43.898266,47.878384,48.772495,43.77377,32.46344,16.81459,14.203933,9.009028,6.677546,9.050528,14.373701,14.373701,17.45971,18.233097,14.237886,5.9494295,3.0709167,6.2323766,14.335975,22.53389,22.21699,9.910686,7.164215,12.419481,18.451908,12.37421,6.820906,6.6586833,6.0739264,3.7348988,2.806833,5.138315,6.7567716,6.9454026,5.5797124,3.127506,1.7014539,1.7655885,1.5920477,0.86770374,0.67152727,0.97710985,1.3015556,0.9997456,0.33576363,0.45648763,0.17731337,0.14335975,0.181086,0.19994913,0.19994913,0.1358145,0.3772625,0.83752275,1.2185578,1.0223814,0.91297525,0.9016574,1.2940104,1.8749946,1.9391292,2.071171,2.7011995,2.8294687,2.1466236,1.0223814,0.814887,0.754525,0.87147635,1.1695137,1.6335466,1.5958204,1.5052774,1.5279131,1.780679,2.305074,2.2183034,1.8749946,1.4373702,0.98465514,0.5357128,0.9997456,0.7922512,0.482896,0.35839936,0.44139713,0.331991,0.20372175,0.39989826,0.7884786,0.76207024,1.4600059,1.7165444,1.81086,1.8599042,1.7995421,0.935611,0.69039035,0.573439,0.4074435,0.32067314,0.30935526,0.20372175,0.094315626,0.030181,0.030181,0.018863125,0.060362,0.10940613,0.10940613,0.0,0.011317875,0.0150905,0.094315626,0.16976812,0.0,0.011317875,0.00754525,0.071679875,0.15467763,0.0452715,0.071679875,0.20372175,0.331991,0.4376245,0.59607476,1.0336993,1.1732863,1.0940613,1.0450171,1.448688,1.3166461,0.7432071,0.35839936,0.29426476,0.18485862,0.10940613,0.14713238,0.23013012,0.29426476,0.26031113,0.18485862,0.120724,0.09808825,0.10940613,0.120724,0.08677038,0.030181,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.02263575,0.02263575,0.0,0.060362,0.24899325,0.2867195,0.13958712,0.030181,0.00754525,0.00754525,0.0150905,0.011317875,0.0,0.0,0.00754525,0.02263575,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.32444575,0.52439487,0.5772116,0.56589377,0.30935526,0.16222288,0.08677038,0.06790725,0.090543,0.150905,0.1056335,0.056589376,0.041498873,0.0150905,0.0150905,0.0150905,0.00754525,0.011317875,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.041498873,0.030181,0.030181,0.090543,0.08677038,0.120724,0.19240387,0.23013012,0.15467763,0.090543,0.049044125,0.030181,0.030181,0.030181,0.041498873,0.056589376,0.07922512,0.090543,0.07922512,0.056589376,0.071679875,0.11317875,0.1358145,0.08677038,0.049044125,0.02263575,0.018863125,0.030181,0.030181,0.049044125,0.06790725,0.07922512,0.090543,0.12826926,0.17354076,0.19240387,0.18485862,0.18485862,0.27917424,0.331991,0.38103512,0.44894236,0.5357128,0.59607476,0.59230214,0.7130261,0.87147635,0.70170826,0.8111144,0.6451189,0.41498876,0.26408374,0.27540162,0.31312788,0.33953625,0.38103512,0.43007925,0.44139713,0.4074435,0.38858038,0.41121614,0.52062225,0.76207024,0.58098423,0.52439487,0.59230214,0.694163,0.65643674,0.6187105,0.6111652,0.573439,0.5357128,0.59607476,0.52062225,0.52062225,0.5885295,0.7092535,0.87147635,0.724344,0.58475685,0.52439487,0.52439487,0.48666862,0.4640329,0.3734899,0.33953625,0.36971724,0.38103512,0.51684964,0.694163,0.7922512,0.784706,0.7469798,0.5772116,0.44139713,0.38103512,0.35085413,0.23013012,0.19240387,0.19240387,0.22258487,0.24522063,0.18485862,0.120724,0.14335975,0.211267,0.2678564,0.24522063,0.2678564,0.26408374,0.25276586,0.2678564,0.36594462,0.32821837,0.32821837,0.32821837,0.32821837,0.36594462,0.40367088,0.40367088,0.42630664,0.4979865,0.59607476,0.6073926,0.59230214,0.58475685,0.58475685,0.55080324,0.52439487,0.573439,0.58098423,0.5319401,0.52062225,0.47157812,0.44894236,0.41121614,0.362172,0.35085413,0.422534,0.55080324,0.5696664,0.5093044,0.59607476,0.77716076,0.8601585,0.87902164,0.845068,0.7469798,0.9318384,0.875249,0.7582976,0.73188925,0.91674787,0.694163,0.52062225,0.44894236,0.44139713,0.38103512,0.392353,0.35085413,0.30935526,0.30181,0.35085413,0.30181,0.29803738,0.27540162,0.241448,0.29049212,0.422534,0.49421388,0.58475685,0.6828451,0.67152727,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08299775,0.41498876,1.3807807,2.2183034,2.8219235,3.7462165,6.2097406,7.3679366,5.8626595,4.564876,4.7874613,6.2814207,6.4436436,5.383536,4.142342,3.5424948,4.1612053,4.798779,5.0138187,4.991183,4.851596,4.6327834,3.3840446,1.9429018,0.8941121,0.39989826,0.20749438,0.041498873,0.06413463,0.06413463,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.003772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.094315626,0.049044125,0.030181,0.030181,0.06790725,0.18485862,0.5319401,1.6675003,2.9351022,4.5422406,7.5792036,12.038446,15.9695215,25.917934,41.472466,55.253864,44.25289,32.101265,25.65385,24.997414,23.401592,18.576405,32.33517,63.961082,91.244705,70.51414,33.236828,20.534397,19.153618,23.933533,37.81302,68.45051,76.56165,66.84337,52.53003,55.397224,52.137676,42.38544,36.65105,40.42745,54.16735,53.63541,38.54491,24.872917,21.941587,32.429485,36.36056,31.041159,28.109829,32.154083,40.733032,37.228264,26.461191,26.570599,36.243607,34.704376,30.290405,23.72981,18.214233,14.981093,13.309821,10.785934,12.245941,14.483108,13.475817,4.3875628,5.05909,7.0510364,6.8925858,4.478106,3.0860074,5.3571277,4.9760923,4.7044635,6.7643166,12.845788,10.250222,6.6322746,4.5233774,5.481624,10.095545,11.1782875,9.725827,7.54525,6.4436436,8.2507305,11.819634,13.890805,15.897841,17.64834,17.346529,20.311813,17.89356,18.346275,22.337713,22.911152,18.414183,18.693357,20.330677,19.915688,14.019074,11.231105,12.034674,15.55076,23.38273,39.574837,67.37154,52.296127,31.93527,25.012505,31.34674,11.355601,7.277394,10.499215,16.060064,22.65084,23.526089,22.820608,25.665169,31.399557,33.565044,37.677204,33.606544,28.1966,24.963459,24.080666,15.886524,11.672502,8.68081,6.156924,5.349582,4.7233267,3.5387223,2.8294687,3.150142,4.5761943,5.9796104,8.929804,13.607859,17.516298,15.482853,14.543469,15.494171,23.103556,42.35903,78.47437,97.462,92.410446,76.39565,60.022465,51.402016,43.51346,51.285065,75.154465,119.52431,192.74718,214.79063,186.52989,149.3205,118.71319,84.45398,56.679916,46.531555,41.62337,35.805984,29.17371,23.16769,17.923742,15.165953,14.332202,12.543978,10.050273,9.748463,16.565596,24.042938,14.324657,18.316093,17.37671,16.286423,17.293713,20.14959,21.78691,23.737356,22.299986,17.342756,12.325166,19.081938,25.419947,28.1966,27.898561,28.664404,34.187527,35.65508,35.032597,34.489338,36.394512,40.725487,49.006397,47.689754,34.040394,16.15438,10.672756,9.446653,14.25675,19.549744,12.483616,14.260523,18.761265,20.1345,16.056292,7.7678347,3.2482302,3.832987,10.159679,18.089737,18.700903,12.166716,9.495697,13.215506,18.878216,15.033911,6.1795597,6.270103,7.858378,8.265821,9.593785,7.492433,7.3415284,6.3644185,4.2102494,2.957738,1.9957186,1.3958713,1.0940613,0.995973,0.97710985,1.0676528,0.95447415,0.67152727,0.38858038,0.43385187,0.241448,0.15467763,0.1961765,0.34330887,0.5281675,0.52439487,0.5093044,0.7205714,1.0072908,0.8526133,0.7922512,0.90920264,1.2298758,1.6071383,1.7655885,1.901403,1.9881734,1.9730829,1.7429527,1.1091517,0.8601585,0.694163,0.69793564,0.91297525,1.327964,1.9730829,2.2447119,1.8674494,1.2411937,1.4260522,1.2902378,1.0978339,1.0676528,1.0525624,0.5357128,0.6187105,0.51684964,0.3055826,0.1358145,0.211267,0.23767537,0.1659955,0.35085413,0.66775465,0.5055317,0.68661773,1.3958713,1.9089483,1.8259505,1.0789708,0.4678055,0.271629,0.21881226,0.18485862,0.18485862,0.18485862,0.11317875,0.056589376,0.049044125,0.06790725,0.026408374,0.02263575,0.033953626,0.033953626,0.011317875,0.0150905,0.030181,0.15467763,0.2678564,0.03772625,0.011317875,0.0,0.049044125,0.120724,0.120724,0.08299775,0.13204187,0.24899325,0.39989826,0.5093044,0.784706,0.9507015,0.98842776,0.97710985,1.1091517,0.98465514,0.56589377,0.26408374,0.18863125,0.15845025,0.1358145,0.10940613,0.14713238,0.211267,0.18485862,0.10186087,0.07922512,0.060362,0.03772625,0.049044125,0.05281675,0.02263575,0.0,0.0,0.003772625,0.003772625,0.003772625,0.00754525,0.0150905,0.0,0.011317875,0.24899325,0.31312788,0.150905,0.041498873,0.00754525,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.011317875,0.1659955,0.33953625,0.5583485,1.0148361,0.91674787,0.41876137,0.07922512,0.041498873,0.056589376,0.1056335,0.17354076,0.150905,0.060362,0.0150905,0.003772625,0.011317875,0.0150905,0.0150905,0.02263575,0.0452715,0.018863125,0.0,0.0,0.0,0.03772625,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.026408374,0.018863125,0.018863125,0.041498873,0.06413463,0.07922512,0.094315626,0.13204187,0.17354076,0.10940613,0.049044125,0.033953626,0.056589376,0.0452715,0.0452715,0.041498873,0.041498873,0.041498873,0.06790725,0.049044125,0.03772625,0.05281675,0.08677038,0.060362,0.03772625,0.02263575,0.0150905,0.018863125,0.018863125,0.030181,0.041498873,0.056589376,0.07922512,0.09808825,0.10940613,0.116951376,0.120724,0.120724,0.181086,0.30935526,0.45648763,0.56212115,0.5583485,0.4640329,0.45648763,0.5998474,0.77338815,0.70170826,0.6451189,0.4678055,0.3055826,0.23013012,0.26408374,0.29803738,0.32067314,0.362172,0.41876137,0.43007925,0.43385187,0.40367088,0.452715,0.60362,0.7997965,0.7130261,0.60362,0.5394854,0.5394854,0.5696664,0.58475685,0.7696155,0.7922512,0.62625575,0.5583485,0.59230214,0.6413463,0.6488915,0.633801,0.68661773,0.65643674,0.58475685,0.5583485,0.5583485,0.452715,0.49421388,0.5281675,0.5093044,0.46026024,0.45648763,0.5319401,0.66020936,0.73188925,0.7205714,0.6752999,0.55080324,0.482896,0.482896,0.5093044,0.4376245,0.30181,0.23390275,0.2263575,0.23767537,0.20749438,0.12826926,0.120724,0.17354076,0.23013012,0.20749438,0.19240387,0.18863125,0.18863125,0.2263575,0.35462674,0.41498876,0.38858038,0.33576363,0.29426476,0.27917424,0.32821837,0.3961256,0.47912338,0.55457586,0.59607476,0.62625575,0.60362,0.59607476,0.6111652,0.58475685,0.59230214,0.62625575,0.6073926,0.52439487,0.44516975,0.45648763,0.44139713,0.41121614,0.362172,0.29049212,0.31312788,0.35839936,0.3961256,0.4376245,0.52062225,0.724344,0.935611,1.0148361,0.9205205,0.73566186,0.7432071,0.694163,0.5998474,0.5394854,0.6828451,0.66775465,0.55457586,0.47912338,0.4640329,0.392353,0.3961256,0.38103512,0.3470815,0.3055826,0.27917424,0.3055826,0.27917424,0.21503963,0.16976812,0.23013012,0.2867195,0.36594462,0.45648763,0.5281675,0.5357128,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.1358145,0.35462674,1.3241913,2.214531,2.9652832,4.0291634,6.3719635,7.9262853,6.6020937,5.4967146,5.696664,6.247467,5.4891696,4.644101,3.953711,3.5802212,3.6141748,3.802806,3.3953626,3.180323,3.270866,3.1312788,2.2711203,1.4826416,0.80356914,0.30935526,0.1056335,0.02263575,0.056589376,0.056589376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.033953626,0.03772625,0.0,0.0,0.0,0.00754525,0.041498873,0.124496624,0.10186087,0.116951376,0.20372175,0.3772625,0.67152727,1.9202662,4.9647746,8.031919,10.876478,14.803781,25.72553,36.292652,51.764187,70.302864,82.95625,65.54936,47.946293,36.96418,32.146538,25.770802,23.639269,41.283836,79.4628,111.82815,84.95574,41.830868,24.054256,19.078165,22.688566,39.02026,86.34784,98.673004,82.99398,58.102196,54.559704,43.132423,32.644524,27.125174,28.030603,34.24789,33.738586,21.65864,12.936331,13.690856,21.217243,26.747911,25.272816,22.454664,22.31885,27.21949,27.99665,21.115381,20.360857,26.634733,27.947605,25.68403,19.444109,12.743927,7.9036493,6.0286546,5.27413,6.609639,9.476834,10.714255,4.5422406,5.1760416,5.824933,5.43258,4.085753,3.0105548,3.6745367,3.2935016,3.9159849,6.530414,11.057564,9.537196,6.8774953,5.621211,6.5341864,8.60913,9.0807085,8.00551,6.33801,5.5268955,7.4999785,9.563604,10.93684,12.208215,13.3626375,13.7851715,17.308804,16.365646,15.313085,15.539442,15.460217,14.332202,15.045229,16.55428,16.731592,12.355347,8.835487,8.360137,11.657412,20.172226,36.05875,56.7931,54.378616,44.682972,37.292397,35.496628,13.804035,6.820906,9.563604,18.549997,31.79191,40.849983,38.710907,33.018013,29.467974,31.799456,35.836166,31.874908,26.879953,24.261751,23.888262,17.399347,13.977575,11.193378,8.420499,6.8661776,4.4630156,3.4330888,3.6594462,4.459243,4.587512,5.6363015,7.4773426,10.431308,13.441863,14.04171,14.520834,15.935568,26.581915,51.070026,90.32419,91.531425,76.16175,59.245304,49.013943,46.89373,46.19202,55.736763,80.93413,125.49637,191.48712,196.62544,173.27667,152.96863,137.07455,96.79047,64.040306,47.42567,37.115086,28.554998,22.473528,21.922724,19.357338,18.52736,19.4592,18.429274,12.377983,10.457717,14.784918,19.564833,11.121698,16.505234,14.034165,13.257004,16.558052,19.17248,26.08393,26.551735,21.862362,16.539188,18.35382,25.446356,33.338688,32.361576,24.695602,24.386248,24.476791,28.796446,30.95816,29.573606,28.234325,36.088932,48.100967,49.72697,36.681232,14.947141,8.820397,14.68683,24.895552,28.200373,9.748463,10.533169,14.694374,18.078419,17.240896,9.405154,4.2102494,2.584248,4.353609,8.6732645,13.996439,18.69713,15.39231,15.131999,18.387774,15.060319,7.598067,6.960493,9.940866,12.487389,9.699419,6.1720147,8.797762,10.552032,8.507269,3.821669,2.335255,1.4637785,0.9922004,0.7696155,0.7130261,0.7809334,0.91297525,0.7507524,0.36594462,0.27917424,0.13958712,0.08677038,0.120724,0.24899325,0.52062225,0.8224323,0.8941121,0.9997456,1.0978339,0.8262049,0.845068,1.116697,1.4222796,1.6071383,1.5882751,1.5543215,1.4298248,1.3732355,1.3355093,1.0638802,0.95447415,0.935611,0.9205205,1.0186088,1.5543215,3.0746894,3.9084394,3.350091,1.8976303,1.2411937,1.0450171,1.0035182,1.0487897,0.9997456,0.5357128,0.3734899,0.3169005,0.20372175,0.060362,0.08677038,0.1358145,0.1056335,0.17354076,0.30181,0.2678564,0.30181,0.8563859,1.4411428,1.6033657,0.94692886,0.32444575,0.14335975,0.20749438,0.36594462,0.5281675,0.36594462,0.211267,0.13958712,0.15845025,0.20372175,0.09808825,0.041498873,0.02263575,0.02263575,0.041498873,0.026408374,0.030181,0.116951376,0.23390275,0.19994913,0.056589376,0.02263575,0.124496624,0.31312788,0.47535074,0.33953625,0.18863125,0.20372175,0.41876137,0.69793564,0.8865669,1.0676528,1.1921495,1.2185578,1.1431054,0.8563859,0.5093044,0.25276586,0.1358145,0.124496624,0.1056335,0.07922512,0.10186087,0.1659955,0.22258487,0.1358145,0.10186087,0.060362,0.00754525,0.011317875,0.030181,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.15467763,0.24522063,0.19240387,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.003772625,0.0,0.0,0.00754525,0.056589376,0.120724,0.2678564,0.633801,0.9393836,0.5093044,0.1358145,0.07922512,0.0452715,0.116951376,0.2678564,0.25276586,0.09808825,0.071679875,0.02263575,0.018863125,0.06790725,0.120724,0.071679875,0.049044125,0.0452715,0.041498873,0.030181,0.0,0.018863125,0.011317875,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.018863125,0.0150905,0.0150905,0.018863125,0.03772625,0.0452715,0.049044125,0.071679875,0.11317875,0.08677038,0.049044125,0.033953626,0.05281675,0.041498873,0.03772625,0.033953626,0.030181,0.030181,0.05281675,0.0452715,0.03772625,0.033953626,0.041498873,0.03772625,0.02263575,0.011317875,0.00754525,0.0150905,0.00754525,0.0150905,0.026408374,0.0452715,0.0754525,0.0754525,0.071679875,0.08299775,0.094315626,0.08677038,0.150905,0.29049212,0.39989826,0.45648763,0.482896,0.3470815,0.33576363,0.4376245,0.5885295,0.663982,0.51684964,0.3734899,0.2565385,0.18863125,0.1961765,0.211267,0.23390275,0.29426476,0.38480774,0.45648763,0.482896,0.41498876,0.44139713,0.59230214,0.7167987,0.7582976,0.7507524,0.6451189,0.4979865,0.5017591,0.5583485,0.66775465,0.7130261,0.6413463,0.47535074,0.5885295,0.8111144,0.90920264,0.8337501,0.694163,0.6073926,0.58475685,0.6413463,0.70170826,0.6073926,0.5885295,0.62248313,0.60362,0.52439487,0.49044126,0.58098423,0.69793564,0.7469798,0.7092535,0.6451189,0.56589377,0.48666862,0.4678055,0.48666862,0.422534,0.32444575,0.27540162,0.24522063,0.21881226,0.18485862,0.14335975,0.12826926,0.150905,0.18863125,0.16976812,0.16222288,0.181086,0.211267,0.26031113,0.34330887,0.42630664,0.41498876,0.38103512,0.35085413,0.29426476,0.29426476,0.35085413,0.41498876,0.44894236,0.43007925,0.51684964,0.59230214,0.6187105,0.6187105,0.66775465,0.62248313,0.6526641,0.663982,0.6073926,0.5093044,0.452715,0.4376245,0.43007925,0.41498876,0.40367088,0.35085413,0.32067314,0.33953625,0.41498876,0.5583485,0.79602385,0.90543,0.995973,1.0336993,0.84129536,0.73188925,0.7469798,0.7054809,0.60362,0.5998474,0.6790725,0.6111652,0.543258,0.52439487,0.52439487,0.44516975,0.41876137,0.3772625,0.3055826,0.24899325,0.241448,0.23767537,0.22258487,0.20749438,0.22258487,0.23767537,0.29803738,0.35085413,0.38480774,0.44894236,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.11317875,0.23013012,1.0827434,1.8976303,2.7917426,3.9612563,5.670255,7.0359454,6.009792,5.160951,5.160951,4.7535076,3.5839937,2.9992368,2.704972,2.5502944,2.5276587,2.7502437,2.4672968,2.3428001,2.4371157,2.1956677,1.5128226,1.0525624,0.6375736,0.24522063,0.03772625,0.00754525,0.02263575,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.033953626,0.03772625,0.0,0.0150905,0.011317875,0.02263575,0.056589376,0.094315626,0.13958712,0.331991,0.8262049,1.569412,2.3013012,5.5457587,11.019837,15.331948,17.25976,17.727566,26.740366,36.062523,48.40278,62.003094,70.62731,59.347164,46.327835,37.069813,32.138992,27.185535,27.823109,36.307743,58.328556,78.98368,62.780254,34.930737,20.175999,13.996439,15.826162,29.071848,66.92259,78.21029,68.182655,49.602474,42.732525,29.24539,21.466236,17.572887,16.70141,18.946123,19.61765,11.955449,8.07719,11.050018,14.875461,18.991394,18.485863,16.16947,14.588741,16.026112,18.289686,17.308804,16.750456,17.742655,18.874443,18.146326,14.124708,9.06939,4.67051,2.052308,1.8561316,2.5125682,4.7648253,6.828451,4.3913355,5.66271,5.836251,5.111907,3.9612563,3.127506,2.2748928,1.8146327,2.595566,4.9421387,8.688355,7.5565677,6.9793563,7.2962565,7.77538,6.6058664,7.194396,7.1868505,6.228604,5.342037,6.9265394,8.186596,9.578695,10.812344,11.570641,11.4838705,12.777881,13.317367,12.396846,10.86516,11.125471,11.59705,12.249713,13.336229,13.800262,11.268831,7.7942433,6.458734,7.7150183,12.51757,22.337713,31.40333,40.906574,47.523758,47.855747,38.435505,15.999702,7.9413757,11.729091,22.571615,33.42923,44.879147,49.6402,44.022762,33.195328,31.184519,32.82561,29.860327,25.559534,22.601797,23.084692,20.017548,17.40312,14.479335,11.18206,8.14887,4.772371,3.9688015,4.4931965,5.168496,4.878004,5.3986263,6.462507,8.013056,10.084227,12.815607,17.165443,23.997667,39.17494,61.765415,84.04654,71.98168,56.114025,43.328598,36.307743,33.51977,34.72324,44.48302,68.269424,104.67902,145.44978,136.6407,126.57534,129.28032,132.21164,96.24344,72.28727,54.79738,38.986305,24.869144,17.248442,21.636003,20.006231,18.731083,20.802254,25.857573,14.551015,11.461235,13.211733,14.969776,10.461489,13.2607765,10.340765,10.193633,14.1926155,16.561823,27.215717,25.631214,20.945614,19.07062,22.703657,25.32186,32.88597,33.783855,27.483574,24.556017,20.228815,26.815819,30.546946,28.087193,26.525326,34.6742,43.837902,43.611546,32.859562,19.738375,12.306303,15.196134,21.915178,23.34123,7.7150183,6.3908267,8.710991,14.102073,17.20317,7.8734684,6.221059,5.247721,3.6368105,3.5990841,10.876478,21.296469,18.467,15.222542,15.562078,14.626467,13.626721,12.2119875,14.086982,16.863634,12.053536,7.786698,10.816116,13.151371,11.491416,7.2396674,3.7537618,2.6823363,2.1692593,1.3920987,0.55080324,0.5998474,0.83752275,0.79602385,0.44894236,0.18485862,0.1056335,0.116951376,0.13958712,0.19240387,0.3772625,0.73188925,0.9318384,1.1996948,1.4298248,1.1883769,1.1355602,1.4109617,1.8448136,2.1390784,1.8485862,1.5656394,1.2298758,1.0827434,1.1431054,1.2185578,1.0978339,1.1242423,1.1280149,1.1732863,1.5467763,3.1576872,4.7572803,4.4441524,2.5502944,1.6524098,1.4147344,1.4977322,1.5618668,1.3694628,0.80734175,0.49421388,0.41498876,0.27917424,0.06790725,0.026408374,0.060362,0.06790725,0.060362,0.06413463,0.12826926,0.16222288,0.43385187,0.90543,1.4411428,1.8184053,0.68661773,0.22258487,0.18863125,0.38480774,0.6375736,0.40367088,0.241448,0.19994913,0.24522063,0.271629,0.15845025,0.071679875,0.02263575,0.026408374,0.06790725,0.06413463,0.056589376,0.09808825,0.1961765,0.34330887,0.120724,0.056589376,0.14335975,0.33953625,0.56212115,0.47535074,0.26408374,0.22258487,0.41498876,0.69793564,0.814887,0.98842776,1.146878,1.20724,1.0751982,0.76207024,0.663982,0.4979865,0.24522063,0.120724,0.090543,0.060362,0.06413463,0.11317875,0.19994913,0.13204187,0.08299775,0.03772625,0.0,0.0,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.120724,0.14335975,0.041498873,0.011317875,0.049044125,0.090543,0.090543,0.00754525,0.0,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.02263575,0.0,0.0,0.00754525,0.003772625,0.003772625,0.0452715,0.18485862,0.5281675,0.35085413,0.150905,0.10186087,0.041498873,0.094315626,0.22258487,0.23013012,0.15467763,0.26031113,0.06413463,0.02263575,0.071679875,0.12826926,0.08299775,0.060362,0.08299775,0.07922512,0.03772625,0.011317875,0.00754525,0.003772625,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.011317875,0.0150905,0.0150905,0.02263575,0.026408374,0.026408374,0.041498873,0.05281675,0.05281675,0.03772625,0.026408374,0.041498873,0.033953626,0.033953626,0.03772625,0.033953626,0.030181,0.049044125,0.05281675,0.041498873,0.026408374,0.0150905,0.02263575,0.0150905,0.00754525,0.00754525,0.00754525,0.0,0.003772625,0.0150905,0.033953626,0.06413463,0.0754525,0.06790725,0.071679875,0.08299775,0.08299775,0.150905,0.25276586,0.34330887,0.3961256,0.40367088,0.29803738,0.271629,0.32444575,0.44139713,0.58475685,0.42630664,0.32067314,0.24522063,0.18485862,0.15845025,0.14335975,0.17731337,0.2565385,0.35462674,0.422534,0.452715,0.35085413,0.34330887,0.45648763,0.4979865,0.59230214,0.694163,0.66020936,0.5281675,0.5357128,0.66775465,0.6187105,0.59230214,0.5998474,0.49421388,0.6073926,0.84884065,0.9808825,0.9242931,0.76207024,0.65643674,0.59230214,0.6111652,0.6828451,0.694163,0.68661773,0.7205714,0.7092535,0.633801,0.5394854,0.63002837,0.7167987,0.73566186,0.694163,0.6451189,0.6187105,0.543258,0.4640329,0.40367088,0.35839936,0.30935526,0.29803738,0.2678564,0.211267,0.16222288,0.15467763,0.14335975,0.15467763,0.18485862,0.18485862,0.17354076,0.181086,0.20749438,0.24522063,0.27540162,0.33576363,0.35085413,0.36971724,0.392353,0.36971724,0.28294688,0.31312788,0.35839936,0.362172,0.31312788,0.42630664,0.49421388,0.513077,0.543258,0.694163,0.66020936,0.65643674,0.6451189,0.5998474,0.5281675,0.4678055,0.47157812,0.47157812,0.45648763,0.4640329,0.38480774,0.331991,0.32067314,0.362172,0.46026024,0.694163,0.7432071,0.8186596,0.90920264,0.7809334,0.6526641,0.6752999,0.66020936,0.58475685,0.58098423,0.62248313,0.5583485,0.4979865,0.5055317,0.6149379,0.49044126,0.41498876,0.35085413,0.29426476,0.2565385,0.20372175,0.19994913,0.20749438,0.21503963,0.22258487,0.21881226,0.26031113,0.2867195,0.29049212,0.32821837,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.00754525,0.011317875,0.0754525,0.26031113,0.9205205,1.539231,2.463524,3.7009451,4.9345937,5.300538,4.478106,3.8065786,3.5160866,2.71629,1.9881734,1.5958204,1.4109617,1.4298248,1.7618159,2.3277097,2.5238862,2.4182527,2.071171,1.5467763,0.9808825,0.5357128,0.24899325,0.09808825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.0150905,0.033953626,0.026408374,0.041498873,0.07922512,0.09808825,0.35085413,0.9205205,2.2220762,3.9273026,4.983638,9.665465,17.199398,21.96045,21.526598,16.659912,16.795727,17.338985,20.153362,25.201136,30.535627,32.425713,29.094484,25.43881,23.952396,24.740875,25.985842,21.073883,18.632996,20.63626,22.398075,18.316093,12.306303,8.805306,10.336992,17.497435,24.548471,28.917171,29.781101,26.721502,19.719511,12.166716,10.397354,9.480607,8.345046,9.81637,10.763299,6.48137,4.8440504,7.6622014,10.672756,12.294985,10.816116,9.107117,8.239413,7.4773426,7.4999785,12.494934,15.079182,13.124963,9.74469,10.178542,8.201687,5.5457587,3.1840954,1.2902378,0.9393836,0.95447415,1.9278114,3.2821836,3.2557755,4.5912848,4.870459,4.22534,3.2331395,2.9237845,1.6410918,1.0676528,1.4637785,3.1727777,6.6549106,5.2137675,6.6586833,8.311093,8.171506,4.878004,5.1156793,5.753253,5.3910813,4.496969,5.409944,6.749226,8.288457,9.646602,10.269085,9.439108,7.5188417,9.159933,9.771099,8.635539,8.941121,9.880505,9.95973,10.18986,10.453944,9.540969,7.0774446,5.2590394,4.4743333,5.583485,9.910686,12.664702,22.115128,36.83591,48.3311,41.06502,21.179516,12.178034,15.769572,25.521809,26.872408,35.104275,49.432705,51.36806,40.291634,33.474503,35.06655,35.95689,33.093468,27.645796,25.012505,24.231571,21.696367,17.693611,12.97783,8.744945,6.2097406,5.379763,5.1571784,5.160951,5.7079816,6.1833324,7.0887623,8.544995,11.004747,15.24895,23.352549,38.41664,59.38112,77.1615,74.69043,59.807423,49.300663,40.276543,31.27506,22.284895,16.886269,23.013012,41.310246,66.122795,85.51786,72.5589,75.98067,93.69314,107.20291,81.62829,73.09461,60.456314,42.660843,23.982576,14.011529,19.681786,17.765291,15.169725,17.240896,27.770292,14.758509,12.359119,13.93985,14.471789,10.544487,9.133525,7.5716586,8.345046,11.510279,14.690601,24.997414,22.424482,22.367893,26.510237,22.790428,20.30804,26.166927,32.96897,34.85528,27.502436,20.922977,25.92548,28.853037,27.411894,30.671442,36.190792,36.530327,30.509218,23.703403,28.438047,20.511763,11.740409,9.265567,11.706455,9.148616,4.4215164,3.9084394,10.110635,16.712729,8.60913,10.589758,14.5132885,14.158662,9.899368,8.741172,18.278368,18.467,15.901614,14.566105,15.8676605,20.843754,18.92726,18.297232,19.478064,15.358356,12.774108,13.626721,13.3626375,11.52537,11.736636,6.0512905,4.5497856,3.8443048,2.4371157,0.6828451,0.84129536,0.72811663,0.67152727,0.6413463,0.25276586,0.1961765,0.241448,0.26031113,0.23013012,0.24522063,0.35839936,0.5772116,1.0978339,1.7240896,1.8523588,1.569412,1.6260014,2.1013522,2.6182017,2.3465726,2.0258996,1.4260522,1.056335,1.1242423,1.5430037,1.3091009,1.177059,1.1506506,1.177059,1.1280149,1.991946,3.8556228,3.9725742,2.4107075,2.022127,1.8976303,2.0296721,2.203213,2.1315331,1.4939595,0.995973,0.83752275,0.60362,0.241448,0.030181,0.03772625,0.07922512,0.090543,0.0754525,0.11317875,0.16222288,0.25276586,0.543258,1.2562841,2.704972,1.1544232,0.35085413,0.090543,0.1659955,0.36594462,0.24522063,0.18863125,0.20372175,0.241448,0.20749438,0.150905,0.06790725,0.018863125,0.02263575,0.06413463,0.08677038,0.08299775,0.09808825,0.17731337,0.35462674,0.181086,0.090543,0.090543,0.16976812,0.31312788,0.38103512,0.28294688,0.241448,0.32821837,0.4640329,0.58475685,0.7394345,0.87147635,0.94315624,0.935611,0.68661773,0.87902164,0.8563859,0.482896,0.14713238,0.10186087,0.056589376,0.03772625,0.05281675,0.094315626,0.060362,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.02263575,0.018863125,0.18863125,0.3169005,0.27540162,0.041498873,0.00754525,0.0,0.0,0.003772625,0.003772625,0.011317875,0.0452715,0.041498873,0.003772625,0.003772625,0.0,0.0,0.00754525,0.011317875,0.00754525,0.030181,0.0754525,0.1056335,0.090543,0.033953626,0.041498873,0.09808825,0.13204187,0.181086,0.41121614,0.09808825,0.018863125,0.018863125,0.033953626,0.056589376,0.10186087,0.1358145,0.10940613,0.0452715,0.030181,0.018863125,0.00754525,0.0,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0150905,0.0150905,0.02263575,0.02263575,0.018863125,0.026408374,0.026408374,0.030181,0.026408374,0.018863125,0.02263575,0.030181,0.041498873,0.0452715,0.041498873,0.033953626,0.05281675,0.056589376,0.0452715,0.026408374,0.0150905,0.018863125,0.0150905,0.0150905,0.011317875,0.0,0.003772625,0.003772625,0.00754525,0.018863125,0.041498873,0.08299775,0.071679875,0.06413463,0.0754525,0.090543,0.150905,0.211267,0.31312788,0.40367088,0.35839936,0.30935526,0.271629,0.29049212,0.36971724,0.45648763,0.35839936,0.27917424,0.23013012,0.20749438,0.1659955,0.124496624,0.16976812,0.24899325,0.3169005,0.34330887,0.35085413,0.24899325,0.211267,0.25276586,0.23390275,0.32067314,0.5017591,0.58475685,0.55457586,0.58475685,0.77716076,0.66020936,0.543258,0.543258,0.5772116,0.62248313,0.7054809,0.76584285,0.77716076,0.76207024,0.7394345,0.6375736,0.55080324,0.543258,0.633801,0.72811663,0.7884786,0.80734175,0.77338815,0.633801,0.694163,0.7092535,0.69039035,0.66775465,0.65643674,0.69793564,0.65643674,0.51684964,0.35085413,0.31312788,0.29049212,0.29049212,0.27540162,0.23013012,0.16222288,0.15845025,0.15845025,0.181086,0.20749438,0.211267,0.18863125,0.16222288,0.16222288,0.18485862,0.1961765,0.23013012,0.26408374,0.3169005,0.392353,0.44516975,0.30935526,0.31312788,0.35462674,0.35839936,0.30935526,0.3772625,0.34330887,0.33576363,0.43007925,0.6451189,0.68661773,0.62625575,0.56212115,0.5394854,0.5281675,0.52439487,0.5319401,0.51684964,0.47157812,0.43385187,0.38103512,0.33953625,0.30181,0.26408374,0.23013012,0.40367088,0.513077,0.5885295,0.63002837,0.60362,0.49044126,0.44139713,0.41121614,0.41498876,0.5281675,0.48666862,0.43007925,0.43385187,0.52439487,0.67152727,0.55080324,0.3961256,0.31312788,0.31312788,0.3055826,0.23013012,0.18863125,0.17354076,0.17731337,0.211267,0.1961765,0.21881226,0.241448,0.23767537,0.1961765,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.041498873,0.060362,0.211267,0.44139713,0.5772116,1.1581959,2.2748928,3.4594972,3.6783094,3.361409,2.987919,2.493705,1.9353566,1.4939595,1.4222796,1.2223305,1.1091517,1.1619685,1.297783,1.9806281,2.1315331,1.871222,1.3505998,0.77716076,0.77716076,0.47535074,0.1659955,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041498873,0.10186087,0.0754525,0.026408374,0.02263575,0.041498873,0.120724,0.36594462,1.1846043,2.3956168,4.798779,7.4735703,7.7678347,9.49947,17.53139,23.277096,23.4695,20.187317,19.210207,15.165953,11.419736,10.310584,13.155144,17.037174,14.335975,10.891568,9.861642,11.7026825,10.801025,9.835234,9.465516,9.982366,11.276376,12.657157,11.846043,12.604341,15.803526,19.440336,11.434827,7.7376537,6.9755836,7.2962565,6.379509,5.168496,5.1873593,4.768598,4.568649,7.5829763,9.1825695,5.0515447,2.2447119,3.2255943,5.873977,6.802043,4.938366,3.308592,2.71629,1.7391801,2.4974778,7.884786,10.510533,8.76758,6.851087,6.6813188,4.4403796,2.4069347,1.3770081,0.65643674,1.2411937,1.3166461,1.2864652,1.2902378,1.20724,1.2298758,1.2713746,1.4373702,1.6675003,1.7391801,1.6675003,1.3543724,1.6184561,2.384299,2.7011995,3.6028569,6.5040054,8.16396,7.0774446,3.4632697,3.0746894,4.08198,4.2064767,3.410453,3.9197574,5.3382645,5.6476197,5.8664317,6.205968,6.058836,5.0439997,6.4021444,6.862405,5.828706,5.402399,7.17176,7.677292,7.786698,7.635793,6.620957,5.975838,4.1197066,2.8143783,3.1124156,5.372218,8.971302,12.162943,19.613878,30.48281,38.390232,35.9003,22.296213,17.176762,23.43932,27.298714,38.929718,48.112286,49.519474,44.166122,39.38243,47.244583,58.343647,61.388153,52.062225,33.018013,25.951887,22.903606,19.644058,15.052773,11.121698,9.205205,7.5112963,6.9869013,7.6131573,8.409182,9.993684,10.408672,12.079946,16.493916,24.186298,31.05625,49.49307,74.38862,92.84053,84.152176,74.275444,65.64368,54.38239,40.189774,26.336695,16.923996,17.833199,26.37065,40.778305,60.214867,47.176674,51.04739,63.50837,71.37807,56.642193,51.907547,43.313507,30.66767,17.610613,11.642321,12.449662,10.672756,9.507015,9.718282,9.646602,9.95973,12.706201,15.524352,15.082954,7.066127,6.175787,6.3719635,8.307321,12.593022,19.806282,27.49489,24.714466,32.282352,43.698315,25.144547,27.14781,31.135473,33.553726,32.67848,28.626678,19.896824,17.670975,19.58747,24.484337,32.39553,39.374886,29.000168,19.017803,18.991394,30.320587,28.536135,15.365902,11.54046,18.4255,18.03692,6.598321,2.987919,7.8961043,17.897333,25.46522,19.644058,32.99915,41.52151,32.30876,3.6028569,14.468017,21.311558,24.929506,25.159636,20.873934,19.87419,17.444618,16.795727,16.014793,8.058327,15.418718,17.999193,15.977067,12.336484,12.849561,7.7678347,5.3458095,3.5877664,1.8561316,0.8526133,1.6373192,0.9242931,0.52062225,0.76584285,0.5357128,0.29049212,0.28294688,0.28294688,0.21881226,0.18485862,0.21881226,0.32821837,0.7432071,1.4977322,2.425798,1.8900851,1.5430037,1.4298248,1.6146835,2.2107582,2.5540671,1.8787673,1.1544232,0.995973,1.6788181,1.629774,1.2789198,1.0336993,0.94692886,0.70170826,0.87147635,1.0450171,1.1053791,1.0940613,1.20724,1.5467763,1.5882751,2.003264,2.6521554,2.5804756,1.7127718,1.4222796,1.2147852,0.8111144,0.150905,0.090543,0.15845025,0.21503963,0.211267,0.19994913,0.24899325,0.22258487,0.32067314,0.6413463,1.1921495,0.7130261,0.32067314,0.120724,0.09808825,0.120724,0.2565385,0.29803738,0.24522063,0.1358145,0.060362,0.02263575,0.00754525,0.0,0.003772625,0.0150905,0.026408374,0.02263575,0.033953626,0.08677038,0.18485862,0.1961765,0.116951376,0.08677038,0.13204187,0.1659955,0.21503963,0.19240387,0.124496624,0.120724,0.36594462,0.7696155,0.91674787,0.9393836,0.9997456,1.267602,0.80356914,0.77716076,0.8337501,0.694163,0.18485862,0.10940613,0.10186087,0.0754525,0.033953626,0.0452715,0.02263575,0.0150905,0.00754525,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.452715,0.663982,0.47912338,0.1358145,0.026408374,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.026408374,0.0150905,0.003772625,0.00754525,0.033953626,0.056589376,0.0452715,0.00754525,0.018863125,0.060362,0.094315626,0.0452715,0.0452715,0.1659955,0.17731337,0.08299775,0.1056335,0.056589376,0.026408374,0.0150905,0.033953626,0.1056335,0.181086,0.19994913,0.19240387,0.150905,0.030181,0.018863125,0.00754525,0.00754525,0.02263575,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.033953626,0.033953626,0.011317875,0.0,0.03772625,0.0452715,0.0452715,0.0452715,0.0452715,0.0452715,0.0452715,0.041498873,0.026408374,0.0150905,0.026408374,0.02263575,0.00754525,0.0,0.0,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.026408374,0.049044125,0.056589376,0.056589376,0.090543,0.13958712,0.20749438,0.24522063,0.26031113,0.32067314,0.331991,0.30935526,0.30935526,0.32444575,0.27540162,0.26408374,0.20372175,0.1659955,0.1659955,0.1659955,0.1056335,0.1358145,0.18485862,0.23390275,0.32067314,0.29426476,0.25276586,0.18485862,0.124496624,0.1358145,0.271629,0.5885295,0.663982,0.47157812,0.41121614,0.5093044,0.543258,0.543258,0.5281675,0.5017591,0.47912338,0.47157812,0.47912338,0.5055317,0.58098423,0.663982,0.7884786,0.7696155,0.62248313,0.55080324,0.633801,0.7092535,0.79602385,0.8526133,0.7922512,0.84129536,0.7809334,0.70170826,0.65643674,0.65643674,0.76584285,0.7582976,0.5998474,0.3734899,0.29049212,0.27917424,0.26408374,0.26031113,0.24899325,0.19994913,0.17354076,0.18485862,0.19240387,0.17354076,0.1358145,0.124496624,0.13204187,0.150905,0.18485862,0.24522063,0.32821837,0.35085413,0.35839936,0.38480774,0.45648763,0.4074435,0.3772625,0.3772625,0.38103512,0.32067314,0.271629,0.2678564,0.32821837,0.452715,0.6111652,0.6111652,0.5470306,0.55080324,0.6488915,0.7469798,0.6752999,0.56589377,0.5093044,0.5055317,0.45648763,0.38480774,0.3470815,0.27917424,0.18485862,0.120724,0.20749438,0.3772625,0.5281675,0.63002837,0.70170826,0.47157812,0.32067314,0.26408374,0.28294688,0.32067314,0.35839936,0.43007925,0.6752999,0.9507015,0.8526133,0.6828451,0.5017591,0.4376245,0.4640329,0.42630664,0.3055826,0.23013012,0.19240387,0.18485862,0.19994913,0.17354076,0.150905,0.1358145,0.14713238,0.18485862,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.0754525,0.07922512,0.060362,0.17354076,0.13204187,0.58475685,1.3732355,2.1277604,2.2598023,2.0108092,2.052308,1.9278114,1.569412,1.2864652,1.1657411,1.0186088,0.9016574,0.8601585,0.90543,1.5430037,1.8561316,1.6788181,1.1317875,0.65643674,0.47157812,0.28294688,0.11317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.0150905,0.0150905,0.018863125,0.060362,0.23767537,0.7092535,2.9728284,5.6061206,7.654656,8.333729,7.0359454,7.91874,10.978339,12.706201,12.249713,11.385782,11.133017,9.774872,9.673011,11.257513,13.019329,15.279131,16.976812,18.28214,19.33093,20.247679,15.301767,15.482853,15.184815,12.310076,8.273367,7.3000293,7.726336,9.669238,13.853079,21.613369,11.359374,4.9345937,3.591539,5.915476,7.8432875,6.428553,6.277648,5.4665337,4.2819295,5.2175403,6.6586833,4.195159,2.305074,2.8143783,4.8855495,4.214022,2.9501927,2.0296721,1.5430037,0.76207024,2.2409391,5.938112,6.6813188,4.45547,4.3724723,4.5535583,3.0181,1.5052774,0.73188925,0.362172,0.59607476,0.9922004,0.9393836,0.5470306,0.65643674,0.7092535,1.0299267,1.2638294,1.2638294,1.0940613,1.2034674,1.146878,1.146878,1.1883769,0.9808825,1.9202662,4.2027044,5.1534057,3.9876647,1.780679,1.6637276,2.1315331,2.3314822,2.2107582,2.5314314,3.078462,3.3576362,3.3236825,3.1539145,3.2520027,4.1008434,4.7120085,4.285702,3.2444575,3.229367,4.821415,5.541986,5.8437963,5.9230213,5.7306175,5.3269467,4.002755,2.7879698,3.5047686,8.741172,12.1252165,10.253995,11.317875,18.94235,32.154083,43.27578,32.45212,21.296469,19.108345,22.88097,27.698612,33.863083,37.75266,38.175194,36.368107,46.474968,66.764145,93.84782,110.44737,85.408455,52.511166,36.168156,28.238098,22.432028,14.27184,15.626213,19.583696,21.605824,19.538425,13.59654,15.230087,21.217243,34.817554,54.725697,75.071465,75.576996,76.64842,77.659485,77.64817,75.31669,62.323765,56.242294,46.56551,32.157856,21.221016,14.739646,17.293713,22.4358,27.502436,33.62541,43.44932,46.614555,44.271755,37.61307,27.860836,25.125683,21.273832,15.633758,9.616421,6.722818,7.9489207,10.378491,9.397609,6.4964604,9.265567,9.476834,8.341274,8.714764,9.484379,5.5759397,11.638548,9.971047,9.5183325,14.136025,22.590479,29.467974,26.71773,28.679495,32.259716,16.920223,23.38273,35.364586,36.126656,24.499426,14.867915,16.346785,17.60684,19.055529,21.205925,24.69183,23.062057,18.663176,18.357594,23.258234,28.709677,16.448645,11.415963,13.302276,18.976303,22.49239,17.810562,10.20495,8.469543,13.298503,17.301258,8.167733,11.2650585,13.656902,11.578186,10.423763,31.765503,41.36306,41.487556,35.225,26.4876,20.760756,20.096773,22.488617,22.281124,10.133271,13.411682,17.229578,16.4411,13.687083,19.353567,22.50748,17.222033,10.4049,6.379509,6.8737226,3.942393,2.444661,1.659955,1.0827434,0.39989826,0.24522063,0.22258487,0.19994913,0.17731337,0.3055826,0.48666862,0.73566186,1.0110635,1.3317367,1.7919968,2.3767538,2.2107582,1.9768555,2.0108092,2.2862108,2.625747,2.6182017,2.0447628,1.2525115,1.1544232,1.1619685,0.8563859,0.65643674,0.6451189,0.55457586,0.68661773,0.91297525,0.9620194,0.80356914,0.6790725,0.90543,1.0412445,1.388326,1.9127209,2.2484846,1.3543724,0.90920264,0.7809334,0.7394345,0.47157812,0.33953625,0.48666862,0.482896,0.2678564,0.150905,0.2263575,0.26031113,0.27540162,0.4074435,0.90920264,0.76584285,0.6073926,0.392353,0.16976812,0.08677038,0.18863125,0.31312788,0.271629,0.1056335,0.060362,0.0150905,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.018863125,0.049044125,0.07922512,0.094315626,0.08677038,0.07922512,0.1056335,0.23390275,0.3734899,0.3772625,0.271629,0.29426476,0.694163,0.9318384,1.0978339,1.267602,1.4977322,1.0148361,0.76584285,0.633801,0.49044126,0.18485862,0.060362,0.060362,0.060362,0.030181,0.02263575,0.0150905,0.03772625,0.060362,0.06413463,0.03772625,0.00754525,0.0,0.00754525,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.27917424,0.58098423,0.6451189,0.18485862,0.0754525,0.018863125,0.0,0.003772625,0.003772625,0.011317875,0.011317875,0.02263575,0.03772625,0.0150905,0.003772625,0.0,0.041498873,0.11317875,0.181086,0.0754525,0.0452715,0.06413463,0.09808825,0.1056335,0.056589376,0.17354076,0.2678564,0.26408374,0.19240387,0.15467763,0.13204187,0.15845025,0.32821837,0.7884786,0.4640329,0.20749438,0.1056335,0.116951376,0.056589376,0.02263575,0.00754525,0.00754525,0.018863125,0.033953626,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.026408374,0.026408374,0.011317875,0.0,0.00754525,0.02263575,0.03772625,0.05281675,0.08299775,0.071679875,0.07922512,0.06790725,0.03772625,0.0150905,0.026408374,0.030181,0.026408374,0.02263575,0.011317875,0.003772625,0.003772625,0.003772625,0.003772625,0.0150905,0.018863125,0.02263575,0.02263575,0.026408374,0.056589376,0.0754525,0.1358145,0.2263575,0.30181,0.29426476,0.29049212,0.29049212,0.31312788,0.33953625,0.29803738,0.24899325,0.20749438,0.1961765,0.1961765,0.15467763,0.094315626,0.08299775,0.090543,0.124496624,0.211267,0.20749438,0.271629,0.24899325,0.13958712,0.11317875,0.29426476,0.59607476,0.90543,1.026154,0.6790725,0.58475685,0.573439,0.55080324,0.4678055,0.34330887,0.41876137,0.46026024,0.4979865,0.52439487,0.482896,0.5583485,0.7054809,0.7167987,0.5772116,0.47535074,0.56212115,0.58475685,0.6073926,0.6828451,0.8526133,1.0110635,1.0186088,0.9280658,0.7922512,0.7054809,0.73566186,0.68661773,0.5583485,0.3961256,0.29049212,0.33576363,0.3169005,0.29049212,0.27540162,0.23390275,0.16976812,0.1659955,0.1659955,0.15845025,0.16222288,0.13958712,0.1358145,0.15845025,0.19994913,0.23013012,0.2678564,0.31312788,0.33576363,0.35085413,0.43385187,0.482896,0.513077,0.48666862,0.41498876,0.331991,0.28294688,0.27917424,0.3169005,0.38480774,0.47535074,0.49421388,0.49421388,0.49044126,0.5093044,0.5772116,0.6413463,0.6451189,0.6451189,0.6375736,0.56589377,0.45648763,0.4376245,0.392353,0.27540162,0.14713238,0.15467763,0.17731337,0.241448,0.331991,0.3961256,0.33953625,0.26408374,0.23013012,0.24522063,0.271629,0.27917424,0.34330887,0.5583485,0.79602385,0.7092535,0.60362,0.56589377,0.49044126,0.40367088,0.4640329,0.46026024,0.3470815,0.26408374,0.24899325,0.22258487,0.17731337,0.1358145,0.11317875,0.120724,0.14713238,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.033953626,0.018863125,0.08677038,0.018863125,0.17731337,0.573439,1.0186088,1.1204696,1.1808317,1.3958713,1.4901869,1.3845534,1.1883769,0.9808825,0.7582976,0.6413463,0.6413463,0.633801,1.0072908,1.2298758,1.0978339,0.7092535,0.47912338,0.32821837,0.15467763,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.00754525,0.049044125,0.2867195,0.77338815,1.50905,2.4220252,3.6707642,4.7610526,5.704209,6.1908774,5.6061206,6.006019,6.8963585,7.786698,8.567632,9.533423,10.186088,11.732863,14.977322,18.99894,21.179516,23.68454,24.141027,25.042685,26.547962,26.476282,19.787418,17.53516,13.585222,8.07719,7.432071,13.536179,14.320885,11.23865,8.801534,14.566105,10.065364,5.0251365,2.6068838,4.0178456,8.484633,6.5945487,5.43258,4.236658,3.1237335,3.0746894,4.085753,2.8822856,1.690136,1.6750455,2.9351022,2.4333432,1.690136,2.6785638,4.5497856,3.6481283,4.3347464,5.330719,4.266839,1.9844007,2.546522,2.9086938,1.720317,0.66775465,0.35085413,0.27917424,0.24522063,0.47157812,0.44139713,0.22258487,0.44516975,0.60362,1.086516,1.9994912,2.5993385,1.297783,0.90543,0.83752275,0.8941121,0.875249,0.58475685,0.94315624,2.0787163,2.7389257,2.305074,0.7997965,0.9280658,1.1808317,1.3430545,1.4109617,1.5769572,1.901403,2.704972,3.2218218,3.1539145,2.674791,3.4972234,3.6179473,3.1576872,2.625747,2.916239,3.0520537,3.4632697,3.8292143,3.9914372,3.953711,3.6481283,2.9803739,2.2975287,2.6936543,5.994701,11.883769,9.805053,8.793989,13.671993,25.046457,33.97626,27.117628,20.526854,19.63274,19.229069,17.53139,22.066084,30.350769,39.386204,45.682716,51.371834,70.54809,103.30956,135.22597,137.35373,98.62019,61.550377,38.654316,29.037895,18.402864,26.959179,39.405067,45.64499,41.20838,27.24967,23.046967,28.875671,45.592175,68.26188,86.170525,89.13958,86.928825,79.65143,73.45301,80.500275,54.933193,45.25641,37.333897,26.536644,17.738882,10.736891,12.079946,14.784918,16.746683,20.734346,34.538383,35.07032,29.32084,22.458437,17.82188,15.565851,13.830443,12.313848,9.831461,4.293247,7.8734684,11.385782,9.442881,4.9044123,8.858124,9.446653,10.533169,9.733373,7.828197,8.756263,14.007756,11.276376,9.378746,12.981603,22.590479,27.200626,23.61286,24.367384,27.061039,14.339747,15.958203,23.356321,22.797974,15.501716,17.652113,17.667202,15.24895,14.479335,17.18808,22.960196,21.42851,20.492899,22.46221,25.291677,22.582933,10.325675,12.525115,16.920223,19.149845,22.764019,24.457928,19.862871,16.124199,14.656648,11.148107,13.147598,16.761772,17.440845,15.580941,16.505234,40.842438,49.50816,44.890465,34.632698,31.599506,25.431265,22.194353,22.137764,21.696367,13.487134,14.260523,20.172226,23.209188,23.914669,31.407103,28.475773,17.712475,8.341274,5.0968165,8.213005,3.9084394,2.9992368,2.474842,1.3166461,0.49421388,0.6149379,0.6488915,0.6828451,0.7582976,0.8865669,1.3958713,1.4637785,1.3015556,1.1091517,1.056335,1.5505489,1.5769572,1.659955,2.003264,2.4786146,2.3654358,2.3956168,2.1202152,1.5920477,1.3430545,1.0374719,0.6413463,0.4376245,0.46026024,0.49044126,0.67152727,1.1091517,1.2411937,0.9205205,0.422534,0.56589377,0.73188925,0.94315624,1.1808317,1.4071891,1.1619685,0.9205205,0.87147635,0.9280658,0.7432071,0.3734899,0.36594462,0.3470815,0.22258487,0.15467763,0.38103512,0.35839936,0.2678564,0.30935526,0.7092535,0.8111144,0.6451189,0.392353,0.17354076,0.049044125,0.08677038,0.14713238,0.12826926,0.049044125,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.011317875,0.0150905,0.060362,0.08299775,0.07922512,0.06790725,0.10186087,0.46026024,0.784706,0.814887,0.63002837,0.62248313,0.965792,1.1544232,1.2789198,1.3656902,1.3656902,1.0299267,0.8601585,0.80356914,0.7167987,0.40367088,0.1961765,0.090543,0.041498873,0.018863125,0.0150905,0.0150905,0.049044125,0.094315626,0.11317875,0.056589376,0.011317875,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.0452715,0.124496624,0.24522063,0.30935526,0.14335975,0.20372175,0.124496624,0.05281675,0.033953626,0.018863125,0.0150905,0.00754525,0.011317875,0.026408374,0.0150905,0.011317875,0.003772625,0.018863125,0.05281675,0.08677038,0.060362,0.08299775,0.120724,0.150905,0.17731337,0.10940613,0.14713238,0.22258487,0.29426476,0.34330887,0.23767537,0.16976812,0.17731337,0.27540162,0.45648763,0.3169005,0.2263575,0.16222288,0.11317875,0.07922512,0.026408374,0.011317875,0.00754525,0.00754525,0.02263575,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.011317875,0.0150905,0.0150905,0.00754525,0.0150905,0.02263575,0.02263575,0.0150905,0.00754525,0.00754525,0.011317875,0.018863125,0.03772625,0.071679875,0.0754525,0.090543,0.090543,0.06413463,0.033953626,0.02263575,0.02263575,0.026408374,0.026408374,0.0150905,0.003772625,0.003772625,0.00754525,0.00754525,0.00754525,0.0150905,0.011317875,0.011317875,0.018863125,0.026408374,0.041498873,0.08677038,0.16976812,0.24522063,0.24522063,0.23013012,0.26031113,0.3169005,0.35462674,0.2867195,0.241448,0.22258487,0.20749438,0.18485862,0.14335975,0.1056335,0.06413463,0.05281675,0.090543,0.18485862,0.24899325,0.43385187,0.3772625,0.116951376,0.07922512,0.19240387,0.33953625,0.5281675,0.784706,1.1317875,0.9507015,0.69039035,0.5017591,0.422534,0.3772625,0.41876137,0.41498876,0.41121614,0.42630664,0.47535074,0.59230214,0.68661773,0.66020936,0.52439487,0.422534,0.482896,0.52439487,0.56212115,0.6451189,0.8224323,0.97710985,0.98842776,0.9280658,0.8526133,0.77338815,0.7469798,0.7809334,0.7432071,0.59607476,0.392353,0.4074435,0.36594462,0.3169005,0.2867195,0.27917424,0.23767537,0.24522063,0.2263575,0.17354076,0.150905,0.16222288,0.14713238,0.14713238,0.1659955,0.19240387,0.20749438,0.24899325,0.29049212,0.331991,0.3734899,0.46026024,0.5470306,0.58098423,0.5357128,0.42630664,0.38480774,0.35839936,0.35839936,0.38858038,0.43385187,0.45648763,0.49421388,0.5319401,0.56212115,0.58098423,0.633801,0.65643674,0.694163,0.7092535,0.5772116,0.4979865,0.43007925,0.36971724,0.29426476,0.16976812,0.14335975,0.11317875,0.124496624,0.1961765,0.29426476,0.23767537,0.19994913,0.1961765,0.21881226,0.24899325,0.271629,0.30181,0.39989826,0.5281675,0.56212115,0.5772116,0.58098423,0.5281675,0.45648763,0.45648763,0.5017591,0.41121614,0.33953625,0.32821837,0.32821837,0.2678564,0.21503963,0.19994913,0.21881226,0.21881226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.03772625,0.03772625,0.0452715,0.00754525,0.0,0.13958712,0.3772625,0.47912338,0.7054809,0.9808825,1.2185578,1.327964,1.2147852,0.8526133,0.513077,0.35839936,0.36971724,0.392353,0.66020936,0.814887,0.7054809,0.47157812,0.5470306,0.29049212,0.090543,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.03772625,0.049044125,0.0754525,0.19994913,0.65643674,1.5580941,2.8219235,4.1498876,4.708236,4.398881,4.459243,5.1269975,5.6363015,5.6815734,6.149379,7.2962565,8.688355,9.1976595,10.699164,12.713746,16.886269,22.541435,26.70264,33.293415,35.47022,34.330887,31.648552,29.882963,27.913652,21.394556,11.717773,4.9157305,11.664956,23.726038,22.873425,14.02662,5.1760416,7.3717093,8.228095,5.696664,2.8898308,2.3616633,6.092789,4.7006907,3.361409,2.3616633,1.780679,1.5015048,1.871222,1.5241405,0.9997456,0.7696155,1.2525115,1.1959221,1.1280149,2.8785129,5.1835866,3.6556737,3.7952607,3.6028569,2.3880715,0.97333723,1.6976813,2.3767538,1.2261031,0.271629,0.27540162,0.7205714,0.56212115,0.3169005,0.14713238,0.1659955,0.4376245,0.58475685,1.5656394,3.1312788,3.8820312,1.267602,0.76207024,0.65643674,0.76207024,0.8563859,0.663982,0.63002837,0.8186596,1.1355602,1.237421,0.55457586,0.69039035,0.95447415,1.1393328,1.1996948,1.2411937,1.5165952,2.6068838,3.451952,3.4670424,2.5314314,3.0633714,2.6634734,2.1768045,2.263575,3.4142256,2.444661,2.2862108,2.5087957,2.704972,2.505023,2.2673476,2.071171,2.173032,2.595566,3.1425967,8.7600355,8.386545,8.175279,11.3820095,18.38023,21.851044,18.881989,17.350302,18.68204,17.833199,14.890551,20.225042,29.090712,39.02026,49.82883,51.85096,64.191216,88.76232,121.78411,153.7986,140.82077,92.49722,52.03959,33.74613,22.93756,36.021023,52.36781,59.792336,54.220165,39.69556,29.928234,30.120638,40.81603,56.22343,64.22894,67.914795,68.68064,63.64041,58.834087,69.23144,43.777542,32.45212,27.90988,24.891779,20.243906,9.167479,8.737399,10.540714,11.495189,13.849306,21.462463,21.145563,18.58395,16.7995,16.143063,13.241914,12.0233555,15.056546,16.859861,3.904667,9.420244,13.038192,10.344538,5.2062225,9.756008,11.0613365,12.898605,11.589504,9.137298,13.223051,16.497688,10.944386,7.232122,10.31813,19.451654,18.116146,17.184307,20.760756,23.997667,13.132507,9.752235,11.506506,10.801025,9.95973,21.217243,18.059555,11.77059,10.601076,15.965749,22.4773,23.212961,23.797718,24.582424,24.178753,19.440336,10.140816,11.695138,16.32792,19.1423,18.104828,22.020813,24.435291,23.518545,18.885761,11.6008215,24.80501,29.769783,27.257215,21.085201,18.112373,40.849983,50.854984,48.89699,41.993088,43.46064,32.425713,24.401339,20.096773,17.723793,13.008011,14.856597,21.4436,25.676485,27.34776,33.14251,28.74363,18.648085,11.291467,10.246449,14.203933,9.933322,5.873977,2.8936033,1.2411937,0.5357128,0.79602385,0.965792,1.086516,1.1808317,1.2638294,1.599593,1.50905,1.3166461,1.1355602,0.86770374,0.8601585,0.87902164,1.056335,1.4524606,2.0636258,2.093807,2.0673985,1.901403,1.7467253,2.003264,1.5958204,0.94692886,0.47912338,0.33576363,0.38858038,0.5696664,1.0299267,1.3091009,1.1280149,0.3961256,0.36971724,0.4640329,0.55457586,0.62625575,0.79602385,1.0374719,1.0676528,1.146878,1.2902378,1.2525115,0.5319401,0.24522063,0.16222288,0.14713238,0.14335975,0.38858038,0.392353,0.29426476,0.25276586,0.44139713,0.58098423,0.5055317,0.3169005,0.120724,0.030181,0.026408374,0.02263575,0.018863125,0.018863125,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.05281675,0.090543,0.094315626,0.07922512,0.094315626,0.63002837,1.0035182,1.056335,0.9318384,1.0789708,1.4939595,1.5807298,1.5354583,1.4260522,1.1921495,0.9922004,0.95824677,0.98465514,0.94315624,0.67152727,0.38480774,0.2263575,0.120724,0.0452715,0.041498873,0.026408374,0.041498873,0.0754525,0.094315626,0.049044125,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.003772625,0.011317875,0.049044125,0.094315626,0.06790725,0.03772625,0.041498873,0.0754525,0.22258487,0.21881226,0.14713238,0.071679875,0.03772625,0.02263575,0.00754525,0.003772625,0.00754525,0.00754525,0.033953626,0.03772625,0.02263575,0.0,0.0,0.026408374,0.06790725,0.09808825,0.120724,0.13958712,0.14713238,0.14713238,0.20749438,0.33953625,0.5319401,0.44139713,0.2867195,0.19240387,0.16976812,0.116951376,0.150905,0.20372175,0.17731337,0.090543,0.06790725,0.033953626,0.018863125,0.00754525,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0150905,0.0150905,0.00754525,0.02263575,0.06413463,0.06413463,0.030181,0.02263575,0.011317875,0.003772625,0.003772625,0.0150905,0.03772625,0.05281675,0.071679875,0.07922512,0.06790725,0.0452715,0.026408374,0.018863125,0.018863125,0.02263575,0.0150905,0.00754525,0.011317875,0.0150905,0.011317875,0.0,0.011317875,0.00754525,0.003772625,0.00754525,0.00754525,0.02263575,0.05281675,0.1056335,0.1659955,0.19994913,0.18863125,0.20749438,0.25276586,0.29426476,0.26408374,0.241448,0.23767537,0.2263575,0.18863125,0.13204187,0.10186087,0.06790725,0.056589376,0.090543,0.18863125,0.29803738,0.46026024,0.3734899,0.090543,0.049044125,0.090543,0.124496624,0.17731337,0.36971724,0.9242931,0.8941121,0.76207024,0.56589377,0.3961256,0.36594462,0.35085413,0.32444575,0.31312788,0.33953625,0.43385187,0.56589377,0.63002837,0.6149379,0.5319401,0.422534,0.43007925,0.51684964,0.5998474,0.6752999,0.7884786,0.9393836,0.9393836,0.8903395,0.8563859,0.8337501,0.7922512,0.814887,0.79602385,0.6752999,0.3961256,0.3734899,0.33953625,0.31312788,0.30935526,0.34330887,0.271629,0.27917424,0.27917424,0.23390275,0.15467763,0.17354076,0.17354076,0.1659955,0.15845025,0.18485862,0.19994913,0.23013012,0.2678564,0.30181,0.32444575,0.41498876,0.5093044,0.58098423,0.5998474,0.513077,0.48666862,0.41498876,0.38480774,0.4074435,0.452715,0.4376245,0.49044126,0.55457586,0.60362,0.63002837,0.633801,0.6413463,0.7054809,0.77338815,0.6790725,0.6752999,0.5772116,0.452715,0.33576363,0.1961765,0.15845025,0.1056335,0.090543,0.12826926,0.20749438,0.14713238,0.1358145,0.150905,0.17354076,0.19994913,0.23390275,0.25276586,0.27540162,0.32067314,0.40367088,0.47912338,0.51684964,0.55080324,0.58475685,0.5696664,0.56212115,0.47912338,0.41876137,0.42630664,0.4640329,0.40367088,0.38858038,0.3734899,0.36594462,0.4074435,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.07922512,0.071679875,0.0,0.011317875,0.00754525,0.05281675,0.15467763,0.24522063,0.392353,0.6451189,0.95824677,1.1996948,1.177059,0.72811663,0.35462674,0.1358145,0.090543,0.15845025,0.48666862,0.67152727,0.6073926,0.4678055,0.7130261,0.2867195,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.018863125,0.003772625,0.011317875,0.03772625,0.060362,0.12826926,0.36594462,0.5696664,1.297783,2.3993895,3.6368105,4.7044635,5.492942,5.0968165,4.9987283,5.7570257,6.9982195,7.5905213,8.688355,10.005001,10.638803,9.046755,11.7026825,16.448645,24.737103,33.1576,33.45941,39.786102,44.845192,41.657326,32.4823,28.800219,34.60629,24.842735,10.993429,4.1800685,15.169725,26.397057,23.982576,13.777626,3.6783094,3.5651307,5.881522,5.2250857,3.138824,1.3958713,2.0145817,1.7316349,1.2185578,0.9242931,0.8903395,0.7469798,0.4979865,0.58475685,0.6413463,0.5319401,0.38103512,0.4074435,0.91674787,2.033445,2.6823363,0.62625575,0.8224323,1.4373702,1.5015048,1.1091517,1.4411428,2.3880715,1.3505998,0.35085413,0.331991,1.1619685,1.026154,0.7432071,0.56212115,0.5772116,0.73188925,0.56212115,2.1466236,3.9914372,4.29702,0.9808825,0.8865669,0.7054809,0.7130261,0.86770374,0.8186596,0.9016574,0.56212115,0.362172,0.48666862,0.7092535,0.8337501,1.1657411,1.4373702,1.5920477,1.7693611,1.6863633,2.6634734,3.3161373,3.078462,2.191895,3.2784111,2.3314822,1.388326,1.7127718,3.7613072,2.505023,1.9881734,2.0862615,2.293756,1.750498,1.539231,1.5430037,2.8747404,4.485651,3.1539145,5.2854476,6.115425,7.3151197,9.57115,12.585477,13.743673,14.049255,14.268067,14.924504,16.286423,16.32792,22.439573,27.46471,31.384468,41.34797,43.709633,47.946293,60.03001,87.55885,139.77953,170.81691,127.40909,73.619,40.774532,27.453392,38.854263,52.122585,57.325035,52.779022,45.05646,33.34246,26.374422,27.027086,32.00695,31.848501,31.995632,34.727013,34.666653,33.331142,39.114574,27.789156,19.68933,19.515789,25.35204,28.645542,11.076427,8.926031,12.37421,14.264296,10.072908,9.378746,9.846551,11.3669195,13.426772,15.0905,12.113899,11.272603,17.384256,22.232079,4.5950575,11.000975,14.694374,11.989402,6.8963585,11.114153,13.0646,12.287439,10.695392,11.057564,17.014538,18.991394,9.786189,4.666737,8.311093,14.807553,7.6018395,10.416218,17.25976,20.568352,11.185833,8.544995,8.062099,7.383027,9.027891,20.394812,16.358103,8.722309,9.0957985,17.037174,20.055275,22.337713,26.091475,25.917934,21.835953,19.296976,11.857361,9.001483,13.483362,19.927006,14.84528,14.252977,23.016785,26.778091,21.915178,15.55076,33.365097,37.141495,30.03764,20.006231,19.783646,39.589928,50.409817,55.797123,57.84943,57.21563,36.786865,24.955914,18.02183,13.317367,9.190115,13.671993,18.670721,20.711712,20.68153,23.812809,25.15209,22.454664,20.311813,20.383493,21.379465,17.746428,9.6051035,3.289729,0.9318384,0.42630664,0.6073926,0.9016574,1.0638802,1.0789708,1.1657411,0.9808825,0.8563859,0.9997456,1.2940104,1.2902378,1.0940613,0.94315624,0.8186596,0.8262049,1.1959221,1.8787673,1.961765,1.7014539,1.5920477,2.3993895,2.5087957,1.6637276,0.7922512,0.3470815,0.29426476,0.38858038,0.6828451,1.0450171,1.1732863,0.58098423,0.482896,0.36971724,0.3169005,0.39989826,0.70170826,0.95824677,1.1242423,1.3392819,1.6033657,1.7882242,0.94692886,0.41498876,0.16222288,0.09808825,0.116951376,0.22258487,0.331991,0.33953625,0.2565385,0.18863125,0.18485862,0.2867195,0.2565385,0.09808825,0.056589376,0.02263575,0.011317875,0.02263575,0.049044125,0.049044125,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.033953626,0.094315626,0.124496624,0.1056335,0.090543,0.58098423,0.845068,0.9205205,0.965792,1.2525115,1.7014539,1.6939086,1.5203679,1.3128735,1.0638802,1.0148361,1.0827434,1.1280149,1.086516,0.95824677,0.62248313,0.4376245,0.26408374,0.094315626,0.08299775,0.05281675,0.041498873,0.03772625,0.030181,0.030181,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.011317875,0.00754525,0.02263575,0.11317875,0.09808825,0.05281675,0.018863125,0.02263575,0.11317875,0.20749438,0.19240387,0.090543,0.056589376,0.041498873,0.0150905,0.0,0.0,0.0,0.049044125,0.06790725,0.0452715,0.003772625,0.0,0.011317875,0.0150905,0.018863125,0.018863125,0.030181,0.13204187,0.16222288,0.23767537,0.40367088,0.6187105,0.633801,0.43385187,0.23390275,0.13204187,0.094315626,0.09808825,0.124496624,0.10186087,0.0452715,0.026408374,0.03772625,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.011317875,0.011317875,0.03772625,0.10940613,0.116951376,0.060362,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.018863125,0.033953626,0.041498873,0.041498873,0.0452715,0.033953626,0.02263575,0.0150905,0.0150905,0.011317875,0.011317875,0.011317875,0.0150905,0.011317875,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.011317875,0.030181,0.06413463,0.1056335,0.1659955,0.15467763,0.1358145,0.150905,0.19994913,0.23767537,0.23767537,0.24522063,0.241448,0.21503963,0.14335975,0.09808825,0.08677038,0.090543,0.116951376,0.19994913,0.29426476,0.31312788,0.22258487,0.07922512,0.033953626,0.041498873,0.056589376,0.071679875,0.10186087,0.1961765,0.38480774,0.6375736,0.6111652,0.35085413,0.271629,0.23013012,0.21503963,0.23767537,0.2867195,0.3169005,0.41498876,0.5055317,0.5696664,0.56589377,0.44516975,0.41121614,0.51684964,0.63002837,0.694163,0.72811663,0.90543,0.9318384,0.86770374,0.7997965,0.845068,0.8299775,0.72811663,0.6451189,0.56212115,0.331991,0.331991,0.32821837,0.32067314,0.32821837,0.41498876,0.28294688,0.25276586,0.27917424,0.29049212,0.18863125,0.17354076,0.1961765,0.1961765,0.17354076,0.20372175,0.20749438,0.23767537,0.24899325,0.2565385,0.29803738,0.392353,0.46026024,0.5319401,0.59607476,0.5885295,0.5772116,0.48666862,0.43007925,0.4376245,0.47535074,0.40367088,0.4640329,0.5357128,0.59230214,0.663982,0.63002837,0.6149379,0.6790725,0.784706,0.77338815,0.814887,0.7507524,0.5998474,0.40367088,0.23013012,0.17354076,0.10940613,0.08299775,0.08677038,0.10186087,0.07922512,0.08299775,0.10186087,0.120724,0.1358145,0.16222288,0.18863125,0.21503963,0.23767537,0.271629,0.331991,0.39989826,0.5093044,0.62625575,0.6790725,0.59230214,0.5055317,0.46026024,0.47535074,0.52439487,0.52062225,0.5696664,0.5696664,0.543258,0.63002837,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.060362,0.0,0.060362,0.030181,0.0,0.0,0.0,0.0,0.1358145,0.3772625,0.6149379,0.70170826,0.55457586,0.34330887,0.1358145,0.0,0.0,0.18485862,0.3772625,0.46026024,0.43385187,0.3961256,0.21503963,0.06790725,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.0754525,0.0754525,0.06790725,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.08677038,0.08677038,0.0150905,0.0150905,0.02263575,0.060362,0.3169005,1.1581959,1.2940104,2.746471,3.9008942,3.983892,3.0671442,3.3953626,3.4783602,3.9725742,5.2288585,7.277394,11.121698,13.5663595,14.641558,14.18507,11.84227,16.931541,38.756176,67.6658,84.408714,60.11678,43.505913,40.36709,34.89301,24.612606,20.402355,26.05375,18.03692,7.183078,0.94692886,3.3878171,6.270103,7.594294,5.27413,1.1846043,1.1581959,2.3918443,2.4522061,1.8787673,1.2449663,1.1581959,0.633801,0.59607476,0.80356914,1.0148361,0.9922004,0.51684964,0.6073926,0.8563859,0.8563859,0.19994913,0.1358145,0.4074435,1.3091009,2.1013522,0.9922004,0.80734175,2.674791,3.3764994,2.1466236,0.67152727,1.1581959,1.0638802,0.573439,0.10186087,0.26031113,0.211267,1.599593,2.354118,2.003264,1.6486372,0.6451189,2.052308,3.7499893,4.0103,1.4939595,1.4939595,0.97333723,0.7432071,0.9507015,1.0978339,1.6712729,0.90920264,0.24522063,0.23013012,0.55080324,1.267602,1.4864142,1.780679,2.4408884,3.4783602,2.233394,3.169005,3.5349495,2.71629,2.2296214,5.2665844,4.032936,2.1881225,1.7467253,3.0520537,1.659955,1.6976813,2.2220762,2.335255,1.1732863,0.80734175,0.88279426,4.496969,8.986393,5.934339,5.9984736,5.6363015,5.783434,6.541732,7.201941,9.484379,12.657157,13.822898,12.038446,8.314865,8.477088,9.431562,10.687846,13.894578,22.843245,28.64177,27.823109,37.760204,72.0345,140.42842,195.47856,169.68135,112.67322,59.713108,31.678732,34.730785,40.593445,44.113304,43.69077,41.2612,31.76173,23.759993,20.89657,23.280869,27.46471,25.427492,22.371666,19.56106,17.486116,15.886524,13.162688,10.925522,13.392818,22.594252,38.37514,14.290704,9.405154,18.504726,27.07613,11.306557,7.594294,6.458734,6.349328,7.0359454,9.597558,10.099318,11.385782,11.996947,10.382264,4.9119577,12.238396,15.690348,13.422999,8.710991,9.918231,11.747954,8.782671,6.8774953,9.87296,19.57615,18.040693,8.737399,5.5080323,10.11818,12.268577,9.009028,7.462252,11.2650585,15.871433,8.560086,15.041456,13.117417,9.767326,10.751981,20.613623,16.048746,8.031919,8.586494,15.845025,14.037937,17.91997,33.12742,35.60226,23.005466,14.694374,7.432071,11.631002,18.38023,23.26955,26.381968,13.211733,21.334194,25.484081,18.674494,12.193124,29.049213,32.29367,25.272816,19.444109,34.345978,53.537323,53.043106,56.449787,64.65902,55.90653,30.041412,19.655376,14.871688,10.925522,8.179051,10.7557535,12.51757,12.668475,12.985375,17.80679,18.297232,22.160398,23.639269,20.37972,13.460726,10.382264,8.001738,4.515832,0.7696155,0.24522063,0.3169005,0.52062225,0.573439,0.52062225,0.70170826,0.663982,0.482896,0.56212115,1.0450171,1.8146327,2.354118,2.1579416,1.6825907,1.2223305,0.91674787,1.539231,1.8599042,1.6222287,1.1431054,1.3128735,2.7879698,2.2786655,1.3204187,0.694163,0.42630664,0.41498876,0.66775465,0.8262049,0.83752275,0.94692886,1.3958713,0.91674787,0.52062225,0.60362,0.94692886,1.0072908,1.0487897,1.2449663,1.5316857,1.6184561,1.5580941,1.0110635,0.4376245,0.116951376,0.150905,0.150905,0.2263575,0.3734899,0.47157812,0.27540162,0.1056335,0.1056335,0.19994913,0.26408374,0.150905,0.041498873,0.02263575,0.06790725,0.1358145,0.18485862,0.09808825,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.03772625,0.10940613,0.17731337,0.150905,0.24899325,0.32821837,0.44516975,0.56589377,0.58098423,0.5319401,0.482896,0.482896,0.573439,0.7922512,1.1959221,1.388326,1.448688,1.4335974,1.3732355,1.0072908,0.6413463,0.32444575,0.120724,0.1056335,0.1056335,0.08677038,0.056589376,0.030181,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.02263575,0.011317875,0.0,0.049044125,0.09808825,0.08677038,0.02263575,0.0,0.0,0.0,0.02263575,0.06790725,0.090543,0.06790725,0.02263575,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.018863125,0.02263575,0.018863125,0.030181,0.056589376,0.116951376,0.20749438,0.30181,0.35085413,0.422534,0.3772625,0.26408374,0.13204187,0.0452715,0.02263575,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.06413463,0.0754525,0.07922512,0.090543,0.018863125,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.02263575,0.0452715,0.033953626,0.02263575,0.0150905,0.011317875,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.011317875,0.02263575,0.056589376,0.090543,0.090543,0.090543,0.08299775,0.13204187,0.21503963,0.21503963,0.21503963,0.21503963,0.2263575,0.241448,0.23013012,0.15467763,0.12826926,0.13958712,0.17354076,0.19994913,0.23390275,0.18863125,0.12826926,0.08299775,0.0452715,0.033953626,0.030181,0.030181,0.03772625,0.060362,0.08677038,0.15467763,0.20372175,0.22258487,0.26031113,0.19994913,0.1659955,0.15845025,0.16976812,0.18485862,0.23013012,0.362172,0.45648763,0.45648763,0.3961256,0.422534,0.45648763,0.5357128,0.60362,0.52062225,0.69039035,0.814887,0.784706,0.6752999,0.7469798,0.7582976,0.6526641,0.513077,0.41876137,0.44139713,0.5772116,0.56589377,0.422534,0.3055826,0.48666862,0.36594462,0.27917424,0.24522063,0.23767537,0.21503963,0.17731337,0.15845025,0.15845025,0.1659955,0.1659955,0.14335975,0.15467763,0.181086,0.21503963,0.27540162,0.3961256,0.5017591,0.573439,0.6375736,0.7469798,0.73566186,0.694163,0.63002837,0.5357128,0.42630664,0.36594462,0.43385187,0.56212115,0.6752999,0.68661773,0.62625575,0.56589377,0.5772116,0.5998474,0.44139713,0.41876137,0.4678055,0.49044126,0.4376245,0.29049212,0.15467763,0.1056335,0.07922512,0.06413463,0.0754525,0.06413463,0.071679875,0.08677038,0.10940613,0.120724,0.15845025,0.1659955,0.19240387,0.23390275,0.26031113,0.30935526,0.31312788,0.31312788,0.32444575,0.33576363,0.3470815,0.35085413,0.35839936,0.36594462,0.36594462,0.48666862,0.59230214,0.694163,0.76584285,0.7167987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.1358145,0.1659955,0.06790725,0.018863125,0.05281675,0.060362,0.011317875,0.094315626,0.21881226,0.3169005,0.33576363,0.27540162,0.20749438,0.16976812,0.150905,0.071679875,0.17731337,0.26408374,0.30935526,0.3169005,0.31312788,0.090543,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.0754525,0.094315626,0.049044125,0.026408374,0.03772625,0.0,0.12826926,0.06413463,0.0,0.0,0.0,0.0,0.060362,0.13204187,0.16976812,0.124496624,0.15467763,0.27917424,1.1280149,2.7502437,4.6252384,2.7087448,3.2972744,4.164978,4.1272516,3.0671442,4.1272516,4.9421387,5.6589375,7.284939,11.695138,22.631977,28.415411,30.61108,28.207916,17.603067,11.706455,27.600525,47.38417,58.283283,52.66207,35.549446,28.449366,24.510744,19.63274,12.491161,11.23865,6.8359966,2.5616124,0.3961256,1.0299267,1.6184561,3.0558262,2.5993385,0.633801,0.694163,1.0223814,1.1996948,1.0487897,0.76584285,0.9016574,0.55457586,0.5055317,0.56212115,0.7205714,1.1732863,0.52439487,0.5055317,1.3505998,2.2296214,1.2487389,0.29049212,0.35462674,1.1619685,2.142851,2.4672968,2.0108092,1.9730829,2.0372176,1.7731338,0.66020936,0.845068,1.0902886,0.9280658,0.4678055,0.392353,0.6073926,1.1846043,1.5958204,1.6486372,1.4901869,0.6752999,1.9429018,3.6066296,4.2027044,2.5087957,2.1843498,1.2902378,0.70170826,0.6526641,0.73188925,1.0336993,0.8111144,0.46026024,0.2867195,0.48666862,1.7165444,2.0145817,1.50905,0.95824677,1.780679,3.338773,2.916239,2.1353056,1.8599042,2.191895,3.0935526,3.0369632,2.354118,1.6675003,1.8787673,0.90920264,0.8299775,1.1506506,1.3958713,1.1129243,0.7582976,1.418507,4.5309224,7.914967,5.7909794,4.67051,4.504514,5.010046,5.8400235,6.56814,7.092535,8.137552,8.371455,7.6810646,7.1793056,8.492179,9.910686,12.494934,15.746937,17.60684,21.187061,19.930779,27.242125,51.417107,95.65491,173.52943,185.32643,142.77122,77.252045,39.78233,35.22877,37.48103,41.340424,42.19304,36.024796,30.05273,26.90636,23.511,20.794708,23.695858,28.977533,28.822855,24.491882,18.561316,14.920732,11.348056,8.348819,12.936331,23.673222,30.69785,13.166461,6.7680893,7.779153,10.9594755,9.559832,8.68081,6.971811,6.692637,7.9489207,8.6581745,8.103599,11.02361,12.095036,9.265567,3.7650797,11.374464,18.448135,15.897841,7.484888,9.797507,10.759526,5.987156,4.08198,8.303548,16.561823,11.996947,6.349328,7.5263867,13.570132,12.6345215,9.590013,7.6697464,9.110889,10.989656,5.240176,10.03141,11.744182,8.7600355,5.3609,11.729091,8.45068,7.149124,10.106862,14.173752,10.767072,15.546988,24.205162,25.261497,18.648085,15.69412,10.208723,13.521088,18.731083,20.304268,14.04171,12.804289,27.792929,31.686277,20.402355,13.072145,29.588697,33.236828,29.068075,26.404602,38.839176,52.590393,57.611755,62.77648,64.82501,48.387688,28.28337,16.784409,11.3820095,9.374973,7.8508325,10.182315,10.714255,11.589504,14.898096,22.688566,25.650078,27.313805,26.325377,22.65084,17.584206,12.513797,6.9567204,2.806833,0.84129536,0.694163,0.3961256,0.30935526,0.2867195,0.32444575,0.55457586,0.2565385,0.14713238,0.21881226,0.4640329,0.8639311,1.177059,1.358145,1.3732355,1.3204187,1.4147344,1.5618668,1.7844516,1.841041,1.6222287,1.1280149,1.267602,1.1846043,1.2185578,1.3317367,1.1091517,0.77716076,0.80356914,1.026154,1.1732863,0.87147635,1.4411428,1.2223305,0.845068,0.7205714,1.0299267,1.0223814,0.7507524,0.5998474,0.69793564,0.9205205,1.388326,1.4713237,1.1959221,0.70170826,0.24899325,0.27917424,0.2565385,0.3169005,0.43007925,0.4074435,0.19994913,0.1056335,0.11317875,0.15467763,0.1056335,0.041498873,0.0452715,0.090543,0.16222288,0.21881226,0.22258487,0.124496624,0.03772625,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.003772625,0.0,0.02263575,0.05281675,0.06790725,0.041498873,0.08299775,0.14713238,0.18485862,0.18485862,0.17731337,0.15845025,0.14713238,0.17354076,0.27540162,0.47535074,0.73188925,1.1355602,1.4034165,1.3958713,1.1431054,1.0487897,0.8299775,0.513077,0.22258487,0.181086,0.16222288,0.15845025,0.1056335,0.02263575,0.030181,0.0150905,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.011317875,0.060362,0.07922512,0.060362,0.0150905,0.0,0.011317875,0.011317875,0.011317875,0.02263575,0.056589376,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.00754525,0.049044125,0.08299775,0.011317875,0.011317875,0.00754525,0.003772625,0.00754525,0.018863125,0.0150905,0.05281675,0.10940613,0.1659955,0.21503963,0.24899325,0.1961765,0.11317875,0.0452715,0.00754525,0.0150905,0.00754525,0.003772625,0.003772625,0.003772625,0.003772625,0.011317875,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.041498873,0.041498873,0.0452715,0.06790725,0.02263575,0.003772625,0.0,0.0,0.0,0.011317875,0.0150905,0.011317875,0.003772625,0.00754525,0.0150905,0.0150905,0.0150905,0.011317875,0.0,0.011317875,0.011317875,0.00754525,0.003772625,0.0,0.003772625,0.0,0.0,0.003772625,0.011317875,0.003772625,0.018863125,0.0452715,0.06413463,0.056589376,0.0452715,0.049044125,0.08299775,0.13204187,0.150905,0.16222288,0.14335975,0.14713238,0.17731337,0.20372175,0.16222288,0.16222288,0.16976812,0.1659955,0.150905,0.18485862,0.19240387,0.1659955,0.10940613,0.033953626,0.02263575,0.026408374,0.026408374,0.018863125,0.02263575,0.049044125,0.0754525,0.094315626,0.120724,0.18485862,0.1659955,0.116951376,0.1056335,0.1358145,0.15845025,0.2263575,0.362172,0.4074435,0.35462674,0.3734899,0.3470815,0.331991,0.4074435,0.5394854,0.59230214,0.68661773,0.84884065,0.8526133,0.7054809,0.663982,0.65643674,0.60362,0.5093044,0.41498876,0.36971724,0.38480774,0.38103512,0.331991,0.30181,0.42630664,0.44139713,0.3961256,0.35085413,0.31312788,0.24899325,0.23390275,0.1961765,0.16976812,0.16222288,0.19240387,0.1961765,0.1961765,0.20372175,0.23767537,0.29803738,0.32444575,0.3734899,0.46026024,0.59230214,0.77338815,0.83752275,0.84884065,0.80356914,0.73566186,0.6828451,0.6526641,0.6451189,0.68661773,0.77716076,0.90543,0.814887,0.69039035,0.633801,0.6488915,0.6375736,0.51684964,0.5394854,0.62625575,0.68661773,0.6073926,0.49421388,0.32821837,0.20749438,0.15467763,0.1358145,0.124496624,0.10186087,0.090543,0.09808825,0.10940613,0.14713238,0.124496624,0.116951376,0.14335975,0.19994913,0.2565385,0.29803738,0.32444575,0.3169005,0.24899325,0.25276586,0.25276586,0.27917424,0.31312788,0.3055826,0.35839936,0.46026024,0.56212115,0.6526641,0.7432071,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.06790725,0.11317875,0.049044125,0.030181,0.06790725,0.030181,0.08677038,0.071679875,0.09808825,0.14713238,0.09808825,0.25276586,0.28294688,0.28294688,0.2565385,0.1358145,0.25276586,0.27917424,0.28294688,0.27917424,0.23390275,0.1056335,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.041498873,0.018863125,0.030181,0.06413463,0.0,0.06413463,0.030181,0.026408374,0.05281675,0.0,0.030181,0.090543,0.14335975,0.23767537,0.5093044,0.5093044,0.52439487,1.1959221,2.746471,4.961002,4.640329,4.478106,4.5196047,4.617693,4.4139714,5.6287565,6.296511,7.5188417,12.566614,26.864862,36.545418,41.28761,38.80522,29.252934,15.226315,7.888559,12.808062,21.90386,29.671696,33.202873,24.51829,18.49718,16.252468,15.041456,8.2507305,4.447925,2.1541688,0.8299775,0.18863125,0.23013012,0.23767537,1.448688,1.4977322,0.3772625,0.46026024,0.5055317,0.52439487,0.49421388,0.47912338,0.6451189,0.58475685,0.44516975,0.34330887,0.44894236,0.9922004,0.7922512,0.6526641,1.056335,1.7580433,1.8033148,2.071171,1.0789708,0.7092535,1.569412,3.0218725,3.5085413,3.3764994,2.7200627,1.8297231,1.177059,2.071171,1.7844516,1.1619685,0.724344,0.65643674,0.965792,1.358145,1.7240896,1.9278114,1.7882242,1.1581959,1.8372684,2.969056,3.6858547,3.0822346,2.1881225,1.2638294,0.84129536,0.8526133,0.62248313,0.68661773,0.6828451,0.59230214,0.44516975,0.3169005,1.5241405,2.7540162,2.6295197,1.4449154,1.1732863,2.1353056,2.2409391,2.505023,2.9501927,2.584248,3.6254926,3.9650288,3.0143273,1.5203679,1.569412,1.1619685,0.87147635,0.91297525,1.1732863,1.1996948,0.97710985,1.7429527,4.3196554,6.673774,3.904667,3.4179983,3.4783602,4.1008434,4.8327327,4.768598,4.9723196,5.4967146,5.3910813,4.859141,5.2665844,6.56814,7.575431,9.574923,12.336484,14.136025,14.996184,16.546734,24.574879,42.638206,72.09109,130.35928,158.25784,134.03381,76.00707,42.577847,35.247635,35.387222,38.190285,38.880672,32.735065,28.75872,28.419184,24.857826,18.791445,18.51227,21.922724,19.772327,16.105335,13.59654,13.517315,10.201178,10.18986,14.102073,19.383747,20.300495,14.739646,10.367173,7.360391,5.8136153,5.745708,7.17176,7.605612,8.707218,9.929549,8.503497,7.541477,12.50248,12.90615,7.8244243,5.885295,9.691874,10.733118,9.239159,7.635793,10.56335,10.910432,5.587258,3.5160866,7.515069,14.305794,10.412445,6.330465,6.960493,11.514051,13.494679,10.121953,8.907167,9.454198,9.288202,3.8405323,8.710991,11.800771,9.910686,6.4436436,11.41219,6.507778,8.627994,12.981603,14.7736,9.216523,9.740918,14.286931,17.652113,17.91997,16.475054,10.993429,11.887542,15.690348,17.20317,9.480607,11.306557,30.060276,35.51549,23.695858,16.859861,24.333431,27.834427,27.144037,26.374422,33.964943,47.025772,54.189987,59.320755,59.44148,44.750877,28.532362,16.429781,10.359629,9.020347,7.9036493,10.510533,11.2801485,12.66093,16.320375,23.133736,23.163918,20.153362,16.233604,13.004238,11.529142,8.477088,4.074435,1.2298758,0.67152727,0.94692886,0.5319401,0.24522063,0.10940613,0.120724,0.21503963,0.071679875,0.0452715,0.12826926,0.35462674,0.7922512,1.1657411,1.358145,1.2940104,1.1506506,1.3656902,1.7655885,1.991946,2.4031622,2.7426984,2.1277604,1.418507,0.9242931,0.88279426,1.2110126,1.5015048,1.0714256,1.1355602,1.2751472,1.1959221,0.73566186,0.995973,1.0638802,1.0186088,0.98465514,1.0978339,1.2298758,1.0601076,0.8941121,0.84129536,0.84884065,1.2487389,1.7655885,1.7693611,1.1657411,0.40367088,0.29426476,0.2263575,0.26408374,0.38858038,0.51684964,0.392353,0.23390275,0.15467763,0.15467763,0.15467763,0.1659955,0.1358145,0.13204187,0.15845025,0.17354076,0.19240387,0.13958712,0.0754525,0.033953626,0.018863125,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.00754525,0.0150905,0.018863125,0.02263575,0.120724,0.181086,0.18863125,0.16222288,0.15845025,0.116951376,0.1056335,0.1358145,0.23767537,0.46026024,0.5696664,0.814887,1.0676528,1.2147852,1.1393328,0.90920264,0.62625575,0.36971724,0.19994913,0.181086,0.18485862,0.18863125,0.12826926,0.030181,0.02263575,0.0150905,0.02263575,0.0150905,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.033953626,0.094315626,0.120724,0.090543,0.018863125,0.00754525,0.00754525,0.003772625,0.003772625,0.018863125,0.0150905,0.003772625,0.0,0.0,0.00754525,0.02263575,0.026408374,0.094315626,0.181086,0.124496624,0.0452715,0.026408374,0.026408374,0.02263575,0.00754525,0.0,0.0150905,0.041498873,0.07922512,0.120724,0.14335975,0.11317875,0.0754525,0.06790725,0.10186087,0.0452715,0.0150905,0.0,0.0,0.00754525,0.00754525,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.026408374,0.041498873,0.041498873,0.03772625,0.033953626,0.041498873,0.02263575,0.00754525,0.0,0.0,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.003772625,0.00754525,0.00754525,0.003772625,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.018863125,0.026408374,0.033953626,0.041498873,0.03772625,0.030181,0.0452715,0.06413463,0.08299775,0.10186087,0.12826926,0.1056335,0.10186087,0.13204187,0.150905,0.17354076,0.21503963,0.21503963,0.17354076,0.1659955,0.20749438,0.19994913,0.17354076,0.13204187,0.0754525,0.049044125,0.030181,0.018863125,0.0150905,0.0150905,0.033953626,0.06790725,0.08299775,0.08299775,0.11317875,0.116951376,0.08677038,0.08677038,0.124496624,0.16222288,0.23390275,0.33953625,0.38480774,0.3734899,0.392353,0.35085413,0.3734899,0.452715,0.5470306,0.6187105,0.633801,0.8262049,0.91674787,0.8186596,0.6488915,0.5583485,0.4979865,0.452715,0.41121614,0.38858038,0.35462674,0.33953625,0.3169005,0.29803738,0.31312788,0.2867195,0.2565385,0.23767537,0.23767537,0.26031113,0.24899325,0.18485862,0.1358145,0.124496624,0.16222288,0.181086,0.20372175,0.20372175,0.18863125,0.20372175,0.241448,0.33576363,0.452715,0.58475685,0.7432071,0.87147635,0.9242931,0.875249,0.7696155,0.7582976,0.8111144,0.7884786,0.7922512,0.875249,0.9997456,0.9507015,0.84129536,0.7130261,0.6187105,0.62248313,0.482896,0.4640329,0.52062225,0.5885295,0.58475685,0.63002837,0.47535074,0.30935526,0.20749438,0.16222288,0.12826926,0.09808825,0.08299775,0.08299775,0.07922512,0.10940613,0.10186087,0.1056335,0.13204187,0.15467763,0.20749438,0.23767537,0.24899325,0.23767537,0.18485862,0.18863125,0.20372175,0.23013012,0.2565385,0.25276586,0.27540162,0.35085413,0.43007925,0.5093044,0.6375736,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.056589376,0.1056335,0.15467763,0.060362,0.16222288,0.1961765,0.211267,0.21503963,0.150905,0.31312788,0.35462674,0.38103512,0.38480774,0.23390275,0.30935526,0.32067314,0.2867195,0.22258487,0.120724,0.08299775,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.0452715,0.0,0.0,0.0,0.026408374,0.09808825,0.20749438,0.124496624,0.17731337,0.28294688,0.47535074,0.90543,1.3015556,1.7580433,2.5427492,3.7914882,5.534441,6.115425,5.4778514,5.323174,6.1833324,7.4169807,7.798016,8.959985,13.200415,22.911152,40.5859,39.789875,38.526047,32.357803,20.956932,8.084735,4.255521,3.3312278,5.6476197,10.887795,18.074646,15.354584,11.359374,10.355856,10.868933,5.670255,2.2107582,0.8978847,0.4640329,0.2565385,0.2263575,0.18863125,0.98465514,1.0035182,0.24522063,0.35085413,0.48666862,0.3169005,0.2263575,0.3055826,0.35839936,0.41876137,0.36971724,0.4376245,0.6451189,0.80734175,1.297783,1.2487389,0.9808825,0.8941121,1.4864142,2.9200118,1.7542707,0.86770374,1.569412,3.6330378,4.5950575,5.0025005,4.0706625,2.535204,2.6295197,4.3724723,3.3576362,1.7240896,0.754525,0.8865669,1.4373702,1.7316349,2.2069857,2.7653341,2.7540162,1.9466745,1.9844007,2.425798,2.9011486,3.1199608,2.233394,1.2562841,1.0110635,1.2298758,0.5357128,0.513077,0.5998474,0.69039035,0.6375736,0.27540162,1.1959221,3.0709167,3.8367596,2.969056,1.4675511,1.6712729,1.7127718,2.161714,2.6710186,1.9881734,3.8141239,4.293247,3.1161883,1.4600059,2.033445,1.7052265,1.2940104,1.3091009,1.690136,1.8146327,1.2751472,2.214531,4.217795,5.613666,3.4632697,3.983892,4.044254,4.255521,4.459243,3.7499893,3.610402,4.032936,3.8254418,3.4745877,5.149633,5.1043615,5.111907,6.187105,8.2507305,10.167224,10.763299,14.950912,23.1526,37.009453,59.392437,91.76156,117.211685,106.49366,66.458565,40.065277,33.463184,31.803228,32.391758,33.13119,32.49739,28.136238,28.377686,24.782373,17.157898,13.555041,15.83748,12.759018,9.265567,8.231868,10.453944,9.42779,11.3820095,12.883514,13.072145,13.679539,14.611377,12.642066,9.87296,7.3075747,4.82896,5.534441,7.2170315,9.129752,10.11818,8.6581745,10.940613,12.593022,10.816116,7.0548086,6.9680386,8.00551,5.406172,5.6363015,9.484379,12.057309,10.47658,5.458988,3.108643,5.836251,12.366665,12.955194,8.971302,6.5756855,8.507269,14.086982,10.38981,9.122208,9.035437,8.14887,3.7575345,8.718536,12.551523,11.570641,8.299775,11.465008,5.5080323,9.6201935,14.498198,14.373701,6.983129,6.0362,12.332711,17.101309,17.640795,17.30503,11.117926,9.107117,12.879742,17.727566,12.642066,11.989402,27.257215,31.184519,21.236107,19.60256,18.202915,20.756983,23.09601,24.337204,26.898817,40.838665,49.991055,54.389935,52.66207,42.060997,29.052984,17.38803,10.495442,8.371455,7.5792036,12.506252,13.656902,14.494425,17.13149,22.356575,20.934296,17.13149,12.581704,8.59404,6.1531515,4.0706625,1.750498,0.55457586,0.6488915,0.995973,0.62248313,0.271629,0.07922512,0.049044125,0.056589376,0.030181,0.026408374,0.116951376,0.39989826,0.9922004,1.7769064,2.3956168,2.1805773,1.3845534,1.1732863,1.6675003,1.720317,2.0070364,2.5238862,2.5729303,2.0258996,1.2298758,0.7884786,0.9280658,1.478869,1.3656902,1.6561824,1.7580433,1.4071891,0.66775465,0.7507524,1.026154,1.2034674,1.2034674,1.177059,1.3091009,1.3091009,1.3204187,1.3430545,1.2261031,1.2034674,1.5845025,1.690136,1.2751472,0.513077,0.3055826,0.23767537,0.24522063,0.30935526,0.4678055,0.4640329,0.362172,0.271629,0.23767537,0.241448,0.27540162,0.26031113,0.23013012,0.211267,0.211267,0.18863125,0.1659955,0.120724,0.06413463,0.030181,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.0150905,0.0150905,0.011317875,0.02263575,0.060362,0.17731337,0.27540162,0.3169005,0.29803738,0.24522063,0.17731337,0.15845025,0.18863125,0.29426476,0.5357128,0.6149379,0.724344,0.8639311,0.97333723,0.8941121,0.56212115,0.31312788,0.17731337,0.1358145,0.13204187,0.124496624,0.124496624,0.08677038,0.026408374,0.0150905,0.011317875,0.0150905,0.011317875,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.018863125,0.0150905,0.06790725,0.10940613,0.10186087,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.08299775,0.08299775,0.14713238,0.2678564,0.29049212,0.1056335,0.041498873,0.033953626,0.030181,0.0,0.0,0.0,0.011317875,0.03772625,0.08299775,0.1358145,0.150905,0.12826926,0.10940613,0.1358145,0.10186087,0.041498873,0.00754525,0.00754525,0.00754525,0.0150905,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.041498873,0.0452715,0.041498873,0.033953626,0.02263575,0.02263575,0.018863125,0.011317875,0.00754525,0.003772625,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.00754525,0.011317875,0.0150905,0.033953626,0.033953626,0.033953626,0.041498873,0.056589376,0.049044125,0.060362,0.06790725,0.06790725,0.06413463,0.090543,0.08299775,0.07922512,0.09808825,0.1056335,0.150905,0.19994913,0.20372175,0.17354076,0.18485862,0.19240387,0.17354076,0.15467763,0.14335975,0.11317875,0.090543,0.049044125,0.026408374,0.02263575,0.02263575,0.03772625,0.08299775,0.10186087,0.07922512,0.06413463,0.071679875,0.06413463,0.06790725,0.09808825,0.13204187,0.20749438,0.27540162,0.32821837,0.36971724,0.3734899,0.32821837,0.3772625,0.452715,0.52062225,0.58475685,0.56212115,0.68661773,0.7922512,0.77716076,0.6073926,0.4979865,0.41498876,0.362172,0.3470815,0.362172,0.331991,0.30181,0.271629,0.241448,0.2263575,0.17354076,0.15467763,0.150905,0.1659955,0.21503963,0.21503963,0.15845025,0.11317875,0.11317875,0.150905,0.15467763,0.19994913,0.21881226,0.19994913,0.16222288,0.20372175,0.29426476,0.39989826,0.5017591,0.62625575,0.76584285,0.8601585,0.8601585,0.7997965,0.7922512,0.8526133,0.8601585,0.8941121,0.98465514,1.0940613,1.0827434,0.9922004,0.84129536,0.6828451,0.56589377,0.44894236,0.38858038,0.38858038,0.42630664,0.4376245,0.5470306,0.52062225,0.3961256,0.24899325,0.19994913,0.15845025,0.116951376,0.09808825,0.10940613,0.116951376,0.13204187,0.116951376,0.116951376,0.13958712,0.15467763,0.17354076,0.21881226,0.241448,0.21881226,0.14713238,0.16976812,0.18863125,0.211267,0.23013012,0.211267,0.21881226,0.271629,0.32067314,0.362172,0.4376245,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.15467763,0.3470815,0.44139713,0.28294688,0.30181,0.3961256,0.44139713,0.43007925,0.48666862,0.41121614,0.38480774,0.42630664,0.46026024,0.32067314,0.32444575,0.29803738,0.241448,0.150905,0.026408374,0.003772625,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.00754525,0.0,0.00754525,0.10940613,0.46026024,0.29803738,0.6187105,1.2034674,1.8259505,2.2560298,3.218049,4.6818275,6.5832305,8.216777,8.2507305,6.8359966,6.092789,6.828451,8.843033,10.944386,10.450171,12.491161,20.560806,33.346233,44.747105,30.860073,22.17549,15.716756,9.1976595,1.0336993,1.0827434,0.91297525,1.4675511,4.4630156,12.370438,9.7296,6.832224,6.4511886,7.2283497,3.6971724,2.082489,1.2223305,0.8111144,0.6375736,0.56589377,0.7130261,0.86770374,0.6149379,0.15845025,0.29803738,0.59607476,0.35085413,0.181086,0.21503963,0.09808825,0.10940613,0.26031113,0.694163,1.1204696,0.80734175,1.6788181,2.093807,1.5958204,0.66775465,0.7205714,2.2560298,2.1088974,1.8033148,2.3201644,4.112161,4.889322,5.828706,5.372218,3.9348478,3.9008942,6.2889657,4.9421387,2.4182527,0.6488915,0.91674787,1.8448136,1.9504471,2.7351532,3.99521,3.832987,2.674791,2.4672968,2.335255,2.1843498,2.6898816,2.4069347,1.3619176,1.0789708,1.3807807,0.392353,0.392353,0.56212115,0.8111144,0.90543,0.47535074,1.1506506,3.0105548,4.561104,4.5912848,2.2069857,3.059599,2.1843498,1.3920987,1.2336484,1.0110635,2.71629,3.169005,2.4408884,1.599593,2.7313805,2.191895,1.720317,2.0183544,2.8445592,3.0331905,1.5543215,2.5616124,4.2027044,5.4363527,6.047518,7.77538,6.722818,5.191132,4.142342,3.2142766,3.127506,3.2633207,2.8558772,2.8143783,5.7117543,4.738417,3.7160356,3.9650288,5.330719,6.2135134,8.586494,12.804289,18.791445,28.841719,47.636936,66.798096,84.20122,80.52291,56.81573,34.489338,30.184772,26.597006,24.699375,26.231062,33.708405,27.543936,26.359331,22.57916,15.131999,9.446653,13.008011,11.77059,8.296002,5.492942,6.6058664,8.341274,10.133271,9.639057,8.360137,11.653639,11.012292,10.20495,10.280403,10.235131,7.0359454,5.028909,5.511805,6.677546,7.84706,9.480607,14.713238,9.805053,6.3116016,6.990674,5.798525,6.043745,5.7004366,7.6508837,12.249713,17.323895,9.344792,5.2552667,3.6066296,4.534695,9.763554,15.62244,11.849815,6.828451,6.4134626,13.951167,10.642575,8.201687,7.213259,6.752999,4.406426,7.605612,11.476325,11.857361,9.378746,9.461743,4.5422406,10.359629,14.84528,12.551523,4.606375,6.4474163,16.127972,19.376202,15.384765,16.81459,11.276376,7.383027,11.578186,20.175999,19.357338,16.018566,24.431519,25.906616,19.911915,24.046711,20.628714,27.415667,33.380184,33.006695,26.27256,36.243607,46.158066,49.94201,46.37688,39.09194,27.698612,17.836971,11.019837,7.7829256,7.673519,15.165953,16.309057,16.233604,17.882242,22.009495,21.496418,20.089228,16.852316,11.634775,5.0741806,2.3465726,1.1506506,0.995973,1.2864652,1.3091009,0.7507524,0.35085413,0.1659955,0.16222288,0.23013012,0.08299775,0.018863125,0.090543,0.3734899,0.97333723,2.0560806,3.2972744,3.4066803,2.3805263,1.5052774,1.6033657,1.3091009,1.056335,1.1883769,1.9542197,2.1843498,1.5656394,0.94315624,0.76584285,1.086516,1.4034165,1.9579924,2.2107582,1.8259505,0.70170826,0.8563859,1.2223305,1.3656902,1.2600567,1.2525115,1.2411937,1.2864652,1.4826416,1.7014539,1.599593,1.1619685,1.0336993,1.056335,0.9922004,0.513077,0.32444575,0.27917424,0.23767537,0.1961765,0.27540162,0.35085413,0.36594462,0.3470815,0.31312788,0.29803738,0.3169005,0.35462674,0.3470815,0.30935526,0.3169005,0.2678564,0.25276586,0.21503963,0.14335975,0.08677038,0.033953626,0.00754525,0.003772625,0.011317875,0.0150905,0.041498873,0.03772625,0.030181,0.041498873,0.094315626,0.1659955,0.32067314,0.41876137,0.40367088,0.27917424,0.20372175,0.17354076,0.21503963,0.33576363,0.5357128,0.6790725,0.7696155,0.784706,0.69793564,0.482896,0.2565385,0.14335975,0.1358145,0.16976812,0.1358145,0.049044125,0.018863125,0.00754525,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.003772625,0.018863125,0.041498873,0.018863125,0.00754525,0.0150905,0.03772625,0.041498873,0.018863125,0.018863125,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.120724,0.13958712,0.181086,0.2867195,0.43385187,0.28294688,0.10186087,0.0150905,0.02263575,0.003772625,0.0,0.0,0.003772625,0.026408374,0.07922512,0.18485862,0.22258487,0.18485862,0.10940613,0.07922512,0.124496624,0.06413463,0.011317875,0.011317875,0.0,0.011317875,0.003772625,0.003772625,0.011317875,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.03772625,0.033953626,0.02263575,0.0150905,0.011317875,0.011317875,0.011317875,0.0150905,0.011317875,0.003772625,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.0150905,0.00754525,0.003772625,0.0150905,0.033953626,0.03772625,0.041498873,0.06413463,0.10940613,0.090543,0.0754525,0.071679875,0.06790725,0.049044125,0.060362,0.06790725,0.07922512,0.090543,0.08677038,0.1056335,0.12826926,0.14335975,0.14713238,0.16976812,0.12826926,0.12826926,0.13958712,0.13958712,0.11317875,0.10940613,0.071679875,0.03772625,0.026408374,0.030181,0.056589376,0.10186087,0.120724,0.10186087,0.060362,0.056589376,0.056589376,0.056589376,0.060362,0.0754525,0.15467763,0.19994913,0.26031113,0.32444575,0.331991,0.30181,0.32067314,0.36971724,0.43385187,0.5017591,0.5017591,0.49421388,0.5281675,0.5772116,0.52439487,0.47535074,0.362172,0.271629,0.23390275,0.26408374,0.29803738,0.2565385,0.19994913,0.17354076,0.19994913,0.16976812,0.15845025,0.14713238,0.1358145,0.1358145,0.14335975,0.124496624,0.1056335,0.116951376,0.150905,0.13204187,0.16976812,0.22258487,0.24899325,0.21503963,0.20749438,0.2263575,0.271629,0.35462674,0.48666862,0.58098423,0.6828451,0.76584285,0.8224323,0.84129536,0.8262049,0.8526133,0.9242931,1.0336993,1.1883769,1.2600567,1.2147852,1.0940613,0.8941121,0.5885295,0.45648763,0.35839936,0.34330887,0.3734899,0.33953625,0.362172,0.46026024,0.4376245,0.29803738,0.25276586,0.21503963,0.15467763,0.12826926,0.14713238,0.17731337,0.181086,0.14713238,0.124496624,0.1358145,0.16976812,0.14713238,0.21881226,0.26408374,0.23013012,0.1358145,0.16976812,0.181086,0.1961765,0.20749438,0.1659955,0.1659955,0.20372175,0.23013012,0.23013012,0.23013012,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.060362,0.0,0.0,0.40367088,0.87147635,1.1016065,0.80734175,0.7092535,0.4376245,0.33576363,0.52439487,0.91674787,0.62248313,0.5583485,0.45648763,0.28294688,0.26031113,0.331991,0.13958712,0.071679875,0.17354076,0.1358145,0.026408374,0.0,0.030181,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.1659955,0.033953626,0.0,0.018863125,0.08299775,0.23013012,0.5470306,1.9429018,4.032936,6.013564,6.696409,7.405663,9.680555,13.88326,17.18808,13.551269,7.201941,6.7039547,9.159933,11.883769,12.419481,13.324911,14.558559,21.643549,32.07486,35.308,19.83269,10.012547,4.61392,2.0598533,0.41121614,0.1056335,0.0754525,0.6451189,3.1425967,9.918231,6.0248823,3.6594462,3.572676,4.3196554,2.2598023,2.625747,2.5502944,2.093807,1.4826416,1.1280149,2.252257,1.2789198,0.29426476,0.116951376,0.27540162,0.482896,0.29426476,0.20372175,0.24522063,0.0,0.060362,0.11317875,0.5017591,1.0374719,0.97710985,1.2449663,2.5767028,2.8181508,1.6863633,0.73188925,1.478869,2.4220252,2.9351022,2.9766011,3.1124156,4.29702,5.692891,6.571913,5.9003854,2.3503454,5.353355,4.5837393,2.4295704,0.6828451,0.55080324,1.6712729,1.6863633,3.218049,5.372218,3.7235808,2.757789,3.1954134,2.8596497,1.750498,2.0296721,2.1390784,1.3958713,0.9280658,0.845068,0.26031113,0.19994913,0.49421388,1.0299267,1.4034165,0.91674787,1.7467253,3.3161373,4.9534564,5.3684454,2.6710186,5.4665337,4.7912335,3.2633207,2.3390274,2.305074,1.50905,1.4147344,1.6146835,1.9881734,2.6710186,2.6597006,1.8938577,2.565385,4.3875628,4.606375,1.7995421,1.8749946,3.874486,7.194396,11.627231,15.863888,11.080199,5.13077,1.7618159,0.62625575,3.2746384,2.8822856,1.8787673,1.5580941,2.1202152,4.3422914,3.0935526,1.9089483,2.6597006,5.553304,7.9451485,8.141325,9.7220545,15.460217,27.298714,47.818024,74.51689,76.81819,53.031788,30.365858,27.385485,22.035902,18.87067,21.390783,32.05977,25.468992,21.45869,17.006994,11.314102,5.783434,6.405917,7.213259,6.9793563,5.775889,4.961002,5.873977,7.907422,9.114662,9.175024,9.382519,4.7950063,3.8669407,5.873977,8.499724,7.828197,5.715527,3.0369632,2.071171,4.659192,12.193124,9.14107,4.402653,3.9876647,6.72659,4.274384,2.4182527,5.2137675,8.201687,14.064346,32.606796,9.012801,6.417235,8.578949,7.809334,4.991183,10.751981,9.846551,5.873977,4.3913355,12.925014,11.631002,7.956466,5.9532022,6.092789,5.247721,2.8332415,4.2894745,8.6581745,12.272349,8.744945,6.507778,14.181297,17.1164,11.747954,5.583485,9.454198,12.298758,11.668729,9.480607,11.993175,11.555551,8.733627,10.710483,17.380484,21.345512,22.481071,32.55021,39.887962,40.8198,39.672924,45.592175,73.94722,87.32872,72.84939,42.189266,33.644268,37.745113,41.60828,40.20109,36.33038,21.915178,15.343266,11.69891,9.469289,10.544487,15.720529,16.70141,17.57666,19.787418,22.156626,19.836462,16.22606,12.759018,9.408927,4.6856003,3.5990841,2.2107582,2.2220762,3.2482302,2.8219235,1.1996948,0.44516975,0.27540162,0.42630664,0.67152727,0.21881226,0.041498873,0.030181,0.13204187,0.35085413,0.63002837,1.4901869,2.9652832,4.1762958,3.3123648,2.7389257,2.1994405,1.6373192,1.146878,0.97710985,1.3053282,1.1581959,0.9016574,0.7092535,0.55080324,0.62248313,1.2638294,1.9278114,1.9957186,0.76207024,0.95824677,1.2713746,1.2902378,1.0940613,1.267602,1.2902378,1.2525115,1.3807807,1.539231,1.2223305,0.8903395,0.633801,0.513077,0.47535074,0.36594462,0.2565385,0.23767537,0.18485862,0.090543,0.090543,0.12826926,0.1659955,0.19994913,0.23767537,0.27540162,0.32444575,0.33576363,0.32444575,0.3055826,0.3055826,0.35462674,0.43007925,0.45648763,0.40367088,0.3055826,0.14713238,0.041498873,0.0,0.003772625,0.0150905,0.041498873,0.03772625,0.02263575,0.02263575,0.0452715,0.1056335,0.22258487,0.30935526,0.31312788,0.23013012,0.14335975,0.11317875,0.17354076,0.29049212,0.35085413,0.4979865,0.47157812,0.3961256,0.38480774,0.52062225,0.52062225,0.34330887,0.34330887,0.48666862,0.36594462,0.1358145,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.003772625,0.0150905,0.05281675,0.08677038,0.071679875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.07922512,0.10940613,0.1659955,0.45648763,0.72811663,0.34330887,0.033953626,0.0150905,0.0150905,0.003772625,0.0,0.0,0.00754525,0.030181,0.1659955,0.14335975,0.08299775,0.041498873,0.030181,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.018863125,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.00754525,0.003772625,0.0150905,0.0150905,0.033953626,0.06413463,0.10940613,0.18485862,0.1358145,0.0754525,0.05281675,0.060362,0.060362,0.071679875,0.094315626,0.124496624,0.150905,0.1358145,0.124496624,0.11317875,0.10186087,0.09808825,0.120724,0.10940613,0.150905,0.15845025,0.11317875,0.0754525,0.06413463,0.05281675,0.033953626,0.018863125,0.030181,0.056589376,0.116951376,0.1659955,0.16976812,0.120724,0.09808825,0.10186087,0.08299775,0.05281675,0.0754525,0.124496624,0.19240387,0.271629,0.34330887,0.38103512,0.43007925,0.38858038,0.331991,0.331991,0.44139713,0.47912338,0.41498876,0.3961256,0.452715,0.48666862,0.42630664,0.29426476,0.18863125,0.15467763,0.1659955,0.32821837,0.31312788,0.24899325,0.21503963,0.21503963,0.150905,0.120724,0.094315626,0.0754525,0.0754525,0.06413463,0.05281675,0.0452715,0.05281675,0.0754525,0.08677038,0.08299775,0.10186087,0.1659955,0.27540162,0.18863125,0.1659955,0.181086,0.2565385,0.48666862,0.513077,0.5017591,0.56212115,0.7092535,0.8526133,0.8186596,0.754525,0.7582976,0.8865669,1.1280149,1.5316857,1.7240896,1.5958204,1.1996948,0.7469798,0.4678055,0.34330887,0.392353,0.4979865,0.41121614,0.32821837,0.331991,0.362172,0.362172,0.29049212,0.19240387,0.13204187,0.10186087,0.090543,0.090543,0.116951376,0.120724,0.1056335,0.08677038,0.120724,0.09808825,0.08299775,0.08677038,0.11317875,0.1358145,0.16222288,0.13958712,0.120724,0.120724,0.1056335,0.094315626,0.10186087,0.11317875,0.13204187,0.1659955,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.10186087,0.071679875,0.0150905,0.060362,0.09808825,0.07922512,0.0,0.049044125,0.17731337,0.38480774,0.5772116,0.5772116,1.3204187,1.3656902,1.0148361,0.62248313,0.62248313,0.49421388,0.4376245,0.34330887,0.241448,0.29426476,0.48666862,0.35462674,0.18485862,0.094315626,0.026408374,0.003772625,0.0,0.026408374,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.071679875,0.071679875,0.06413463,0.116951376,0.45648763,1.4600059,2.9200118,4.22534,4.515832,4.221567,5.062863,5.5268955,5.409944,6.983129,9.7220545,10.303039,10.8576145,9.876732,9.318384,9.322156,8.209232,6.779407,6.485142,8.171506,11.578186,15.339493,11.883769,7.9828744,5.1798143,3.3878171,0.9016574,0.28294688,0.07922512,0.38103512,1.6486372,4.6931453,3.62172,3.308592,3.2067313,2.867195,1.9655377,1.4411428,1.7618159,1.7391801,1.2940104,1.4600059,1.0601076,1.2261031,0.97710985,0.35462674,0.44516975,0.62248313,0.5017591,0.35462674,0.2867195,0.2565385,0.06413463,0.0754525,0.19994913,0.3470815,0.40367088,0.58475685,1.8334957,2.282438,1.5467763,0.7205714,0.94692886,1.1129243,1.3317367,1.8184053,2.8822856,2.5804756,3.531177,5.553304,7.2358947,5.938112,5.1232247,4.4705606,3.6066296,2.6710186,2.282438,2.6446102,2.2069857,3.229367,4.8930945,3.2821836,2.897376,2.9501927,2.8898308,2.6219745,2.4823873,3.1576872,2.595566,2.1353056,1.8184053,0.392353,0.41121614,0.66775465,0.9808825,1.2562841,1.4901869,2.493705,3.2520027,4.0895257,4.538468,3.3538637,3.610402,4.146115,3.5764484,2.6408374,4.195159,3.0331905,1.8825399,1.1996948,1.2713746,2.2183034,1.7467253,1.0035182,1.9278114,4.014073,4.2894745,3.5349495,5.028909,5.9532022,6.013564,7.466025,6.9755836,5.2665844,4.7044635,5.413717,5.2779026,7.2623034,8.586494,11.517824,16.143063,20.357084,10.9594755,5.4438977,5.20245,7.3905725,4.930821,4.3347464,4.9119577,6.6549106,11.7555,24.601288,53.458096,82.17155,80.61345,50.36077,24.665422,21.179516,20.673985,22.424482,24.069347,21.636003,19.810055,16.731592,14.120935,12.6345215,11.898859,8.926031,8.130007,7.5527954,6.828451,7.1793056,9.337247,8.484633,7.0510364,6.300284,6.319147,4.659192,4.8742313,6.790725,8.246958,5.1043615,5.534441,5.1269975,5.674028,7.3905725,8.956212,5.4665337,4.7120085,6.9944468,10.408672,10.86516,3.7273536,2.4672968,6.1003346,14.418973,28.030603,12.196897,15.426264,18.440592,13.513543,4.4516973,7.0510364,10.408672,9.178797,6.066381,11.827179,10.502988,7.3188925,6.458734,7.8017883,6.9227667,3.0218725,6.0248823,11.668729,15.128226,11.027383,7.462252,13.008011,14.260523,8.60913,4.2404304,8.461998,10.03141,8.941121,7.4811153,10.26154,13.238141,11.676274,12.770335,17.16167,18.94235,21.073883,26.11411,33.610317,40.09923,39.099487,56.5441,97.30732,116.03463,98.19011,60.082825,42.574074,35.44004,31.241108,26.366877,21.013521,17.033401,15.23386,13.29473,11.7894535,14.181297,18.79899,21.1682,21.496418,22.156626,27.649569,22.760246,17.082445,11.92904,8.213005,6.428553,4.055572,2.161714,2.1843498,3.4029078,2.9464202,1.0487897,0.3734899,0.39989826,0.6752999,0.7809334,0.4678055,0.19994913,0.17731337,0.32444575,0.29049212,0.38480774,0.6526641,1.2034674,1.9579924,2.6634734,3.663219,3.270866,2.6106565,2.2975287,2.4295704,1.7316349,1.0902886,0.80734175,0.84129536,0.7696155,0.6451189,0.8299775,1.2751472,1.6788181,1.4713237,1.7919968,1.750498,1.6071383,1.5316857,1.5845025,1.5203679,1.5769572,1.6486372,1.5354583,0.91674787,0.7130261,0.6187105,0.6790725,0.80356914,0.7809334,0.6413463,0.5281675,0.33576363,0.10940613,0.041498873,0.049044125,0.049044125,0.08677038,0.16976812,0.27540162,0.3055826,0.29049212,0.27540162,0.27917424,0.2678564,0.3169005,0.4074435,0.5319401,0.6111652,0.52439487,0.3470815,0.15845025,0.05281675,0.030181,0.003772625,0.018863125,0.033953626,0.056589376,0.0754525,0.071679875,0.08299775,0.11317875,0.1358145,0.124496624,0.071679875,0.06413463,0.060362,0.124496624,0.25276586,0.362172,0.47157812,0.38103512,0.241448,0.1659955,0.24899325,0.513077,0.42630664,0.2678564,0.16222288,0.10940613,0.0452715,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041498873,0.033953626,0.0150905,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.030181,0.049044125,0.056589376,0.05281675,0.049044125,0.030181,0.011317875,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.033953626,0.1056335,0.15845025,0.10186087,0.056589376,0.0452715,0.026408374,0.026408374,0.011317875,0.0,0.0,0.00754525,0.05281675,0.0754525,0.09808825,0.10186087,0.030181,0.0754525,0.033953626,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.0150905,0.00754525,0.011317875,0.02263575,0.011317875,0.003772625,0.00754525,0.00754525,0.003772625,0.0150905,0.011317875,0.003772625,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.018863125,0.02263575,0.0150905,0.0150905,0.033953626,0.08299775,0.14335975,0.14713238,0.116951376,0.10186087,0.1056335,0.11317875,0.071679875,0.0754525,0.116951376,0.181086,0.2263575,0.17354076,0.14335975,0.14713238,0.15467763,0.15467763,0.16976812,0.18863125,0.17354076,0.15467763,0.13958712,0.11317875,0.10940613,0.071679875,0.03772625,0.026408374,0.018863125,0.041498873,0.15467763,0.20372175,0.16222288,0.1358145,0.090543,0.0754525,0.06413463,0.060362,0.0754525,0.08677038,0.11317875,0.17354076,0.24899325,0.29426476,0.2867195,0.2565385,0.24899325,0.26031113,0.28294688,0.29049212,0.30935526,0.35462674,0.42630664,0.513077,0.38480774,0.2678564,0.18863125,0.14713238,0.13204187,0.181086,0.241448,0.28294688,0.29049212,0.24899325,0.19994913,0.16222288,0.1358145,0.10940613,0.05281675,0.041498873,0.033953626,0.033953626,0.033953626,0.041498873,0.060362,0.071679875,0.1056335,0.16976812,0.24899325,0.23390275,0.20749438,0.18485862,0.18863125,0.2565385,0.36971724,0.5093044,0.6488915,0.7696155,0.87902164,0.8337501,0.875249,0.9242931,0.9808825,1.1280149,1.3543724,1.4600059,1.5505489,1.5354583,1.1016065,0.59607476,0.4376245,0.4074435,0.41121614,0.47157812,0.38858038,0.3734899,0.362172,0.331991,0.29049212,0.211267,0.16976812,0.14335975,0.12826926,0.12826926,0.150905,0.1659955,0.17731337,0.17731337,0.14713238,0.11317875,0.07922512,0.08299775,0.116951376,0.150905,0.19240387,0.17731337,0.13958712,0.1056335,0.08299775,0.060362,0.06413463,0.06790725,0.06413463,0.08299775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05281675,0.124496624,0.120724,0.11317875,0.26408374,0.32444575,0.22258487,0.090543,0.10186087,0.116951376,0.181086,0.3169005,0.5281675,1.1657411,1.237421,1.0336993,0.754525,0.5017591,0.59230214,0.513077,0.36594462,0.2678564,0.331991,0.52439487,0.38103512,0.1659955,0.030181,0.0,0.0,0.071679875,0.08299775,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.120724,0.32821837,0.5093044,0.6828451,1.0148361,2.5691576,1.6410918,0.7167987,0.9318384,2.0636258,3.1916409,3.500996,3.4670424,3.6066296,4.4818783,7.986647,8.379,7.726336,7.8206515,10.159679,10.38981,9.593785,8.311093,6.952948,5.802297,3.742444,2.5616124,2.323937,3.1010978,4.9534564,5.855114,5.2590394,4.2517486,3.0369632,0.9318384,0.26408374,0.056589376,0.26408374,0.8865669,1.9881734,1.6561824,1.8297231,2.3013012,2.4371157,1.1695137,0.62248313,0.8299775,1.026154,1.0186088,1.2034674,0.90543,1.0525624,0.935611,0.5055317,0.35839936,0.43007925,0.4376245,0.33576363,0.2263575,0.33953625,0.23013012,0.211267,0.21881226,0.21881226,0.1961765,0.2867195,1.3241913,1.8863125,1.5618668,0.97333723,0.62625575,0.6073926,0.6828451,0.91674787,1.6976813,1.8674494,2.5993385,3.9650288,5.3344917,5.372218,4.7648253,4.847823,4.610148,3.9084394,3.4481792,3.2821836,3.531177,4.0706625,4.353609,3.3953626,3.3689542,3.5123138,3.3236825,2.806833,2.4672968,2.7351532,2.2484846,2.1202152,2.1579416,0.86770374,1.2487389,1.3845534,1.3091009,1.2751472,1.7316349,3.0256453,5.323174,6.405917,6.485142,8.175279,6.4134626,6.168242,4.678055,2.2899833,2.463524,2.7653341,1.659955,0.8978847,0.98465514,1.20724,1.0412445,0.7696155,1.9806281,3.9688015,3.772625,3.4557245,4.293247,4.4516973,4.236658,6.085244,5.481624,5.836251,6.3455553,6.3342376,5.247721,6.270103,7.0548086,8.552541,10.672756,12.283667,6.8699503,4.9345937,5.2137675,5.764571,3.953711,2.565385,2.535204,3.9348478,8.699674,20.613623,43.879402,67.39795,69.71811,49.06676,23.329912,17.271078,17.538933,21.353058,23.910898,18.387774,15.150862,12.664702,11.627231,11.812089,12.064855,8.371455,7.303802,7.515069,8.224322,9.239159,9.175024,6.379509,3.9876647,3.259548,3.5877664,4.4743333,5.6061206,7.1679873,7.865923,4.9119577,6.4247804,7.8696957,11.283921,13.445636,5.8513412,4.821415,7.273621,10.299266,12.381755,13.392818,4.402653,1.841041,6.507778,16.648594,27.966469,13.70972,18.229324,22.239624,17.255987,5.6098933,6.33801,11.050018,11.151879,7.5490227,10.653893,10.955703,8.412953,7.254758,7.865923,6.790725,3.2557755,6.530414,12.174261,14.392565,6.0211096,9.435335,16.158154,15.697892,8.529905,6.085244,13.219278,11.197151,8.107371,7.9791017,10.789707,11.61214,11.676274,12.536433,14.181297,15.026365,17.20317,18.587723,25.39354,36.46242,43.268234,51.52274,72.08732,84.238945,77.36522,50.956844,35.304226,27.144037,22.149082,18.09351,14.837734,14.109617,14.622695,14.354838,13.890805,16.399601,22.01704,22.530117,21.319103,21.594505,26.412148,23.020557,19.010258,14.056801,9.382519,7.752744,5.824933,4.9987283,4.5761943,3.9499383,2.5993385,1.1242423,0.49421388,0.44894236,0.6526641,0.6790725,0.43007925,0.22258487,0.2263575,0.38103512,0.43007925,0.35462674,0.31312788,0.43007925,0.77338815,1.3656902,2.1277604,2.0447628,1.8070874,1.8146327,2.161714,1.6976813,1.1091517,0.9016574,1.1393328,1.418507,1.2110126,1.1280149,1.3732355,1.841041,2.0862615,2.142851,2.1088974,2.0372176,1.9768555,1.991946,1.6071383,1.6863633,1.8070874,1.629774,0.9016574,0.80734175,0.875249,0.95447415,0.9922004,1.0487897,1.1959221,1.2034674,0.9695646,0.543258,0.120724,0.041498873,0.018863125,0.0452715,0.12826926,0.2565385,0.27917424,0.27540162,0.271629,0.2678564,0.241448,0.28294688,0.36971724,0.5357128,0.6488915,0.422534,0.29049212,0.181086,0.090543,0.02263575,0.0,0.011317875,0.033953626,0.06413463,0.090543,0.094315626,0.06413463,0.049044125,0.049044125,0.049044125,0.02263575,0.018863125,0.02263575,0.06790725,0.17354076,0.33953625,0.43007925,0.36594462,0.2263575,0.11317875,0.15467763,0.40367088,0.3961256,0.27540162,0.14335975,0.056589376,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.030181,0.026408374,0.018863125,0.0150905,0.00754525,0.0,0.0,0.0150905,0.030181,0.0,0.011317875,0.0150905,0.033953626,0.071679875,0.1056335,0.060362,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.03772625,0.071679875,0.07922512,0.056589376,0.041498873,0.0452715,0.026408374,0.003772625,0.0,0.0,0.011317875,0.041498873,0.06790725,0.071679875,0.02263575,0.0452715,0.02263575,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.0150905,0.018863125,0.00754525,0.00754525,0.011317875,0.00754525,0.003772625,0.0150905,0.0150905,0.011317875,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.018863125,0.0150905,0.02263575,0.030181,0.06790725,0.124496624,0.15467763,0.1659955,0.1659955,0.16222288,0.150905,0.1056335,0.09808825,0.124496624,0.19240387,0.26031113,0.21881226,0.1961765,0.18863125,0.1659955,0.14713238,0.18485862,0.22258487,0.1961765,0.1659955,0.1659955,0.18485862,0.15845025,0.120724,0.120724,0.14335975,0.116951376,0.10940613,0.16222288,0.17731337,0.14713238,0.12826926,0.08677038,0.060362,0.071679875,0.1056335,0.13204187,0.13958712,0.1659955,0.19994913,0.241448,0.28294688,0.30935526,0.3055826,0.28294688,0.25276586,0.21503963,0.20372175,0.23013012,0.25276586,0.271629,0.32821837,0.28294688,0.21881226,0.1659955,0.13204187,0.120724,0.13204187,0.16976812,0.19994913,0.20749438,0.18485862,0.181086,0.181086,0.16222288,0.120724,0.056589376,0.033953626,0.030181,0.026408374,0.02263575,0.02263575,0.030181,0.041498873,0.071679875,0.120724,0.16976812,0.19994913,0.23390275,0.23390275,0.19994913,0.181086,0.24899325,0.36971724,0.482896,0.58475685,0.7205714,0.7884786,0.95447415,1.0751982,1.0940613,1.056335,1.0714256,1.1431054,1.2864652,1.3807807,1.1808317,0.7507524,0.58475685,0.5772116,0.62248313,0.5885295,0.5093044,0.47912338,0.44516975,0.38858038,0.34330887,0.29426476,0.22258487,0.181086,0.181086,0.19994913,0.1961765,0.17731337,0.17354076,0.17731337,0.14335975,0.1358145,0.14713238,0.14335975,0.12826926,0.1358145,0.14713238,0.12826926,0.094315626,0.06790725,0.06790725,0.049044125,0.0452715,0.041498873,0.03772625,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05281675,0.12826926,0.13204187,0.38103512,0.91674787,1.026154,0.60362,0.13958712,0.10940613,0.1358145,0.1659955,0.24899325,0.5017591,0.8903395,0.8865669,0.77716076,0.67152727,0.47912338,0.55457586,0.47912338,0.35462674,0.26031113,0.24899325,0.34330887,0.27540162,0.1659955,0.08677038,0.049044125,0.011317875,0.071679875,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.16976812,0.36971724,0.79602385,1.1431054,1.2487389,1.2789198,1.7127718,3.2520027,2.1390784,0.95824677,0.91297525,1.8297231,2.5993385,3.270866,3.7386713,3.9650288,3.9612563,8.054554,9.593785,8.560086,6.8473144,8.280911,7.118943,6.7680893,6.0550632,4.9421387,4.52715,2.6295197,1.4071891,1.1053791,1.3694628,1.2223305,2.1164427,2.6031113,2.6068838,2.0145817,0.694163,0.18863125,0.03772625,0.1659955,0.44516975,0.7092535,0.5017591,0.59230214,2.4899325,4.2706113,0.5583485,0.23013012,0.35462674,0.5357128,0.6149379,0.6526641,0.84884065,0.77338815,0.62248313,0.47157812,0.31312788,0.3055826,0.35839936,0.32067314,0.2263575,0.28294688,0.46026024,0.6187105,0.65643674,0.5281675,0.21881226,0.2867195,0.7922512,1.3543724,1.6448646,1.3807807,0.724344,0.6413463,0.69039035,0.72811663,0.87902164,1.5203679,2.1390784,2.7426984,3.3840446,4.1800685,5.243949,5.6061206,5.119452,4.3121104,4.376245,4.3875628,4.6327834,4.4931965,3.92353,3.4557245,3.7575345,4.3422914,4.2291126,3.3727267,2.6597006,2.4069347,1.7655885,1.6184561,1.8033148,1.1091517,1.6863633,1.6524098,1.388326,1.3053282,1.8297231,3.821669,5.9984736,7.3415284,7.8961043,8.793989,7.0359454,5.8928404,3.953711,1.7165444,1.6071383,2.9464202,1.750498,0.77716076,0.7922512,0.58098423,0.6149379,0.6526641,1.7165444,3.259548,3.1539145,3.0105548,3.3915899,3.169005,2.9464202,5.040227,5.8513412,7.3000293,7.432071,6.1342883,5.1269975,5.1873593,5.836251,5.6287565,4.561104,4.085753,4.6742826,6.432326,6.2021956,4.08198,3.3953626,3.0709167,2.2598023,2.7125173,6.541732,16.21097,30.203636,44.037853,48.697044,41.43097,25.770802,17.787928,15.784663,17.003222,17.984104,14.547242,14.698147,12.0082655,9.7296,9.416472,10.940613,8.239413,6.851087,6.6586833,7.232122,7.809334,6.1041074,3.5990841,1.8938577,1.6222287,2.4333432,4.508287,5.696664,6.72659,7.0510364,4.847823,6.9982195,10.906659,14.679284,14.754736,5.915476,6.156924,8.967529,11.725319,12.860879,11.861133,4.104616,1.7731338,5.9494295,15.309312,26.117884,13.577678,17.040947,21.23988,18.21046,7.3113475,7.7942433,11.959221,11.996947,8.695901,11.415963,12.332711,9.310839,7.3377557,7.462252,6.809588,4.9459114,7.598067,11.091517,11.02361,2.2296214,9.880505,18.738628,18.150099,10.4049,10.736891,17.052265,12.151625,7.9262853,8.718536,11.32542,10.521852,15.448899,18.79899,17.527617,12.853333,15.494171,19.519562,27.815563,40.70285,55.93671,59.592384,58.977448,56.02348,49.549656,35.262726,24.631468,19.08571,16.063837,14.003984,12.336484,12.253486,14.305794,15.984612,16.999449,19.304522,23.465727,23.246916,22.658386,23.688313,26.310287,24.918188,22.028357,15.965749,9.031664,7.484888,6.7643166,6.609639,5.775889,4.0103,2.0636258,1.2034674,0.6752999,0.49044126,0.5281675,0.4979865,0.27540162,0.18485862,0.23767537,0.38103512,0.47912338,0.3169005,0.18863125,0.17354076,0.29803738,0.52439487,1.0148361,1.1921495,1.4373702,1.7919968,1.9466745,1.7429527,1.2110126,1.0072908,1.3317367,1.8938577,1.5618668,1.3996439,1.6788181,2.191895,2.252257,2.191895,2.3465726,2.293756,2.04099,2.0296721,1.7769064,1.9957186,2.0485353,1.6788181,1.026154,1.0450171,1.2261031,1.3430545,1.3091009,1.177059,1.2185578,1.2034674,1.0186088,0.66775465,0.29426476,0.23013012,0.15467763,0.09808825,0.09808825,0.17731337,0.211267,0.24899325,0.271629,0.26408374,0.21503963,0.24899325,0.3169005,0.47535074,0.58475685,0.34330887,0.211267,0.19240387,0.14335975,0.05281675,0.0,0.00754525,0.026408374,0.049044125,0.06413463,0.08299775,0.049044125,0.02263575,0.011317875,0.0150905,0.00754525,0.0,0.003772625,0.026408374,0.08299775,0.21503963,0.2867195,0.28294688,0.20372175,0.1056335,0.10186087,0.23390275,0.24899325,0.1961765,0.124496624,0.060362,0.018863125,0.003772625,0.003772625,0.011317875,0.030181,0.00754525,0.0,0.003772625,0.0150905,0.041498873,0.018863125,0.011317875,0.0150905,0.026408374,0.049044125,0.03772625,0.049044125,0.060362,0.060362,0.026408374,0.011317875,0.003772625,0.0150905,0.030181,0.0,0.0,0.0,0.0150905,0.0452715,0.08299775,0.049044125,0.026408374,0.011317875,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.00754525,0.030181,0.05281675,0.05281675,0.033953626,0.026408374,0.033953626,0.02263575,0.011317875,0.003772625,0.0,0.0,0.018863125,0.033953626,0.030181,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.00754525,0.011317875,0.011317875,0.00754525,0.0150905,0.011317875,0.011317875,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0150905,0.026408374,0.041498873,0.07922512,0.14335975,0.19994913,0.18863125,0.16222288,0.13958712,0.10940613,0.1056335,0.120724,0.20749438,0.31312788,0.3055826,0.26031113,0.241448,0.20749438,0.17354076,0.17731337,0.211267,0.20372175,0.19994913,0.21881226,0.25276586,0.20372175,0.17731337,0.20372175,0.25276586,0.21881226,0.18485862,0.1961765,0.19240387,0.1659955,0.150905,0.120724,0.08299775,0.0754525,0.09808825,0.13204187,0.17354076,0.21881226,0.25276586,0.28294688,0.331991,0.35085413,0.33576363,0.30181,0.26408374,0.241448,0.22258487,0.23390275,0.21503963,0.16976812,0.15467763,0.1659955,0.14713238,0.124496624,0.10940613,0.10940613,0.11317875,0.116951376,0.124496624,0.13958712,0.14335975,0.14335975,0.14335975,0.12826926,0.09808825,0.056589376,0.033953626,0.026408374,0.018863125,0.011317875,0.0150905,0.0150905,0.02263575,0.041498873,0.06413463,0.08677038,0.124496624,0.19240387,0.21881226,0.20372175,0.19994913,0.23390275,0.25276586,0.29049212,0.38103512,0.55457586,0.69793564,0.87902164,1.0487897,1.1204696,0.995973,0.91297525,0.9808825,1.1355602,1.2525115,1.1242423,0.80356914,0.6790725,0.69039035,0.73188925,0.6488915,0.62625575,0.58475685,0.513077,0.44139713,0.43007925,0.4074435,0.32067314,0.2565385,0.24522063,0.24522063,0.21503963,0.18485862,0.16976812,0.16222288,0.1358145,0.150905,0.1961765,0.211267,0.17731337,0.14713238,0.124496624,0.094315626,0.06413463,0.049044125,0.06790725,0.049044125,0.0452715,0.049044125,0.05281675,0.041498873,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05281675,0.1358145,0.15845025,0.8111144,1.841041,2.0145817,1.1619685,0.15467763,0.07922512,0.15467763,0.21881226,0.24522063,0.36594462,0.66020936,0.62625575,0.47535074,0.3734899,0.43385187,0.41498876,0.33576363,0.271629,0.2263575,0.11317875,0.090543,0.1358145,0.18485862,0.18863125,0.09808825,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.17731337,0.4979865,0.7884786,1.3807807,1.6524098,1.5203679,1.2487389,1.4449154,1.4713237,1.1657411,0.76207024,0.6073926,1.1619685,2.293756,4.063117,4.745962,4.0480266,3.078462,4.5988297,6.48137,6.541732,5.0138187,4.557331,3.4632697,3.3236825,3.31991,3.3312278,3.9574835,2.6144292,1.7165444,1.8448136,2.3088465,1.1506506,0.5998474,0.77338815,1.0487897,0.9997456,0.40367088,0.13204187,0.033953626,0.060362,0.13958712,0.15845025,0.10940613,0.1056335,2.9916916,5.934339,0.4074435,0.27540162,0.3961256,0.39989826,0.23390275,0.17354076,0.5319401,0.45648763,0.32067314,0.29049212,0.31312788,0.32444575,0.3772625,0.3734899,0.29049212,0.181086,0.55457586,0.935611,1.0374719,0.7809334,0.27917424,0.3470815,0.2565385,0.6828451,1.4524606,1.5430037,0.995973,0.77338815,0.91674787,1.1959221,1.0902886,1.4298248,2.1013522,2.5087957,2.9124665,4.425289,6.2663302,6.228604,5.2628117,4.644101,5.9984736,6.488915,5.6815734,4.8063245,4.3007927,3.8254418,3.9914372,4.8968673,5.194905,4.478106,3.240685,2.6408374,1.8485862,1.3430545,1.177059,0.97710985,1.4600059,1.4109617,1.3468271,1.50905,1.8599042,5.1345425,4.938366,6.006019,8.073418,5.873977,4.6214657,3.4972234,2.5427492,2.1881225,3.2218218,5.100589,3.9650288,2.1768045,1.0412445,0.80734175,0.90543,0.8337501,1.2034674,2.0108092,2.6672459,2.7351532,3.2784111,2.9841464,2.305074,3.470815,5.3910813,7.0284004,7.043491,5.96452,6.1720147,5.7494807,6.571913,5.96452,4.214022,4.5988297,7.0057645,8.959985,7.756517,4.6214657,4.719554,5.783434,4.0178456,3.0445085,5.372218,12.385528,20.77962,24.982323,26.981813,27.8797,27.864609,22.424482,17.493662,13.29473,10.386037,9.669238,17.761518,14.864142,9.771099,7.805561,10.785934,8.850578,6.8133607,5.323174,4.429062,3.5953116,2.214531,1.5958204,1.4600059,1.7618159,2.7011995,4.2102494,4.9232755,5.7419353,6.1078796,3.99521,6.319147,11.744182,13.283413,10.193633,7.967784,8.145098,8.869441,10.79348,11.853588,7.303802,3.1124156,1.9429018,4.429062,10.54826,19.60256,11.974312,13.970031,16.980585,15.705438,8.156415,9.435335,12.377983,11.91395,9.457971,12.898605,13.494679,10.152134,7.865923,7.726336,6.9152217,6.809588,8.492179,9.084481,7.0849895,2.372981,8.367682,16.912678,17.463482,12.057309,15.32063,16.214743,10.585986,7.33021,8.854351,11.087745,11.012292,22.854563,29.849009,25.574625,13.973803,18.900852,30.098001,40.336906,50.051414,67.36399,75.0941,66.63965,50.062733,33.297188,24.125937,16.72782,13.807808,13.422999,13.347548,11.0613365,12.31762,15.513034,18.218006,20.036411,22.60557,23.910898,25.10682,26.796955,28.464457,28.502182,27.027086,23.503454,15.75071,7.0774446,6.2663302,6.560595,6.228604,5.43258,4.074435,1.7919968,1.267602,0.8639311,0.5772116,0.3961256,0.32067314,0.14713238,0.15467763,0.29803738,0.452715,0.422534,0.23013012,0.124496624,0.120724,0.20372175,0.34330887,0.965792,1.4826416,2.191895,2.8898308,2.8558772,2.4484336,1.6410918,1.177059,1.3355093,1.9202662,1.4071891,1.2713746,1.7731338,2.4522061,2.1277604,2.0258996,2.3616633,2.3654358,1.9994912,1.9504471,2.305074,2.7615614,2.6672459,2.0070364,1.4222796,1.478869,1.5958204,1.7089992,1.6561824,1.1846043,0.8186596,0.62625575,0.47912338,0.36971724,0.40367088,0.5093044,0.38103512,0.20372175,0.08299775,0.071679875,0.10940613,0.181086,0.23767537,0.24899325,0.20372175,0.22258487,0.271629,0.38480774,0.48666862,0.392353,0.2263575,0.21503963,0.19240387,0.1056335,0.00754525,0.0,0.0150905,0.018863125,0.018863125,0.03772625,0.026408374,0.011317875,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.049044125,0.08677038,0.120724,0.11317875,0.0754525,0.03772625,0.06413463,0.06413463,0.0452715,0.03772625,0.06413463,0.026408374,0.00754525,0.011317875,0.03772625,0.08677038,0.018863125,0.0,0.00754525,0.033953626,0.1056335,0.056589376,0.03772625,0.03772625,0.056589376,0.10940613,0.094315626,0.116951376,0.14713238,0.14713238,0.09808825,0.0452715,0.018863125,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.011317875,0.0150905,0.033953626,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.011317875,0.0,0.0,0.00754525,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.011317875,0.0150905,0.0150905,0.0150905,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.02263575,0.033953626,0.10186087,0.16976812,0.15845025,0.12826926,0.10940613,0.094315626,0.10186087,0.12826926,0.23767537,0.3772625,0.3772625,0.29803738,0.27917424,0.2678564,0.24522063,0.20372175,0.23767537,0.25276586,0.2678564,0.29049212,0.3055826,0.28294688,0.24899325,0.26408374,0.30935526,0.29426476,0.26031113,0.30181,0.30181,0.23767537,0.19240387,0.16222288,0.116951376,0.0754525,0.060362,0.08677038,0.15845025,0.21881226,0.26408374,0.3055826,0.3734899,0.362172,0.33953625,0.31312788,0.29049212,0.31312788,0.29049212,0.27540162,0.23013012,0.15467763,0.08677038,0.0754525,0.06790725,0.071679875,0.08299775,0.07922512,0.090543,0.08677038,0.09808825,0.12826926,0.1358145,0.1056335,0.0754525,0.060362,0.056589376,0.041498873,0.033953626,0.02263575,0.011317875,0.00754525,0.018863125,0.0150905,0.02263575,0.026408374,0.026408374,0.030181,0.056589376,0.1056335,0.14335975,0.17354076,0.2263575,0.26408374,0.20372175,0.17731337,0.25276586,0.42630664,0.5772116,0.73188925,0.90920264,1.0374719,0.95824677,0.90543,0.9507015,1.1204696,1.2638294,1.0751982,0.77716076,0.694163,0.6752999,0.6488915,0.6375736,0.68661773,0.65643674,0.5696664,0.49421388,0.543258,0.5394854,0.452715,0.3772625,0.331991,0.27917424,0.23013012,0.211267,0.1961765,0.16976812,0.13958712,0.15467763,0.211267,0.24899325,0.241448,0.19994913,0.1659955,0.116951376,0.0754525,0.056589376,0.0754525,0.05281675,0.06413463,0.090543,0.1056335,0.0754525,0.1659955,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.1358145,0.3055826,1.267602,2.3993895,2.595566,1.6561824,0.29049212,0.056589376,0.10940613,0.16976812,0.120724,0.0,0.14713238,0.23013012,0.19240387,0.116951376,0.21503963,0.60362,0.4074435,0.24522063,0.271629,0.19994913,0.1358145,0.11317875,0.094315626,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.3961256,0.7884786,0.33576363,0.12826926,0.1056335,0.12826926,0.12826926,0.090543,0.21503963,0.5093044,0.814887,1.0148361,1.0525624,3.3463185,3.4255435,2.4559789,1.5882751,1.9693103,2.1013522,2.9049213,3.3689542,3.361409,3.6179473,2.9313297,2.1956677,1.7240896,2.052308,3.9197574,3.651901,2.2748928,2.203213,3.0558262,1.6637276,0.80734175,0.5017591,0.392353,0.3169005,0.3055826,0.120724,0.030181,0.0,0.0,0.0,0.0,0.0,0.6149379,1.3505998,0.58098423,0.70170826,0.5017591,0.29426476,0.211267,0.19994913,0.18485862,0.19240387,0.181086,0.13958712,0.090543,0.19994913,0.4376245,0.47535074,0.29049212,0.1659955,0.19240387,0.34330887,0.32067314,0.13204187,0.1056335,0.056589376,0.026408374,0.1358145,0.4074435,0.76207024,0.7130261,0.4074435,0.7696155,1.750498,2.335255,2.04099,3.1312788,3.5764484,3.802806,6.6813188,6.270103,5.80607,5.6061206,6.5002327,9.857869,9.869187,8.039464,6.881268,6.741681,5.8136153,4.3611546,4.640329,5.3344917,5.3646727,3.874486,2.8256962,2.5087957,2.0070364,1.1959221,0.73188925,1.0487897,1.5241405,2.0787163,2.372981,1.7995421,6.9755836,4.9647746,5.20245,8.914713,9.110889,4.3121104,4.3196554,5.372218,5.7872066,5.9796104,10.0465,10.906659,7.6848373,2.7879698,1.9089483,2.6898816,2.2598023,1.5769572,1.4713237,2.655928,2.263575,2.1579416,1.8523588,1.5430037,2.0900342,4.274384,5.251494,5.9494295,6.515323,6.3342376,6.5530496,4.9949555,3.3425457,3.0369632,5.292993,6.541732,5.7079816,4.7836885,5.6476197,10.038955,10.137043,6.40969,3.893349,5.1458607,10.223814,21.19838,22.14531,18.87067,16.98813,21.941587,28.449366,23.68454,16.693865,12.208215,10.63503,19.791191,18.674494,14.268067,11.136789,11.442371,7.3415284,5.172269,4.3800178,3.731126,1.3128735,0.995973,1.2826926,2.0636258,2.8596497,2.8219235,2.214531,3.187868,5.040227,5.934339,2.8822856,3.9084394,5.723072,6.1908774,5.587258,6.5756855,9.163706,8.246958,8.722309,9.159933,1.7844516,2.3578906,3.289729,5.451443,8.114917,8.956212,9.201432,11.012292,11.268831,9.220296,6.485142,8.145098,10.601076,11.072655,9.918231,10.650121,12.811834,13.140053,12.15917,9.7220545,5.036454,4.90064,5.975838,6.56814,5.7570257,3.3878171,6.598321,7.884786,8.605357,10.253995,14.464244,9.914458,5.50426,5.406172,8.975075,10.7557535,11.306557,26.887499,33.48582,25.997158,18.233097,28.705904,43.155056,49.27048,48.150013,54.291847,57.623074,51.647236,39.601246,26.54419,19.319613,11.140562,10.174769,13.385274,16.014793,11.59705,16.87118,19.87419,20.036411,19.606333,23.620405,26.770548,29.241617,30.675215,30.403585,27.44962,22.19058,18.16519,12.781653,7.24344,6.5455046,6.752999,6.428553,6.477597,6.0286546,2.425798,1.5241405,1.1053791,0.7092535,0.28294688,0.19994913,0.16222288,0.2263575,0.5017591,0.77716076,0.5357128,0.241448,0.11317875,0.11317875,0.15845025,0.120724,0.41498876,1.780679,3.2255943,4.3347464,5.247721,4.432834,2.897376,1.6788181,1.2487389,1.5430037,0.9318384,0.73188925,1.3619176,2.3578906,2.3956168,1.6033657,1.961765,2.516341,2.7804246,2.7313805,3.5236318,4.1083884,4.0706625,3.410453,2.5314314,2.323937,2.0183544,1.780679,1.5618668,1.0978339,0.9393836,0.7167987,0.422534,0.16976812,0.18485862,0.513077,0.45648763,0.2678564,0.1056335,0.0452715,0.0452715,0.06413463,0.13204187,0.21503963,0.23013012,0.21503963,0.26031113,0.33953625,0.41876137,0.44139713,0.34330887,0.23767537,0.150905,0.090543,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.030181,0.041498873,0.0754525,0.041498873,0.011317875,0.02263575,0.071679875,0.120724,0.02263575,0.00754525,0.02263575,0.041498873,0.090543,0.090543,0.06413463,0.06413463,0.120724,0.24522063,0.21881226,0.1961765,0.23767537,0.3169005,0.3055826,0.14713238,0.060362,0.02263575,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.1056335,0.0452715,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.0754525,0.08677038,0.12826926,0.16976812,0.181086,0.1056335,0.094315626,0.17354076,0.27917424,0.34330887,0.3055826,0.29426476,0.25276586,0.26031113,0.31312788,0.35085413,0.46026024,0.452715,0.392353,0.34330887,0.36594462,0.452715,0.3734899,0.3169005,0.34330887,0.38103512,0.392353,0.51684964,0.51684964,0.35085413,0.1659955,0.120724,0.08677038,0.08299775,0.10186087,0.1358145,0.150905,0.181086,0.211267,0.241448,0.29049212,0.41121614,0.47157812,0.452715,0.38480774,0.33576363,0.27540162,0.22258487,0.1659955,0.11317875,0.0754525,0.05281675,0.03772625,0.03772625,0.041498873,0.030181,0.030181,0.041498873,0.056589376,0.0754525,0.0754525,0.06413463,0.060362,0.060362,0.056589376,0.030181,0.030181,0.030181,0.02263575,0.018863125,0.030181,0.018863125,0.00754525,0.00754525,0.018863125,0.030181,0.06790725,0.094315626,0.120724,0.13958712,0.150905,0.150905,0.124496624,0.120724,0.15845025,0.24522063,0.4640329,0.77338815,0.9280658,0.8978847,0.8865669,0.8601585,0.8262049,0.9318384,1.1242423,1.1581959,0.8526133,0.694163,0.6111652,0.5772116,0.62625575,0.6752999,0.73188925,0.7130261,0.6526641,0.70170826,0.6790725,0.58098423,0.48666862,0.4376245,0.41121614,0.32821837,0.2678564,0.23013012,0.19994913,0.150905,0.17731337,0.21881226,0.23767537,0.23390275,0.26031113,0.24899325,0.181086,0.11317875,0.0754525,0.0754525,0.06413463,0.09808825,0.150905,0.18485862,0.1358145,0.056589376,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.1358145,0.52439487,0.935611,1.2336484,1.3807807,1.448688,0.875249,0.36594462,0.10186087,0.05281675,0.0,0.030181,0.0452715,0.03772625,0.02263575,0.041498873,0.120724,0.08299775,0.049044125,0.05281675,0.041498873,0.026408374,0.08299775,0.07922512,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.10940613,0.19240387,0.1056335,0.06413463,0.10186087,0.33576363,0.5470306,0.17731337,0.24899325,0.84884065,1.2411937,1.1619685,0.80734175,1.3355093,1.7655885,1.8938577,1.720317,1.4562333,2.7615614,7.798016,8.401636,4.666737,4.9345937,11.77059,9.359882,4.4441524,1.8485862,4.459243,3.651901,2.3918443,1.3920987,0.83752275,0.38103512,0.21881226,0.13958712,0.094315626,0.06413463,0.060362,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.10186087,1.0412445,1.9466745,0.3470815,0.18863125,0.10186087,0.10186087,0.12826926,0.041498873,0.03772625,0.03772625,0.1056335,0.20749438,0.23767537,0.3169005,0.32821837,0.23390275,0.124496624,0.21503963,0.41498876,0.3772625,0.27540162,0.21503963,0.241448,0.11317875,0.041498873,0.10940613,0.35839936,0.8111144,1.2600567,1.0223814,1.6222287,2.7351532,2.1881225,2.071171,2.9766011,3.6707642,4.689373,8.345046,6.1908774,5.983383,7.5112963,9.718282,10.710483,10.93684,9.442881,7.8244243,6.79827,6.205968,4.5950575,4.9647746,6.187105,6.9189944,5.583485,4.3686996,4.183841,3.942393,3.240685,2.354118,1.7844516,2.04099,2.806833,3.3915899,2.727608,4.6214657,3.4632697,3.338773,5.409944,7.888559,4.7421894,4.327201,4.508287,4.2102494,3.429316,5.824933,10.0465,9.303293,5.040227,6.9227667,5.753253,3.2633207,1.4449154,1.4600059,3.6179473,3.0709167,2.1956677,1.7278622,2.4823873,5.323174,4.715781,4.8855495,4.8553686,5.010046,7.115171,8.084735,6.066381,4.323428,4.6516466,7.3679366,6.428553,4.3800178,3.8292143,5.5457587,8.465771,8.526133,7.405663,5.847569,5.383536,8.345046,14.151116,15.803526,13.702174,11.593277,16.558052,21.817091,23.307278,20.655123,14.852824,8.265821,17.569115,14.803781,9.42779,6.4210076,6.319147,4.919503,4.8930945,5.2665844,4.9345937,2.655928,1.9957186,2.3088465,2.9426475,3.3764994,3.2142766,3.7160356,4.644101,6.360646,7.062354,2.7992878,4.6931453,7.3679366,8.424272,8.805306,12.800517,15.086727,13.441863,10.084227,6.820906,5.032682,12.577931,15.807299,14.434063,9.612649,3.953711,8.669493,10.001229,8.737399,6.2927384,4.689373,9.348565,9.81637,8.952439,9.469289,13.920986,14.2944765,15.878979,15.671484,12.830698,8.661947,5.040227,6.8699503,8.428044,8.0206,7.9753294,14.596286,16.075155,13.690856,9.488152,6.2889657,5.934339,5.938112,7.2170315,9.156161,9.608876,15.207452,24.412657,28.038149,27.19308,33.28587,48.825314,69.929375,87.74371,93.70446,79.53448,57.494804,45.279045,36.164383,27.434528,20.353312,13.690856,14.143571,15.663939,15.120681,12.291212,18.72731,21.537916,22.42071,24.823872,33.94608,31.531599,31.358059,32.45212,32.142765,26.08393,19.727057,13.826671,8.956212,6.33801,7.828197,6.1229706,7.375482,6.900131,4.074435,2.3767538,1.8561316,1.4600059,0.86770374,0.241448,0.23390275,0.23767537,0.38480774,0.58475685,0.7696155,0.875249,0.513077,0.24522063,0.094315626,0.0452715,0.03772625,0.17354076,0.70170826,1.448688,2.3013012,3.199186,5.311856,5.1760416,3.9725742,2.7615614,2.516341,2.052308,1.6146835,1.7995421,2.4333432,2.5804756,1.7655885,2.1805773,3.361409,4.2291126,3.0860074,3.9386206,4.727099,4.768598,4.3121104,4.534695,4.08198,3.127506,2.5238862,2.3201644,1.7580433,1.7052265,1.1581959,0.543258,0.1358145,0.060362,0.14713238,0.13204187,0.08677038,0.041498873,0.02263575,0.011317875,0.018863125,0.049044125,0.10940613,0.23013012,0.27540162,0.28294688,0.32821837,0.41121614,0.45648763,0.47535074,0.331991,0.18863125,0.10186087,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.026408374,0.011317875,0.003772625,0.003772625,0.0150905,0.02263575,0.0150905,0.00754525,0.00754525,0.026408374,0.056589376,0.08299775,0.08677038,0.08299775,0.09808825,0.16976812,0.12826926,0.11317875,0.1358145,0.18485862,0.23013012,0.11317875,0.03772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.00754525,0.003772625,0.011317875,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.026408374,0.041498873,0.06413463,0.09808825,0.124496624,0.13204187,0.14713238,0.17731337,0.20749438,0.241448,0.29426476,0.35085413,0.35462674,0.38480774,0.4640329,0.5696664,0.41498876,0.38480774,0.40367088,0.41876137,0.41498876,0.3734899,0.35839936,0.362172,0.40367088,0.5281675,0.40367088,0.331991,0.32067314,0.35839936,0.39989826,0.271629,0.22258487,0.181086,0.150905,0.19994913,0.23013012,0.2565385,0.331991,0.40367088,0.32821837,0.38103512,0.44139713,0.452715,0.422534,0.422534,0.47912338,0.47535074,0.4074435,0.27917424,0.124496624,0.060362,0.030181,0.02263575,0.033953626,0.030181,0.030181,0.041498873,0.049044125,0.05281675,0.06413463,0.041498873,0.0452715,0.0452715,0.033953626,0.030181,0.02263575,0.026408374,0.030181,0.026408374,0.018863125,0.026408374,0.018863125,0.0150905,0.0150905,0.018863125,0.026408374,0.03772625,0.056589376,0.090543,0.150905,0.16222288,0.1659955,0.15467763,0.1358145,0.1358145,0.2565385,0.4640329,0.6451189,0.8224323,1.1544232,1.0223814,0.8299775,0.72811663,0.72811663,0.694163,0.5281675,0.513077,0.52062225,0.5017591,0.49044126,0.6375736,0.6752999,0.663982,0.66020936,0.7394345,0.7432071,0.66775465,0.56212115,0.4678055,0.422534,0.4074435,0.3961256,0.35085413,0.27917424,0.24899325,0.21503963,0.19240387,0.18863125,0.19240387,0.19994913,0.20749438,0.22258487,0.241448,0.24899325,0.24899325,0.23390275,0.20372175,0.181086,0.18485862,0.22258487,0.011317875,0.003772625,0.0,0.0,0.011317875,0.056589376,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.1358145,0.23013012,0.58098423,1.1393328,1.539231,0.90920264,0.42630664,0.17731337,0.116951376,0.06413463,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.090543,0.124496624,0.08299775,0.08299775,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06790725,0.3470815,0.22258487,0.1056335,0.05281675,0.056589376,0.06413463,0.049044125,0.06790725,0.2263575,0.4376245,0.41876137,0.62625575,1.0450171,1.1846043,1.026154,1.0148361,1.1996948,1.8070874,2.0145817,1.6939086,1.4298248,2.7200627,9.144843,9.442881,3.663219,3.138824,12.185578,10.574668,5.1760416,1.327964,2.8709676,2.5238862,2.0296721,1.2261031,0.3734899,0.116951376,0.06413463,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05281675,0.46026024,0.87147635,0.27917424,0.2263575,0.19994913,0.16976812,0.10940613,0.0,0.0,0.026408374,0.08299775,0.15845025,0.23013012,0.573439,0.49044126,0.35085413,0.362172,0.56589377,0.6375736,0.331991,0.16222288,0.2867195,0.52062225,0.27917424,0.10940613,0.241448,0.7809334,1.7014539,2.1315331,2.0560806,2.1768045,2.3654358,1.6675003,1.9957186,2.9200118,3.519859,4.7044635,9.208978,6.507778,6.722818,9.288202,12.411936,13.075918,10.653893,8.186596,6.330465,5.4740787,5.7419353,4.08198,3.5274043,4.821415,6.673774,5.7381625,4.606375,4.7874613,4.587512,3.572676,2.5616124,1.599593,2.5729303,3.8895764,4.4177437,3.500996,4.002755,3.2746384,3.3425457,4.7233267,6.4210076,3.8707132,3.7575345,3.8782585,3.4859054,3.2859564,4.2328854,6.7114997,6.85486,5.13077,6.375736,7.7338815,5.081726,2.263575,1.5618668,3.6971724,3.2331395,2.335255,1.9768555,2.5616124,3.9273026,5.089271,4.9157305,4.3611546,4.534695,6.696409,9.042982,7.7904706,7.1793056,9.012801,12.657157,10.231359,6.983129,7.0510364,10.495442,13.27964,10.401127,6.488915,3.893349,4.4705606,9.593785,11.766817,11.480098,9.906913,10.502988,19.002712,42.951336,34.45161,19.583696,11.046246,8.160188,13.487134,12.596795,9.544742,7.118943,6.828451,8.650629,8.582722,7.2887115,5.1873593,2.4597516,1.9429018,2.5427492,3.4029078,4.5535583,6.888813,7.6282477,9.156161,10.401127,9.646602,4.515832,5.6853456,9.510788,10.502988,9.74469,14.916959,17.455936,17.040947,11.902632,5.783434,7.911195,16.15438,18.206688,13.675766,5.8928404,1.8938577,8.307321,10.4049,8.91094,5.9720654,5.1647234,11.136789,11.393328,9.533423,9.903141,17.57666,16.18456,15.47908,14.298248,12.00072,8.458225,9.0807085,12.2270775,12.064855,8.993938,9.654147,17.610613,18.463226,14.268067,8.269594,4.8930945,9.235386,9.544742,8.341274,7.3981175,7.748972,21.794455,40.74435,46.09016,41.00466,50.36077,62.76139,79.50807,93.21024,94.915474,74.15472,51.647236,44.169895,39.789875,32.41062,21.78691,19.108345,19.398838,19.813826,19.334703,18.772581,23.661903,24.054256,25.163408,29.479292,36.768,33.1991,32.9652,34.312023,34.108303,27.875927,19.281887,12.559069,7.3868,4.798779,7.1604424,6.6813188,8.182823,6.9265394,3.1765501,2.1805773,2.0975795,1.6410918,0.935611,0.28294688,0.16976812,0.2565385,0.36594462,0.49044126,0.66020936,0.94315624,0.69793564,0.7167987,0.513077,0.20749438,0.5470306,1.7731338,1.2185578,0.69793564,0.9016574,1.4034165,2.7540162,3.3010468,3.6292653,3.8141239,3.4217708,2.8634224,2.1956677,2.1881225,2.7200627,2.7804246,1.8297231,2.1805773,3.259548,4.123479,3.440634,3.9461658,4.7912335,4.9534564,4.5761943,4.9534564,4.8742313,4.1536603,3.3915899,2.806833,2.2447119,1.7882242,0.9997456,0.3734899,0.094315626,0.049044125,0.0452715,0.033953626,0.02263575,0.011317875,0.00754525,0.0,0.00754525,0.02263575,0.056589376,0.12826926,0.181086,0.23767537,0.28294688,0.31312788,0.3470815,0.35462674,0.2678564,0.16976812,0.09808825,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.033953626,0.041498873,0.018863125,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.00754525,0.018863125,0.049044125,0.09808825,0.1056335,0.071679875,0.08677038,0.05281675,0.05281675,0.06413463,0.08299775,0.094315626,0.041498873,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.00754525,0.011317875,0.030181,0.056589376,0.08677038,0.120724,0.18863125,0.19240387,0.17731337,0.181086,0.21503963,0.24522063,0.30181,0.36594462,0.422534,0.47157812,0.41876137,0.38480774,0.43007925,0.52062225,0.5357128,0.543258,0.4640329,0.3961256,0.3961256,0.482896,0.3961256,0.35839936,0.3734899,0.41121614,0.422534,0.3055826,0.23013012,0.20372175,0.20372175,0.1961765,0.18863125,0.19994913,0.27540162,0.3961256,0.44516975,0.4376245,0.44894236,0.47157812,0.5055317,0.52439487,0.51684964,0.44894236,0.35085413,0.23767537,0.120724,0.060362,0.026408374,0.018863125,0.02263575,0.02263575,0.030181,0.030181,0.026408374,0.030181,0.041498873,0.041498873,0.033953626,0.033953626,0.041498873,0.049044125,0.0452715,0.041498873,0.041498873,0.03772625,0.02263575,0.030181,0.02263575,0.0150905,0.0150905,0.0150905,0.0150905,0.018863125,0.030181,0.049044125,0.07922512,0.09808825,0.1056335,0.120724,0.1358145,0.1358145,0.20372175,0.30935526,0.43385187,0.59607476,0.8639311,0.87902164,0.77338815,0.7167987,0.7130261,0.6073926,0.4376245,0.422534,0.4678055,0.52062225,0.56589377,0.694163,0.73188925,0.7167987,0.67152727,0.6111652,0.66775465,0.67152727,0.6073926,0.5017591,0.45648763,0.46026024,0.4678055,0.44139713,0.41498876,0.48666862,0.4074435,0.35839936,0.34330887,0.35085413,0.35839936,0.29426476,0.35085413,0.43007925,0.49044126,0.52062225,0.5281675,0.4376245,0.32067314,0.23767537,0.21503963,0.08677038,0.030181,0.00754525,0.0,0.011317875,0.056589376,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.23767537,0.663982,0.9393836,0.49421388,0.25276586,0.14335975,0.10186087,0.06413463,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.10186087,0.10940613,0.124496624,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.094315626,0.40367088,0.27540162,0.124496624,0.041498873,0.05281675,0.120724,0.056589376,0.033953626,0.08677038,0.24522063,0.5357128,0.79602385,0.965792,0.97710985,1.0186088,1.5316857,1.7542707,2.5729303,2.4559789,1.4071891,0.9393836,2.0070364,6.960493,7.0057645,2.1692593,1.2864652,9.265567,8.786444,4.727099,1.2449663,1.7354075,1.569412,1.4449154,1.056335,0.49421388,0.23767537,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041498873,0.20749438,0.29803738,0.35839936,0.36594462,0.29049212,0.09808825,0.06790725,0.21881226,0.21881226,0.124496624,0.41121614,0.87902164,0.7507524,0.6526641,0.7809334,0.87147635,0.6526641,0.23767537,0.10940613,0.36971724,0.76584285,0.5583485,0.42630664,0.56589377,1.1393328,2.3088465,2.7917426,3.270866,3.0256453,2.214531,1.8674494,1.9278114,2.9426475,3.5349495,4.7572803,10.061591,7.5829763,7.152897,9.574923,13.030646,13.072145,8.567632,6.688864,5.7306175,5.0025005,4.8100967,3.6028569,2.9237845,4.2706113,6.3644185,5.168496,4.45547,4.447925,4.085753,3.2142766,2.6144292,1.9202662,2.6898816,3.5839937,4.032936,4.2328854,4.8742313,4.055572,3.8669407,5.5193505,9.344792,7.175533,5.987156,5.5570765,6.043745,7.9753294,6.477597,6.1229706,5.485397,4.357382,3.712263,6.1418333,4.617693,2.3956168,1.7391801,3.8971217,3.6556737,3.0407357,2.6785638,2.674791,2.5917933,6.1078796,4.98741,3.9801195,5.2099953,8.171506,8.43559,7.786698,8.518587,10.812344,12.721292,9.454198,6.7114997,7.3981175,10.627484,11.714001,8.379,4.696918,2.9954643,4.727099,10.431308,10.099318,8.729855,8.899622,11.544232,15.9695215,45.33941,31.780594,13.932304,7.8696957,7.1038527,8.201687,10.691619,10.967021,8.643084,6.560595,9.242931,9.061845,6.960493,4.085753,1.780679,1.81086,2.7917426,4.2291126,6.5530496,11.114153,13.45318,14.4152,13.238141,9.937095,5.2854476,5.7607985,9.891823,11.476325,11.012292,15.724301,17.550251,15.743164,11.208468,7.484888,10.7557535,12.811834,13.483362,10.242677,4.478106,1.5052774,6.8435416,10.148361,9.5183325,6.462507,5.885295,10.963248,10.355856,9.0957985,11.46878,20.98334,19.319613,14.8339615,11.34051,10.054046,9.574923,13.404137,16.29774,14.015302,8.597813,8.386545,15.286676,15.120681,10.982111,6.590776,6.3153744,13.370183,13.166461,10.178542,8.82417,13.460726,38.118603,62.93493,65.70404,52.53003,57.838116,64.040306,72.076004,78.3876,77.45953,61.806915,46.716415,43.094696,40.778305,34.583652,24.299479,26.00093,26.012249,25.71044,25.89907,26.812046,28.702131,28.766266,30.245134,33.10856,34.093212,32.055996,32.55398,32.301216,29.581152,24.254206,17.255987,11.378237,6.651138,4.1498876,6.017337,7.1038527,7.8319697,6.039973,2.6710186,1.8033148,1.9051756,1.4335974,0.8111144,0.34330887,0.19994913,0.27540162,0.30181,0.43385187,0.66775465,0.8563859,0.7884786,0.97333723,0.77338815,0.32821837,0.55080324,1.7618159,1.0789708,0.30935526,0.18863125,0.35462674,0.6073926,1.1506506,2.2371666,3.5462675,4.2064767,3.7613072,2.957738,2.7200627,3.0218725,2.8709676,1.961765,2.0598533,2.584248,2.9916916,2.7879698,3.1312788,3.9310753,4.346064,4.4101987,5.0439997,5.149633,4.90064,4.29702,3.4217708,2.41448,1.3920987,0.6149379,0.20749438,0.13204187,0.150905,0.09808825,0.041498873,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.03772625,0.071679875,0.14335975,0.18863125,0.1961765,0.21881226,0.211267,0.19240387,0.16222288,0.11317875,0.049044125,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.003772625,0.003772625,0.02263575,0.08677038,0.13204187,0.06790725,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.071679875,0.08677038,0.05281675,0.0452715,0.026408374,0.06790725,0.12826926,0.15467763,0.0754525,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.018863125,0.030181,0.05281675,0.08677038,0.1961765,0.18863125,0.1659955,0.1659955,0.1659955,0.1659955,0.24899325,0.32821837,0.36594462,0.392353,0.44516975,0.39989826,0.41876137,0.52062225,0.59230214,0.6149379,0.56589377,0.513077,0.5055317,0.58098423,0.4640329,0.44516975,0.452715,0.42630664,0.3169005,0.2678564,0.24522063,0.2565385,0.2867195,0.2565385,0.24522063,0.241448,0.28294688,0.362172,0.4640329,0.48666862,0.47535074,0.4979865,0.55080324,0.58098423,0.4979865,0.4074435,0.3169005,0.23013012,0.15467763,0.08299775,0.033953626,0.0150905,0.0150905,0.0150905,0.02263575,0.018863125,0.018863125,0.030181,0.049044125,0.03772625,0.02263575,0.026408374,0.041498873,0.049044125,0.05281675,0.0452715,0.041498873,0.041498873,0.041498873,0.033953626,0.026408374,0.02263575,0.02263575,0.02263575,0.0150905,0.0150905,0.018863125,0.02263575,0.02263575,0.049044125,0.060362,0.08299775,0.11317875,0.120724,0.16222288,0.20749438,0.27540162,0.3734899,0.51684964,0.59607476,0.60362,0.6451189,0.7092535,0.62625575,0.513077,0.44139713,0.422534,0.46026024,0.56589377,0.66020936,0.663982,0.6451189,0.6073926,0.482896,0.543258,0.62248313,0.63002837,0.58475685,0.5885295,0.5470306,0.5055317,0.47157812,0.47535074,0.5696664,0.5281675,0.48666862,0.47157812,0.482896,0.51684964,0.482896,0.5319401,0.573439,0.59230214,0.6413463,0.7432071,0.65643674,0.5093044,0.38103512,0.31312788,0.23013012,0.0754525,0.0150905,0.0,0.0,0.0,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06790725,0.10186087,0.06413463,0.0,0.0,0.0,0.030181,0.1056335,0.23390275,0.09808825,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.056589376,0.08677038,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.06790725,0.18863125,0.3055826,0.19240387,0.06413463,0.041498873,0.150905,0.05281675,0.03772625,0.094315626,0.241448,0.5055317,0.7809334,0.7884786,0.95824677,1.5505489,2.6408374,2.505023,3.0256453,2.5502944,1.0412445,0.090543,0.935611,2.9086938,2.9200118,1.0789708,0.7092535,6.085244,5.9230213,3.470815,1.3392819,1.5241405,1.1091517,0.814887,0.62625575,0.49421388,0.3470815,0.116951376,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.08677038,0.19240387,0.31312788,0.44139713,0.4678055,0.1961765,0.1358145,0.43385187,0.4376245,0.26031113,0.784706,1.0336993,0.90920264,0.8903395,1.0110635,0.87902164,0.48666862,0.26031113,0.271629,0.5017591,0.87147635,0.77716076,1.0336993,1.2525115,1.4750963,2.1390784,2.9766011,4.063117,3.893349,2.7502437,2.7238352,2.11267,3.1048703,3.7914882,5.1156793,10.868933,8.843033,7.183078,8.59404,11.631002,10.687846,5.9305663,5.938112,6.4964604,5.726845,4.074435,3.8480775,4.1272516,5.4740787,6.598321,4.349837,4.1197066,3.5236318,2.9652832,2.6483827,2.5880208,2.535204,2.323937,2.1390784,2.6106565,4.821415,6.485142,5.3194013,4.4516973,6.8397694,15.260268,12.721292,9.578695,8.620448,10.423763,13.355092,9.329701,7.6886096,6.119198,3.9008942,1.9089483,2.8332415,2.704972,2.082489,2.1353056,4.6629643,4.485651,4.1574326,3.6368105,3.0860074,2.8747404,6.651138,4.983638,4.466788,7.0963078,10.269085,6.462507,6.1720147,7.7187905,8.99771,7.496206,4.515832,3.8254418,4.7535076,5.6287565,3.783943,3.180323,3.5538127,4.504514,6.19465,9.337247,7.9262853,8.145098,10.691619,12.536433,6.900131,21.794455,14.543469,8.16396,8.635539,4.919503,3.4368613,8.273367,11.415963,9.669238,4.640329,5.6287565,5.753253,4.5950575,2.6898816,1.5354583,2.0145817,3.0520537,4.870459,7.9791017,13.177779,17.780382,16.188334,11.736636,7.1604424,4.5799665,4.9119577,8.503497,11.7026825,13.558814,15.82239,14.766054,9.922004,8.224322,10.578441,11.864905,6.066381,7.0359454,8.66572,7.375482,2.1315331,5.032682,9.246704,9.963503,7.224577,5.9230213,8.888305,7.069899,7.5301595,12.996693,21.866135,20.417446,13.4644985,8.616675,8.627994,11.404645,14.264296,15.773345,12.849561,7.383027,6.25124,10.997202,10.495442,7.726336,5.802297,7.9715567,14.683057,14.634012,12.755245,14.569878,26.1707,56.49506,75.19596,70.46132,52.26972,52.394215,54.32203,55.182186,57.177906,58.49832,53.33737,43.521004,40.031322,37.669662,33.693314,27.815563,32.029587,32.26349,31.376923,31.097748,32.014496,31.633461,34.632698,37.299942,36.469967,29.524563,29.569836,30.592216,27.789156,21.696367,18.176508,15.207452,10.431308,6.436098,4.610148,5.1345425,7.3717093,6.983129,4.7346444,2.1013522,1.2864652,1.3091009,0.90920264,0.5470306,0.3961256,0.36594462,0.4678055,0.3961256,0.52062225,0.77338815,0.6790725,0.754525,0.84129536,0.6828451,0.32067314,0.0754525,0.08677038,0.06413463,0.030181,0.011317875,0.05281675,0.15845025,0.33953625,0.9242931,2.1805773,4.304565,4.52715,3.8292143,3.361409,3.361409,3.138824,2.4672968,2.0862615,1.8334957,1.6071383,1.3619176,1.8184053,2.6144292,3.3878171,4.142342,5.2628117,5.3684454,5.383536,5.0213637,4.032936,2.214531,0.86770374,0.30935526,0.17731337,0.22258487,0.27917424,0.18485862,0.06790725,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.041498873,0.071679875,0.094315626,0.116951376,0.12826926,0.150905,0.15845025,0.1358145,0.08299775,0.033953626,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0452715,0.03772625,0.02263575,0.0150905,0.0452715,0.150905,0.24899325,0.15845025,0.056589376,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.03772625,0.03772625,0.03772625,0.030181,0.11317875,0.23767537,0.31312788,0.18485862,0.071679875,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.011317875,0.026408374,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.0150905,0.0150905,0.0150905,0.026408374,0.06413463,0.1659955,0.15845025,0.14713238,0.1659955,0.15467763,0.16222288,0.241448,0.31312788,0.35839936,0.41121614,0.45648763,0.3961256,0.3772625,0.4376245,0.52439487,0.5093044,0.5772116,0.633801,0.69039035,0.845068,0.63002837,0.5281675,0.46026024,0.36971724,0.20372175,0.24522063,0.29049212,0.32067314,0.32821837,0.34330887,0.38480774,0.38858038,0.38480774,0.38103512,0.35839936,0.4640329,0.5093044,0.52062225,0.5319401,0.5696664,0.48666862,0.44139713,0.3772625,0.27917424,0.20372175,0.10940613,0.0452715,0.018863125,0.0150905,0.0150905,0.011317875,0.0150905,0.026408374,0.049044125,0.06790725,0.026408374,0.0150905,0.018863125,0.026408374,0.030181,0.041498873,0.03772625,0.033953626,0.03772625,0.056589376,0.03772625,0.033953626,0.033953626,0.033953626,0.026408374,0.018863125,0.0150905,0.0150905,0.0150905,0.011317875,0.030181,0.049044125,0.06413463,0.07922512,0.08677038,0.10940613,0.14335975,0.18485862,0.24522063,0.32821837,0.33953625,0.38103512,0.46026024,0.543258,0.5583485,0.5772116,0.49044126,0.38103512,0.3470815,0.48666862,0.5470306,0.47912338,0.452715,0.47912338,0.422534,0.44516975,0.52062225,0.58098423,0.62625575,0.7205714,0.6413463,0.52062225,0.44894236,0.44894236,0.46026024,0.48666862,0.482896,0.49044126,0.52439487,0.5583485,0.62625575,0.65643674,0.6187105,0.56212115,0.5998474,0.845068,0.83752275,0.724344,0.5998474,0.52439487,0.3055826,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23767537,0.40367088,0.32821837,0.0,0.0,0.0,0.0,0.041498873,0.19994913,0.29426476,0.12826926,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.090543,0.3961256,0.9205205,0.6790725,0.2867195,0.06413463,0.0150905,0.0150905,0.1358145,0.32821837,0.52062225,0.58098423,1.177059,1.0148361,1.5052774,3.0445085,5.036454,3.6556737,2.11267,1.3166461,1.0676528,0.030181,0.090543,0.27917424,0.31312788,0.35462674,1.0374719,3.712263,2.9237845,1.2940104,0.36594462,0.6111652,0.48666862,0.23013012,0.08299775,0.12826926,0.27540162,0.13958712,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041498873,0.08677038,0.0,0.0,0.24899325,0.5093044,0.724344,0.9922004,0.724344,0.7582976,0.72811663,0.55080324,0.42630664,0.36594462,0.67152727,0.8111144,0.72811663,0.8224323,0.59230214,1.780679,2.6219745,2.384299,1.358145,2.6634734,3.5047686,3.6669915,3.31991,2.9916916,2.916239,3.5387223,3.9989824,5.3873086,10.7557535,8.793989,7.5037513,8.145098,9.880505,9.797507,5.6815734,5.515578,6.2399216,6.0776987,4.5007415,5.4288073,6.4474163,7.277394,6.862405,3.3727267,3.0558262,2.5993385,2.1654868,1.780679,1.3430545,1.5618668,1.7731338,1.7957695,2.3314822,4.9421387,7.605612,6.428553,5.515578,8.13378,16.739138,11.174516,8.296002,9.14107,11.25374,8.729855,5.1043615,5.0213637,5.4212623,4.847823,3.4330888,4.0178456,4.1197066,3.410453,3.0897799,5.8588867,5.1156793,4.9459114,4.3724723,3.4368613,3.2029586,3.7650797,5.0213637,7.816879,10.182315,7.3415284,4.508287,5.5759397,6.911449,6.7756343,5.311856,4.772371,5.643847,5.934339,4.749735,2.3201644,3.6368105,5.093044,6.1418333,6.63982,6.8359966,6.749226,11.351829,13.917213,11.306557,3.983892,4.4705606,6.6058664,10.763299,12.879742,4.45547,1.9768555,5.0477724,10.005001,12.14408,5.7381625,4.9685473,4.719554,4.323428,3.5236318,2.4861598,2.3880715,2.4823873,3.4255435,5.855114,10.4049,14.275613,8.303548,3.561358,3.531177,4.104616,4.2517486,7.6093845,12.864652,16.663685,13.626721,6.6322746,3.6292653,6.3945994,10.93684,7.5075235,3.2105038,6.6322746,10.948157,11.091517,3.7688525,5.66271,9.8239155,11.314102,8.975075,5.4476705,7.5829763,7.2472124,8.322411,11.9064045,16.31283,12.102581,7.533932,6.458734,8.20546,7.5829763,7.779153,9.778644,9.159933,6.519096,7.4471617,11.853588,13.404137,11.664956,8.616675,8.66572,12.291212,12.759018,14.7321005,21.790682,36.436012,54.506886,58.920856,49.485523,36.14552,39.001396,43.37387,43.75868,44.62261,46.64851,46.78432,37.05472,36.179474,37.23581,36.104023,31.478783,33.94608,34.632698,32.961426,30.26777,29.815056,30.988342,38.194054,43.622864,41.53283,28.230553,28.411638,29.52079,27.44962,23.450638,24.107073,19.859098,12.985375,7.5603404,5.0854983,4.5007415,8.786444,7.9451485,4.538468,1.2223305,0.7469798,0.724344,0.452715,0.34330887,0.4640329,0.55080324,1.0978339,0.90543,0.7432071,0.7394345,0.3961256,0.543258,0.5055317,0.42630664,0.35839936,0.26031113,0.06413463,0.00754525,0.0,0.003772625,0.0150905,0.16222288,0.19994913,0.362172,1.0110635,2.6106565,4.304565,4.217795,3.8895764,3.9801195,4.2706113,3.8065786,2.6936543,1.6524098,0.995973,0.6413463,1.0789708,2.142851,3.2670932,4.247976,5.247721,5.9796104,5.8437963,5.20245,3.983892,1.6788181,0.70170826,0.32821837,0.24522063,0.24522063,0.24522063,0.15845025,0.071679875,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.041498873,0.06413463,0.0754525,0.08299775,0.1056335,0.056589376,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0452715,0.1056335,0.120724,0.094315626,0.056589376,0.056589376,0.150905,0.33576363,0.29049212,0.17354076,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.13204187,0.2565385,0.24522063,0.071679875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.02263575,0.0754525,0.1358145,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.02263575,0.041498873,0.0754525,0.10186087,0.116951376,0.120724,0.120724,0.1056335,0.14335975,0.20749438,0.27540162,0.32821837,0.35085413,0.3734899,0.362172,0.38103512,0.41498876,0.36594462,0.42630664,0.47912338,0.5281675,0.6488915,0.9922004,0.845068,0.633801,0.422534,0.26408374,0.23013012,0.32821837,0.2867195,0.20749438,0.16976812,0.24522063,0.35462674,0.39989826,0.43007925,0.422534,0.27540162,0.35839936,0.5017591,0.5357128,0.48666862,0.5357128,0.4979865,0.452715,0.34330887,0.19240387,0.1056335,0.071679875,0.041498873,0.02263575,0.0150905,0.0150905,0.003772625,0.00754525,0.02263575,0.030181,0.030181,0.030181,0.02263575,0.0150905,0.018863125,0.030181,0.030181,0.041498873,0.0452715,0.0452715,0.0452715,0.0452715,0.0452715,0.0452715,0.041498873,0.0150905,0.026408374,0.02263575,0.0150905,0.011317875,0.0,0.0,0.018863125,0.049044125,0.08677038,0.120724,0.14713238,0.16976812,0.18863125,0.20372175,0.23013012,0.29049212,0.32444575,0.29803738,0.25276586,0.29049212,0.33953625,0.35839936,0.35462674,0.38858038,0.59607476,0.5583485,0.43007925,0.362172,0.38858038,0.41121614,0.41121614,0.36594462,0.35462674,0.41498876,0.55080324,0.6451189,0.52439487,0.4376245,0.4376245,0.35085413,0.33953625,0.38103512,0.47157812,0.5470306,0.47157812,0.47157812,0.5357128,0.5998474,0.62248313,0.6111652,0.965792,1.0789708,0.995973,0.80734175,0.67152727,0.120724,0.10186087,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.030181,0.011317875,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3470815,0.47535074,0.28294688,0.15845025,0.95824677,0.9997456,0.5357128,0.030181,0.150905,0.21881226,0.094315626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.181086,0.8865669,1.1280149,0.8639311,0.422534,0.08299775,0.06413463,0.3470815,0.9997456,2.1202152,3.3048196,3.6179473,4.6554193,3.8782585,2.5804756,2.1805773,4.2291126,3.682082,1.8448136,0.6375736,0.43007925,0.06790725,0.041498873,1.0072908,1.0601076,0.2867195,0.7432071,1.0450171,0.7922512,0.452715,0.25276586,0.18485862,0.120724,0.056589376,0.030181,0.033953626,0.056589376,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.0,0.06790725,0.18485862,0.422534,0.84884065,1.5165952,1.1619685,1.1355602,1.1355602,0.9393836,0.42630664,0.482896,0.7432071,1.4939595,2.022127,0.6149379,0.754525,1.9164935,2.8747404,3.0935526,2.7615614,3.169005,3.85185,4.2291126,4.002755,3.138824,2.7615614,3.0897799,3.7160356,4.7346444,6.719045,6.432326,6.25124,7.6508837,9.35611,7.3679366,4.9232755,5.3194013,5.775889,5.0062733,3.2067313,5.666483,6.63982,6.488915,5.2967653,2.8709676,2.1654868,1.7429527,1.6222287,1.5279131,0.9016574,0.9280658,1.1129243,1.2713746,1.5505489,2.4031622,6.4738245,5.2665844,3.9461658,6.1229706,13.8719425,10.216269,7.99042,8.103599,8.756263,5.406172,4.1083884,4.9119577,5.304311,4.9232755,5.5683947,6.888813,5.3269467,3.1350515,2.2371666,4.236658,4.9157305,5.828706,5.50426,4.164978,3.7160356,5.2364035,4.044254,4.112161,5.907931,6.4134626,4.9157305,7.515069,8.548768,7.2698483,7.835742,8.137552,7.816879,7.541477,7.322665,6.4926877,4.8138695,5.2137675,6.72659,8.82417,11.41219,13.328684,13.430545,10.461489,5.692891,2.9200118,4.5799665,11.140562,14.128481,10.982111,5.040227,2.3578906,2.9841464,7.5490227,12.185578,8.518587,5.1043615,3.9197574,3.6594462,3.6179473,3.682082,5.481624,5.0968165,5.1534057,6.2361493,6.903904,7.7640624,5.764571,5.172269,6.3229194,5.617439,6.692637,10.386037,12.679792,12.166716,10.072908,10.167224,10.665211,10.242677,7.960239,3.270866,3.9763467,8.827943,12.132762,10.495442,2.8294687,3.482133,3.9348478,6.881268,10.853842,10.242677,9.22784,8.952439,8.186596,6.9454026,6.511551,4.6818275,5.9532022,9.042982,11.6008215,10.197406,5.926794,9.374973,10.303039,6.466279,3.6254926,10.336992,13.479589,12.73261,9.6201935,7.5188417,9.359882,9.876732,11.646093,15.716756,21.594505,27.155355,28.868126,26.317833,22.409393,23.34123,29.799965,27.906107,25.623669,26.676231,30.550716,33.60277,38.2016,42.694798,44.633926,40.766987,37.979015,36.66614,35.08164,33.236828,32.889744,37.1679,40.204865,41.019753,38.62036,32.010723,27.56657,27.027086,26.910133,25.914162,24.903097,19.247932,13.3626375,10.20495,9.337247,6.907676,9.031664,6.187105,2.584248,0.5394854,0.45648763,0.7432071,0.58475685,0.43385187,0.46026024,0.58475685,1.4298248,1.4864142,0.9507015,0.2867195,0.23767537,0.3055826,0.30935526,0.30181,0.29803738,0.26031113,0.0754525,0.018863125,0.018863125,0.05281675,0.16222288,0.3961256,0.33576363,0.28294688,0.5093044,1.2789198,2.3993895,2.8407867,3.0822346,3.561358,4.6742826,4.5912848,3.4632697,2.0108092,0.87902164,0.6413463,0.9620194,1.659955,2.323937,2.8785129,3.5764484,3.5877664,3.4594972,3.078462,2.2711203,0.8111144,0.41121614,0.2867195,0.23767537,0.181086,0.120724,0.06413463,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.018863125,0.033953626,0.041498873,0.0452715,0.03772625,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.05281675,0.14335975,0.14713238,0.17731337,0.1659955,0.14335975,0.24899325,1.1544232,0.95447415,0.482896,0.18863125,0.14713238,0.116951376,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.026408374,0.05281675,0.049044125,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.003772625,0.060362,0.26031113,0.10186087,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.03772625,0.090543,0.18485862,0.13204187,0.1358145,0.1358145,0.11317875,0.08299775,0.09808825,0.1358145,0.181086,0.241448,0.362172,0.41498876,0.45648763,0.44516975,0.38480774,0.3169005,0.6526641,0.69039035,0.5885295,0.5583485,0.87147635,0.7432071,0.7997965,0.754525,0.5394854,0.33953625,0.32067314,0.26408374,0.35085413,0.77338815,1.7467253,1.4147344,0.88279426,0.49044126,0.3169005,0.19994913,0.2565385,0.32444575,0.3772625,0.43385187,0.5696664,0.52439487,0.44516975,0.34330887,0.23013012,0.14335975,0.08677038,0.049044125,0.030181,0.026408374,0.0150905,0.003772625,0.0,0.003772625,0.00754525,0.00754525,0.0150905,0.02263575,0.026408374,0.026408374,0.030181,0.030181,0.041498873,0.0452715,0.0452715,0.0452715,0.03772625,0.041498873,0.0452715,0.0452715,0.041498873,0.033953626,0.02263575,0.0150905,0.011317875,0.0,0.0,0.011317875,0.026408374,0.0452715,0.071679875,0.09808825,0.11317875,0.12826926,0.13958712,0.15467763,0.2263575,0.29803738,0.30935526,0.2565385,0.21503963,0.2565385,0.33953625,0.40367088,0.43007925,0.46026024,0.5017591,0.49044126,0.422534,0.32821837,0.25276586,0.331991,0.35085413,0.33576363,0.331991,0.3772625,0.42630664,0.43385187,0.40367088,0.35839936,0.30181,0.30935526,0.32821837,0.4376245,0.5696664,0.48666862,0.4074435,0.47535074,0.55080324,0.5772116,0.58475685,0.7054809,0.9242931,1.0299267,0.9393836,0.694163,0.34330887,0.5319401,0.5055317,0.331991,0.120724,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.1961765,0.331991,0.29049212,0.10186087,0.071679875,0.026408374,0.00754525,0.026408374,0.060362,0.026408374,0.00754525,0.003772625,0.00754525,0.0,0.0,0.0,0.018863125,0.03772625,0.00754525,0.0,0.150905,0.1961765,0.10940613,0.07922512,1.7391801,1.9768555,1.146878,0.08677038,0.10186087,0.08677038,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.116951376,0.5017591,0.56589377,0.5055317,0.31312788,0.15467763,0.3772625,0.7922512,0.9922004,1.569412,2.293756,2.1013522,2.9766011,2.8219235,1.841041,0.9808825,1.9693103,2.5578396,1.3920987,0.39989826,0.181086,0.030181,0.011317875,0.4979865,0.5885295,0.2867195,0.5055317,0.22258487,0.1358145,0.13958712,0.1358145,0.049044125,0.0150905,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.06790725,0.271629,0.63002837,0.9507015,0.91674787,0.8337501,0.7809334,0.80734175,0.9318384,0.9280658,0.8941121,1.0714256,1.2600567,0.80356914,2.3390274,3.0030096,2.7125173,1.9844007,1.9240388,2.493705,3.451952,4.0216184,4.025391,3.8971217,4.4630156,5.1345425,4.9723196,4.496969,5.7079816,6.156924,6.2323766,7.2962565,8.167733,5.13077,3.893349,4.5799665,5.0062733,4.4630156,3.7084904,5.3156285,5.5570765,4.7912335,3.4217708,1.9051756,1.3166461,1.1204696,1.3468271,1.5769572,0.95824677,1.1317875,1.6260014,1.9353566,1.9429018,1.9353566,6.477597,5.1269975,3.3689542,4.044254,7.356619,6.3531003,6.4474163,8.469543,10.170997,6.2436943,4.8930945,5.1269975,4.9119577,4.187614,4.8855495,6.790725,5.3759904,3.640583,3.048281,3.5387223,3.9801195,4.727099,4.851596,4.395108,4.349837,5.081726,3.6254926,3.4859054,5.2364035,6.5266414,5.3684454,6.145606,6.432326,6.0248823,6.94163,6.719045,6.168242,6.2399216,6.507778,5.1571784,4.3309736,6.6850915,10.582213,14.886778,18.976303,18.368912,11.7894535,5.704209,2.776652,1.8938577,4.183841,9.989911,11.019837,7.122716,6.296511,4.1536603,3.1048703,4.357382,6.5945487,6.013564,3.8254418,2.704972,2.463524,2.848332,3.5424948,4.6856003,4.889322,6.485142,8.82417,8.269594,7.5905213,6.5643673,7.2094865,8.854351,8.167733,8.805306,12.012038,13.019329,10.774617,7.9225125,15.384765,17.96524,14.377474,7.2283497,3.0105548,7.4584794,10.536942,10.008774,6.4738245,3.3727267,5.221313,5.27413,7.3151197,11.747954,15.580941,11.563096,8.379,6.009792,4.8138695,5.523123,5.8928404,8.043237,10.001229,10.170997,7.3415284,4.1197066,6.349328,7.073672,5.0175915,4.564876,10.140816,13.060828,11.98563,8.541223,7.333983,9.201432,9.544742,10.680302,13.041965,15.181043,15.362129,16.120426,16.365646,15.916705,15.497944,19.527107,21.42851,25.370903,34.051712,48.697044,60.939213,67.933655,71.178116,69.39744,58.55114,43.083378,35.534355,31.810774,29.679241,28.788902,37.190536,38.68827,37.111313,34.255436,29.90937,27.457165,25.902843,26.05375,27.44962,28.339958,22.062311,16.505234,12.525115,9.548513,5.5495315,6.145606,4.1272516,1.8372684,0.5998474,0.7205714,0.66775465,0.573439,0.6451189,0.8978847,1.1732863,1.5241405,1.3958713,0.83752275,0.2867195,0.573439,0.32821837,0.30181,0.36971724,0.46026024,0.55080324,0.3772625,0.21503963,0.1056335,0.094315626,0.23390275,0.43385187,0.56589377,0.5998474,0.58475685,0.67152727,1.297783,1.9089483,2.2107582,2.293756,2.6144292,3.0143273,2.8445592,2.142851,1.3015556,1.0336993,0.80734175,1.0072908,1.2940104,1.5165952,1.720317,1.5807298,1.4411428,1.2449663,0.91297525,0.35839936,0.25276586,0.211267,0.16976812,0.1056335,0.0452715,0.018863125,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.02263575,0.0150905,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.056589376,0.124496624,0.17731337,0.31312788,0.38103512,0.3734899,0.392353,1.0487897,1.1808317,1.0751982,0.83752275,0.41121614,0.22258487,0.1358145,0.06790725,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.116951376,0.049044125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.17731337,0.25276586,0.25276586,0.1961765,0.120724,0.10186087,0.10186087,0.10186087,0.08677038,0.090543,0.124496624,0.15845025,0.19994913,0.30181,0.422534,0.5319401,0.5357128,0.42630664,0.2867195,0.5583485,0.6488915,0.7130261,0.8262049,0.98465514,0.7167987,0.77716076,0.73566186,0.52062225,0.43007925,0.543258,0.573439,0.94692886,1.9391292,3.6783094,2.1315331,1.0148361,0.4376245,0.30181,0.2565385,0.20372175,0.24899325,0.32444575,0.392353,0.44139713,0.55457586,0.52439487,0.43385187,0.331991,0.25276586,0.21503963,0.17731337,0.13204187,0.07922512,0.02263575,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.0150905,0.02263575,0.02263575,0.026408374,0.033953626,0.049044125,0.056589376,0.049044125,0.05281675,0.049044125,0.041498873,0.056589376,0.049044125,0.033953626,0.02263575,0.02263575,0.00754525,0.00754525,0.011317875,0.018863125,0.026408374,0.05281675,0.09808825,0.12826926,0.16222288,0.181086,0.1659955,0.18863125,0.22258487,0.23013012,0.20372175,0.16976812,0.19994913,0.23767537,0.28294688,0.3169005,0.33576363,0.40367088,0.47157812,0.48666862,0.43007925,0.29426476,0.32821837,0.3734899,0.3772625,0.35462674,0.362172,0.38480774,0.38480774,0.3734899,0.362172,0.3734899,0.39989826,0.38103512,0.41876137,0.49044126,0.47157812,0.5055317,0.6488915,0.66020936,0.5281675,0.452715,0.4979865,0.69039035,0.87147635,0.9205205,0.7469798,0.9695646,1.1619685,0.87147635,0.452715,0.1358145,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.38103512,0.6375736,0.5357128,0.10186087,0.071679875,0.056589376,0.030181,0.011317875,0.056589376,0.011317875,0.00754525,0.0150905,0.011317875,0.0,0.0,0.0,0.018863125,0.03772625,0.00754525,0.0,0.116951376,0.17731337,0.116951376,0.0,1.2600567,1.4750963,0.87902164,0.0754525,0.0452715,0.049044125,0.018863125,0.0,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.094315626,0.094315626,0.026408374,0.011317875,0.00754525,0.02263575,0.05281675,0.094315626,0.16222288,0.124496624,0.20749438,0.22258487,0.23390275,0.5319401,0.7582976,0.56212115,0.55080324,0.7205714,0.48666862,1.2525115,1.3204187,0.8186596,0.23390275,0.41876137,1.3468271,0.845068,0.2678564,0.10940613,0.018863125,0.003772625,0.026408374,0.094315626,0.18863125,0.2678564,0.090543,0.041498873,0.05281675,0.06413463,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.15467763,0.36971724,0.5696664,0.48666862,0.5772116,0.513077,0.47535074,0.5998474,0.98465514,0.91674787,0.8526133,0.633801,0.43007925,0.7432071,2.6672459,3.1916409,2.4107075,1.1581959,0.9997456,1.4449154,2.5767028,3.4859054,3.9688015,4.5120597,5.523123,6.598321,6.258785,5.1269975,5.8966126,6.7077274,6.375736,6.3153744,6.138061,3.6707642,2.7917426,3.6858547,4.745962,4.9760923,4.025391,3.99521,3.8254418,3.218049,2.214531,1.1959221,1.1317875,1.1053791,1.3430545,1.6222287,1.2751472,1.50905,2.0372176,2.565385,2.9086938,3.0030096,6.247467,5.168496,3.5651307,3.2444575,4.006528,4.1197066,4.776143,7.183078,9.616421,7.4396167,5.3382645,5.534441,4.8100967,3.2029586,4.006528,5.617439,4.9949555,4.644101,5.081726,4.847823,3.470815,3.904667,4.5309224,4.6290107,4.3724723,3.983892,3.048281,3.259548,4.606375,5.3759904,4.798779,4.4894238,4.2894745,4.164978,4.168751,3.7575345,3.5802212,3.863168,4.349837,4.285702,7.213259,9.680555,11.578186,13.343775,15.984612,14.200161,7.466025,2.7653341,2.1202152,2.584248,4.112161,8.695901,8.790216,5.036454,6.247467,4.187614,2.7540162,2.022127,2.0183544,2.7351532,2.354118,1.6939086,1.4826416,2.093807,3.5538127,4.8063245,6.7944975,9.476834,11.729091,11.321648,9.076936,7.201941,7.5792036,9.623966,10.272858,9.616421,10.287949,10.269085,8.963757,7.201941,14.0907545,15.78089,12.155397,6.2399216,4.236658,8.956212,9.039209,6.719045,4.3686996,4.5120597,8.820397,8.224322,7.779153,10.140816,15.565851,10.93684,7.356619,5.5193505,5.534441,6.903904,7.4018903,8.209232,9.005256,8.567632,4.768598,2.704972,4.6629643,5.987156,6.043745,8.182823,13.664448,13.894578,11.065109,8.09228,8.60913,10.438853,10.736891,11.23865,12.095036,11.861133,10.446399,11.32542,12.193124,12.170488,11.812089,13.819125,20.360857,30.920435,45.96189,66.93768,94.3194,100.54046,96.575424,86.442154,67.23195,44.31325,34.11585,30.826118,30.101774,29.071848,37.907337,38.97876,35.847485,31.4901,28.309778,27.804247,26.755457,27.400576,29.671696,31.192064,25.78212,19.353567,13.287186,8.5563135,5.726845,4.5007415,3.4330888,2.4672968,1.6712729,1.2525115,0.814887,0.6790725,1.0412445,1.6788181,1.9278114,1.5618668,1.1431054,0.7394345,0.56212115,0.95824677,0.42630664,0.3169005,0.36971724,0.46026024,0.6149379,0.55080324,0.362172,0.18863125,0.116951376,0.19994913,0.43007925,0.9242931,1.1016065,0.8865669,0.6790725,0.814887,1.1544232,1.4034165,1.4675511,1.4750963,2.4522061,3.3764994,3.3463185,2.3805263,1.4373702,0.7469798,0.7432071,0.8262049,0.7696155,0.7130261,0.6451189,0.47535074,0.32821837,0.24899325,0.241448,0.20749438,0.15845025,0.10940613,0.060362,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.0452715,0.094315626,0.18485862,0.3734899,0.52062225,0.5772116,0.58475685,0.8186596,1.0902886,1.3392819,1.3732355,0.9016574,0.5055317,0.35839936,0.21503963,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08299775,0.21503963,0.29426476,0.27917424,0.16976812,0.12826926,0.094315626,0.08299775,0.090543,0.08677038,0.090543,0.116951376,0.13958712,0.1659955,0.23390275,0.36594462,0.51684964,0.573439,0.49044126,0.32444575,0.5055317,0.62248313,0.79602385,0.995973,1.0412445,0.7507524,0.7469798,0.633801,0.42630664,0.5394854,0.87147635,0.7809334,1.0148361,1.9278114,3.451952,2.0070364,0.8978847,0.33576363,0.241448,0.2263575,0.14713238,0.18863125,0.26408374,0.30935526,0.29426476,0.48666862,0.5583485,0.5357128,0.47157812,0.44894236,0.40367088,0.32444575,0.23767537,0.15467763,0.071679875,0.03772625,0.0150905,0.00754525,0.003772625,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.00754525,0.011317875,0.026408374,0.041498873,0.049044125,0.060362,0.056589376,0.049044125,0.041498873,0.060362,0.060362,0.049044125,0.041498873,0.033953626,0.0150905,0.018863125,0.018863125,0.0150905,0.018863125,0.033953626,0.0754525,0.11317875,0.15845025,0.19240387,0.16976812,0.19240387,0.23013012,0.23390275,0.20749438,0.19994913,0.22258487,0.19994913,0.18863125,0.211267,0.24522063,0.31312788,0.3961256,0.49044126,0.5357128,0.422534,0.3734899,0.39989826,0.392353,0.33576363,0.32821837,0.33953625,0.35085413,0.35462674,0.362172,0.3961256,0.422534,0.38480774,0.362172,0.3961256,0.47535074,0.543258,0.6526641,0.6451189,0.51684964,0.392353,0.35839936,0.4678055,0.65643674,0.7997965,0.724344,1.50905,1.50905,0.83752275,0.24522063,0.03772625,0.071679875,0.0150905,0.0,0.0,0.0,0.0,0.011317875,0.41498876,0.66775465,0.52062225,0.0,0.0,0.060362,0.060362,0.003772625,0.02263575,0.00754525,0.0150905,0.018863125,0.011317875,0.0150905,0.003772625,0.0,0.011317875,0.02263575,0.0,0.049044125,0.39989826,0.6073926,0.4640329,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.07922512,0.049044125,0.00754525,0.0,0.0,0.0,0.0,0.033953626,0.07922512,0.049044125,0.011317875,0.0,0.0,0.003772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.13204187,0.32821837,0.33953625,0.15467763,0.026408374,0.02263575,0.094315626,0.21503963,0.3169005,0.2867195,0.150905,0.33953625,0.5583485,0.6752999,0.7205714,0.7054809,0.30935526,0.026408374,0.056589376,0.27917424,0.98842776,0.6828451,0.24522063,0.0754525,0.124496624,0.5394854,0.331991,0.10940613,0.07922512,0.0452715,0.00754525,0.00754525,0.011317875,0.026408374,0.0754525,0.0452715,0.018863125,0.018863125,0.033953626,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18485862,0.43385187,0.63002837,0.67152727,0.47157812,0.3470815,0.38480774,0.44894236,0.47912338,0.4640329,0.38480774,0.5281675,0.46026024,0.24522063,0.44894236,1.4071891,2.0862615,2.0183544,1.4298248,1.2449663,0.83752275,1.6071383,2.7125173,3.7009451,4.538468,5.0515447,6.3719635,6.828451,6.319147,6.2889657,7.1793056,6.2135134,5.0854983,4.38379,3.5764484,1.9127209,2.8936033,5.036454,6.205968,3.6292653,2.2899833,2.2975287,2.4333432,2.0749438,1.1883769,1.4298248,1.4713237,1.5316857,1.7014539,1.931584,1.9579924,2.1503963,2.757789,3.6707642,4.4215164,5.3948536,5.2628117,4.2517486,3.3123648,4.1083884,4.293247,3.85185,4.4931965,6.1795597,7.1000805,5.100589,6.1078796,5.2326307,2.6672459,3.6971724,4.4441524,4.610148,5.3986263,6.5568223,6.349328,3.3953626,3.85185,4.817642,4.847823,3.9688015,2.9916916,2.4786146,2.637065,3.127506,3.0558262,3.3576362,3.591539,3.3651814,2.5880208,1.4864142,1.4562333,1.8184053,2.1843498,2.897376,5.0251365,10.325675,10.555805,7.91874,5.0062733,4.8063245,4.3347464,3.2633207,2.5276587,2.6823363,3.9197574,3.8556228,8.080963,8.60913,5.0025005,4.353609,2.3013012,1.4675511,1.0110635,0.7092535,0.9695646,1.4034165,1.1544232,1.0374719,1.8334957,4.255521,7.111398,10.831206,13.551269,14.796235,15.448899,10.653893,7.149124,7.333983,10.555805,13.151371,9.982366,7.0849895,6.398372,7.54525,7.8319697,7.5565677,7.164215,6.2135134,5.062863,4.8629136,7.462252,5.704209,4.3611546,4.9345937,5.613666,11.593277,9.763554,7.254758,7.605612,10.785934,7.6395655,6.696409,6.937857,7.443389,7.3868,6.541732,5.7872066,6.4964604,7.2660756,3.9197574,2.2484846,5.802297,8.228095,8.431817,10.616167,17.350302,14.400109,10.016319,8.288457,9.144843,10.370946,10.880251,10.993429,10.465261,8.473316,8.213005,10.552032,11.144334,9.684328,9.910686,12.709973,22.49239,36.036114,51.97923,70.82726,116.07236,120.22979,106.26353,86.86469,64.44398,44.633926,36.711414,36.251152,38.895763,40.35577,44.501884,43.483276,37.801704,30.701622,28.158873,27.943834,28.449366,29.924461,31.512737,31.263742,28.60027,21.398329,13.687083,8.635539,8.552541,5.6325293,4.4894238,3.9612563,3.2067313,1.6939086,1.237421,1.1581959,1.7467253,2.6031113,2.6408374,1.8599042,1.2638294,1.0035182,1.0487897,1.1996948,0.5319401,0.3961256,0.35462674,0.28294688,0.3734899,0.47912338,0.482896,0.38858038,0.23767537,0.090543,0.38103512,1.0827434,1.3656902,1.1129243,0.8903395,0.8903395,0.6526641,0.73188925,1.20724,1.690136,2.9501927,4.3686996,4.5912848,3.4179983,1.81086,0.9695646,0.97710985,1.0487897,0.94315624,0.935611,0.76207024,0.4979865,0.27917424,0.18485862,0.26031113,0.18863125,0.13204187,0.08299775,0.0452715,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.08677038,0.18485862,0.3470815,0.52439487,0.67152727,0.77716076,0.8262049,0.9016574,1.1242423,1.3770081,1.327964,0.97333723,0.7092535,0.452715,0.19994913,0.030181,0.00754525,0.003772625,0.003772625,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05281675,0.08677038,0.120724,0.150905,0.14713238,0.14713238,0.124496624,0.1056335,0.09808825,0.08677038,0.10186087,0.11317875,0.116951376,0.13958712,0.19994913,0.27540162,0.4074435,0.5017591,0.5017591,0.38858038,0.58098423,0.6828451,0.8111144,0.94692886,0.9318384,0.7809334,0.7432071,0.56589377,0.35462674,0.56212115,0.97333723,0.663982,0.47912338,0.76207024,1.3505998,1.7354075,0.94315624,0.271629,0.14335975,0.116951376,0.090543,0.120724,0.16222288,0.18485862,0.18863125,0.33576363,0.5017591,0.6187105,0.66020936,0.6488915,0.59607476,0.46026024,0.33576363,0.24522063,0.15467763,0.0754525,0.033953626,0.018863125,0.011317875,0.0,0.003772625,0.00754525,0.011317875,0.011317875,0.003772625,0.0,0.00754525,0.018863125,0.026408374,0.026408374,0.049044125,0.049044125,0.0452715,0.049044125,0.056589376,0.060362,0.06413463,0.060362,0.0452715,0.026408374,0.033953626,0.026408374,0.018863125,0.0150905,0.018863125,0.026408374,0.049044125,0.094315626,0.13958712,0.150905,0.22258487,0.29049212,0.29803738,0.2565385,0.25276586,0.26408374,0.22258487,0.18485862,0.16976812,0.18485862,0.23767537,0.29426476,0.39989826,0.51684964,0.5093044,0.40367088,0.392353,0.35085413,0.2678564,0.24522063,0.25276586,0.3055826,0.331991,0.32821837,0.34330887,0.35839936,0.3169005,0.2867195,0.32067314,0.46026024,0.47157812,0.45648763,0.47157812,0.4979865,0.43385187,0.3169005,0.331991,0.47535074,0.6375736,0.59607476,0.94692886,0.7997965,0.34330887,0.041498873,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.23390275,0.29426476,0.16976812,0.0,0.0,0.0,0.0,0.02263575,0.1056335,0.033953626,0.00754525,0.0,0.0150905,0.0754525,0.0150905,0.0,0.056589376,0.10940613,0.0,0.24522063,0.83752275,1.2826926,1.1544232,0.090543,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0452715,0.0452715,0.0,0.0,0.0,0.0,0.049044125,0.09808825,0.0,0.0,0.0,0.0,0.02263575,0.1056335,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.090543,0.422534,0.7130261,0.76207024,0.5017591,0.0150905,0.041498873,0.29426476,0.6828451,0.9808825,0.8224323,0.43385187,1.0487897,1.8561316,2.233394,1.7693611,2.1353056,0.95447415,0.06413463,0.0,0.0,0.071679875,0.06413463,0.033953626,0.0150905,0.0150905,0.026408374,0.02263575,0.0150905,0.02263575,0.0452715,0.00754525,0.0,0.0,0.0150905,0.0754525,0.026408374,0.0150905,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48666862,0.6375736,0.56589377,0.422534,0.41121614,0.08299775,0.18485862,0.34330887,0.32821837,0.060362,0.011317875,0.0,0.0,0.120724,0.59607476,0.5470306,0.72811663,1.3845534,2.3428001,2.9916916,1.4901869,1.0487897,1.4109617,2.3767538,3.8292143,3.7575345,5.342037,6.6850915,7.020855,6.730363,7.0359454,5.885295,5.149633,5.311856,5.43258,1.6486372,2.305074,5.1534057,6.9491754,3.4330888,1.7240896,2.0560806,2.7351532,2.7992878,2.0296721,1.2487389,1.3920987,1.7391801,2.1994405,3.3123648,2.9464202,2.8709676,2.938875,3.2859564,4.349837,4.5196047,5.9909286,5.070408,2.093807,1.4335974,3.874486,4.3121104,3.9386206,3.8895764,5.2175403,5.6325293,6.937857,6.0626082,3.4142256,2.8521044,3.5236318,4.3422914,4.708236,4.346064,3.2972744,2.5880208,3.2633207,4.134797,4.5196047,4.22534,3.531177,2.9728284,2.71629,2.5917933,2.0900342,2.384299,2.5125682,2.4031622,1.9994912,1.267602,0.97333723,1.5430037,2.9086938,4.191386,3.6934,2.3616633,1.8372684,2.1541688,2.9992368,3.7084904,3.440634,3.783943,3.6443558,2.8332415,2.0900342,1.5656394,4.255521,5.4438977,3.8254418,1.4939595,1.3505998,0.9922004,0.65643674,0.5319401,0.76207024,1.177059,1.0148361,1.0525624,2.142851,5.2175403,9.35611,12.113899,15.494171,19.598787,22.613113,13.822898,8.8618965,10.650121,17.01831,20.704166,12.577931,8.329956,8.975075,11.653639,9.627739,6.5266414,7.9489207,8.499724,6.33801,3.187868,5.704209,5.994701,5.0062733,4.346064,6.2851934,10.242677,9.491924,8.5563135,8.782671,8.329956,5.938112,6.1908774,6.960493,7.194396,6.911449,6.349328,5.0666356,3.6745367,2.5804756,1.9693103,3.519859,8.793989,9.650374,6.0739264,6.19465,11.653639,9.65792,7.2698483,6.4474163,4.044254,4.983638,5.832478,5.8513412,5.0175915,4.0291634,8.986393,15.286676,15.316857,9.982366,8.710991,15.011275,27.351532,41.178204,54.076805,65.79458,115.604546,120.27883,101.16294,76.82196,63.063198,54.94451,49.03658,48.6065,54.34466,64.3308,60.509132,51.688736,40.178455,29.611334,24.94837,26.8045,28.08342,29.034122,29.20389,27.41944,29.422703,24.67674,17.346529,11.472552,10.970794,8.224322,6.3945994,5.1232247,3.8178966,1.6335466,1.7429527,2.2748928,2.9200118,3.361409,3.2482302,2.8709676,2.3465726,1.9881734,1.7731338,1.358145,0.7092535,0.77716076,0.663982,0.25276586,0.23013012,0.35085413,0.8224323,1.0223814,0.7130261,0.030181,0.116951376,0.33953625,0.7432071,1.0374719,0.6111652,1.5882751,0.8224323,0.23767537,0.44516975,0.76207024,1.2525115,1.8787673,2.516341,2.8709676,2.4559789,1.7240896,1.3770081,1.5731846,2.0485353,2.1202152,1.1921495,0.6790725,0.38480774,0.19994913,0.0754525,0.06413463,0.07922512,0.056589376,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.120724,0.21881226,0.32821837,0.47157812,0.66775465,0.9016574,0.98465514,0.935611,0.7432071,0.63002837,1.0223814,1.448688,1.0902886,0.80356914,0.69039035,0.090543,0.030181,0.0150905,0.0150905,0.018863125,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.0452715,0.09808825,0.120724,0.1358145,0.12826926,0.12826926,0.1358145,0.1358145,0.16222288,0.15845025,0.13958712,0.13958712,0.21503963,0.23767537,0.26408374,0.29426476,0.32821837,0.35085413,0.58475685,0.694163,0.8299775,0.9318384,0.7469798,0.6752999,0.65643674,0.5093044,0.27917424,0.24522063,0.3055826,0.23767537,0.1659955,0.21503963,0.52062225,3.1916409,1.8636768,0.3734899,0.13958712,0.150905,0.06790725,0.056589376,0.060362,0.06790725,0.090543,0.23767537,0.41121614,0.69793564,0.9318384,0.68661773,0.7092535,0.62625575,0.5017591,0.3734899,0.23013012,0.120724,0.06413463,0.033953626,0.011317875,0.0,0.011317875,0.00754525,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.003772625,0.0150905,0.026408374,0.030181,0.041498873,0.056589376,0.0452715,0.056589376,0.071679875,0.0754525,0.0754525,0.0754525,0.06413463,0.05281675,0.033953626,0.018863125,0.030181,0.018863125,0.0150905,0.041498873,0.08677038,0.1358145,0.211267,0.21881226,0.19994913,0.181086,0.1659955,0.1659955,0.17731337,0.17731337,0.16222288,0.1358145,0.150905,0.18863125,0.23767537,0.30181,0.41121614,0.32821837,0.29426476,0.28294688,0.2678564,0.24522063,0.23013012,0.23013012,0.24899325,0.28294688,0.32067314,0.34330887,0.3055826,0.24899325,0.23013012,0.29049212,0.38858038,0.392353,0.35839936,0.3470815,0.45648763,0.422534,0.32821837,0.38480774,0.52062225,0.41121614,1.0450171,0.5470306,0.18485862,0.0452715,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0452715,0.094315626,0.10186087,0.0,0.0,0.0,0.0,0.011317875,0.056589376,0.0150905,0.0,0.0,0.003772625,0.0150905,0.02263575,0.08299775,0.181086,0.29803738,0.40367088,0.31312788,0.33953625,0.38480774,0.32821837,0.018863125,0.003772625,0.0,0.018863125,0.056589376,0.08677038,0.018863125,0.00754525,0.00754525,0.011317875,0.049044125,0.1056335,0.094315626,0.05281675,0.018863125,0.0,0.0,0.0,0.0150905,0.033953626,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.0150905,0.02263575,0.08677038,0.18863125,0.20749438,0.5885295,0.55457586,0.1358145,0.17354076,0.73566186,0.66020936,0.62248313,1.3770081,3.7763977,1.7580433,1.3656902,1.7165444,2.516341,4.063117,1.6675003,0.6073926,0.19240387,0.02263575,0.011317875,0.026408374,0.018863125,0.00754525,0.003772625,0.003772625,0.026408374,0.030181,0.026408374,0.02263575,0.00754525,0.011317875,0.003772625,0.033953626,0.071679875,0.0150905,0.003772625,0.003772625,0.00754525,0.011317875,0.003772625,0.030181,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09808825,0.38480774,0.4979865,0.3772625,0.27917424,0.211267,0.211267,0.23013012,0.2565385,0.27917424,0.26031113,0.34330887,0.241448,0.24899325,1.2525115,0.754525,0.5470306,0.6790725,1.2826926,2.565385,1.5807298,1.116697,1.3543724,2.3126192,3.8405323,3.6896272,4.4403796,5.2665844,5.541986,4.8365054,4.3611546,3.92353,4.1008434,5.3344917,7.9451485,3.3915899,1.8485862,3.863168,6.9982195,5.824933,3.832987,2.8785129,2.916239,3.2369123,2.4672968,1.6976813,1.871222,2.5201135,3.1727777,3.3953626,2.463524,2.848332,3.289729,3.3689542,3.5424948,5.73439,4.304565,1.991946,0.94692886,2.7389257,4.304565,4.2706113,4.2706113,5.0138187,6.304056,4.7950063,5.624984,5.481624,4.1272516,4.4139714,5.27413,4.8629136,3.8895764,3.3312278,4.432834,2.6106565,2.5389767,3.0181,3.0633714,1.8825399,2.1843498,2.8256962,2.7502437,1.9164935,1.3091009,1.6410918,1.9051756,1.9994912,1.9655377,1.9881734,1.6448646,2.463524,3.097325,2.9464202,2.1541688,1.9466745,1.901403,1.6675003,1.297783,1.2411937,1.1996948,1.358145,1.418507,1.2185578,0.7469798,0.6149379,2.1390784,2.8634224,2.1353056,1.1431054,1.0035182,0.9997456,0.8903395,0.68661773,0.6526641,1.2449663,2.2107582,2.6483827,3.0520537,5.3269467,7.805561,9.525878,12.15917,14.78869,13.898351,10.080454,10.9594755,13.992666,16.11288,13.736128,8.303548,5.59103,6.4964604,8.465771,5.4891696,10.718028,15.131999,12.468526,4.8742313,2.897376,6.964266,6.790725,5.2062225,5.0553174,9.190115,9.144843,7.3679366,8.318638,11.193378,9.929549,6.952948,7.745199,8.793989,8.314865,6.2663302,5.1571784,4.13857,3.150142,2.3993895,2.3465726,4.357382,7.152897,6.519096,3.9084394,6.4511886,7.454707,7.809334,9.344792,11.555551,11.61214,8.29223,6.7379084,6.356873,6.009792,4.002755,12.015811,17.440845,16.739138,12.989148,15.890297,23.888262,34.059258,43.9209,53.009155,62.88966,98.42024,120.90508,114.35581,86.11394,66.847145,62.742527,63.0217,67.069725,74.27921,84.03145,67.26968,50.870075,39.804966,34.040394,28.49841,24.556017,21.711456,21.534143,23.646814,25.721758,28.468227,23.246916,16.746683,12.774108,12.264804,11.8045435,9.424017,7.020855,5.2326307,3.4255435,3.9273026,4.1083884,4.002755,3.7575345,3.6292653,3.3689542,3.048281,2.6710186,2.1315331,1.1996948,1.0223814,0.7205714,0.44516975,0.28294688,0.27917424,0.38103512,0.7997965,1.0072908,0.77338815,0.18863125,0.1659955,0.181086,0.27540162,0.41498876,0.47535074,0.7582976,0.7809334,0.513077,0.19240387,0.33576363,0.69793564,0.87902164,1.0223814,1.3468271,2.1654868,2.7502437,2.173032,1.7655885,2.203213,3.5236318,2.0296721,0.9393836,0.35085413,0.150905,0.041498873,0.03772625,0.049044125,0.40367088,0.76584285,0.11317875,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.150905,0.38103512,0.63002837,0.8186596,0.8639311,1.0676528,1.1846043,0.935611,0.513077,0.58475685,1.3430545,1.8485862,2.0108092,1.8184053,1.3505998,0.4074435,0.08677038,0.026408374,0.026408374,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.03772625,0.11317875,0.1961765,0.14713238,0.11317875,0.10940613,0.124496624,0.11317875,0.1358145,0.14713238,0.14713238,0.13958712,0.1659955,0.15845025,0.13958712,0.14713238,0.19240387,0.26408374,0.44894236,0.49044126,0.58475685,0.7582976,0.87147635,0.66020936,0.5470306,0.40367088,0.22258487,0.14713238,0.14713238,0.124496624,0.10186087,0.11317875,0.21503963,0.7469798,0.47535074,0.3055826,0.4640329,0.5055317,0.56589377,0.271629,0.056589376,0.060362,0.1056335,0.19240387,0.40367088,0.633801,0.7394345,0.51684964,0.58098423,0.5772116,0.5319401,0.44894236,0.30181,0.23013012,0.16976812,0.1056335,0.0452715,0.011317875,0.0150905,0.00754525,0.003772625,0.018863125,0.041498873,0.026408374,0.018863125,0.00754525,0.0,0.003772625,0.0150905,0.026408374,0.03772625,0.049044125,0.0452715,0.056589376,0.06413463,0.06413463,0.060362,0.05281675,0.060362,0.05281675,0.041498873,0.03772625,0.030181,0.026408374,0.018863125,0.0150905,0.026408374,0.06413463,0.15845025,0.16976812,0.1961765,0.26031113,0.32821837,0.23013012,0.17731337,0.17354076,0.18863125,0.17354076,0.116951376,0.124496624,0.18485862,0.33953625,0.694163,0.52062225,0.422534,0.35839936,0.29426476,0.23013012,0.21881226,0.21503963,0.2263575,0.24899325,0.29426476,0.331991,0.2867195,0.20749438,0.15467763,0.20372175,0.32067314,0.3470815,0.3055826,0.24899325,0.24899325,0.38858038,0.35085413,0.35462674,0.452715,0.5093044,1.4901869,0.9393836,0.41121614,0.22258487,0.26408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.049044125,0.071679875,0.2263575,0.1056335,0.0,0.003772625,0.018863125,0.011317875,0.003772625,0.0,0.0,0.0,0.03772625,0.20372175,0.392353,0.47912338,0.33953625,0.241448,0.12826926,0.06413463,0.060362,0.06413463,0.049044125,0.02263575,0.0150905,0.026408374,0.041498873,0.00754525,0.0,0.0,0.003772625,0.02263575,0.05281675,0.0452715,0.02263575,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.056589376,0.026408374,0.00754525,0.0150905,0.05281675,0.1056335,0.08677038,0.24522063,0.21881226,0.06413463,0.241448,0.84129536,0.59607476,0.5394854,1.2638294,2.9426475,1.4071891,0.8224323,0.7922512,1.5203679,3.7952607,1.2336484,0.38858038,0.1659955,0.033953626,0.0150905,0.00754525,0.003772625,0.0,0.003772625,0.026408374,0.08677038,0.060362,0.026408374,0.018863125,0.00754525,0.00754525,0.003772625,0.02263575,0.041498873,0.00754525,0.00754525,0.003772625,0.003772625,0.003772625,0.0,0.0150905,0.011317875,0.003772625,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12826926,0.19240387,0.14713238,0.09808825,0.09808825,0.24522063,0.5696664,0.8262049,0.5017591,0.28294688,0.211267,0.120724,0.24899325,1.2525115,0.46026024,0.2678564,0.41121614,0.83752275,1.6675003,1.0487897,0.8639311,1.2600567,2.191895,3.4066803,3.3312278,4.478106,5.3986263,5.304311,4.0895257,3.7273536,3.6707642,3.7499893,4.3083377,6.19465,5.7607985,3.2331395,3.0256453,5.59103,7.413208,3.9197574,2.897376,2.8822856,3.0331905,3.138824,1.7957695,1.4901869,2.1579416,3.338773,4.195159,3.451952,3.6594462,3.610402,3.0822346,2.8558772,5.2552667,3.500996,1.2525115,0.5696664,1.9429018,2.5804756,2.5427492,3.1765501,4.38379,4.5912848,3.3689542,3.9008942,4.221567,3.7198083,3.1124156,3.942393,3.5424948,3.0143273,3.218049,4.7874613,3.1576872,2.293756,2.1088974,2.1277604,1.4977322,3.169005,3.572676,3.1539145,2.4069347,1.8825399,2.4371157,2.263575,2.1503963,2.2484846,2.0749438,2.0296721,2.5427492,2.5993385,2.071171,1.7316349,1.6976813,1.5505489,1.3053282,1.056335,0.965792,0.9016574,0.8111144,0.7507524,0.70170826,0.55080324,0.543258,1.1959221,1.50905,1.2411937,0.935611,0.7997965,0.77338815,0.7507524,0.69039035,0.6451189,1.901403,3.6745367,4.459243,4.3422914,4.979865,6.6549106,7.5188417,8.186596,8.616675,8.103599,9.137298,10.303039,10.216269,8.560086,6.1078796,4.508287,3.9386206,6.1229706,8.914713,6.2663302,9.646602,11.446144,8.850578,4.7950063,7.960239,14.86037,12.151625,6.971811,4.6026025,8.461998,7.0963078,5.828706,7.2057137,10.080454,9.635284,7.7338815,8.088508,8.152642,6.7944975,4.3196554,3.8782585,6.462507,9.258021,10.208723,8.024373,5.587258,5.7419353,5.7909794,5.772116,8.439363,7.5301595,7.7301087,8.741172,10.284176,12.083718,10.631257,7.4811153,5.3609,5.111907,5.7192993,15.528125,16.833452,15.973294,17.13149,22.36412,29.709421,36.8095,43.309734,48.810223,52.835613,77.09737,108.60633,121.42948,108.225296,80.25505,62.946247,61.214615,67.560165,76.86723,86.404434,71.96659,58.083336,46.55419,37.824337,30.973251,26.05375,22.413166,21.405874,22.77911,24.669195,25.948114,20.979568,15.437581,12.694883,13.822898,14.600059,11.649866,8.356364,6.217286,4.8365054,5.4288073,5.119452,4.293247,3.5236318,3.5839937,3.1199608,2.8030603,2.5880208,2.282438,1.5354583,1.2525115,0.80734175,0.422534,0.23390275,0.29803738,0.35462674,0.6149379,0.6752999,0.4678055,0.2565385,0.43385187,0.331991,0.17731337,0.12826926,0.2678564,0.452715,0.6111652,0.63002837,0.52062225,0.45648763,1.2336484,1.1280149,1.1355602,1.5656394,2.0447628,2.7917426,2.4786146,1.9730829,1.8863125,2.5767028,1.871222,1.0110635,0.39989826,0.14335975,0.0754525,0.026408374,0.033953626,0.24899325,0.4640329,0.090543,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.13958712,0.40367088,0.7167987,0.95824677,0.965792,1.0223814,1.1129243,1.1393328,1.1129243,1.1506506,1.3204187,1.5128226,1.7655885,1.9127209,1.599593,0.80734175,0.29426476,0.056589376,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.049044125,0.1056335,0.14713238,0.19240387,0.20372175,0.16976812,0.1358145,0.150905,0.1961765,0.18485862,0.10940613,0.07922512,0.08299775,0.0754525,0.08677038,0.120724,0.16976812,0.35462674,0.46026024,0.5319401,0.59230214,0.633801,0.573439,0.4376245,0.33576363,0.29426476,0.22258487,0.10940613,0.06413463,0.056589376,0.060362,0.071679875,0.071679875,0.07922512,0.30935526,0.6828451,0.8337501,0.8224323,0.40367088,0.09808825,0.060362,0.08677038,0.16222288,0.3055826,0.5017591,0.6451189,0.52062225,0.452715,0.4678055,0.5470306,0.6526641,0.7432071,0.76207024,0.6451189,0.5055317,0.3961256,0.29803738,0.116951376,0.033953626,0.011317875,0.018863125,0.026408374,0.030181,0.02263575,0.00754525,0.0,0.0,0.011317875,0.018863125,0.02263575,0.026408374,0.026408374,0.041498873,0.041498873,0.0452715,0.05281675,0.056589376,0.05281675,0.049044125,0.0452715,0.0452715,0.041498873,0.033953626,0.02263575,0.011317875,0.011317875,0.026408374,0.06790725,0.1056335,0.1659955,0.23013012,0.26408374,0.23013012,0.20749438,0.1961765,0.181086,0.15467763,0.14713238,0.15467763,0.16222288,0.21881226,0.41498876,0.43385187,0.44894236,0.40367088,0.31312788,0.27540162,0.20372175,0.19240387,0.19240387,0.19994913,0.23390275,0.26408374,0.26031113,0.21503963,0.150905,0.12826926,0.241448,0.3055826,0.28294688,0.20749438,0.16222288,0.26408374,0.27540162,0.33953625,0.513077,0.77338815,1.2525115,0.9318384,0.5281675,0.33576363,0.29803738,0.0,0.0,0.0,0.00754525,0.0150905,0.0,0.0,0.0,0.0,0.02263575,0.10940613,0.23390275,0.1358145,0.030181,0.00754525,0.03772625,0.0150905,0.003772625,0.0,0.0,0.0,0.030181,0.16222288,0.32444575,0.38103512,0.15467763,0.11317875,0.041498873,0.0,0.011317875,0.06413463,0.049044125,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.00754525,0.0,0.0452715,0.2263575,0.1659955,0.060362,0.003772625,0.018863125,0.049044125,0.05281675,0.090543,0.14713238,0.27540162,0.59607476,1.3996439,0.90920264,0.49421388,0.6828451,1.146878,0.59230214,0.271629,0.15467763,0.5357128,2.0258996,0.67152727,0.2263575,0.11317875,0.049044125,0.0150905,0.003772625,0.0,0.0,0.003772625,0.026408374,0.116951376,0.0754525,0.02263575,0.00754525,0.00754525,0.0,0.0,0.00754525,0.018863125,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.06790725,0.0,0.0,0.15845025,0.49044126,0.73188925,0.36594462,0.15467763,0.041498873,0.0,0.150905,0.754525,0.150905,0.15467763,0.30935526,0.44894236,0.68661773,0.4074435,1.4222796,2.474842,3.0520537,3.361409,2.9313297,4.1762958,4.9044123,4.357382,3.240685,3.4783602,3.7575345,3.4066803,2.806833,3.399135,5.093044,3.4896781,2.7879698,5.2892203,11.385782,7.1868505,3.863168,2.305074,2.4371157,3.199186,2.1503963,1.4524606,1.7769064,3.0897799,4.659192,4.055572,3.8480775,3.3236825,2.7653341,3.440634,5.4967146,3.5160866,1.3920987,0.98842776,2.1051247,1.8900851,1.6939086,2.323937,3.31991,2.9539654,2.4371157,2.7011995,2.9313297,2.8106055,2.5201135,2.4974778,2.323937,2.5087957,3.2369123,4.38379,3.2105038,2.093807,1.7278622,1.9806281,1.9240388,3.7235808,3.663219,2.9351022,2.4786146,3.0256453,3.1161883,2.372981,1.9881734,2.071171,1.659955,2.6144292,2.565385,2.0636258,1.5958204,1.569412,1.4335974,1.1506506,1.026154,1.1053791,1.177059,1.0336993,0.8601585,0.73566186,0.694163,0.73188925,0.6752999,0.83752275,0.95447415,0.9280658,0.8111144,0.67152727,0.784706,0.8865669,1.0223814,1.5467763,2.5993385,4.376245,5.0477724,4.5422406,4.52715,6.085244,6.379509,6.247467,6.4511886,7.673519,9.491924,8.228095,5.9192486,4.772371,7.1566696,6.8397694,6.4511886,11.159425,17.391802,12.815607,8.099826,5.8626595,5.1156793,7.0812173,15.16218,23.767538,16.644821,7.8734684,4.610148,7.0849895,7.8432875,9.880505,10.231359,8.578949,7.273621,6.2361493,6.688864,6.9227667,5.832478,2.897376,3.9122121,10.084227,14.830189,14.637785,9.0957985,4.9459114,5.455216,6.907676,7.5075235,7.3717093,7.1906233,6.8963585,6.515323,6.771862,9.107117,9.450426,6.6020937,4.432834,4.768598,7.3868,18.38023,17.757746,16.293968,18.62545,23.246916,27.943834,32.19181,36.71896,40.67644,41.6611,61.346657,98.09957,129.67644,139.15327,114.9632,76.85214,61.61074,61.173115,67.82048,74.16226,68.284515,61.158024,51.688736,41.355515,34.187527,29.517017,25.66894,24.363613,24.933279,24.314568,23.914669,20.862616,16.87118,13.913441,14.222796,15.237633,12.626976,9.891823,8.201687,6.3945994,6.1229706,5.292993,4.2517486,3.4330888,3.3538637,2.8106055,2.2786655,2.1088974,2.1843498,1.9429018,1.3053282,0.7582976,0.36594462,0.18485862,0.2565385,0.31312788,0.44894236,0.452715,0.331991,0.32444575,0.48666862,0.34330887,0.14335975,0.049044125,0.12826926,0.29803738,0.4074435,0.5281675,0.6111652,0.5017591,1.3355093,1.3958713,1.3430545,1.448688,1.5731846,1.9051756,1.8561316,1.5203679,1.146878,1.1280149,1.0978339,0.8186596,0.47912338,0.21503963,0.120724,0.071679875,0.06413463,0.08677038,0.1056335,0.049044125,0.0150905,0.018863125,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.033953626,0.09808825,0.2867195,0.5772116,0.8941121,1.1053791,1.0223814,1.0487897,1.2940104,1.7769064,2.4182527,1.8297231,1.3996439,1.4147344,1.6675003,1.4335974,0.8903395,0.3961256,0.1056335,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.094315626,0.16222288,0.17354076,0.1358145,0.120724,0.18863125,0.23013012,0.181086,0.0754525,0.030181,0.041498873,0.05281675,0.06413463,0.07922512,0.10940613,0.30181,0.44516975,0.4979865,0.4640329,0.4074435,0.44139713,0.32067314,0.26408374,0.30181,0.30935526,0.124496624,0.049044125,0.033953626,0.03772625,0.02263575,0.02263575,0.03772625,0.20749438,0.49421388,0.6752999,0.7205714,0.42630664,0.16976812,0.094315626,0.10186087,0.18863125,0.26031113,0.35462674,0.4376245,0.4074435,0.3169005,0.33576363,0.4376245,0.62248313,0.90543,1.0412445,0.97710985,0.84129536,0.7092535,0.5998474,0.331991,0.16222288,0.07922512,0.049044125,0.0452715,0.05281675,0.049044125,0.03772625,0.02263575,0.011317875,0.0150905,0.0150905,0.011317875,0.011317875,0.0150905,0.02263575,0.026408374,0.03772625,0.049044125,0.06790725,0.056589376,0.05281675,0.049044125,0.0452715,0.05281675,0.041498873,0.030181,0.026408374,0.018863125,0.0150905,0.0150905,0.05281675,0.10940613,0.1659955,0.21503963,0.26031113,0.26031113,0.23013012,0.18485862,0.1358145,0.150905,0.16222288,0.16976812,0.16976812,0.1961765,0.30181,0.40367088,0.41121614,0.33953625,0.31312788,0.23013012,0.1961765,0.181086,0.17354076,0.20372175,0.22258487,0.241448,0.21881226,0.16222288,0.10940613,0.1961765,0.27540162,0.27917424,0.211267,0.150905,0.18485862,0.18863125,0.24899325,0.41498876,0.724344,0.573439,0.482896,0.3961256,0.29049212,0.16222288,0.011317875,0.003772625,0.0,0.0150905,0.030181,0.0,0.0,0.0,0.011317875,0.03772625,0.071679875,0.0150905,0.07922512,0.07922512,0.0150905,0.071679875,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.0754525,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.030181,0.0,0.07922512,0.38858038,0.3734899,0.14713238,0.0,0.0150905,0.08299775,0.1056335,0.27540162,0.44516975,0.6451189,1.086516,2.2711203,1.5543215,0.5319401,0.018863125,0.02263575,0.0452715,0.056589376,0.08677038,0.13204187,0.17731337,0.116951376,0.09808825,0.09808825,0.08677038,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.07922512,0.05281675,0.0150905,0.0,0.0,0.0,0.0,0.011317875,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.17731337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026408374,0.1358145,0.026408374,0.17731337,0.19994913,0.049044125,0.0,0.0,2.2107582,3.8367596,3.9348478,3.4179983,2.3578906,3.0520537,3.2746384,2.535204,2.0749438,2.7653341,3.2859564,2.7313805,1.5354583,1.4675511,2.1579416,2.3126192,2.6521554,5.3571277,14.056801,11.740409,5.5495315,1.6976813,1.8070874,2.8936033,2.9766011,2.0787163,1.9957186,3.048281,4.06689,3.640583,3.138824,2.4974778,2.4710693,4.636556,6.126743,3.6556737,1.4939595,1.4750963,3.0105548,2.938875,2.2371666,2.033445,2.4333432,2.5389767,2.493705,2.4559789,2.3805263,2.5578396,3.591539,2.3805263,2.335255,2.9766011,3.7084904,3.8141239,2.5201135,1.7391801,1.7844516,2.3088465,2.293756,3.3048196,3.199186,2.4672968,2.2447119,4.304565,3.2520027,2.0447628,1.4977322,1.5618668,1.3128735,3.180323,2.6408374,1.8259505,1.5958204,1.5543215,1.2449663,0.94692886,0.9242931,1.1204696,1.1431054,0.9620194,0.875249,0.8337501,0.8224323,0.87147635,0.73566186,0.8941121,1.1506506,1.2751472,0.9922004,1.0714256,1.2940104,1.3770081,1.6410918,3.0143273,3.0030096,4.0178456,4.2630663,3.832987,4.696918,6.5455046,6.851087,7.575431,9.137298,10.412445,9.122208,5.7381625,3.7650797,5.80607,13.562587,11.668729,9.922004,16.893814,26.672459,18.885761,7.273621,3.0445085,4.2291126,9.559832,18.489635,24.903097,15.618668,7.3905725,6.470052,8.624221,10.487898,15.030138,13.853079,7.175533,3.7952607,3.3651814,4.9044123,6.4964604,6.398372,3.0407357,4.7648253,11.536687,15.124454,12.37421,5.20245,4.1762958,6.862405,8.548768,7.1679873,3.2935016,5.6476197,5.594803,4.587512,4.134797,5.794752,5.9494295,4.6214657,4.323428,6.0776987,9.4013815,18.1086,18.293459,16.618414,16.550507,18.372684,20.006231,22.582933,26.64605,31.44483,34.93451,55.18973,93.21402,133.60751,159.9593,154.88889,105.17701,74.222626,60.897713,59.245304,58.430416,58.241783,55.898983,50.598446,43.622864,38.307236,33.365097,28.78513,27.732567,28.739857,25.714212,23.95617,22.92247,20.028866,15.788436,13.7851715,14.317112,12.774108,11.521597,10.680302,8.103599,6.5341864,5.4703064,4.727099,4.123479,3.4896781,2.8596497,1.9278114,1.569412,1.8636768,2.0673985,1.1959221,0.59230214,0.2678564,0.17354076,0.19994913,0.30181,0.3772625,0.42630664,0.4376245,0.3734899,0.27540162,0.17731337,0.116951376,0.10940613,0.14713238,0.18485862,0.241448,0.3055826,0.33576363,0.29426476,0.69039035,1.116697,1.0223814,0.60362,0.8262049,0.70170826,0.7884786,0.724344,0.4678055,0.26408374,0.3470815,0.5583485,0.573439,0.3961256,0.32821837,0.181086,0.10940613,0.07922512,0.08677038,0.14713238,0.049044125,0.041498873,0.041498873,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.011317875,0.011317875,0.026408374,0.09808825,0.27917424,0.6073926,1.1016065,1.1016065,1.177059,1.4713237,2.123988,3.2746384,2.3465726,1.6033657,1.3053282,1.3091009,1.0789708,0.62248313,0.35839936,0.19240387,0.0754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.011317875,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.026408374,0.026408374,0.026408374,0.03772625,0.071679875,0.1961765,0.20372175,0.14335975,0.06413463,0.033953626,0.041498873,0.049044125,0.05281675,0.06413463,0.1056335,0.271629,0.38103512,0.41876137,0.3961256,0.35085413,0.331991,0.24522063,0.18485862,0.19994913,0.2867195,0.15845025,0.071679875,0.033953626,0.026408374,0.0150905,0.018863125,0.026408374,0.033953626,0.071679875,0.18485862,0.38858038,0.362172,0.25276586,0.1659955,0.150905,0.26408374,0.3055826,0.2565385,0.17354076,0.181086,0.1961765,0.23767537,0.27540162,0.36594462,0.63002837,0.84884065,0.91297525,0.86770374,0.7922512,0.7809334,0.62625575,0.42630664,0.24899325,0.13204187,0.094315626,0.11317875,0.13204187,0.116951376,0.071679875,0.0452715,0.030181,0.018863125,0.00754525,0.003772625,0.0150905,0.0150905,0.02263575,0.03772625,0.05281675,0.071679875,0.06413463,0.060362,0.056589376,0.049044125,0.056589376,0.049044125,0.049044125,0.041498873,0.030181,0.02263575,0.0150905,0.02263575,0.049044125,0.1056335,0.20749438,0.2867195,0.29803738,0.2678564,0.211267,0.150905,0.11317875,0.120724,0.16222288,0.19994913,0.19994913,0.22258487,0.31312788,0.3734899,0.362172,0.32067314,0.28294688,0.23013012,0.18863125,0.18485862,0.21881226,0.23767537,0.23013012,0.19994913,0.15845025,0.1358145,0.181086,0.24522063,0.26031113,0.21503963,0.1659955,0.1659955,0.12826926,0.11317875,0.17354076,0.35462674,0.97710985,0.573439,0.26408374,0.150905,0.16976812,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.120724,0.0,0.0,0.10940613,0.10940613,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15845025,0.07922512,0.0,0.0452715,0.23013012,0.30181,0.12826926,0.0,0.02263575,0.1056335,0.27917424,0.694163,0.935611,0.9393836,1.0374719,2.1353056,1.6222287,0.663982,0.011317875,0.0,0.0,0.00754525,0.08299775,0.150905,0.030181,0.030181,0.041498873,0.11317875,0.17731337,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09808825,0.1961765,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.049044125,0.0,0.0,0.9507015,1.6863633,1.8938577,2.1353056,1.0751982,1.4034165,1.6675003,1.4524606,1.4034165,1.539231,1.81086,1.750498,1.3355093,0.9922004,2.1503963,2.093807,1.4939595,1.7278622,4.851596,8.601585,5.7570257,2.3993895,1.6222287,3.5387223,4.112161,2.7917426,2.916239,4.0517993,2.0145817,2.7728794,2.4559789,1.8599042,1.961765,3.953711,4.025391,2.625747,1.1581959,0.5319401,1.1280149,3.9612563,2.637065,1.3128735,1.6373192,2.746471,3.440634,3.048281,3.4632697,4.6554193,4.6554193,3.531177,3.8707132,5.172269,6.047518,4.2404304,1.629774,1.2789198,1.780679,2.1843498,2.0145817,3.6028569,3.92353,3.5160866,3.5085413,5.643847,3.6669915,2.1466236,1.539231,1.7278622,2.0447628,2.7879698,2.1956677,1.8749946,2.1994405,2.335255,1.4675511,1.0676528,1.2562841,1.5958204,1.0827434,0.9507015,0.8865669,0.9016574,0.9318384,0.87147635,0.8337501,1.6373192,2.4371157,2.6521554,1.9693103,2.9464202,2.3390274,1.7014539,1.9881734,3.5387223,2.9916916,3.0256453,3.2331395,4.014073,6.5756855,8.737399,10.11818,11.955449,12.989148,9.461743,5.50426,3.5274043,2.4484336,3.31991,9.337247,6.126743,4.847823,10.570895,17.91997,11.11038,4.7610526,3.3576362,4.6327834,6.9152217,9.125979,6.330465,5.2175403,6.9227667,11.359374,17.240896,9.529651,7.2698483,5.96452,3.7198083,1.267602,2.9766011,6.0022464,7.7678347,7.254758,5.0213637,4.055572,5.8211603,7.8206515,8.171506,5.5683947,9.035437,10.178542,8.620448,5.0251365,1.0827434,6.013564,6.900131,5.775889,4.5007415,4.745962,5.0741806,4.0404816,4.949684,8.816625,14.358611,10.902886,10.314357,11.487643,12.830698,12.268577,13.268322,16.120426,20.734346,27.596752,37.763977,56.95532,86.85715,114.93302,136.78784,156.1565,128.03157,101.06863,81.59811,69.6087,58.74732,52.190495,46.10525,42.807976,42.215675,41.823322,36.194565,30.878935,30.429993,33.11233,30.91289,27.2044,24.21648,19.425245,14.358611,14.603831,14.43029,13.400364,12.294985,11.193378,9.461743,7.8017883,7.3377557,6.94163,6.089017,4.8666863,3.440634,1.9844007,1.3015556,1.418507,1.6033657,1.0638802,0.6451189,0.33576363,0.17731337,0.27540162,0.33576363,0.34330887,0.3470815,0.3470815,0.27540162,0.13958712,0.20749438,0.29426476,0.32821837,0.36594462,0.2565385,0.18485862,0.19994913,0.24522063,0.120724,0.20749438,0.40367088,0.42630664,0.32821837,0.47157812,0.33953625,0.663982,0.8941121,0.76207024,0.27540162,0.5055317,0.70170826,0.7130261,0.694163,1.0978339,0.3055826,0.07922512,0.060362,0.16976812,0.6111652,0.16976812,0.041498873,0.03772625,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.018863125,0.03772625,0.0,0.02263575,0.0754525,0.13204187,0.271629,0.68661773,1.1242423,1.539231,1.8863125,2.04099,1.7844516,1.3468271,0.98842776,0.76207024,0.6149379,0.3961256,0.24899325,0.35085413,0.35085413,0.17731337,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.0452715,0.094315626,0.1358145,0.13958712,0.1056335,0.0452715,0.0452715,0.06413463,0.08299775,0.1056335,0.150905,0.24899325,0.29426476,0.34330887,0.39989826,0.41121614,0.362172,0.2678564,0.1659955,0.090543,0.090543,0.17731337,0.116951376,0.049044125,0.026408374,0.0150905,0.026408374,0.030181,0.030181,0.049044125,0.120724,0.16976812,0.26408374,0.31312788,0.28294688,0.19994913,0.331991,0.3470815,0.27540162,0.1659955,0.1056335,0.14335975,0.26408374,0.31312788,0.26408374,0.21503963,0.38480774,0.4376245,0.48666862,0.6111652,0.8526133,0.9016574,0.80734175,0.55457586,0.25276586,0.1056335,0.19240387,0.29426476,0.271629,0.14335975,0.1056335,0.08299775,0.041498873,0.00754525,0.003772625,0.0150905,0.0150905,0.02263575,0.03772625,0.049044125,0.060362,0.060362,0.060362,0.060362,0.056589376,0.0452715,0.056589376,0.060362,0.056589376,0.0452715,0.0452715,0.02263575,0.0150905,0.02263575,0.03772625,0.060362,0.16976812,0.26408374,0.29426476,0.26031113,0.19994913,0.11317875,0.071679875,0.071679875,0.1056335,0.150905,0.1659955,0.1961765,0.26408374,0.331991,0.32067314,0.28294688,0.23767537,0.20749438,0.20749438,0.24522063,0.27917424,0.23390275,0.181086,0.14713238,0.120724,0.15845025,0.17731337,0.17731337,0.1659955,0.150905,0.1056335,0.090543,0.090543,0.09808825,0.120724,0.41498876,0.17731337,0.18863125,0.4640329,0.7922512,0.7205714,0.14335975,0.0,0.0,0.0,0.0,0.0,0.27917424,0.8337501,1.2789198,0.8526133,0.16976812,0.02263575,0.060362,0.07922512,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.0452715,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.10940613,0.14335975,0.17731337,0.2263575,0.241448,0.13204187,0.23390275,0.35839936,0.47912338,0.513077,0.32821837,0.44894236,0.43007925,0.31312788,0.19240387,0.23013012,0.452715,0.35839936,0.15845025,0.02263575,0.049044125,0.018863125,0.00754525,0.0150905,0.030181,0.00754525,0.00754525,0.0452715,0.07922512,0.0754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.094315626,0.0452715,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.11317875,0.16976812,0.38480774,0.17731337,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.08677038,0.25276586,0.33576363,0.3169005,0.31312788,0.5998474,0.2263575,0.3961256,0.6073926,0.77338815,1.2223305,0.84129536,1.146878,1.4109617,1.4449154,1.5618668,1.3845534,1.2261031,1.2147852,1.5882751,2.7125173,4.4894238,3.1916409,1.3543724,0.6790725,2.0447628,5.9984736,6.3908267,5.3344917,4.093298,3.1010978,4.006528,3.874486,5.081726,6.56814,3.8556228,2.425798,1.6675003,1.2411937,1.2789198,2.3880715,2.5125682,2.214531,1.4335974,0.7809334,1.5430037,4.825187,2.806833,1.1883769,1.81086,2.637065,3.8292143,3.7801702,4.5761943,5.994701,5.4967146,3.610402,4.172523,5.8136153,6.628502,4.168751,2.5125682,1.4260522,1.6675003,2.7615614,2.9916916,4.168751,4.036709,3.802806,3.8480775,3.731126,3.127506,3.4632697,3.5500402,3.0369632,2.3880715,2.4371157,2.6898816,2.806833,2.746471,2.7615614,2.1503963,2.3616633,4.45547,6.1644692,1.901403,1.2298758,1.4750963,2.1503963,2.5767028,1.8825399,1.7014539,4.4516973,5.511805,3.983892,2.7238352,3.651901,3.31991,2.8256962,2.9049213,3.9197574,4.3649273,4.6742826,5.5797124,7.0774446,8.431817,7.8206515,7.907422,8.14887,7.6886096,5.372218,4.4516973,3.712263,3.1614597,4.2291126,9.7296,7.6697464,5.5080323,5.794752,6.9680386,3.3689542,2.987919,8.590267,11.291467,9.171251,7.2698483,5.323174,4.006528,7.77538,14.634012,16.143063,6.952948,6.511551,6.458734,4.1800685,2.7917426,6.092789,11.106608,12.340257,9.318384,6.6058664,5.4476705,6.511551,8.903395,10.695392,8.914713,8.8769865,7.0472636,4.4743333,2.425798,2.3880715,9.673011,10.597303,7.273621,3.0860074,2.6936543,4.90064,4.7950063,6.3531003,11.974312,22.4773,10.008774,7.5301595,8.707218,10.197406,11.657412,14.173752,16.324148,19.48561,25.001186,34.202618,47.980244,61.874825,73.03047,85.476364,110.13047,112.63549,104.252716,91.87851,79.34585,67.38663,59.075535,49.749607,42.69857,39.26548,38.846718,37.42821,34.66288,34.670425,35.77203,30.4979,28.24187,25.985842,21.692595,16.51278,14.7736,15.803526,14.362384,12.989148,12.415709,11.570641,11.563096,11.212241,9.948412,8.265821,7.748972,5.243949,3.1614597,2.0258996,1.6675003,1.237421,0.91297525,0.7696155,0.56589377,0.34330887,0.422534,0.69793564,0.56589377,0.543258,0.663982,0.49421388,0.1358145,0.10186087,0.17354076,0.24899325,0.35462674,0.56589377,0.3961256,0.41121614,0.67152727,0.7432071,0.5470306,0.5319401,0.3961256,0.17354076,0.241448,0.41121614,0.6752999,0.6488915,0.331991,0.12826926,0.23390275,0.2867195,0.26031113,0.20372175,0.2565385,0.07922512,0.026408374,0.0452715,0.11317875,0.27917424,0.49421388,0.3470815,0.1358145,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.00754525,0.018863125,0.02263575,0.011317875,0.033953626,0.060362,0.090543,0.1056335,0.060362,0.056589376,0.041498873,0.049044125,0.12826926,0.36971724,1.2298758,1.6637276,1.5052774,0.9808825,0.73566186,0.5093044,0.331991,0.21881226,0.15467763,0.090543,0.05281675,0.1056335,0.120724,0.06790725,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.011317875,0.0150905,0.018863125,0.033953626,0.05281675,0.094315626,0.11317875,0.09808825,0.0452715,0.056589376,0.08299775,0.1056335,0.13958712,0.23767537,0.3055826,0.27540162,0.31312788,0.4074435,0.35085413,0.28294688,0.26408374,0.20372175,0.13204187,0.19994913,0.150905,0.09808825,0.120724,0.20749438,0.271629,0.18485862,1.4373702,1.6750455,0.6413463,0.20749438,0.120724,0.1056335,0.1358145,0.181086,0.22258487,0.23013012,0.20749438,0.17354076,0.14713238,0.14335975,0.19994913,0.27917424,0.31312788,0.2867195,0.23767537,0.22258487,0.20749438,0.2263575,0.32067314,0.52439487,0.69039035,0.7394345,0.69039035,0.55080324,0.32821837,0.20749438,0.23767537,0.271629,0.24899325,0.19240387,0.14713238,0.094315626,0.05281675,0.033953626,0.0150905,0.0150905,0.018863125,0.02263575,0.03772625,0.049044125,0.049044125,0.056589376,0.060362,0.060362,0.056589376,0.060362,0.060362,0.060362,0.056589376,0.0452715,0.030181,0.026408374,0.03772625,0.060362,0.08677038,0.12826926,0.18863125,0.23013012,0.24522063,0.22258487,0.20749438,0.14713238,0.08677038,0.060362,0.07922512,0.150905,0.2263575,0.28294688,0.33576363,0.43007925,0.43385187,0.3470815,0.2678564,0.23013012,0.21881226,0.18863125,0.15467763,0.13958712,0.13958712,0.1358145,0.120724,0.120724,0.116951376,0.1056335,0.1056335,0.08299775,0.071679875,0.071679875,0.07922512,0.08677038,0.24899325,0.116951376,0.18863125,0.62625575,1.1619685,1.0789708,0.21503963,0.0,0.0,0.018863125,0.090543,0.21503963,1.1016065,2.354118,3.0218725,1.5882751,0.4074435,0.14713238,0.181086,0.15467763,0.0,0.0,0.0,0.0,0.0,0.0,0.05281675,0.03772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.056589376,0.056589376,0.07922512,0.13958712,0.1961765,0.18863125,0.5772116,0.66775465,0.6149379,0.5583485,0.5998474,1.2449663,0.69793564,0.16222288,0.06413463,0.030181,0.02263575,0.018863125,0.0150905,0.011317875,0.033953626,0.026408374,0.011317875,0.0,0.0,0.0,0.0452715,0.06413463,0.049044125,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.049044125,0.02263575,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.03772625,0.08677038,0.19240387,0.15467763,0.06413463,0.0,0.0,0.0,0.0,0.030181,0.07922512,0.1056335,0.13958712,0.16976812,0.15467763,0.23013012,0.6828451,0.482896,0.29803738,0.34330887,0.83752275,2.0258996,1.0072908,1.1431054,1.5807298,1.9768555,2.516341,1.448688,0.8601585,0.875249,1.4373702,2.3201644,3.399135,2.372981,1.327964,1.3807807,2.6597006,4.6818275,6.115425,6.692637,5.9607477,3.3123648,2.2862108,2.3805263,4.6554193,7.149124,4.878004,2.2107582,1.3241913,1.1280149,1.1808317,1.6675003,1.7957695,1.9391292,1.5165952,0.9242931,1.5015048,3.187868,2.252257,2.093807,3.4179983,4.221567,3.9725742,3.6783094,4.063117,4.708236,4.0480266,2.9124665,3.6368105,4.90064,5.2552667,3.1350515,1.7467253,1.2261031,1.9240388,3.270866,3.7763977,4.036709,4.0895257,4.636556,5.0251365,3.259548,4.3007927,5.1232247,4.870459,3.5424948,2.003264,1.9994912,1.9768555,2.161714,2.5578396,2.9313297,3.240685,2.8256962,3.7235808,5.0779533,3.169005,1.871222,2.3993895,3.3161373,3.5349495,2.3013012,2.233394,3.0218725,3.4330888,3.31991,3.6028569,4.398881,3.7348988,2.655928,2.3578906,4.195159,6.2399216,6.1606965,6.126743,6.5455046,6.047518,6.360646,8.152642,8.00551,5.560849,3.4783602,2.7841973,2.3993895,3.9763467,7.779153,12.683565,9.016574,7.0849895,5.7306175,4.0103,1.2223305,4.38379,10.072908,10.631257,6.326692,5.323174,5.9192486,5.138315,6.6322746,9.865415,10.121953,10.808571,15.656394,14.958458,8.084735,3.5047686,7.2887115,10.084227,9.371201,6.330465,5.80607,5.3948536,6.670001,9.0543,10.20495,6.0248823,4.67051,3.229367,3.4217708,5.5797124,8.627994,10.065364,7.7112455,4.398881,2.3578906,3.218049,6.4738245,6.1644692,5.6400743,7.360391,12.879742,8.284684,8.605357,10.125726,12.555296,19.029121,15.886524,15.275358,17.859608,22.865881,28.08342,34.489338,39.672924,44.0039,52.15654,73.13233,87.879524,90.38455,86.19316,78.621506,68.76363,59.086853,49.29689,42.102493,37.903564,34.787376,33.527317,34.213936,34.13094,31.512737,25.506718,27.227036,26.283878,23.703403,20.96825,20.006231,17.293713,15.147089,13.841762,13.091009,12.045992,12.193124,12.483616,11.966766,10.506761,8.778898,5.847569,3.7499893,2.927557,2.9011486,2.2711203,1.5467763,1.1695137,0.95447415,0.7696155,0.55080324,0.6451189,0.6752999,0.76207024,0.77716076,0.33953625,0.1358145,0.09808825,0.12826926,0.1961765,0.331991,0.60362,0.5696664,0.63002837,0.87147635,1.0638802,0.88279426,0.91674787,0.8865669,0.7432071,0.66775465,0.663982,0.91674787,0.8978847,0.66775465,0.87902164,1.3619176,1.5543215,1.0676528,0.2565385,0.23013012,0.13204187,0.05281675,0.02263575,0.041498873,0.08677038,0.24899325,0.26031113,0.2263575,0.1659955,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.02263575,0.0150905,0.00754525,0.02263575,0.026408374,0.026408374,0.033953626,0.041498873,0.090543,0.1056335,0.15467763,0.21503963,0.1961765,0.124496624,0.06790725,0.0452715,0.1056335,0.33576363,0.7054809,0.86770374,0.7130261,0.38103512,0.25276586,0.16222288,0.08299775,0.033953626,0.0150905,0.00754525,0.0,0.018863125,0.030181,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.00754525,0.018863125,0.026408374,0.030181,0.041498873,0.09808825,0.10940613,0.06413463,0.0452715,0.071679875,0.116951376,0.13204187,0.14713238,0.2867195,0.31312788,0.25276586,0.25276586,0.32821837,0.3734899,0.32067314,0.38103512,0.31312788,0.1659955,0.26408374,0.3055826,0.43007925,0.6526641,1.1053791,2.0560806,1.4562333,1.4034165,1.2110126,0.7394345,0.41121614,0.20372175,0.1056335,0.07922512,0.090543,0.12826926,0.116951376,0.10940613,0.120724,0.150905,0.19994913,0.47912338,0.8299775,1.0110635,0.90920264,0.5357128,0.30935526,0.18863125,0.150905,0.18485862,0.2678564,0.3470815,0.41876137,0.48666862,0.5394854,0.56589377,0.39989826,0.29803738,0.2565385,0.24522063,0.21503963,0.19994913,0.181086,0.13958712,0.090543,0.041498873,0.02263575,0.0150905,0.018863125,0.02263575,0.026408374,0.026408374,0.03772625,0.049044125,0.06413463,0.07922512,0.071679875,0.0754525,0.08299775,0.08677038,0.08299775,0.07922512,0.071679875,0.07922512,0.1056335,0.1358145,0.17731337,0.19994913,0.22258487,0.24522063,0.24899325,0.211267,0.1659955,0.11317875,0.06790725,0.05281675,0.10186087,0.16222288,0.23390275,0.30935526,0.35839936,0.3772625,0.362172,0.3169005,0.24899325,0.20372175,0.14713238,0.116951376,0.1056335,0.116951376,0.1358145,0.1358145,0.11317875,0.090543,0.07922512,0.071679875,0.060362,0.049044125,0.05281675,0.0754525,0.1056335,0.44139713,0.1659955,0.1358145,0.41498876,0.7922512,0.77338815,0.15467763,0.0,0.011317875,0.08677038,0.34330887,1.2713746,2.837014,3.85185,3.5047686,1.358145,0.35839936,0.14713238,0.16222288,0.116951376,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.18485862,0.094315626,0.07922512,0.0754525,0.07922512,0.14713238,0.49044126,0.543258,0.6375736,0.8337501,0.9242931,1.3053282,0.72811663,0.31312788,0.30181,0.049044125,0.02263575,0.00754525,0.0,0.0,0.00754525,0.0150905,0.00754525,0.0,0.0,0.0,0.0452715,0.0452715,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06413463,0.08677038,0.0452715,0.0,0.0,0.0,0.060362,0.16222288,0.19240387,0.1358145,0.24899325,0.32444575,0.41876137,0.87147635,0.6790725,0.33576363,0.41121614,1.237421,2.9313297,1.9693103,2.022127,2.3013012,2.5880208,3.2821836,1.7995421,1.1657411,1.0186088,1.1393328,1.4335974,1.6637276,1.6448646,2.3654358,3.8367596,5.100589,4.0291634,4.2328854,5.111907,5.5797124,4.08198,1.5128226,1.2185578,3.4859054,6.1795597,4.7308717,2.2107582,1.7618159,1.8863125,1.9089483,1.9881734,1.7655885,1.8523588,1.4675511,0.8224323,1.1053791,1.5845025,2.897376,4.847823,6.2436943,4.8742313,3.4859054,3.2557755,3.270866,3.048281,2.5125682,2.1881225,2.7879698,3.4557245,3.4859054,2.335255,1.1657411,1.146878,2.8294687,5.1534057,5.4363527,4.587512,4.961002,6.2135134,6.828451,4.1197066,5.2967653,5.7419353,5.2288585,3.7386713,1.4600059,2.0673985,2.1994405,2.474842,2.9124665,2.9464202,3.5651307,2.7992878,2.584248,3.3915899,4.255521,2.5314314,2.9049213,3.5047686,3.361409,2.4220252,2.546522,2.4220252,2.5767028,3.2029586,4.1574326,5.0138187,4.187614,2.8106055,2.3013012,4.3724723,6.6813188,6.6360474,5.8098426,4.938366,3.9122121,6.934085,9.635284,9.035437,5.7419353,3.953711,2.6597006,1.9429018,3.832987,7.707473,10.26154,6.7680893,6.730363,6.3832817,4.3385186,1.5580941,5.4288073,10.416218,10.578441,6.4926877,5.2552667,6.5040054,6.647365,6.537959,6.3531003,5.6023483,11.234878,16.097792,14.7321005,8.284684,4.504514,7.164215,7.424526,5.643847,3.742444,5.198677,6.0701537,7.4811153,8.959985,8.737399,3.7348988,3.361409,5.2175403,7.54525,9.307066,10.174769,7.383027,4.2706113,3.3274553,4.4441524,4.9421387,6.0776987,5.745708,4.636556,3.8103511,4.6742826,16.21097,13.517315,10.774617,14.332202,22.692339,17.757746,14.871688,15.150862,18.070873,21.436056,24.042938,26.597006,29.988596,36.669914,50.624855,64.855194,71.30639,74.68666,75.34686,69.28049,63.217876,54.69929,46.82582,40.646263,35.160866,31.686277,32.29367,32.199356,29.5472,25.401085,26.412148,25.834936,24.888006,24.20139,23.77131,18.719765,16.45619,15.513034,14.532151,12.264804,12.630749,13.347548,13.245687,11.910177,9.665465,6.7454534,4.817642,4.6026025,5.093044,3.519859,2.8822856,2.3390274,1.7655885,1.2147852,0.9205205,0.87147635,1.0223814,1.1808317,1.0751982,0.38858038,0.41498876,0.4074435,0.33953625,0.27917424,0.39989826,0.7507524,0.965792,1.0638802,1.2034674,1.6750455,1.6637276,1.6712729,1.6561824,1.5203679,1.1129243,0.94315624,0.98465514,0.8941121,0.7582976,1.1053791,1.6863633,1.9579924,1.4034165,0.41498876,0.27917424,0.14713238,0.094315626,0.05281675,0.00754525,0.0150905,0.018863125,0.090543,0.1659955,0.1659955,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.030181,0.033953626,0.041498873,0.041498873,0.03772625,0.049044125,0.1056335,0.15845025,0.16222288,0.18863125,0.25276586,0.27917424,0.211267,0.12826926,0.071679875,0.090543,0.23767537,0.23390275,0.21881226,0.16976812,0.10186087,0.06413463,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.003772625,0.011317875,0.018863125,0.02263575,0.02263575,0.06413463,0.116951376,0.1056335,0.0452715,0.0452715,0.06790725,0.10940613,0.12826926,0.16222288,0.31312788,0.35839936,0.33953625,0.32444575,0.33953625,0.38480774,0.3772625,0.452715,0.41876137,0.32067314,0.422534,0.49421388,1.0827434,1.7052265,2.233394,2.9124665,1.9693103,1.2562841,0.995973,0.98465514,0.6073926,0.44516975,0.31312788,0.181086,0.071679875,0.056589376,0.060362,0.071679875,0.120724,0.21503963,0.33953625,1.0450171,1.8184053,2.191895,1.9466745,1.1242423,0.6413463,0.362172,0.23013012,0.18485862,0.14713238,0.14713238,0.181086,0.24899325,0.35839936,0.51684964,0.44894236,0.38480774,0.32067314,0.2565385,0.18863125,0.19240387,0.211267,0.21881226,0.1961765,0.14713238,0.090543,0.056589376,0.03772625,0.018863125,0.0150905,0.011317875,0.018863125,0.033953626,0.05281675,0.071679875,0.071679875,0.08677038,0.10940613,0.12826926,0.120724,0.120724,0.120724,0.1358145,0.1659955,0.19240387,0.22258487,0.20749438,0.20372175,0.21881226,0.24899325,0.20749438,0.16976812,0.12826926,0.08299775,0.0452715,0.060362,0.08299775,0.13958712,0.21503963,0.25276586,0.3169005,0.36594462,0.35462674,0.2867195,0.21503963,0.17354076,0.12826926,0.1358145,0.18485862,0.19994913,0.16976812,0.1358145,0.09808825,0.06790725,0.056589376,0.049044125,0.033953626,0.03772625,0.06790725,0.120724,0.62625575,0.1659955,0.026408374,0.00754525,0.018863125,0.09808825,0.018863125,0.0,0.018863125,0.18485862,0.7205714,2.8332415,4.5309224,4.304565,2.3163917,0.392353,0.10940613,0.049044125,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.36594462,0.41121614,0.3961256,0.2678564,0.08677038,0.02263575,0.018863125,0.10940613,0.573439,1.1846043,1.1959221,0.70170826,0.44516975,0.45648763,0.5583485,0.35462674,0.21881226,0.094315626,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0754525,0.15845025,0.041498873,0.00754525,0.0,0.06413463,0.17731337,0.2565385,0.24522063,0.55457586,0.7394345,0.80356914,1.1883769,0.80734175,0.39989826,0.5017591,1.3204187,2.757789,2.7200627,2.886058,2.867195,2.746471,3.1048703,2.0900342,1.6712729,1.2487389,0.80734175,0.9242931,0.935611,1.8938577,3.9197574,6.0626082,6.2851934,3.440634,1.7354075,1.9278114,3.5387223,4.851596,2.0108092,1.2525115,2.637065,4.6252384,4.0970707,2.5125682,2.4861598,2.776652,2.8558772,2.8936033,2.123988,1.9164935,1.4109617,0.66775465,0.65643674,1.0110635,4.1612053,7.1566696,7.6018395,3.6896272,2.916239,3.3048196,3.048281,2.0145817,1.7429527,1.9240388,2.2899833,2.5012503,2.4899325,2.4672968,1.5241405,1.267602,3.5538127,6.960493,6.7680893,5.1345425,5.5457587,6.990674,7.6697464,4.9647746,4.927048,4.9044123,4.6856003,3.8178966,1.5958204,2.9200118,3.7499893,4.115934,3.9650288,3.180323,3.0935526,2.5314314,2.354118,2.9766011,4.3649273,3.0181,3.097325,3.1350515,2.7426984,2.6106565,3.108643,3.893349,4.1800685,4.014073,4.293247,4.979865,4.4403796,3.572676,3.361409,4.8742313,5.975838,6.368191,5.624984,4.346064,4.142342,8.688355,10.137043,8.793989,6.2436943,5.330719,4.4139714,3.7235808,3.6783094,4.002755,3.7462165,3.6896272,6.217286,6.930312,4.7648253,2.003264,5.0439997,10.3634,12.14408,9.457971,6.258785,6.541732,7.360391,7.3113475,6.006019,4.0517993,6.224831,6.3719635,6.1116524,6.5643673,8.341274,7.805561,6.530414,4.9044123,4.0216184,5.674028,8.631766,9.665465,9.110889,7.17176,3.9197574,6.006019,11.249968,13.008011,9.922004,5.9230213,4.3649273,4.074435,6.0248823,8.3525915,6.3832817,3.772625,4.5460134,5.089271,4.485651,4.5422406,29.709421,19.836462,10.978339,15.049001,19.817598,17.904879,14.460471,12.15917,12.626976,16.444872,19.591242,23.02433,26.883726,31.882454,39.32207,47.795387,53.084606,60.788307,69.167305,69.1409,71.70628,66.60947,57.362762,47.13895,38.782585,31.878681,29.845236,30.309269,30.875162,29.139755,26.189562,25.778347,26.07261,25.887753,24.66165,20.670212,18.546225,17.437073,16.26756,13.766309,14.535924,14.675511,13.6833105,11.944131,10.718028,8.228095,6.8699503,7.115171,7.4584794,4.402653,4.6327834,4.187614,3.0558262,1.871222,1.9089483,1.7882242,1.81086,1.8900851,1.7429527,0.8865669,0.935611,0.8903395,0.694163,0.5055317,0.7054809,1.388326,1.901403,1.9579924,1.9164935,2.7804246,2.9954643,2.7502437,2.4710693,2.1768045,1.4750963,1.2336484,0.9997456,0.77716076,0.6111652,0.5998474,0.8262049,1.0487897,0.935611,0.5281675,0.23013012,0.11317875,0.14335975,0.116951376,0.0150905,0.011317875,0.003772625,0.003772625,0.0150905,0.026408374,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0,0.003772625,0.011317875,0.033953626,0.06413463,0.06413463,0.05281675,0.049044125,0.056589376,0.090543,0.18863125,0.23767537,0.21881226,0.1961765,0.20749438,0.27917424,0.2678564,0.16976812,0.08299775,0.0452715,0.03772625,0.060362,0.056589376,0.03772625,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.011317875,0.011317875,0.0150905,0.0150905,0.0150905,0.08677038,0.11317875,0.090543,0.0452715,0.0452715,0.0452715,0.060362,0.10186087,0.18485862,0.32821837,0.48666862,0.5696664,0.573439,0.51684964,0.41876137,0.43385187,0.4640329,0.5055317,0.5583485,0.663982,0.6073926,1.539231,2.463524,2.8030603,2.3993895,1.6109109,1.6033657,1.7014539,1.4713237,0.7394345,0.7205714,0.6790725,0.452715,0.13204187,0.049044125,0.056589376,0.06413463,0.13204187,0.27540162,0.45648763,1.5052774,2.6332922,3.1916409,2.8822856,1.7542707,1.0374719,0.6073926,0.3772625,0.2565385,0.150905,0.1358145,0.124496624,0.13204187,0.16222288,0.2263575,0.29049212,0.38858038,0.41121614,0.32821837,0.18863125,0.150905,0.18485862,0.24899325,0.30181,0.29426476,0.2263575,0.15467763,0.10186087,0.06413463,0.026408374,0.011317875,0.011317875,0.018863125,0.030181,0.041498873,0.056589376,0.08677038,0.13204187,0.1659955,0.150905,0.14713238,0.16222288,0.18863125,0.211267,0.22258487,0.22258487,0.18863125,0.1659955,0.1659955,0.20372175,0.1961765,0.16222288,0.124496624,0.08299775,0.049044125,0.0452715,0.033953626,0.041498873,0.08677038,0.1659955,0.271629,0.32444575,0.32821837,0.29426476,0.23390275,0.23390275,0.17731337,0.1961765,0.27540162,0.26408374,0.19994913,0.1659955,0.116951376,0.060362,0.0452715,0.041498873,0.02263575,0.02263575,0.056589376,0.120724,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21881226,1.0978339,3.6141748,3.893349,2.4182527,0.44139713,0.0,0.15845025,0.24522063,0.1659955,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1091517,1.177059,0.8299775,0.4376245,0.120724,0.09808825,0.10186087,0.25276586,0.62248313,1.2223305,0.9507015,0.4640329,0.15845025,0.392353,1.4637785,0.97710985,0.452715,0.10940613,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15845025,0.35839936,0.19994913,0.041498873,0.0,0.0,0.0,0.0,0.0,0.27540162,0.47157812,0.5998474,1.0525624,0.95447415,0.58475685,0.44894236,0.633801,0.7922512,0.84129536,1.3015556,1.7354075,1.8448136,1.478869,1.5430037,0.9808825,0.47157812,0.41121614,0.9016574,1.7316349,2.8709676,3.9763467,4.0895257,1.6486372,2.3088465,1.3091009,1.1996948,2.6785638,4.606375,1.8749946,1.3166461,2.3993895,4.0480266,4.6856003,3.2067313,2.1503963,1.9693103,2.565385,3.2972744,2.3805263,1.9957186,1.5505489,0.9620194,0.65643674,0.91297525,2.9615107,3.5990841,2.3465726,1.478869,3.7273536,4.881777,3.7160356,1.3505998,1.267602,2.3277097,2.9501927,3.048281,3.0181,3.7386713,2.4823873,1.2864652,2.161714,4.3385186,4.304565,2.9124665,2.746471,3.6858547,4.5761943,3.218049,2.6936543,3.1765501,3.62172,3.6481283,3.5236318,4.52715,5.270357,5.311856,4.768598,4.304565,2.9464202,2.1692593,2.1315331,2.5201135,2.5314314,3.2670932,3.92353,3.9688015,3.500996,3.2821836,4.745962,4.82896,4.353609,3.9876647,4.255521,3.440634,3.4179983,3.8895764,4.8365054,6.5455046,6.643593,6.760544,6.6360474,6.3908267,6.5002327,7.356619,6.405917,4.8968673,3.9386206,4.5007415,6.5530496,8.171506,6.4511886,2.9426475,3.663219,8.692128,11.970539,9.725827,3.651901,0.9318384,4.606375,8.756263,9.408927,6.673774,4.745962,6.541732,6.888813,5.5570765,3.31991,1.9542197,1.6373192,2.2069857,6.5040054,13.641812,19.010258,12.811834,9.684328,7.8621507,6.6360474,6.3945994,13.230596,13.483362,9.778644,5.240176,3.4934506,7.7678347,11.314102,10.065364,5.2288585,3.3123648,6.300284,8.661947,10.246449,9.997457,5.9192486,3.4066803,6.9869013,8.646856,6.8850408,6.7152724,30.165909,22.733839,16.335466,19.31584,16.448645,13.238141,10.853842,11.18206,13.698401,15.456445,19.462973,23.38273,24.333431,23.710949,27.17799,34.03662,36.01725,41.212154,51.454834,62.31622,74.022675,76.391884,68.89945,54.13717,37.779068,26.842226,25.985842,27.962696,28.27205,25.148317,25.061548,27.675978,29.471746,28.898308,26.381968,24.48811,21.217243,17.810562,16.048746,18.233097,18.28214,15.99593,12.823153,10.461489,10.86516,9.348565,9.831461,9.967276,8.431817,4.927048,6.319147,6.0550632,4.67051,3.361409,3.983892,3.5424948,3.059599,2.886058,2.7540162,1.7391801,1.3505998,1.0487897,0.80734175,0.80356914,1.448688,2.916239,3.7386713,3.5839937,3.1576872,4.195159,4.636556,3.9499383,3.1199608,2.5729303,2.1805773,1.6561824,1.5807298,1.5618668,1.2600567,0.38103512,0.23390275,0.482896,0.72811663,0.7432071,0.47157812,0.32821837,0.2263575,0.116951376,0.011317875,0.0,0.0,0.026408374,0.056589376,0.07922512,0.090543,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.011317875,0.05281675,0.124496624,0.17354076,0.0754525,0.06413463,0.060362,0.09808825,0.17731337,0.27540162,0.32444575,0.25276586,0.181086,0.1659955,0.23013012,0.23013012,0.120724,0.026408374,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.041498873,0.05281675,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.026408374,0.041498873,0.0452715,0.0452715,0.0452715,0.0452715,0.0452715,0.0754525,0.16976812,0.36594462,0.67152727,0.875249,0.9242931,0.8224323,0.62625575,0.55080324,0.5696664,0.6187105,0.68661773,0.80734175,0.5885295,0.7809334,1.2261031,1.7391801,2.1051247,2.0183544,2.3277097,2.323937,1.750498,0.8224323,0.7394345,1.0751982,0.8978847,0.23013012,0.060362,0.049044125,0.0452715,0.071679875,0.1358145,0.26031113,1.0299267,2.1277604,2.867195,2.8407867,1.9391292,1.1317875,0.7092535,0.4678055,0.29426476,0.19994913,0.124496624,0.116951376,0.120724,0.116951376,0.090543,0.12826926,0.211267,0.34330887,0.44516975,0.33576363,0.19994913,0.18485862,0.21503963,0.271629,0.38103512,0.36971724,0.29426476,0.24522063,0.211267,0.0754525,0.041498873,0.02263575,0.0150905,0.018863125,0.030181,0.041498873,0.08299775,0.13204187,0.17354076,0.19994913,0.18485862,0.18485862,0.18863125,0.19994913,0.19994913,0.19994913,0.181086,0.150905,0.120724,0.1056335,0.1056335,0.1056335,0.10186087,0.08677038,0.060362,0.03772625,0.02263575,0.02263575,0.033953626,0.0452715,0.071679875,0.1056335,0.1358145,0.16222288,0.19994913,0.23390275,0.2263575,0.16976812,0.116951376,0.150905,0.18863125,0.16222288,0.11317875,0.071679875,0.0452715,0.02263575,0.00754525,0.011317875,0.0452715,0.1056335,0.17354076,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0754525,0.3772625,1.478869,1.5731846,0.9695646,0.26408374,0.34330887,0.66775465,0.543258,0.24522063,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30935526,0.6375736,0.8337501,0.8526133,0.7809334,1.4901869,1.3732355,0.86770374,0.36971724,0.2565385,0.19240387,0.094315626,0.030181,0.10186087,0.40367088,0.724344,0.724344,0.47535074,0.14713238,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.11317875,0.24899325,0.049044125,0.0,0.03772625,0.10186087,0.10940613,0.02263575,0.056589376,0.29803738,0.68661773,0.9922004,0.543258,0.21503963,0.12826926,0.2565385,0.41498876,0.452715,0.5696664,0.80734175,1.0072908,0.80734175,0.995973,1.0450171,0.754525,0.32067314,0.33953625,0.7884786,1.297783,1.6976813,1.9278114,2.0636258,1.0525624,0.5017591,1.1808317,2.6144292,3.0709167,1.478869,1.1883769,3.1124156,6.0324273,6.587003,4.3875628,3.240685,2.8747404,2.9841464,3.199186,3.1425967,2.4069347,1.7618159,1.4864142,1.3770081,1.388326,1.539231,1.3430545,1.0676528,1.7240896,5.2892203,5.828706,3.863168,1.1317875,0.6073926,3.3576362,3.6481283,2.9803739,2.425798,2.6408374,2.505023,3.138824,3.7877154,4.0782075,4.0216184,3.3840446,2.746471,2.6483827,2.8294687,2.2560298,2.3767538,2.584248,3.2067313,3.62172,2.2786655,1.9240388,2.9652832,3.4859054,3.2255943,3.5839937,2.655928,2.4031622,2.7087448,3.0633714,2.5578396,2.4597516,3.9499383,4.8138695,4.3875628,3.572676,3.8556228,3.3425457,3.0520537,3.3764994,4.074435,4.1536603,4.1083884,4.115934,4.3083377,4.776143,6.0248823,6.0286546,6.643593,7.7301087,7.145352,5.0515447,4.1800685,4.4743333,5.198677,4.927048,4.938366,5.081726,3.640583,2.123988,5.2854476,13.019329,13.381501,8.575176,3.863168,7.54525,9.258021,7.6886096,6.017337,5.696664,6.4549613,9.273112,7.696155,5.666483,5.726845,9.009028,8.933576,11.6008215,17.316349,21.790682,16.16947,7.3717093,4.9647746,5.13077,5.1760416,3.5236318,4.5988297,5.0251365,4.032936,2.8294687,4.5799665,8.122461,10.042727,9.42779,7.413208,7.2057137,8.213005,8.76758,9.092027,9.235386,9.046755,7.564113,9.948412,9.310839,6.9491754,12.366665,30.52431,24.801237,16.524097,13.947394,12.249713,11.332966,13.124963,14.792462,15.445127,16.127972,17.074902,19.53088,21.949133,23.216734,22.658386,22.469755,24.586197,32.357803,46.373108,64.45152,80.94544,78.3876,66.4397,52.13013,39.85401,30.852528,27.37794,25.484081,22.865881,18.874443,20.964478,23.039421,23.371412,22.382984,22.658386,24.095757,23.560043,21.42851,19.421474,20.590988,22.77911,20.511763,16.35433,12.638294,11.487643,10.091772,11.472552,11.959221,10.212496,7.2358947,8.0206,7.4509344,5.798525,4.1083884,4.2027044,3.7537618,3.440634,3.7499893,4.0103,2.4107075,1.5920477,1.2223305,1.1431054,1.3770081,2.1315331,3.3048196,3.4029078,2.9049213,2.3465726,2.3390274,2.625747,2.5578396,2.263575,1.9957186,2.1315331,1.5316857,1.0751982,0.7582976,0.5357128,0.32067314,0.18485862,0.27917424,0.7922512,1.5241405,1.8900851,1.4411428,0.8978847,0.4074435,0.08299775,0.011317875,0.071679875,0.05281675,0.094315626,0.18863125,0.19994913,0.10186087,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0,0.02263575,0.071679875,0.22258487,0.42630664,0.51684964,0.2678564,0.1358145,0.08299775,0.090543,0.13958712,0.15845025,0.13204187,0.09808825,0.07922512,0.071679875,0.060362,0.041498873,0.018863125,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.03772625,0.06790725,0.08677038,0.10186087,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.003772625,0.003772625,0.0452715,0.049044125,0.0452715,0.049044125,0.056589376,0.049044125,0.05281675,0.08299775,0.18863125,0.452715,0.6111652,0.7054809,0.84129536,0.9620194,0.845068,0.95824677,1.3430545,1.2110126,0.68661773,0.80734175,0.84129536,0.7997965,1.50905,2.674791,2.8747404,2.1353056,1.6561824,1.358145,1.1431054,0.90920264,1.177059,1.539231,1.3241913,0.59230214,0.15845025,0.09808825,0.060362,0.071679875,0.1659955,0.4074435,0.6073926,0.94315624,1.1657411,1.177059,1.0336993,0.8526133,0.6187105,0.44139713,0.35462674,0.29426476,0.23390275,0.2263575,0.24522063,0.26031113,0.2263575,0.26408374,0.26408374,0.30935526,0.3961256,0.43385187,0.42630664,0.28294688,0.1961765,0.241448,0.36971724,0.4074435,0.392353,0.34330887,0.27540162,0.19994913,0.11317875,0.05281675,0.026408374,0.026408374,0.030181,0.06413463,0.1056335,0.14713238,0.16976812,0.17354076,0.150905,0.18485862,0.20749438,0.19994913,0.150905,0.15845025,0.1659955,0.15845025,0.1358145,0.094315626,0.0754525,0.071679875,0.06790725,0.06413463,0.049044125,0.0452715,0.041498873,0.041498873,0.041498873,0.0452715,0.030181,0.041498873,0.05281675,0.060362,0.08677038,0.14335975,0.18485862,0.17731337,0.13958712,0.12826926,0.14713238,0.14335975,0.11317875,0.071679875,0.056589376,0.02263575,0.0150905,0.0150905,0.02263575,0.033953626,0.116951376,0.02263575,0.0,0.0,0.0,0.0,0.0,0.08677038,0.116951376,0.0754525,0.07922512,0.3772625,0.3961256,0.29049212,0.28294688,0.663982,0.77338815,0.42630664,0.1056335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.29049212,0.47535074,0.663982,1.237421,1.5958204,1.1695137,0.8224323,0.663982,0.07922512,0.02263575,0.00754525,0.003772625,0.011317875,0.056589376,0.271629,0.32821837,0.25276586,0.116951376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12826926,0.6451189,0.12826926,0.10940613,0.18485862,0.15845025,0.056589376,0.011317875,0.0,0.10186087,0.28294688,0.392353,0.2263575,0.1961765,0.15467763,0.094315626,0.12826926,0.29049212,0.40367088,0.55080324,0.6526641,0.45648763,0.814887,1.4637785,1.2223305,0.2565385,0.07922512,0.22258487,0.41876137,1.1204696,2.1164427,2.5314314,1.0450171,0.32821837,0.5017591,1.1242423,1.2034674,0.9205205,0.9242931,2.4861598,5.1458607,6.7077274,5.1760416,4.568649,4.085753,3.8141239,4.7120085,4.798779,4.2102494,3.5160866,2.9351022,2.3616633,1.6524098,1.056335,0.6488915,0.7092535,1.7127718,4.919503,5.4363527,3.7499893,1.5731846,1.8146327,3.240685,2.9652832,2.5767028,2.8106055,3.5651307,3.1840954,3.6292653,4.3083377,4.9044123,5.406172,4.38379,3.1237335,2.444661,2.5389767,2.9954643,3.9763467,3.187868,2.8143783,3.2331395,2.9841464,2.9841464,3.1652324,3.2859564,3.308592,3.4029078,2.8785129,2.4899325,2.584248,2.9200118,2.6823363,2.2598023,3.127506,4.1612053,4.538468,3.7575345,3.2670932,3.0709167,3.138824,3.4557245,3.983892,4.6742826,4.055572,3.983892,5.458988,8.627994,9.031664,6.379509,5.2628117,6.175787,5.515578,4.4403796,4.949684,5.938112,6.40969,5.4665337,5.198677,4.82896,5.119452,5.987156,6.515323,9.0807085,8.307321,6.4210076,6.692637,13.411682,12.51757,8.975075,7.5263867,8.76758,9.178797,8.469543,6.304056,5.2967653,7.1038527,12.419481,10.710483,10.33322,12.989148,15.30554,8.865668,3.62172,4.2592936,5.6551647,5.3269467,3.4557245,3.0633714,2.8294687,3.7914882,6.145606,9.246704,8.341274,7.798016,7.466025,7.232122,7.0246277,7.6697464,6.907676,6.7944975,7.779153,8.699674,8.98262,9.590013,9.073163,9.869187,18.28214,30.414904,22.439573,13.539951,10.963248,10.020092,11.170743,12.996693,13.9888935,14.022847,14.320885,16.984358,21.296469,22.541435,20.915434,21.511507,22.26226,24.929506,33.798946,48.878128,65.919075,74.96206,68.14115,55.60472,43.31728,33.04065,27.362848,24.012758,21.96045,20.175999,17.63325,18.651857,19.512016,19.74592,19.855326,21.307787,20.730574,20.300495,21.669958,24.21648,25.05023,27.098766,25.71044,21.115381,15.196134,11.506506,9.895596,10.201178,10.227587,9.235386,7.9489207,8.971302,8.560086,6.8699503,4.870459,4.3196554,3.9574835,3.7386713,4.0970707,4.4215164,3.0633714,2.2748928,1.6712729,1.4600059,1.6260014,1.9089483,2.2484846,2.161714,1.8485862,1.5920477,1.7391801,2.444661,2.0787163,1.569412,1.3732355,1.4449154,0.98842776,0.56589377,0.41498876,0.44516975,0.20372175,0.23767537,0.32067314,0.76207024,1.5920477,2.5729303,2.7011995,1.5430037,0.59607476,0.30935526,0.09808825,0.25276586,0.18863125,0.150905,0.1961765,0.19240387,0.1056335,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.06413463,0.10940613,0.23013012,0.41498876,0.5696664,0.33953625,0.1659955,0.071679875,0.0452715,0.05281675,0.06413463,0.05281675,0.041498873,0.030181,0.02263575,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.05281675,0.08299775,0.15845025,0.03772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.0150905,0.00754525,0.0150905,0.056589376,0.12826926,0.090543,0.05281675,0.03772625,0.03772625,0.041498873,0.05281675,0.09808825,0.1659955,0.27917424,0.47157812,0.55080324,0.663982,0.7997965,0.9016574,0.8639311,1.0223814,1.3128735,1.2298758,0.83752275,0.7997965,0.9922004,1.3355093,2.305074,3.591539,4.1008434,3.0143273,2.5540671,2.252257,1.8485862,1.2525115,1.2449663,1.4147344,1.1619685,0.5281675,0.17354076,0.10940613,0.06790725,0.06413463,0.10940613,0.22258487,0.26031113,0.35462674,0.41121614,0.41876137,0.452715,0.51684964,0.45648763,0.3961256,0.38103512,0.38480774,0.33953625,0.30181,0.28294688,0.271629,0.241448,0.211267,0.19994913,0.241448,0.33576363,0.43007925,0.46026024,0.33576363,0.24522063,0.25276586,0.28294688,0.33953625,0.41121614,0.41121614,0.331991,0.2565385,0.181086,0.10940613,0.071679875,0.06790725,0.06790725,0.09808825,0.12826926,0.13958712,0.18863125,0.422534,0.2678564,0.21881226,0.22258487,0.21881226,0.1659955,0.21503963,0.20749438,0.1659955,0.116951376,0.08299775,0.056589376,0.056589376,0.056589376,0.049044125,0.03772625,0.030181,0.026408374,0.030181,0.03772625,0.0452715,0.03772625,0.026408374,0.02263575,0.02263575,0.033953626,0.06413463,0.09808825,0.124496624,0.12826926,0.11317875,0.10186087,0.10186087,0.094315626,0.07922512,0.05281675,0.03772625,0.026408374,0.02263575,0.0150905,0.0150905,0.06790725,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.08677038,0.116951376,0.06413463,0.03772625,0.0452715,0.018863125,0.1056335,0.5093044,1.5015048,1.2600567,0.58098423,0.120724,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.08677038,0.26408374,0.84129536,1.6637276,2.161714,1.1996948,0.5772116,0.48666862,0.6073926,0.10940613,0.03772625,0.02263575,0.030181,0.03772625,0.018863125,0.011317875,0.00754525,0.026408374,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10940613,0.5394854,0.10940613,0.10940613,0.1659955,0.10940613,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.21881226,0.22258487,0.071679875,0.0,0.14713238,0.2678564,0.38103512,0.4376245,0.32821837,0.4979865,1.0412445,0.8941121,0.14713238,0.041498873,0.0754525,0.09808825,0.845068,1.9202662,1.7693611,0.77338815,0.20749438,0.030181,0.094315626,0.16976812,0.5357128,0.8903395,2.0485353,3.8669407,5.2326307,5.243949,5.2854476,4.9232755,4.5988297,5.613666,6.330465,5.704209,4.6818275,3.7386713,2.867195,2.0183544,1.539231,1.6675003,2.033445,1.6561824,3.4557245,4.6290107,4.055572,2.4861598,2.5616124,2.7087448,2.3013012,2.2598023,2.8256962,3.5387223,3.350091,3.6443558,4.7308717,6.0626082,6.273875,4.402653,3.1124156,2.7011995,3.169005,4.221567,5.194905,4.327201,3.5047686,3.4972234,3.953711,4.0103,3.7160356,3.6481283,3.8480775,3.8292143,3.2255943,2.8445592,2.6483827,2.5578396,2.4333432,2.04099,2.1013522,2.8634224,3.731126,3.2821836,3.0709167,3.2520027,3.2784111,3.2520027,3.9197574,5.617439,4.8553686,4.7120085,6.7944975,11.234878,9.64283,6.7114997,5.96452,7.6848373,8.903395,8.296002,7.8961043,7.375482,6.8397694,6.8397694,5.6363015,7.537705,11.400873,13.604086,8.054554,4.9760923,4.032936,4.447925,6.579458,11.925267,10.744436,7.8998766,7.183078,8.718536,8.941121,7.1378064,7.964011,8.677037,8.929804,10.774617,9.193887,7.118943,6.7152724,7.122716,4.4516973,5.9494295,8.967529,9.491924,7.2057137,5.5004873,5.093044,5.0251365,6.4247804,8.733627,9.710737,7.062354,6.3719635,6.541732,6.4247804,4.8327327,5.3458095,4.504514,4.2404304,5.0741806,6.1003346,7.2358947,7.677292,8.288457,10.585986,16.716501,21.262514,14.649103,9.480607,9.937095,11.759273,12.925014,13.004238,12.7477,12.468526,12.0233555,15.199906,18.92726,18.776354,16.048746,17.765291,20.677757,24.329659,32.674706,45.395996,57.924885,62.429398,58.74732,50.621082,40.55949,29.83769,24.646559,22.04722,20.677757,19.606333,18.334957,17.984104,17.437073,17.60684,18.704676,20.22127,18.41041,17.40689,18.904623,21.911406,22.7527,26.1707,26.502691,22.322622,15.62244,11.796998,10.61994,9.0807085,7.9413757,7.7602897,8.914713,10.970794,10.114408,8.009283,5.8928404,4.5761943,4.0216184,3.6028569,3.7688525,4.1989317,3.8141239,2.9766011,2.1202152,1.6788181,1.5958204,1.3430545,1.2261031,1.2261031,1.2034674,1.1544232,1.237421,2.191895,1.841041,1.4147344,1.3204187,1.1242423,0.67152727,0.33953625,0.2867195,0.38103512,0.20372175,0.44894236,0.8337501,1.2185578,1.7995421,3.108643,3.108643,2.161714,1.2336484,0.694163,0.32821837,0.845068,1.2525115,1.0035182,0.35085413,0.362172,0.18863125,0.06790725,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.1056335,0.22258487,0.30181,0.33953625,0.38858038,0.25276586,0.13204187,0.05281675,0.02263575,0.0150905,0.018863125,0.011317875,0.00754525,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.0452715,0.120724,0.041498873,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.02263575,0.0150905,0.011317875,0.033953626,0.10186087,0.18863125,0.09808825,0.0452715,0.026408374,0.030181,0.030181,0.049044125,0.13204187,0.2867195,0.45648763,0.51684964,0.5357128,0.65643674,0.80356914,0.90920264,0.91297525,0.94315624,1.0148361,0.9695646,0.80734175,0.69039035,0.9318384,1.8976303,3.2482302,4.247976,3.772625,4.217795,4.678055,4.187614,2.776652,1.4524606,1.0827434,1.1883769,1.0638802,0.59230214,0.22258487,0.13204187,0.090543,0.0754525,0.07922512,0.10186087,0.13958712,0.19994913,0.24522063,0.24522063,0.1961765,0.271629,0.30935526,0.33953625,0.3734899,0.392353,0.40367088,0.3961256,0.35839936,0.30181,0.24899325,0.16976812,0.14335975,0.1659955,0.21881226,0.28294688,0.331991,0.29426476,0.26408374,0.2565385,0.23013012,0.26031113,0.33576363,0.3734899,0.35085413,0.32444575,0.30181,0.21881226,0.15845025,0.13204187,0.1056335,0.11317875,0.12826926,0.120724,0.15845025,0.38103512,0.23013012,0.19240387,0.20749438,0.241448,0.3055826,0.3734899,0.2565385,0.1358145,0.08299775,0.06413463,0.049044125,0.049044125,0.0452715,0.03772625,0.030181,0.026408374,0.026408374,0.030181,0.033953626,0.0452715,0.049044125,0.041498873,0.030181,0.026408374,0.0150905,0.02263575,0.03772625,0.06413463,0.090543,0.08677038,0.08299775,0.0754525,0.0754525,0.07922512,0.071679875,0.120724,0.10940613,0.06790725,0.018863125,0.0150905,0.071679875,0.02263575,0.003772625,0.011317875,0.0754525,0.26031113,0.3470815,0.14713238,0.0,0.0150905,0.071679875,0.094315626,0.03772625,0.11317875,0.62625575,2.0145817,1.6033657,0.80734175,0.23767537,0.071679875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.2263575,0.62248313,0.392353,0.48666862,1.6373192,3.1124156,2.7200627,0.7167987,0.18863125,0.16222288,0.13958712,0.07922512,0.0452715,0.030181,0.056589376,0.19994913,0.59230214,0.116951376,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0754525,0.08299775,0.018863125,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.018863125,0.14335975,0.17731337,0.090543,0.018863125,0.03772625,0.08299775,0.14713238,0.20749438,0.2565385,0.05281675,0.0,0.0,0.030181,0.150905,0.24522063,0.20749438,0.44894236,0.77338815,0.4074435,0.14713238,0.071679875,0.05281675,0.06413463,0.18485862,0.47535074,1.0148361,1.9466745,2.9200118,3.0633714,4.587512,5.0138187,4.8440504,4.7535076,5.572167,7.624475,6.8435416,5.1269975,3.6783094,3.0181,2.5578396,2.505023,3.2972744,3.9084394,1.8599042,2.1881225,3.9763467,4.395108,3.097325,2.2371666,2.5238862,2.5012503,2.5427492,2.6672459,2.516341,2.886058,3.572676,4.9157305,6.1720147,5.5382137,3.2784111,2.6823363,2.9916916,3.7273536,4.689373,5.1798143,5.13077,4.6026025,4.006528,4.1197066,3.7688525,3.6745367,3.7914882,4.032936,4.255521,3.308592,3.270866,3.006782,2.3126192,1.901403,1.7391801,1.5731846,2.022127,2.746471,2.4220252,3.169005,3.3878171,3.0407357,2.757789,3.8103511,6.802043,6.470052,5.907931,6.8435416,9.654147,6.9491754,7.1793056,9.454198,12.668475,15.513034,13.675766,10.3634,7.462252,6.4549613,8.394091,5.4967146,10.050273,16.991903,19.48938,8.956212,4.025391,3.712263,4.0291634,3.9612563,5.455216,6.802043,5.2288585,4.1536603,4.7421894,5.926794,7.0585814,12.457208,14.237886,10.574668,5.696664,6.126743,5.772116,4.7535076,3.8707132,4.606375,10.702937,13.830443,12.551523,8.941121,8.59404,8.416726,8.590267,8.492179,7.5263867,5.13077,4.508287,5.587258,6.485142,6.006019,3.6556737,4.2064767,4.5007415,4.353609,4.1612053,4.908185,5.515578,7.039718,8.311093,8.83926,8.801534,7.7678347,6.432326,6.7643166,9.491924,14.0907545,13.992666,12.985375,12.276122,11.691365,9.669238,10.638803,11.18206,10.993429,10.770844,12.200669,15.32063,20.243906,27.743885,36.986816,45.554447,53.46187,57.981472,55.60472,46.173157,32.8822,24.903097,22.56407,21.522825,20.040184,19.006485,18.806536,17.840744,17.369165,17.625704,17.818108,17.123945,16.31283,15.147089,14.483108,16.286423,22.930016,24.846508,21.122927,14.724555,12.498707,11.812089,9.0543,7.1679873,7.696155,10.816116,13.336229,11.732863,9.35611,7.4735703,5.2779026,4.1989317,3.429316,3.3236825,3.783943,4.2894745,3.2746384,2.3465726,1.7580433,1.4147344,0.87902164,0.7997965,0.97333723,1.1242423,1.0487897,0.6375736,1.3770081,1.5241405,1.5430037,1.5241405,1.1883769,0.68661773,0.38480774,0.3055826,0.3734899,0.44139713,0.9507015,1.5165952,1.750498,2.071171,3.6896272,2.8558772,2.7879698,2.354118,1.4826416,1.1242423,1.9655377,2.7841973,2.2447119,0.8337501,0.875249,0.41121614,0.12826926,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.033953626,0.16222288,0.35462674,0.3961256,0.2678564,0.14713238,0.094315626,0.056589376,0.030181,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.02263575,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.03772625,0.02263575,0.02263575,0.05281675,0.10940613,0.1358145,0.060362,0.026408374,0.02263575,0.030181,0.030181,0.041498873,0.12826926,0.331991,0.5696664,0.6111652,0.5583485,0.62625575,0.7922512,0.965792,0.98842776,0.8337501,0.7696155,0.7205714,0.663982,0.6451189,0.8337501,2.214531,3.821669,4.4177437,2.4861598,4.9685473,6.277648,5.4363527,3.078462,1.4600059,0.94315624,1.1016065,1.1506506,0.8111144,0.29426476,0.16976812,0.120724,0.1056335,0.10186087,0.12826926,0.17354076,0.23390275,0.29426476,0.29803738,0.1659955,0.18863125,0.23013012,0.29049212,0.33953625,0.33953625,0.41876137,0.47535074,0.4640329,0.392353,0.3169005,0.23767537,0.18863125,0.14335975,0.10940613,0.10186087,0.15467763,0.20749438,0.241448,0.25276586,0.24899325,0.23390275,0.241448,0.271629,0.32067314,0.3772625,0.41876137,0.33576363,0.2565385,0.211267,0.150905,0.15845025,0.12826926,0.09808825,0.08677038,0.0754525,0.06413463,0.120724,0.17354076,0.241448,0.422534,0.4640329,0.241448,0.0754525,0.056589376,0.0452715,0.049044125,0.041498873,0.033953626,0.030181,0.030181,0.041498873,0.041498873,0.03772625,0.033953626,0.041498873,0.049044125,0.05281675,0.049044125,0.03772625,0.018863125,0.0150905,0.02263575,0.033953626,0.0452715,0.056589376,0.08299775,0.0754525,0.06790725,0.0754525,0.10186087,0.19240387,0.18485862,0.11317875,0.03772625,0.02263575,0.0452715,0.00754525,0.0,0.060362,0.38103512,1.297783,1.7354075,0.7394345,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24899325,1.0751982,2.867195,1.086516,0.66020936,1.20724,1.7316349,0.59607476,0.20372175,0.1056335,0.08299775,0.041498873,0.030181,0.056589376,0.02263575,0.030181,0.6149379,2.776652,0.55457586,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3734899,0.4074435,0.08677038,0.1358145,0.0754525,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.090543,0.18863125,0.241448,0.15467763,0.0,0.0,0.0,0.0,0.0,0.06413463,0.32067314,0.45648763,0.62625575,0.47912338,0.29426476,0.9922004,0.5281675,0.35839936,0.26031113,0.23013012,0.48666862,0.73188925,0.8111144,0.9393836,1.2562841,1.8297231,3.5387223,3.8593953,3.429316,3.5462675,6.1342883,9.454198,9.250477,6.700182,3.8858037,3.7990334,3.1161883,2.9615107,3.1765501,3.3274553,2.71629,2.837014,3.6745367,3.3463185,2.0296721,1.9693103,3.4557245,3.8556228,4.0291634,4.0782075,3.3576362,2.7238352,3.3048196,3.561358,3.2067313,3.218049,2.2183034,2.546522,2.8256962,2.7615614,3.127506,4.5422406,4.496969,3.7009451,2.9351022,3.0218725,3.5085413,3.3010468,3.218049,3.410453,3.3878171,2.71629,2.9426475,2.9426475,2.3880715,1.7542707,1.8749946,2.3013012,2.9916916,3.361409,2.2899833,3.2784111,3.2142766,2.9086938,2.916239,3.5387223,7.273621,7.2472124,5.5570765,4.1612053,4.8666863,5.1232247,9.205205,13.687083,15.999702,14.449154,11.910177,7.8432875,5.481624,5.9192486,8.103599,4.9760923,5.9192486,10.374719,13.59654,6.6360474,4.7836885,6.349328,6.7152724,5.2628117,5.372218,10.0465,7.24344,3.519859,2.4220252,4.485651,8.771353,14.079436,14.618922,9.322156,1.8787673,2.7426984,5.20245,6.417235,5.8626595,5.3269467,6.1795597,6.934085,6.590776,6.688864,11.291467,12.012038,9.371201,5.753253,2.837014,1.6033657,2.505023,3.2972744,4.5761943,6.2323766,7.4773426,9.491924,11.378237,12.102581,11.695138,11.246195,10.612394,11.570641,11.506506,9.156161,4.5761943,7.911195,8.805306,8.130007,7.2924843,8.254503,8.986393,10.076681,11.02361,10.450171,6.1041074,5.1534057,5.3458095,7.213259,10.137043,12.359119,14.128481,20.330677,29.407612,39.36357,47.776524,61.935184,68.29583,64.55716,51.9,34.95714,24.265524,21.553007,20.949387,19.825144,18.79899,20.922977,22.443346,20.866388,16.618414,13.030646,12.785426,13.905896,14.053028,14.418973,19.73083,28.336185,29.743376,24.582424,16.663685,13.000465,10.729345,8.963757,8.873214,10.582213,13.181552,12.902377,11.917723,11.080199,9.955957,6.8058157,5.1081343,4.353609,4.036709,3.8405323,3.6330378,2.7540162,2.1579416,1.7052265,1.2940104,0.8526133,0.5998474,0.9280658,1.1581959,1.0299267,0.68661773,0.91674787,1.1506506,1.0638802,0.7394345,0.6413463,0.60362,0.392353,0.59607476,1.0789708,0.9922004,1.9693103,1.5543215,0.97333723,1.4298248,4.104616,3.3123648,3.5047686,3.500996,3.1237335,3.2331395,3.5387223,3.0407357,2.2899833,1.7429527,1.7542707,0.7432071,0.21503963,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.071679875,0.1056335,0.30181,0.35839936,0.27540162,0.120724,0.060362,0.03772625,0.02263575,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.060362,0.049044125,0.0452715,0.056589376,0.0754525,0.0754525,0.041498873,0.030181,0.030181,0.030181,0.030181,0.041498873,0.056589376,0.12826926,0.32821837,0.73188925,0.56212115,0.5357128,0.633801,0.7809334,0.8563859,0.7092535,0.7092535,0.77338815,0.8903395,1.0978339,1.146878,2.2409391,3.3689542,3.8782585,3.4632697,4.146115,4.1800685,3.361409,2.1315331,1.5731846,1.2298758,1.1431054,1.0035182,0.68661773,0.26031113,0.17354076,0.1358145,0.116951376,0.1056335,0.090543,0.07922512,0.13958712,0.18485862,0.181086,0.1659955,0.23013012,0.271629,0.29426476,0.31312788,0.35085413,0.41121614,0.42630664,0.44516975,0.47535074,0.48666862,0.4376245,0.3734899,0.27917424,0.18485862,0.1358145,0.16222288,0.21503963,0.26408374,0.29803738,0.33576363,0.29803738,0.27917424,0.26408374,0.2565385,0.3055826,0.35462674,0.3470815,0.31312788,0.27540162,0.27540162,0.35839936,0.20749438,0.08677038,0.08677038,0.1358145,0.124496624,0.120724,0.150905,0.18863125,0.150905,0.12826926,0.08677038,0.056589376,0.0452715,0.0452715,0.056589376,0.05281675,0.041498873,0.030181,0.030181,0.030181,0.030181,0.030181,0.026408374,0.0150905,0.0150905,0.02263575,0.030181,0.030181,0.030181,0.00754525,0.00754525,0.02263575,0.033953626,0.0452715,0.08299775,0.090543,0.090543,0.08677038,0.0754525,0.05281675,0.03772625,0.049044125,0.071679875,0.060362,0.00754525,0.0,0.0,0.011317875,0.0754525,0.26031113,0.3470815,0.14713238,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1657411,2.1390784,2.3201644,1.8674494,0.633801,1.0374719,1.5618668,1.358145,0.241448,0.13204187,0.09808825,0.0754525,0.041498873,0.018863125,0.0150905,0.003772625,0.00754525,0.20749438,0.9695646,0.271629,0.03772625,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0754525,0.08299775,0.018863125,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.07922512,0.211267,0.27540162,0.12826926,0.09808825,0.060362,0.02263575,0.120724,0.26031113,0.15467763,0.03772625,0.094315626,0.4678055,0.5017591,0.422534,0.392353,0.7696155,2.0900342,0.97333723,0.754525,0.91297525,0.935611,0.35462674,0.422534,0.59607476,0.8224323,1.3128735,2.5502944,3.5575855,3.5387223,3.169005,3.7160356,7.0246277,7.77538,7.3415284,5.9532022,4.4403796,4.2404304,3.3878171,3.4972234,3.7198083,3.4179983,2.1541688,2.7728794,2.7087448,2.0975795,1.4864142,1.8448136,4.146115,6.1418333,7.066127,6.617184,4.919503,3.591539,3.2029586,2.7691069,2.3956168,3.2670932,3.99521,4.1310244,3.500996,2.7087448,3.1652324,3.7990334,3.2482302,2.7502437,2.886058,3.5462675,3.0369632,2.4069347,2.2409391,2.6483827,3.229367,3.4255435,3.904667,3.8556228,3.078462,1.9730829,1.6863633,1.8825399,2.6182017,3.4896781,3.6556737,4.557331,4.7912335,4.647874,4.689373,5.7607985,6.9869013,5.783434,5.379763,6.8246784,8.967529,8.296002,8.956212,8.616675,6.6624556,4.183841,6.4210076,6.651138,5.221313,3.8895764,5.8211603,5.040227,4.564876,4.949684,5.3571277,3.572676,4.0895257,5.587258,5.704209,5.3194013,8.544995,10.38981,6.6134114,4.044254,5.8513412,11.529142,8.254503,6.9755836,6.8699503,6.63982,4.478106,7.394345,7.5188417,6.5756855,5.6891184,5.3873086,5.119452,4.515832,4.112161,4.90064,8.299775,8.239413,7.17176,5.485397,4.402653,5.9720654,8.213005,7.877241,7.564113,8.812852,12.079946,11.7894535,8.688355,6.039973,5.2590394,5.9003854,6.398372,9.031664,10.076681,8.9788475,8.326183,14.109617,13.845533,10.121953,6.1418333,5.7419353,6.881268,6.802043,6.5756855,6.017337,3.663219,5.4740787,8.627994,10.925522,12.15917,14.117163,16.463736,20.749437,25.887753,31.705141,38.974987,45.626125,42.072315,34.485565,26.061293,17.025856,13.023102,13.015556,14.811326,17.28994,20.43631,23.507227,24.00144,22.013268,18.599041,15.788436,14.452927,12.494934,12.7477,16.780636,24.891779,43.988808,48.27451,38.90708,22.813063,12.706201,12.283667,11.336739,11.465008,12.494934,12.487389,11.895086,12.00072,12.668475,12.370438,8.197914,5.9418845,5.643847,5.3344917,4.323428,3.180323,2.897376,2.4069347,1.8485862,1.3166461,0.87902164,0.90543,1.2336484,1.6561824,2.0787163,2.516341,2.0070364,2.9124665,3.8707132,4.0782075,3.2784111,2.9200118,1.5505489,0.7696155,0.8978847,0.965792,1.991946,1.5958204,1.1280149,1.2261031,1.81086,1.2600567,0.97333723,1.0186088,1.4562333,2.3692086,3.7575345,6.2097406,5.8588867,2.7917426,1.0450171,0.6111652,0.21881226,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.150905,0.21503963,0.21503963,0.18863125,0.150905,0.120724,0.09808825,0.033953626,0.02263575,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.03772625,0.05281675,0.06413463,0.14713238,0.24899325,0.19994913,0.06413463,0.02263575,0.018863125,0.018863125,0.018863125,0.02263575,0.03772625,0.071679875,0.15845025,0.36594462,0.35085413,0.513077,0.6488915,0.6752999,0.62248313,0.573439,0.58475685,0.7432071,1.0902886,1.599593,1.2487389,1.3543724,2.3163917,3.712263,4.293247,3.9122121,3.3727267,2.6710186,2.3465726,3.4745877,2.0900342,1.2826926,1.0035182,0.8903395,0.26031113,0.1358145,0.08677038,0.0754525,0.07922512,0.06790725,0.06413463,0.1056335,0.1358145,0.124496624,0.094315626,0.1659955,0.15845025,0.17731337,0.2565385,0.35085413,0.34330887,0.39989826,0.48666862,0.56589377,0.5998474,0.6451189,0.6187105,0.5281675,0.39989826,0.271629,0.2263575,0.2263575,0.27917424,0.3734899,0.47157812,0.482896,0.42630664,0.34330887,0.2867195,0.3055826,0.29426476,0.3169005,0.3470815,0.362172,0.3734899,0.45648763,0.38480774,0.26408374,0.1659955,0.1358145,0.1056335,0.090543,0.10186087,0.124496624,0.12826926,0.06413463,0.049044125,0.049044125,0.0452715,0.0452715,0.03772625,0.026408374,0.018863125,0.02263575,0.030181,0.030181,0.030181,0.030181,0.026408374,0.0150905,0.026408374,0.03772625,0.041498873,0.049044125,0.06790725,0.041498873,0.02263575,0.0150905,0.02263575,0.033953626,0.07922512,0.11317875,0.150905,0.19994913,0.24899325,0.19240387,0.1358145,0.08677038,0.060362,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.094315626,0.1961765,0.03772625,0.00754525,0.0,0.0,0.00754525,0.0452715,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.573439,1.6750455,2.625747,2.2258487,1.7655885,1.8372684,2.1164427,1.3958713,1.0450171,1.3204187,1.3996439,0.9620194,0.18863125,0.124496624,0.08677038,0.06413463,0.060362,0.124496624,0.033953626,0.003772625,0.003772625,0.05281675,0.23390275,0.1358145,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.1056335,0.12826926,0.10940613,0.056589376,0.090543,0.23390275,0.39989826,0.66020936,0.4979865,0.28294688,0.29426476,0.73188925,0.7884786,0.5885295,0.5093044,0.9242931,2.2107582,1.4826416,1.3468271,1.3656902,1.1883769,0.513077,0.56589377,0.83752275,1.1506506,1.720317,3.1614597,4.093298,3.4896781,2.9841464,3.893349,7.194396,6.488915,5.451443,4.561104,4.1083884,4.183841,4.1197066,4.466788,4.881777,4.6252384,2.5540671,3.3727267,2.7992878,1.931584,1.5543215,2.1353056,4.112161,6.7341356,8.401636,8.262049,6.2361493,3.8178966,3.0671442,2.9954643,3.2067313,3.904667,3.832987,3.7348988,3.410453,3.1237335,3.5839937,3.7386713,2.9954643,2.3428001,2.3918443,3.3651814,2.9766011,2.625747,2.7200627,3.180323,3.4444065,3.5236318,3.640583,3.2972744,2.4899325,1.7089992,1.961765,2.1805773,2.8898308,4.164978,5.643847,6.0701537,6.092789,6.5228686,7.0585814,6.270103,6.6058664,7.001992,7.4094353,7.8244243,8.29223,6.647365,5.802297,4.406426,2.6898816,2.4672968,9.348565,9.039209,5.621211,3.2218218,6.0286546,7.194396,5.541986,4.1197066,4.036709,4.45547,5.4212623,8.130007,8.141325,6.096562,7.7376537,6.8661776,5.100589,6.40969,11.465008,17.64834,7.798016,3.7763977,4.074435,6.273875,7.0585814,8.922258,8.084735,6.571913,5.7079816,6.1078796,5.6589375,4.9232755,5.0779533,6.119198,6.8850408,5.4288073,4.564876,4.6516466,5.7872066,7.8244243,8.805306,7.5829763,6.058836,5.6815734,7.462252,6.6322746,4.98741,3.9084394,3.731126,3.731126,4.538468,6.3417826,7.250985,7.454707,9.190115,12.434572,10.223814,6.643593,4.2894745,4.2328854,4.8855495,5.3156285,6.0362,6.903904,7.1340337,9.514561,11.740409,12.679792,12.96274,14.977322,16.874952,18.765038,21.171972,24.974777,31.437284,34.62138,29.056757,20.75321,13.543724,9.073163,8.156415,9.042982,11.793225,15.671484,19.130981,20.711712,20.447628,19.225298,18.8254,21.926497,21.669958,17.154125,14.362384,16.399601,23.48459,42.653297,51.74155,46.705097,31.105293,16.120426,13.030646,12.525115,13.004238,13.102326,11.68382,10.899114,11.589504,12.419481,12.049765,9.110889,7.4018903,6.8397694,5.828706,4.402653,4.247976,3.712263,2.6182017,1.7655885,1.4411428,1.4260522,1.4071891,3.1312788,4.315883,4.221567,3.663219,2.584248,3.3312278,3.9574835,3.7462165,3.187868,4.425289,2.7502437,1.3166461,1.2336484,1.5845025,1.4864142,1.2826926,1.5128226,1.7995421,0.8865669,0.6488915,0.7130261,0.9016574,1.1959221,1.7127718,4.134797,4.9685473,3.7009451,1.3958713,0.7054809,0.784706,0.43385187,0.11317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.090543,0.1358145,0.120724,0.09808825,0.07922512,0.06790725,0.071679875,0.018863125,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.00754525,0.0,0.0,0.011317875,0.026408374,0.041498873,0.06413463,0.06790725,0.09808825,0.1358145,0.10940613,0.03772625,0.018863125,0.0150905,0.0150905,0.0150905,0.0150905,0.026408374,0.049044125,0.08299775,0.14713238,0.19994913,0.36971724,0.52062225,0.5583485,0.4376245,0.49421388,0.55080324,0.80356914,1.4335974,2.6219745,2.6823363,1.8146327,1.5165952,2.0975795,2.6785638,6.507778,4.3611546,2.282438,2.463524,3.2369123,2.3013012,1.4109617,0.8978847,0.7167987,0.44139713,0.17731337,0.0754525,0.056589376,0.06413463,0.060362,0.05281675,0.071679875,0.08299775,0.071679875,0.056589376,0.10186087,0.094315626,0.1056335,0.1659955,0.241448,0.23013012,0.30181,0.40367088,0.49044126,0.5357128,0.5772116,0.6073926,0.60362,0.5583485,0.47912338,0.34330887,0.28294688,0.29049212,0.3470815,0.41121614,0.5017591,0.5394854,0.5357128,0.4979865,0.422534,0.36971724,0.3734899,0.39989826,0.43007925,0.44139713,0.49044126,0.4640329,0.36594462,0.23767537,0.14713238,0.116951376,0.1056335,0.10940613,0.10940613,0.0754525,0.033953626,0.026408374,0.030181,0.03772625,0.03772625,0.03772625,0.030181,0.02263575,0.018863125,0.030181,0.02263575,0.02263575,0.02263575,0.018863125,0.0150905,0.018863125,0.026408374,0.026408374,0.030181,0.049044125,0.03772625,0.030181,0.02263575,0.026408374,0.030181,0.056589376,0.090543,0.1358145,0.19240387,0.25276586,0.24522063,0.21503963,0.18863125,0.16976812,0.13204187,0.00754525,0.0,0.018863125,0.018863125,0.0,0.0,0.018863125,0.17731337,0.6828451,1.086516,0.3055826,0.14335975,0.06790725,0.026408374,0.00754525,0.0452715,0.041498873,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38480774,1.6373192,2.4031622,2.6521554,3.6707642,3.0256453,1.7052265,1.0638802,1.3920987,1.8976303,1.1996948,1.0035182,0.8299775,0.5017591,0.18485862,0.10186087,0.060362,0.060362,0.09808825,0.1659955,0.06413463,0.041498873,0.030181,0.018863125,0.026408374,0.2678564,0.13204187,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.124496624,0.09808825,0.0,0.0,0.17731337,0.15467763,0.3055826,0.6187105,0.7167987,1.1921495,1.1091517,0.8526133,0.6828451,0.73188925,0.633801,0.67152727,0.83752275,1.3656902,2.7389257,2.3880715,2.0975795,1.7240896,1.2336484,0.7394345,1.0902886,1.6033657,1.8184053,2.1164427,3.7160356,4.98741,4.304565,3.5123138,4.146115,7.435844,6.934085,5.2552667,4.006528,3.8065786,4.2894745,5.138315,6.0701537,6.2851934,5.3194013,3.0407357,3.2067313,2.463524,1.8221779,1.7731338,2.3088465,3.1048703,5.794752,7.960239,8.228095,6.247467,3.663219,3.1199608,3.4594972,3.9650288,4.353609,3.5462675,3.5123138,3.6481283,3.663219,3.5990841,3.2784111,2.8634224,2.6219745,2.7653341,3.4217708,3.078462,2.8709676,3.138824,3.712263,3.874486,3.2482302,2.938875,2.6672459,2.3993895,2.3314822,3.2633207,3.0935526,3.029418,3.7160356,5.2175403,5.59103,5.560849,6.1795597,6.990674,6.0512905,6.6850915,8.631766,9.767326,9.163706,7.1000805,5.2326307,4.0517993,2.8709676,2.3126192,4.2819295,11.117926,8.929804,4.727099,2.938875,5.409944,7.2660756,5.349582,4.2592936,5.13077,5.6098933,6.3455553,10.808571,11.057564,6.7944975,5.3571277,4.2027044,3.8480775,5.975838,10.03141,13.223051,5.0515447,2.5238862,3.4632697,5.5495315,6.277648,6.8171334,6.1305156,5.168496,5.010046,6.8737226,6.349328,5.7004366,6.017337,6.820906,6.0626082,4.055572,3.259548,4.5007415,6.9189944,7.9300575,6.749226,5.945657,5.3684454,5.247721,6.217286,7.960239,10.355856,11.185833,10.223814,9.235386,9.993684,9.322156,7.888559,6.9454026,8.329956,8.695901,6.0701537,4.357382,4.5837393,4.8968673,4.353609,4.666737,6.3531003,8.669493,9.601331,9.831461,10.929295,11.544232,11.891314,13.7700815,15.437581,16.135517,17.274849,20.398582,27.19308,30.131956,25.020048,17.45971,11.246195,8.3525915,7.284939,8.024373,10.133271,12.691111,14.27184,14.86037,15.667711,16.569368,18.568861,23.763765,25.676485,22.771564,18.821627,16.863634,19.191343,31.803228,41.525284,42.532574,33.80649,19.1423,12.849561,11.725319,12.694883,13.460726,12.487389,10.748209,11.083972,11.706455,11.246195,8.763808,8.028146,7.745199,6.85486,5.6061206,5.5193505,3.7499893,2.7653341,2.4672968,2.584248,2.6634734,3.651901,4.644101,4.6856003,4.006528,3.9989824,4.3309736,5.3948536,5.353355,3.9122121,2.293756,6.0286546,4.1989317,1.750498,0.9242931,1.2600567,0.724344,0.6790725,1.1581959,1.539231,0.55080324,0.80734175,1.146878,1.4826416,1.6410918,1.358145,3.6971724,3.361409,1.8825399,0.663982,0.965792,0.69039035,0.35462674,0.1056335,0.0,0.00754525,0.0,0.0,0.003772625,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.041498873,0.049044125,0.0452715,0.033953626,0.018863125,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0150905,0.011317875,0.0150905,0.02263575,0.033953626,0.041498873,0.05281675,0.05281675,0.0452715,0.033953626,0.02263575,0.018863125,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.03772625,0.05281675,0.060362,0.10940613,0.23013012,0.35462674,0.44139713,0.4678055,0.52439487,0.62248313,0.91297525,1.6486372,3.2067313,3.7160356,2.7087448,1.5807298,1.2713746,2.2598023,5.745708,4.191386,3.4670424,4.557331,3.5500402,2.6408374,1.5128226,0.8337501,0.66020936,0.43007925,0.16976812,0.0754525,0.060362,0.06413463,0.060362,0.049044125,0.05281675,0.05281675,0.0452715,0.05281675,0.071679875,0.08299775,0.090543,0.10186087,0.124496624,0.150905,0.24899325,0.35839936,0.43385187,0.44139713,0.47157812,0.51684964,0.5696664,0.60362,0.58475685,0.55457586,0.5017591,0.43385187,0.3734899,0.36971724,0.4640329,0.56589377,0.6375736,0.6526641,0.6073926,0.5583485,0.55080324,0.55457586,0.5470306,0.52062225,0.51684964,0.5319401,0.49044126,0.38103512,0.24899325,0.19994913,0.15467763,0.116951376,0.08299775,0.041498873,0.018863125,0.0150905,0.02263575,0.03772625,0.03772625,0.0452715,0.03772625,0.026408374,0.02263575,0.030181,0.02263575,0.018863125,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.018863125,0.030181,0.026408374,0.030181,0.03772625,0.03772625,0.03772625,0.0452715,0.06790725,0.10186087,0.13958712,0.19240387,0.22258487,0.21503963,0.21503963,0.21503963,0.19240387,0.041498873,0.026408374,0.0452715,0.041498873,0.011317875,0.0,0.094315626,0.45648763,1.2449663,1.780679,0.5583485,0.331991,0.16222288,0.05281675,0.00754525,0.041498873,0.056589376,0.033953626,0.011317875,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,1.0035182,3.7009451,3.9914372,2.071171,2.4522061,2.1202152,1.3468271,0.69039035,1.0336993,3.572676,1.4373702,0.52062225,0.21503963,0.1358145,0.150905,0.06790725,0.030181,0.05281675,0.11317875,0.11317875,0.116951376,0.11317875,0.071679875,0.011317875,0.0,0.4678055,0.23767537,0.018863125,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.06790725,0.10940613,0.24522063,0.21503963,0.030181,0.0,0.23013012,0.33576363,0.56589377,0.87147635,0.8865669,1.4977322,1.5467763,1.3619176,1.0487897,0.48666862,0.18485862,0.56212115,1.1846043,2.1315331,3.9989824,3.3727267,2.8106055,2.1390784,1.4335974,1.0072908,1.6675003,2.5540671,2.7653341,2.7238352,4.1762958,5.7607985,5.43258,4.3083377,4.274384,8.00551,8.601585,6.802043,4.919503,4.146115,4.5912848,6.217286,8.058327,7.9753294,5.836251,3.5387223,2.5993385,1.9089483,1.7165444,1.9089483,2.022127,1.6260014,3.731126,5.6891184,6.0701537,4.6554193,3.2746384,3.2331395,3.5953116,3.9122121,4.2102494,3.4972234,3.9725742,4.4894238,4.395108,3.5274043,2.584248,2.4823873,2.9011486,3.3953626,3.4255435,2.969056,2.6106565,2.848332,3.5990841,4.1989317,2.806833,2.2069857,2.282438,2.8181508,3.5236318,4.587512,4.08198,3.4632697,3.500996,4.304565,4.561104,4.0216184,4.0404816,4.817642,5.413717,6.9189944,9.242931,10.70671,10.091772,6.620957,5.4363527,4.515832,3.6141748,3.5538127,6.2135134,8.60913,5.481624,2.867195,2.8332415,3.4444065,4.5799665,3.8367596,4.8742313,7.284939,6.587003,5.934339,10.355856,10.797253,6.145606,3.2331395,4.617693,4.304565,3.8971217,3.7801702,3.138824,1.8636768,2.233394,3.2105038,3.92353,3.6594462,4.3649273,4.183841,3.8254418,4.4441524,7.643338,7.224577,6.3832817,6.039973,6.1342883,5.6023483,4.5912848,4.1762958,5.4740787,7.5263867,7.284939,5.617439,6.462507,7.911195,9.092027,10.137043,14.219024,18.621677,19.357338,16.927769,16.331694,18.048239,15.569623,11.204697,7.352846,6.507778,5.783434,4.5535583,5.093044,7.0812173,7.594294,5.572167,4.496969,5.726845,8.186596,8.360137,5.9796104,6.9454026,8.488406,9.635284,11.200924,12.826925,13.396591,14.403882,17.37671,23.861853,26.925224,22.258488,16.603323,13.268322,12.132762,9.544742,9.2844305,9.623966,9.5032425,8.533678,9.012801,11.857361,15.098045,17.852062,20.30804,22.982832,23.80149,21.817091,18.184053,16.161926,20.394812,25.74062,29.588697,28.819082,19.794964,12.936331,10.555805,11.2650585,13.132507,13.679539,11.106608,10.955703,11.917723,11.812089,7.5829763,7.0170827,7.647111,7.937603,7.254758,5.8890676,3.229367,2.806833,3.2746384,3.651901,3.3425457,5.5985756,4.606375,2.8521044,2.3805263,4.7535076,6.530414,7.488661,6.9793563,4.949684,1.9579924,6.587003,4.938366,1.9693103,0.392353,0.65643674,0.5998474,0.49044126,0.46026024,0.49044126,0.4074435,1.1581959,1.3392819,2.1202152,3.1425967,2.5087957,2.8294687,2.7728794,2.1579416,1.4373702,1.7240896,0.59230214,0.13204187,0.10186087,0.23390275,0.22258487,0.06413463,0.0150905,0.026408374,0.049044125,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.026408374,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.026408374,0.03772625,0.03772625,0.030181,0.030181,0.026408374,0.026408374,0.033953626,0.033953626,0.018863125,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.03772625,0.056589376,0.071679875,0.13958712,0.2263575,0.35085413,0.60362,0.56589377,0.69039035,1.0072908,1.6222287,2.7011995,3.3425457,2.9841464,2.0372176,1.4939595,2.9351022,1.901403,2.6446102,4.930821,6.749226,4.3196554,2.8521044,1.4411428,0.77716076,0.70170826,0.20372175,0.124496624,0.08299775,0.071679875,0.0754525,0.06413463,0.05281675,0.049044125,0.049044125,0.05281675,0.060362,0.06790725,0.090543,0.090543,0.06790725,0.06790725,0.120724,0.23767537,0.35462674,0.41876137,0.392353,0.43385187,0.45648763,0.513077,0.58475685,0.6111652,0.7809334,0.79602385,0.68661773,0.543258,0.51684964,0.5319401,0.6149379,0.68661773,0.7432071,0.83752275,0.8299775,0.8337501,0.8337501,0.8111144,0.72811663,0.66020936,0.694163,0.6828451,0.58475685,0.46026024,0.36594462,0.23767537,0.124496624,0.05281675,0.03772625,0.02263575,0.0150905,0.026408374,0.041498873,0.0452715,0.0452715,0.03772625,0.030181,0.030181,0.033953626,0.030181,0.02263575,0.0150905,0.018863125,0.018863125,0.0150905,0.0150905,0.0150905,0.018863125,0.026408374,0.018863125,0.033953626,0.041498873,0.041498873,0.041498873,0.0452715,0.0754525,0.10186087,0.116951376,0.150905,0.19240387,0.18863125,0.18485862,0.19994913,0.20372175,0.1358145,0.124496624,0.049044125,0.030181,0.060362,0.0,0.2678564,0.5017591,0.36594462,0.02263575,0.1056335,0.29049212,0.1358145,0.0,0.041498873,0.19994913,0.041498873,0.00754525,0.02263575,0.030181,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.1659955,1.1695137,2.1164427,1.6637276,0.59607476,1.8146327,2.6106565,1.5430037,0.72811663,1.8900851,6.3945994,3.572676,1.2223305,0.16976812,0.23390275,0.19994913,0.08677038,0.033953626,0.0150905,0.026408374,0.0754525,0.23390275,0.18485862,0.071679875,0.0,0.0,0.23013012,0.14335975,0.041498873,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.17731337,0.33576363,0.06790725,0.0,0.07922512,0.15845025,0.0,0.03772625,0.45648763,0.56212115,0.3772625,0.65643674,0.875249,0.8865669,0.935611,0.9280658,0.42630664,0.42630664,0.49044126,1.1317875,2.6710186,5.2326307,3.5123138,3.1010978,2.8445592,2.252257,1.4939595,1.7165444,2.9313297,3.9650288,4.357382,4.395108,5.6287565,5.1760416,3.8443048,3.8065786,8.590267,9.125979,8.537451,7.0963078,5.43258,4.515832,7.0812173,9.74469,10.419991,8.484633,4.7610526,3.6141748,3.006782,2.5314314,1.9353566,1.1280149,0.9205205,1.2261031,1.5430037,1.7127718,1.9089483,2.674791,2.916239,3.0256453,3.1954134,3.4029078,2.584248,3.953711,5.413717,5.7872066,4.821415,3.0746894,2.0070364,1.6486372,1.7655885,1.8787673,2.1315331,1.8863125,2.0447628,2.867195,3.9688015,2.3692086,1.4939595,1.3694628,1.9881734,3.2821836,3.3651814,4.191386,5.828706,7.9451485,9.812597,8.103599,4.6629643,3.3161373,4.2404304,3.9989824,6.145606,8.258276,8.631766,7.0963078,5.0213637,4.961002,4.5309224,4.014073,4.2102494,6.470052,5.1760416,3.0860074,2.6446102,3.482133,2.3956168,1.9693103,4.2328854,8.620448,12.30253,10.178542,4.7572803,3.3953626,2.9916916,2.4371157,2.6106565,7.8319697,8.262049,7.115171,6.375736,6.790725,4.2630663,2.9464202,2.4371157,3.0105548,5.5985756,8.650629,8.096053,6.741681,6.6020937,8.91094,9.80128,8.495952,6.809588,5.8588867,6.043745,7.4811153,7.466025,7.1981683,7.164215,7.1264887,10.069136,12.570387,13.211733,11.970539,10.223814,8.356364,7.3415284,5.8928404,5.093044,8.36391,14.2944765,14.43029,10.770844,6.115425,4.0895257,3.6971724,3.8858037,5.881522,9.046755,10.880251,7.7414265,5.062863,3.5990841,3.62172,4.927048,4.5120597,5.0251365,6.3908267,8.235641,9.857869,10.33322,9.857869,10.93684,13.449409,14.634012,13.290957,9.567377,8.07719,10.925522,17.701157,15.588487,13.083464,11.604594,10.668983,7.8734684,6.9567204,9.540969,12.860879,15.475307,17.25976,15.377219,14.275613,14.807553,16.784409,18.980076,18.848034,19.24416,19.738375,19.68933,18.233097,15.818617,13.060828,10.967021,10.197406,11.076427,10.480352,11.729091,14.464244,15.17727,7.2170315,4.191386,5.3571277,6.771862,6.477597,4.485651,4.032936,2.7125173,1.8146327,1.4977322,0.77716076,1.6222287,2.674791,3.4368613,4.6931453,8.514814,6.058836,3.4142256,2.6446102,3.410453,2.9464202,2.9086938,2.8521044,2.2484846,1.6448646,2.6710186,2.6332922,2.0749438,1.1657411,0.3734899,0.45648763,1.2261031,0.9808825,3.2067313,7.0849895,7.4773426,3.2633207,1.9466745,1.9579924,2.2975287,2.516341,1.6033657,0.58475685,0.5055317,1.1506506,1.0525624,0.30935526,0.06790725,0.08677038,0.14335975,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.0452715,0.071679875,0.056589376,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.060362,0.030181,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.030181,0.030181,0.018863125,0.0150905,0.0150905,0.018863125,0.030181,0.018863125,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.033953626,0.0452715,0.056589376,0.09808825,0.18485862,0.31312788,0.45648763,0.35839936,0.5281675,1.0299267,1.418507,0.7469798,1.2713746,1.4411428,1.3166461,1.056335,0.8865669,1.7165444,2.252257,2.8181508,3.2105038,2.686109,1.6486372,0.9507015,0.5357128,0.30181,0.1056335,0.19240387,0.11317875,0.056589376,0.0754525,0.0754525,0.0754525,0.06790725,0.060362,0.060362,0.060362,0.049044125,0.0452715,0.0452715,0.056589376,0.090543,0.116951376,0.15845025,0.23013012,0.32067314,0.38103512,0.43007925,0.47912338,0.5583485,0.67152727,0.7922512,0.8186596,0.8601585,0.87147635,0.88279426,0.9922004,0.9318384,0.9695646,0.98842776,0.9997456,1.1431054,1.1431054,1.1431054,1.2223305,1.327964,1.267602,1.1091517,1.0789708,0.95447415,0.754525,0.7167987,0.58098423,0.36594462,0.18863125,0.09808825,0.060362,0.03772625,0.02263575,0.0150905,0.02263575,0.0452715,0.0452715,0.03772625,0.02263575,0.02263575,0.0452715,0.033953626,0.02263575,0.02263575,0.030181,0.030181,0.018863125,0.0150905,0.0150905,0.0150905,0.0150905,0.026408374,0.030181,0.030181,0.026408374,0.0150905,0.05281675,0.124496624,0.17354076,0.18863125,0.21503963,0.26408374,0.27540162,0.29426476,0.31312788,0.29049212,0.05281675,0.08677038,0.090543,0.241448,0.38480774,0.0,0.05281675,0.12826926,0.10186087,0.003772625,0.02263575,0.1056335,0.29426476,0.241448,0.011317875,0.05281675,0.018863125,0.00754525,0.003772625,0.00754525,0.00754525,0.041498873,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.08677038,0.00754525,0.033953626,0.23390275,0.6413463,2.7841973,5.5495315,5.2099953,1.7240896,0.8224323,1.659955,3.5651307,6.039973,3.1614597,1.1808317,0.3169005,0.2678564,0.22258487,0.094315626,0.041498873,0.018863125,0.00754525,0.026408374,0.09808825,0.08299775,0.03772625,0.0,0.0,0.0452715,0.041498873,0.026408374,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.094315626,0.14335975,0.120724,0.120724,0.02263575,0.0,0.011317875,0.033953626,0.06790725,0.0150905,0.07922512,0.09808825,0.030181,0.0,0.056589376,0.4074435,0.48666862,0.29049212,0.3772625,0.38103512,0.422534,0.55080324,0.7130261,0.7696155,0.45648763,1.388326,3.1916409,4.98741,5.3910813,2.1579416,2.2296214,3.5236318,4.3007927,3.1916409,2.3956168,2.584248,3.2784111,4.2291126,5.406172,7.001992,5.8513412,4.191386,3.9461658,6.700182,8.348819,8.390318,7.907422,6.971811,4.6516466,5.270357,7.586749,9.371201,9.5183325,8.069645,6.5002327,4.485651,3.0671442,2.4182527,1.8372684,1.599593,2.1013522,2.1654868,1.7655885,2.0296721,3.0331905,2.686109,2.3465726,2.4333432,2.425798,2.625747,3.6481283,4.534695,4.561104,3.2331395,1.871222,1.8863125,2.4861598,2.8106055,1.9240388,1.8900851,2.746471,3.4859054,3.5877664,3.0143273,2.1768045,3.138824,4.8968673,5.7306175,3.2067313,2.5201135,2.7389257,4.38379,6.752999,7.907422,5.4476705,3.7386713,3.3463185,3.9084394,4.146115,4.074435,4.961002,5.6853456,5.3609,3.3236825,4.191386,4.508287,4.719554,4.8930945,4.7120085,3.1916409,2.7841973,3.3312278,4.217795,4.3611546,5.3873086,7.6886096,9.371201,8.873214,4.9421387,3.1237335,2.8445592,3.1539145,3.572676,4.085753,7.533932,7.164215,6.6586833,7.884786,10.929295,9.250477,5.926794,3.6481283,4.014073,7.5301595,14.517061,14.6302395,11.355601,8.231868,8.850578,8.548768,6.9755836,6.273875,7.281166,9.544742,7.364164,5.847569,5.0666356,5.353355,7.3075747,8.756263,8.7600355,8.918486,9.393836,8.918486,5.987156,4.715781,4.7648253,5.8098426,7.567886,9.525878,10.917976,10.299266,7.5188417,3.7348988,2.1051247,1.5430037,2.3654358,4.1800685,5.873977,5.100589,4.236658,3.6971724,3.802806,4.7572803,4.3800178,5.0854983,6.470052,8.043237,9.1976595,8.854351,8.137552,9.122208,11.321648,11.668729,18.184053,16.06761,11.668729,9.378746,11.634775,12.042219,10.174769,7.835742,6.1229706,5.406172,6.1229706,8.7600355,11.4838705,13.841762,16.758,18.606586,17.655886,15.599804,14.219024,15.380992,20.462717,21.145563,18.142553,13.996439,13.072145,12.423254,10.665211,9.880505,11.121698,14.422746,11.461235,10.27663,11.321648,12.174261,7.533932,5.904158,4.636556,3.429316,2.7238352,3.6934,4.90064,4.293247,3.2557755,2.293756,1.0450171,1.177059,1.7429527,2.6521554,3.3915899,3.0218725,2.1692593,2.8822856,3.3915899,3.2784111,3.470815,4.2819295,4.1612053,4.0404816,4.2291126,4.402653,3.4179983,4.0593443,4.82896,4.3196554,1.2034674,2.9766011,3.6707642,6.2927384,10.695392,13.5663595,7.967784,3.5274043,2.0070364,2.8521044,3.187868,2.9464202,2.2975287,1.6939086,1.2298758,0.62625575,0.28294688,0.13204187,0.116951376,0.14713238,0.1056335,0.10940613,0.07922512,0.060362,0.08299775,0.16976812,0.094315626,0.10186087,0.116951376,0.094315626,0.02263575,0.026408374,0.11317875,0.40367088,0.7582976,0.7582976,0.47535074,0.24899325,0.09808825,0.02263575,0.011317875,0.003772625,0.0,0.0,0.003772625,0.02263575,0.026408374,0.030181,0.0452715,0.06413463,0.071679875,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.003772625,0.011317875,0.018863125,0.02263575,0.030181,0.030181,0.018863125,0.0150905,0.0150905,0.0150905,0.018863125,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.124496624,1.1016065,1.0940613,0.10940613,0.033953626,0.056589376,0.12826926,0.25276586,0.36971724,0.35839936,0.33953625,1.0186088,1.8334957,2.033445,0.68661773,0.965792,1.690136,2.0749438,1.7731338,0.84884065,1.2298758,1.50905,1.7580433,2.3956168,4.1762958,2.7087448,1.3958713,1.7052265,2.5578396,0.35085413,0.62248313,0.32444575,0.06413463,0.041498873,0.05281675,0.041498873,0.030181,0.033953626,0.049044125,0.049044125,0.0452715,0.05281675,0.06790725,0.08299775,0.07922512,0.0754525,0.08677038,0.120724,0.17731337,0.24899325,0.3169005,0.4074435,0.5055317,0.6073926,0.7205714,0.73566186,0.7809334,0.83752275,0.8903395,0.94315624,0.98842776,1.086516,1.1732863,1.1695137,0.97333723,1.0412445,1.2713746,1.5203679,1.7014539,1.7655885,1.7052265,1.5769572,1.2789198,0.8978847,0.7054809,0.6375736,0.6828451,0.6413463,0.45648763,0.1961765,0.10186087,0.056589376,0.041498873,0.03772625,0.033953626,0.041498873,0.05281675,0.0452715,0.030181,0.033953626,0.030181,0.030181,0.033953626,0.041498873,0.030181,0.018863125,0.02263575,0.026408374,0.026408374,0.0150905,0.026408374,0.030181,0.030181,0.026408374,0.0150905,0.071679875,0.16976812,0.23013012,0.24522063,0.29803738,0.241448,0.21881226,0.23013012,0.26031113,0.26408374,0.241448,0.120724,0.07922512,0.16222288,0.241448,0.026408374,0.011317875,0.05281675,0.090543,0.08677038,0.0,0.06790725,0.1659955,0.13204187,0.0,0.00754525,0.033953626,0.018863125,0.0,0.0,0.0,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.10940613,0.1056335,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20372175,0.70170826,0.8224323,0.4979865,0.26408374,0.05281675,0.76207024,4.504514,9.163706,8.401636,2.3993895,1.5656394,2.3088465,2.848332,3.2331395,1.7731338,0.8526133,0.38480774,0.23013012,0.17354076,0.08299775,0.041498873,0.02263575,0.011317875,0.0150905,0.033953626,0.060362,0.060362,0.03772625,0.03772625,0.0150905,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.071679875,0.060362,0.060362,0.011317875,0.0,0.0,0.0,0.00754525,0.0,0.041498873,0.041498873,0.0,0.0,0.02263575,0.15845025,0.2565385,0.32821837,0.52439487,0.4678055,0.35839936,0.38858038,0.58475685,0.8186596,0.7130261,1.4864142,3.863168,6.25124,4.7535076,1.9693103,2.897376,4.8025517,5.5797124,3.7537618,3.150142,3.308592,3.229367,3.2520027,5.040227,8.635539,7.937603,5.6513925,4.2781568,6.1531515,7.01331,7.092535,6.934085,6.2323766,3.8141239,3.7650797,5.7079816,7.515069,8.09228,7.4018903,6.0324273,4.1989317,2.8407867,2.2484846,2.0673985,2.082489,2.3013012,2.0598533,1.6788181,2.4710693,3.1237335,2.9237845,2.8634224,2.9426475,2.1654868,2.7540162,2.9841464,3.0105548,2.7804246,2.033445,1.4373702,2.2975287,3.7386713,4.5535583,3.218049,2.704972,3.8405323,5.20245,5.515578,3.6481283,2.625747,4.3611546,6.9189944,7.9262853,4.5799665,2.8747404,2.2975287,3.0105548,4.195159,4.032936,2.9237845,3.6028569,5.2288585,6.5002327,5.6551647,4.1536603,5.081726,6.3229194,6.1833324,3.4029078,4.346064,5.753253,5.8928404,4.5007415,2.7615614,5.1647234,8.145098,8.190369,5.8588867,5.775889,7.967784,7.541477,5.798525,3.942393,3.0822346,4.7308717,5.828706,5.802297,5.3571277,6.4964604,7.220804,5.666483,4.930821,6.017337,7.8244243,6.779407,4.5761943,3.218049,4.025391,7.6622014,13.057055,12.679792,10.137043,8.073418,8.201687,7.2396674,6.620957,7.073672,7.9225125,7.0812173,4.123479,3.5538127,4.032936,5.1043615,7.1981683,7.8206515,7.360391,7.4169807,8.073418,7.9225125,5.6476197,5.764571,7.0284004,8.141325,7.7640624,7.5263867,7.8244243,7.6848373,6.6058664,4.5422406,3.029418,1.8561316,1.6524098,2.4031622,3.470815,3.4179983,3.2935016,3.229367,3.4670424,4.349837,4.1574326,5.492942,7.141579,8.333729,8.710991,7.2170315,6.330465,7.537705,9.997457,10.540714,14.747191,13.879487,11.121698,9.035437,9.548513,9.378746,7.2623034,5.383536,5.040227,6.63982,8.933576,10.978339,11.959221,12.672247,15.524352,19.217752,19.11589,16.399601,13.249459,12.83447,15.871433,15.886524,13.671993,11.219787,11.706455,12.31762,11.589504,10.785934,10.997202,13.117417,9.756008,8.058327,9.650374,12.132762,9.06939,8.4544525,6.651138,4.436607,2.727608,2.5691576,2.8106055,4.4177437,3.8141239,1.4034165,1.5882751,0.91297525,0.9318384,1.297783,1.6410918,1.5580941,1.0110635,2.3465726,2.9954643,2.5880208,2.987919,4.4441524,4.666737,5.6400743,7.0510364,6.3116016,3.2821836,4.9044123,7.145352,7.4697976,4.8402777,5.3873086,4.5761943,5.6325293,8.793989,11.317875,7.1906233,4.5912848,3.832987,4.1008434,3.4594972,3.640583,3.6896272,3.4255435,2.8106055,1.9466745,1.5052774,1.1016065,0.7167987,0.3734899,0.13204187,0.150905,0.11317875,0.116951376,0.16976812,0.17731337,0.13204187,0.13958712,0.124496624,0.0754525,0.041498873,0.09808825,0.116951376,0.4074435,0.95447415,1.4298248,0.91674787,0.5470306,0.29426476,0.13958712,0.071679875,0.030181,0.00754525,0.003772625,0.011317875,0.0150905,0.0150905,0.030181,0.0452715,0.056589376,0.0452715,0.00754525,0.02263575,0.0452715,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.011317875,0.00754525,0.00754525,0.0,0.00754525,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.003772625,0.011317875,0.018863125,0.02263575,0.02263575,0.0150905,0.02263575,0.02263575,0.0150905,0.0150905,0.02263575,0.018863125,0.0150905,0.0150905,0.0150905,0.11317875,0.8337501,0.88279426,0.2263575,0.0754525,0.07922512,0.10186087,0.16222288,0.2565385,0.392353,0.7997965,1.5882751,2.0900342,2.2409391,2.5578396,2.7200627,2.8558772,2.5917933,1.9806281,1.4977322,1.50905,3.4557245,3.6971724,2.41448,3.6141748,3.2255943,2.123988,2.1654868,2.8558772,1.3468271,4.776143,2.8747404,0.6526641,0.071679875,0.0452715,0.026408374,0.011317875,0.011317875,0.018863125,0.018863125,0.026408374,0.20749438,0.5470306,0.7394345,0.17731337,0.09808825,0.071679875,0.0754525,0.094315626,0.13204187,0.20372175,0.36971724,0.49044126,0.543258,0.6375736,0.68661773,0.70170826,0.7092535,0.73566186,0.80356914,0.91297525,1.0638802,1.2034674,1.2487389,1.0789708,1.1846043,1.3505998,1.50905,1.6486372,1.8184053,1.8976303,1.7882242,1.5920477,1.3430545,1.0223814,0.87902164,0.9242931,0.98465514,0.935611,0.66775465,0.36971724,0.18863125,0.10186087,0.06790725,0.041498873,0.03772625,0.041498873,0.03772625,0.033953626,0.041498873,0.041498873,0.041498873,0.041498873,0.041498873,0.030181,0.026408374,0.026408374,0.026408374,0.02263575,0.02263575,0.02263575,0.02263575,0.026408374,0.030181,0.033953626,0.124496624,0.25276586,0.331991,0.35462674,0.392353,0.29426476,0.23013012,0.21881226,0.23767537,0.24899325,0.26031113,0.120724,0.049044125,0.041498873,0.056589376,0.026408374,0.041498873,0.17354076,0.25276586,0.1961765,0.00754525,0.0452715,0.033953626,0.011317875,0.0,0.00754525,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.19240387,0.18863125,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.116951376,0.58475685,1.4901869,2.2786655,2.5125682,2.0749438,1.1506506,0.38480774,1.20724,4.8138695,8.990166,8.09228,3.078462,2.0447628,1.9353566,1.4713237,1.1506506,0.9393836,0.724344,0.44894236,0.17731337,0.11317875,0.06790725,0.03772625,0.02263575,0.0150905,0.00754525,0.00754525,0.041498873,0.05281675,0.041498873,0.060362,0.030181,0.00754525,0.011317875,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.03772625,0.0150905,0.00754525,0.011317875,0.011317875,0.011317875,0.030181,0.00754525,0.0,0.071679875,0.23013012,0.4376245,0.43385187,0.3055826,0.35839936,0.5772116,0.62248313,0.6413463,1.3204187,4.014073,6.722818,4.1083884,2.123988,3.399135,5.4250345,6.1078796,3.7914882,4.055572,4.032936,3.429316,3.1350515,5.2137675,8.835487,8.627994,6.368191,4.429062,5.7570257,6.258785,6.085244,5.7079816,5.1571784,4.0178456,4.3196554,5.572167,6.25124,6.0512905,5.9192486,5.7004366,4.67051,3.5160866,2.637065,2.142851,2.1164427,2.2748928,2.0598533,1.7354075,2.4220252,3.1954134,3.4066803,3.6179473,3.6556737,2.6106565,2.7502437,2.6408374,2.1956677,1.8070874,2.354118,2.293756,2.8822856,4.063117,4.8930945,3.5236318,2.7125173,3.7009451,5.100589,5.5570765,3.7386713,3.0897799,4.2291126,5.847569,6.477597,4.5007415,2.927557,2.444661,2.7615614,3.097325,2.1843498,2.335255,3.8103511,5.696664,6.620957,4.738417,3.7273536,5.1571784,6.651138,6.3531003,2.938875,4.7044635,7.6886096,7.858378,4.9119577,2.2975287,6.5945487,11.23865,10.789707,6.0814714,4.2404304,6.047518,4.606375,2.9652832,3.983892,10.344538,12.083718,9.710737,7.043491,6.2889657,8.024373,5.885295,3.7650797,3.0671442,3.5877664,3.4670424,3.1161883,2.6068838,2.5502944,3.4934506,5.9305663,9.246704,9.061845,7.6848373,6.5266414,6.092789,5.221313,5.3382645,5.7872066,5.617439,3.6179473,2.5767028,4.5497856,5.9909286,5.983383,6.228604,6.360646,6.820906,7.1906233,7.232122,6.85486,6.066381,6.934085,8.028146,8.303548,7.0812173,6.3644185,5.670255,5.3684454,5.534441,5.934339,5.3759904,3.7877154,2.5201135,2.2258487,2.8785129,2.8521044,2.463524,2.1881225,2.335255,3.0558262,3.7952607,5.881522,7.858378,8.835487,8.511042,5.938112,4.557331,5.4174895,8.013056,10.291721,11.796998,11.54046,10.087999,8.537451,8.511042,7.647111,5.4401255,4.432834,6.771862,14.200161,13.275867,13.58145,13.166461,12.294985,13.449409,17.391802,18.372684,16.459963,13.36641,12.453435,13.449409,12.860879,11.548005,10.525623,10.955703,14.6302395,14.916959,12.611885,10.401127,12.879742,13.52486,12.713746,13.981348,16.290195,13.9888935,11.581959,14.418973,14.554788,10.495442,7.201941,6.0550632,6.7341356,5.062863,1.7127718,2.2258487,1.3543724,0.9507015,0.7054809,0.7092535,1.4298248,1.2336484,1.8033148,1.9240388,1.5845025,1.9881734,2.969056,3.2972744,4.4818783,6.085244,5.7079816,3.1199608,4.2064767,5.621211,6.039973,6.1644692,5.8136153,3.9688015,3.7235808,5.311856,6.1116524,4.168751,4.353609,4.7308717,4.395108,3.4594972,3.772625,4.636556,5.070408,4.7572803,4.002755,3.338773,2.637065,1.9278114,1.2562841,0.7092535,0.58475685,0.3961256,0.2867195,0.271629,0.2565385,0.2678564,0.38480774,0.35085413,0.20372175,0.241448,0.24899325,0.13958712,0.24522063,0.7507524,1.6750455,1.9202662,1.569412,1.1317875,0.8299775,0.58098423,0.38858038,0.19994913,0.071679875,0.030181,0.056589376,0.08299775,0.06790725,0.049044125,0.041498873,0.026408374,0.018863125,0.033953626,0.049044125,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.02263575,0.0150905,0.0150905,0.00754525,0.02263575,0.02263575,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.00754525,0.0150905,0.02263575,0.02263575,0.0150905,0.00754525,0.02263575,0.018863125,0.0150905,0.0150905,0.0150905,0.06413463,0.31312788,0.40367088,0.271629,0.15467763,0.181086,0.124496624,0.116951376,0.27917424,0.72811663,1.4637785,1.9844007,2.161714,2.5125682,4.1800685,4.08198,3.078462,2.1654868,1.8523588,2.1503963,1.9429018,3.8367596,4.908185,4.436607,3.893349,3.561358,2.3993895,1.8787673,2.0485353,1.5731846,5.4476705,3.7763977,1.3166461,0.2263575,0.0754525,0.03772625,0.0150905,0.00754525,0.011317875,0.02263575,0.124496624,0.62625575,1.1657411,1.2562841,0.29426476,0.15467763,0.09808825,0.1056335,0.15467763,0.211267,0.3961256,0.55457586,0.59230214,0.5319401,0.5017591,0.6073926,0.62248313,0.62248313,0.6526641,0.7469798,0.80734175,0.97333723,1.1242423,1.1808317,1.1016065,1.2525115,1.3430545,1.4449154,1.5807298,1.720317,1.9353566,1.8976303,1.8297231,1.7580433,1.50905,1.2449663,1.177059,1.146878,1.0978339,1.0638802,0.8224323,0.5470306,0.3169005,0.1659955,0.08677038,0.056589376,0.041498873,0.03772625,0.03772625,0.041498873,0.041498873,0.041498873,0.0452715,0.0452715,0.03772625,0.03772625,0.033953626,0.026408374,0.02263575,0.030181,0.018863125,0.0150905,0.026408374,0.049044125,0.071679875,0.18863125,0.30181,0.35462674,0.35462674,0.362172,0.29803738,0.2565385,0.24522063,0.25276586,0.2565385,0.060362,0.060362,0.041498873,0.018863125,0.003772625,0.02263575,0.06413463,0.271629,0.35462674,0.241448,0.08677038,0.049044125,0.018863125,0.0,0.003772625,0.0150905,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16976812,0.16976812,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06790725,0.1056335,0.32821837,1.2411937,2.6974268,3.440634,3.6254926,3.2255943,2.04099,1.388326,1.8863125,3.6669915,5.4967146,4.745962,2.938875,1.6637276,0.8563859,0.5093044,0.66020936,0.83752275,0.73566186,0.44139713,0.13204187,0.06790725,0.056589376,0.03772625,0.02263575,0.011317875,0.003772625,0.0,0.00754525,0.00754525,0.011317875,0.049044125,0.030181,0.011317875,0.018863125,0.041498873,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.071679875,0.011317875,0.011317875,0.018863125,0.018863125,0.02263575,0.060362,0.011317875,0.0,0.00754525,0.03772625,0.094315626,0.18863125,0.241448,0.4074435,0.6488915,0.72811663,0.331991,1.0751982,3.783943,6.3832817,3.893349,2.082489,2.8747404,4.727099,5.715527,3.5085413,4.304565,4.22534,4.1762958,4.82896,6.63982,7.77538,7.54525,6.221059,5.093044,6.488915,6.5945487,5.715527,4.889322,4.659192,5.081726,5.956975,6.809588,6.296511,4.9345937,5.111907,5.8513412,5.481624,4.606375,3.5500402,2.3578906,1.9994912,2.293756,2.3692086,2.071171,1.961765,3.3161373,4.0782075,4.429062,4.293247,3.31991,2.867195,3.187868,2.8030603,2.1466236,3.5689032,3.3123648,2.8785129,3.0256453,3.361409,2.3428001,1.6788181,2.3277097,3.1954134,3.5538127,3.0558262,3.610402,3.6179473,3.482133,3.4745877,3.7575345,3.308592,3.1727777,3.3425457,3.4330888,2.7011995,2.9728284,3.5047686,4.002755,3.8971217,2.3390274,3.1048703,4.715781,5.873977,5.3646727,2.0598533,4.957229,9.0543,9.435335,5.8664317,2.8256962,5.3759904,8.7751255,8.405409,4.3611546,1.4411428,1.7693611,1.3204187,2.8558772,9.001483,22.243397,20.251451,11.9064045,6.156924,5.8928404,7.9262853,4.1008434,2.505023,2.4899325,2.806833,1.5845025,1.5958204,1.8599042,2.4597516,3.4330888,4.7572803,7.194396,7.3792543,6.3116016,4.8742313,3.874486,3.7198083,3.7235808,3.180323,2.3314822,2.3654358,4.2706113,7.9526935,8.967529,6.862405,5.1835866,5.572167,6.7039547,6.7680893,5.726845,5.304311,5.87775,6.5266414,6.851087,6.722818,6.2851934,6.247467,5.7683434,5.59103,6.0211096,6.9567204,7.2283497,6.013564,4.3800178,3.2142766,3.2331395,3.059599,1.9881734,1.1921495,1.1317875,1.5618668,3.3915899,5.8098426,7.835742,8.635539,7.4999785,4.768598,3.2142766,3.5990841,6.149379,10.54826,12.377983,12.019584,9.861642,7.3490734,6.9793563,6.224831,4.447925,4.085753,8.20546,20.474035,15.690348,15.196134,14.78869,13.264549,12.408164,15.482853,17.4333,17.308804,15.652621,14.48688,15.120681,14.64533,13.400364,11.668729,9.654147,15.430037,16.648594,13.645585,10.38981,14.460471,18.949896,18.463226,18.233097,19.28566,18.470772,13.860624,21.779364,24.371157,18.229324,14.422746,14.25675,11.136789,6.934085,3.4859054,2.5691576,1.9994912,1.6071383,1.1091517,0.8865669,1.9542197,2.5578396,1.9240388,1.4562333,1.5618668,1.6373192,0.9997456,0.965792,1.4524606,2.203213,2.8030603,2.776652,2.7841973,2.5276587,2.5616124,4.2894745,3.92353,2.6182017,2.2711203,2.7917426,2.1164427,1.6335466,2.938875,3.7273536,3.500996,3.5462675,3.7688525,5.032682,5.938112,6.0248823,5.753253,5.036454,4.402653,3.7499893,3.0407357,2.305074,1.9051756,1.3845534,0.9922004,0.8299775,0.83752275,0.8639311,1.1016065,1.0601076,0.7469798,0.6526641,0.513077,0.35462674,0.33576363,0.633801,1.4449154,2.6936543,2.5616124,2.071171,1.6675003,1.2261031,0.80734175,0.41876137,0.14713238,0.03772625,0.09808825,0.16222288,0.10940613,0.06413463,0.056589376,0.056589376,0.05281675,0.033953626,0.0150905,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.02263575,0.018863125,0.0150905,0.02263575,0.041498873,0.041498873,0.03772625,0.030181,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.003772625,0.011317875,0.0,0.011317875,0.0150905,0.0150905,0.011317875,0.003772625,0.011317875,0.0150905,0.0150905,0.018863125,0.018863125,0.030181,0.06790725,0.13958712,0.21503963,0.21503963,0.28294688,0.17354076,0.14713238,0.3772625,0.9808825,1.7919968,1.8938577,2.0900342,2.9615107,4.878004,4.4101987,2.3465726,1.1808317,1.6222287,2.6106565,2.5427492,3.7235808,6.0776987,7.84706,5.587258,4.0706625,2.463524,1.4147344,1.0336993,0.875249,2.2598023,2.7653341,2.071171,0.724344,0.150905,0.08677038,0.0452715,0.071679875,0.16976812,0.29426476,1.1959221,1.8863125,2.0975795,1.6750455,0.59230214,0.45648763,0.5394854,0.663982,0.73566186,0.7432071,0.814887,0.7884786,0.724344,0.633801,0.482896,0.56589377,0.5696664,0.58475685,0.6451189,0.73566186,0.7092535,0.8337501,0.95447415,0.98842776,0.9318384,1.0978339,1.1921495,1.3694628,1.5845025,1.6071383,1.8749946,1.8674494,1.8485862,1.8863125,1.8485862,1.5618668,1.4411428,1.2336484,1.0110635,1.1732863,1.2298758,1.0299267,0.7205714,0.422534,0.21503963,0.120724,0.0754525,0.05281675,0.041498873,0.033953626,0.03772625,0.041498873,0.0452715,0.049044125,0.049044125,0.049044125,0.041498873,0.033953626,0.033953626,0.033953626,0.02263575,0.02263575,0.0452715,0.08299775,0.13204187,0.24899325,0.29426476,0.27917424,0.241448,0.23390275,0.2565385,0.28294688,0.29803738,0.29049212,0.26408374,0.0,0.0,0.090543,0.090543,0.02263575,0.1056335,0.02263575,0.0,0.018863125,0.11317875,0.38103512,0.23390275,0.08677038,0.00754525,0.003772625,0.0150905,0.11317875,0.08299775,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33953625,0.5357128,0.46026024,0.35085413,0.6451189,1.0110635,0.784706,0.392353,1.358145,3.6179473,3.8895764,2.9841464,2.0598533,2.6106565,1.8787673,0.9808825,0.46026024,0.3772625,0.3055826,0.3169005,0.24899325,0.150905,0.06790725,0.030181,0.07922512,0.08299775,0.05281675,0.0150905,0.0150905,0.003772625,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.056589376,0.1056335,0.27917424,0.5017591,0.5093044,0.70170826,2.1654868,0.5319401,0.5998474,2.595566,4.930821,4.2102494,1.599593,1.3015556,2.6634734,4.0216184,2.71629,2.203213,3.904667,6.458734,8.518587,8.790216,7.4811153,6.790725,6.802043,8.050782,11.506506,7.8810134,5.2326307,4.274384,4.5912848,4.6554193,4.9723196,7.2094865,7.6923823,5.96452,4.8063245,3.6707642,3.2859564,3.500996,3.7386713,3.006782,2.565385,2.4484336,2.5880208,2.6597006,2.0598533,3.3651814,5.028909,5.885295,5.3458095,3.4179983,3.8443048,5.0968165,4.927048,3.470815,3.2520027,1.7240896,1.1431054,1.0751982,1.1242423,0.91674787,0.9997456,1.1883769,1.5958204,2.2862108,3.2482302,4.8968673,5.2175403,5.0175915,5.2099953,6.820906,6.7831798,4.8968673,3.1237335,2.323937,2.2748928,1.6260014,1.4449154,1.9353566,2.9728284,4.1197066,5.560849,6.2851934,6.2851934,5.406172,3.3425457,5.2326307,7.884786,7.9225125,4.9760923,1.6788181,1.7769064,2.1013522,2.0673985,2.003264,3.1727777,3.0520537,1.7391801,4.3875628,12.528888,24.061802,16.837225,9.876732,5.572167,4.727099,6.5455046,4.032936,3.9989824,4.908185,5.270357,3.6481283,2.584248,2.3088465,3.187868,5.4288073,9.076936,10.1294985,8.058327,6.0248823,5.2779026,5.142088,5.836251,5.0515447,4.244203,4.146115,4.745962,7.492433,8.013056,7.073672,5.904158,6.2097406,8.737399,7.6923823,4.696918,2.071171,2.837014,3.6066296,4.715781,6.33801,8.039464,8.7751255,9.5183325,10.216269,10.393582,9.374973,6.2851934,5.8211603,6.9227667,7.277394,5.994701,3.6028569,3.2105038,2.1164427,1.478869,1.599593,1.8938577,3.1727777,4.7308717,6.0776987,6.1720147,3.3878171,2.71629,2.9803739,4.515832,7.424526,11.551778,13.758763,12.721292,9.382519,5.73439,4.8063245,3.8178966,2.6936543,2.3805263,3.7499893,7.5829763,11.393328,15.675257,17.286167,16.350557,16.263786,18.010511,20.590988,22.756474,22.748928,18.293459,16.343012,16.999449,17.271078,14.966003,8.66572,7.752744,9.691874,11.559323,12.483616,13.656902,10.216269,6.115425,5.6815734,9.156161,12.694883,12.694883,13.381501,10.287949,6.330465,11.812089,18.35382,13.743673,7.707473,4.327201,2.0447628,1.3015556,1.7919968,1.6335466,1.4637785,4.45547,5.772116,4.044254,3.663219,4.881777,3.783943,1.2336484,0.60362,0.8865669,1.1808317,0.7167987,1.0110635,2.6936543,4.9345937,5.873977,2.6408374,1.7014539,1.8033148,2.1805773,2.384299,2.2748928,1.8221779,1.3996439,1.5882751,2.6068838,4.304565,4.398881,4.8100967,5.2665844,5.6778007,6.119198,5.764571,6.043745,6.145606,5.798525,5.247721,4.6629643,3.682082,2.969056,2.6898816,2.5314314,2.4710693,2.546522,2.4522061,1.9957186,1.1280149,0.9205205,1.0148361,1.2864652,1.4298248,0.9922004,1.0412445,1.327964,1.4864142,1.3505998,0.94692886,0.4074435,0.17354076,0.06413463,0.0,0.0,0.071679875,0.090543,0.09808825,0.1056335,0.1056335,0.08299775,0.056589376,0.041498873,0.026408374,0.0150905,0.0150905,0.02263575,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.02263575,0.02263575,0.0452715,0.0452715,0.026408374,0.026408374,0.05281675,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.030181,0.041498873,0.026408374,0.0452715,0.1056335,0.1659955,0.15467763,0.116951376,0.090543,0.11317875,0.19994913,0.9808825,0.9280658,1.5920477,3.3651814,5.4778514,4.8440504,2.4974778,1.1053791,1.5958204,3.1576872,3.953711,9.552286,12.310076,10.227587,6.94163,5.1232247,3.5047686,1.9542197,0.72811663,0.47157812,1.6825907,3.2935016,3.4330888,1.9202662,0.26031113,0.18485862,0.120724,0.3055826,0.7469798,1.237421,4.8138695,5.028909,4.0291634,2.8634224,1.4939595,1.4600059,2.173032,2.6483827,2.5276587,2.0749438,1.0148361,0.55457586,0.62248313,0.9205205,0.94692886,0.77338815,0.58475685,0.48666862,0.49044126,0.5017591,0.5772116,0.62248313,0.70170826,0.77338815,0.68661773,0.73566186,0.83752275,1.1091517,1.4260522,1.448688,1.6071383,1.4637785,1.4222796,1.5430037,1.5580941,1.5430037,1.6222287,1.5316857,1.2487389,0.9922004,1.1242423,1.2864652,1.2562841,0.9620194,0.47157812,0.241448,0.1358145,0.08299775,0.0452715,0.0452715,0.056589376,0.05281675,0.05281675,0.060362,0.060362,0.060362,0.05281675,0.0452715,0.0452715,0.0452715,0.0452715,0.056589376,0.08677038,0.14335975,0.23013012,0.29049212,0.2678564,0.21503963,0.17354076,0.19994913,0.30935526,0.3734899,0.36594462,0.29803738,0.21503963,0.049044125,0.06790725,0.09808825,0.14713238,0.16222288,0.02263575,0.02263575,0.018863125,0.011317875,0.02263575,0.0754525,0.0452715,0.06790725,0.08299775,0.116951376,0.28294688,0.2263575,0.090543,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.1659955,0.32821837,0.33953625,0.21503963,0.094315626,0.13204187,0.20372175,0.6752999,1.3732355,1.5769572,4.168751,4.142342,2.9841464,1.7354075,0.98465514,0.8865669,0.56589377,0.3470815,0.2867195,0.18485862,0.1358145,0.0754525,0.07922512,0.13958712,0.150905,0.16222288,0.11317875,0.05281675,0.0150905,0.0150905,0.003772625,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0150905,0.0150905,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.0452715,0.0,0.033953626,0.16976812,0.33576363,0.21881226,0.06413463,0.003772625,0.02263575,0.3772625,0.3772625,0.24899325,0.19240387,0.38858038,0.40367088,0.44139713,0.482896,0.6375736,1.1657411,0.7394345,0.80356914,1.8825399,3.6179473,4.772371,2.3767538,2.535204,3.482133,3.7462165,2.1654868,1.81086,2.3201644,4.7421894,8.122461,9.533423,8.186596,7.9036493,7.877241,8.59404,11.834724,6.187105,4.327201,4.889322,6.25124,6.4964604,6.326692,7.696155,7.779153,5.692891,2.5125682,2.5691576,2.7653341,2.969056,3.1010978,3.138824,3.6292653,3.5085413,3.2633207,3.1916409,3.4029078,5.715527,6.25124,5.6476197,4.436607,3.0633714,3.0030096,3.6179473,3.7084904,2.8219235,1.2713746,0.6451189,0.5357128,0.7469798,1.026154,1.0751982,1.2562841,1.4109617,1.4562333,1.5769572,2.1881225,3.953711,4.5724216,4.2027044,3.7273536,4.7836885,5.311856,4.036709,2.7238352,2.3654358,3.1652324,2.8294687,2.2069857,2.2673476,3.0369632,3.6179473,3.663219,3.5424948,3.7613072,3.7877154,2.0485353,3.7952607,4.9949555,4.4818783,2.6144292,1.3015556,3.2142766,4.991183,4.221567,1.8976303,2.4182527,3.0860074,2.5729303,2.584248,4.1498876,7.6207023,5.2854476,3.5387223,3.1916409,3.6858547,3.1048703,3.2557755,5.6815734,6.900131,5.5268955,2.293756,3.0369632,4.4516973,5.9305663,7.281166,8.726082,8.477088,6.790725,5.674028,5.945657,7.2170315,6.749226,5.028909,4.666737,6.300284,8.578949,8.443134,6.304056,4.398881,4.0970707,5.9192486,4.7044635,5.5759397,5.66271,4.376245,3.3878171,5.191132,7.699928,9.148616,9.367428,9.786189,8.880759,9.540969,11.291467,12.823153,12.00072,8.635539,6.330465,5.794752,6.19465,5.149633,2.2598023,1.3543724,1.3430545,1.6109109,2.003264,2.5125682,3.0558262,3.1576872,2.686109,1.8259505,2.4031622,3.1840954,4.4403796,6.2323766,8.424272,8.809079,7.5527954,6.405917,6.307829,7.383027,3.7273536,2.9086938,3.0860074,3.4029078,3.983892,7.0510364,9.97482,11.393328,11.449917,11.823407,13.81158,18.53868,23.631723,26.20088,22.847017,16.569368,17.542706,20.741892,21.371922,14.867915,12.1252165,16.524097,20.689075,21.609596,20.65135,17.237123,13.804035,11.114153,9.869187,10.691619,11.619685,12.268577,10.472807,7.4697976,7.8923316,13.713491,11.038701,11.18206,14.66042,11.234878,7.062354,5.4476705,5.2854476,5.692891,5.9682927,7.2585306,6.273875,6.273875,7.183078,5.613666,7.5075235,5.643847,3.8367596,2.9501927,0.9242931,1.7542707,4.217795,4.7044635,2.6710186,0.62625575,0.7997965,1.6071383,2.7841973,4.006528,4.8742313,4.8025517,3.5953116,2.848332,3.308592,4.889322,3.8141239,3.7537618,3.6368105,3.6971724,5.485397,7.9828744,8.262049,7.466025,6.7039547,7.043491,8.273367,8.537451,8.416726,7.967784,6.7454534,6.6058664,6.7114997,5.7570257,4.014073,3.361409,2.686109,2.093807,1.8938577,1.9957186,1.9089483,1.7127718,1.3091009,0.9242931,0.6790725,0.58098423,0.33576363,0.211267,0.21881226,0.2565385,0.10940613,0.06413463,0.049044125,0.05281675,0.071679875,0.08299775,0.09808825,0.13204187,0.16976812,0.18485862,0.16222288,0.150905,0.14335975,0.14713238,0.14335975,0.08677038,0.03772625,0.03772625,0.060362,0.06413463,0.02263575,0.00754525,0.011317875,0.02263575,0.030181,0.033953626,0.033953626,0.0452715,0.05281675,0.056589376,0.05281675,0.060362,0.03772625,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.011317875,0.003772625,0.0150905,0.003772625,0.011317875,0.0150905,0.018863125,0.018863125,0.02263575,0.018863125,0.026408374,0.05281675,0.094315626,0.090543,0.0754525,0.10186087,0.23390275,0.56589377,1.5430037,2.5276587,3.4896781,3.8971217,2.7200627,2.2107582,1.2789198,0.80356914,1.4034165,3.4632697,5.798525,9.725827,11.480098,9.861642,6.2361493,5.1571784,6.94163,6.356873,2.8596497,0.5696664,1.0940613,1.6939086,2.003264,1.6637276,0.29426476,0.241448,0.211267,0.24522063,0.4074435,0.79602385,2.5087957,2.8445592,3.078462,3.6934,4.376245,3.5764484,2.9652832,2.6710186,2.6144292,2.516341,2.625747,2.686109,2.4522061,1.9655377,1.5807298,1.3204187,1.1695137,1.0336993,0.87147635,0.68661773,0.44894236,0.4376245,0.513077,0.5772116,0.5885295,0.55080324,0.6187105,0.8111144,1.0902886,1.3392819,1.6637276,1.6788181,1.6561824,1.6561824,1.5316857,1.4713237,1.7278622,1.9051756,1.7769064,1.2864652,1.3807807,1.3619176,1.3166461,1.2638294,1.1581959,0.80734175,0.46026024,0.23767537,0.14335975,0.094315626,0.07922512,0.06413463,0.060362,0.06413463,0.071679875,0.08299775,0.1056335,0.12826926,0.13958712,0.120724,0.10940613,0.150905,0.23013012,0.3055826,0.31312788,0.29803738,0.27917424,0.2565385,0.26031113,0.34330887,0.5017591,0.7130261,0.73566186,0.5319401,0.24899325,0.05281675,0.0452715,0.0452715,0.08299775,0.116951376,0.00754525,0.026408374,0.026408374,0.02263575,0.0150905,0.0,0.00754525,0.033953626,0.0452715,0.056589376,0.13958712,0.10186087,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.018863125,0.05281675,0.071679875,0.09808825,0.12826926,0.21503963,0.44139713,0.9280658,0.56589377,0.633801,1.0072908,1.5845025,2.3013012,3.6783094,3.9084394,2.8181508,1.1091517,0.34330887,0.38858038,0.3169005,0.23390275,0.1659955,0.07922512,0.049044125,0.05281675,0.07922512,0.09808825,0.10186087,0.10186087,0.0754525,0.056589376,0.0452715,0.02263575,0.011317875,0.049044125,0.060362,0.030181,0.00754525,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05281675,0.06790725,0.049044125,0.02263575,0.08677038,0.18863125,0.14713238,0.06413463,0.02263575,0.06790725,0.22258487,0.26408374,0.29803738,0.41498876,0.7130261,0.9318384,1.0299267,1.1242423,1.1959221,1.0789708,1.0110635,1.0714256,1.5543215,2.6068838,4.255521,3.651901,3.4255435,4.1083884,4.7874613,3.0746894,2.1466236,2.7691069,5.6891184,9.778644,12.053536,11.234878,11.068882,10.174769,9.152389,10.582213,6.2097406,5.4363527,6.670001,8.314865,8.809079,7.2472124,6.7039547,5.802297,4.093298,2.082489,2.5540671,2.5767028,2.4295704,2.4484336,3.0445085,3.218049,3.0218725,3.218049,3.9273026,4.6252384,6.3908267,6.6360474,5.304311,3.3350005,2.6446102,2.3163917,2.505023,2.4484336,1.841041,0.87147635,1.2223305,1.418507,1.4071891,1.2864652,1.3166461,1.539231,1.4222796,1.327964,1.3204187,1.1619685,1.8674494,2.425798,2.5012503,2.2598023,2.3767538,2.425798,2.0598533,2.1202152,2.637065,2.837014,2.6031113,2.6634734,2.704972,2.6974268,2.8822856,3.0369632,3.4029078,3.712263,3.772625,3.4444065,4.195159,3.6783094,2.7653341,2.2447119,2.8256962,5.20245,6.530414,5.100589,2.123988,1.7240896,3.0897799,4.817642,5.081726,3.9725742,3.4896781,3.1576872,2.5804756,2.5578396,3.0331905,3.0935526,3.8254418,5.7683434,6.247467,4.825187,3.3274553,5.6589375,6.515323,6.0701537,5.081726,4.919503,5.511805,7.0359454,8.643084,9.665465,9.612649,8.182823,6.9152217,6.009792,5.5457587,5.481624,4.8025517,3.6783094,3.169005,3.9914372,6.549277,6.5756855,7.748972,7.786698,6.126743,3.9461658,5.292993,8.065872,9.710737,9.574923,8.914713,8.080963,9.457971,11.895086,13.328684,10.808571,8.91094,8.560086,9.027891,9.473062,8.933576,6.436098,5.1571784,4.7044635,4.357382,3.0369632,2.5616124,2.384299,2.161714,1.991946,2.4333432,3.470815,3.531177,3.6481283,4.285702,5.3194013,5.4740787,4.6214657,5.3986263,7.1302614,5.855114,3.4179983,3.5085413,4.266839,4.432834,3.3576362,4.0103,5.855114,7.3981175,7.9300575,7.515069,8.812852,14.667966,22.526344,27.687294,23.31105,16.497688,18.919714,25.069094,28.102283,19.844007,12.989148,13.88326,17.108854,19.896824,22.107582,22.266033,20.526854,16.373192,11.551778,10.072908,9.167479,9.850324,10.593531,10.306811,8.329956,10.989656,11.431054,13.177779,15.0905,11.355601,7.643338,7.043491,6.651138,6.0550632,7.3453007,8.75249,7.5037513,7.8961043,9.593785,7.6395655,9.937095,10.461489,9.963503,8.699674,6.4134626,2.7200627,4.38379,6.330465,5.8211603,2.4559789,2.335255,2.463524,3.561358,5.221313,5.9003854,6.8699503,6.375736,7.111398,8.616675,7.2962565,4.187614,5.2665844,5.696664,4.45547,4.346064,6.6247296,7.2170315,6.851087,6.5643673,7.7225633,9.382519,11.34051,12.679792,12.804289,11.404645,10.506761,9.507015,7.99042,6.296511,5.5495315,4.949684,4.214022,3.6707642,3.3048196,2.7502437,2.0900342,1.4562333,1.0940613,0.935611,0.5885295,0.5357128,0.43007925,0.49044126,0.6413463,0.49421388,0.32444575,0.25276586,0.271629,0.33576363,0.3772625,0.41876137,0.36971724,0.3169005,0.3169005,0.38103512,0.39989826,0.32067314,0.2678564,0.24522063,0.16976812,0.124496624,0.11317875,0.11317875,0.1056335,0.094315626,0.07922512,0.056589376,0.041498873,0.03772625,0.02263575,0.02263575,0.030181,0.030181,0.026408374,0.03772625,0.060362,0.049044125,0.030181,0.011317875,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.17731337,1.9994912,4.7610526,5.5759397,4.3083377,1.9353566,0.38480774,0.090543,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.00754525,0.00754525,0.00754525,0.011317875,0.011317875,0.011317875,0.02263575,0.018863125,0.0150905,0.018863125,0.026408374,0.049044125,0.056589376,0.05281675,0.14335975,0.452715,1.1581959,2.535204,3.8103511,3.9876647,3.1727777,2.5804756,3.2821836,3.3576362,3.187868,3.0445085,3.0822346,4.323428,6.360646,7.0585814,5.907931,3.9989824,3.399135,6.7756343,6.8435416,2.9652832,1.1355602,1.3128735,1.267602,1.0940613,0.79602385,0.2867195,0.3055826,0.331991,0.35085413,0.38858038,0.52062225,2.0975795,2.7200627,3.7575345,5.617439,7.7602897,5.1081343,2.795515,1.9730829,2.4710693,2.7879698,3.5349495,4.123479,3.9499383,3.2482302,3.0671442,2.916239,2.4333432,1.8863125,1.4298248,1.1242423,0.7432071,0.55457586,0.44894236,0.38480774,0.39989826,0.3772625,0.42630664,0.5394854,0.7205714,0.9808825,1.4298248,1.7127718,1.8863125,1.9466745,1.8448136,1.6637276,2.0975795,2.727608,3.0520537,2.474842,1.9579924,1.5731846,1.3392819,1.2562841,1.2826926,1.1657411,0.90543,0.62248313,0.38858038,0.18863125,0.12826926,0.09808825,0.08299775,0.08299775,0.094315626,0.18863125,0.26031113,0.32821837,0.38480774,0.41121614,0.38480774,0.39989826,0.43385187,0.44516975,0.392353,0.3470815,0.29426476,0.2678564,0.29049212,0.38103512,0.41498876,0.4979865,0.5017591,0.39989826,0.2678564,0.10186087,0.033953626,0.026408374,0.049044125,0.05281675,0.00754525,0.030181,0.041498873,0.033953626,0.0150905,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.17354076,0.35462674,0.3470815,0.2678564,0.59230214,1.0525624,0.59607476,0.5696664,1.6184561,3.6783094,2.2220762,1.2713746,1.1242423,1.8523588,3.31991,3.108643,3.4066803,2.9086938,1.6184561,0.84129536,0.41498876,0.22258487,0.13204187,0.06790725,0.018863125,0.02263575,0.060362,0.06790725,0.033953626,0.026408374,0.041498873,0.041498873,0.056589376,0.06790725,0.018863125,0.02263575,0.06790725,0.09808825,0.08299775,0.02263575,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.056589376,0.0754525,0.049044125,0.00754525,0.02263575,0.03772625,0.03772625,0.041498873,0.116951376,0.06790725,0.15845025,0.3169005,0.55080324,0.9393836,1.3920987,1.6146835,1.7995421,1.780679,1.0487897,0.98842776,0.9620194,1.1883769,1.9202662,3.440634,4.3347464,4.357382,4.534695,4.8327327,4.1612053,3.3463185,4.979865,8.379,12.491161,15.916705,15.886524,14.25675,11.563096,9.110889,8.956212,6.205968,5.753253,6.983129,8.737399,9.333474,7.0359454,5.462761,4.142342,2.886058,1.7844516,1.9051756,1.9504471,1.9164935,1.991946,2.546522,2.3956168,2.293756,2.8294687,4.002755,5.247721,6.2135134,6.326692,4.8629136,2.7917426,2.7804246,2.4031622,2.04099,1.5845025,1.1883769,1.2902378,1.841041,1.8334957,1.5543215,1.3241913,1.478869,1.4977322,1.2525115,1.20724,1.3845534,1.3770081,1.1317875,1.1921495,1.3053282,1.3015556,1.0940613,0.97710985,1.1355602,1.8259505,2.5993385,2.2711203,2.0372176,2.6144292,3.0105548,3.138824,3.8405323,4.274384,4.640329,4.5460134,4.1197066,4.006528,3.9801195,3.0897799,2.4899325,2.7313805,3.7763977,4.919503,5.281675,4.025391,1.9466745,1.4750963,3.9763467,6.356873,6.2021956,4.055572,3.440634,4.002755,3.4783602,3.138824,3.4594972,4.1197066,3.9273026,4.4177437,4.436607,4.3347464,5.945657,9.261794,8.914713,6.5341864,4.025391,3.5839937,4.881777,7.383027,9.842778,11.076427,9.955957,7.884786,7.0887623,6.205968,5.0138187,4.429062,3.9122121,3.7198083,3.6896272,4.274384,6.541732,8.058327,8.488406,7.326438,5.05909,3.1350515,4.8440504,7.281166,8.850578,8.941121,7.91874,7.3000293,8.718536,10.601076,11.261286,8.922258,7.8432875,9.152389,10.31813,10.359629,9.869187,8.303548,7.956466,7.488661,6.1229706,3.6481283,2.8294687,2.2560298,1.9542197,2.11267,3.097325,3.953711,3.6066296,3.0520537,2.8747404,3.218049,4.1989317,3.6066296,4.0593443,5.1269975,3.3123648,2.5993385,3.6141748,5.2326307,5.987156,4.0593443,2.6634734,3.410453,4.772371,5.621211,5.247721,6.1116524,11.944131,21.719002,29.641514,25.170954,20.643805,24.156118,30.320587,32.814293,24.382475,17.206944,16.022339,16.825907,17.976559,20.209951,24.208935,24.755966,21.97554,17.742655,15.701665,13.0646,14.93205,17.512526,17.95015,14.298248,13.272095,14.505743,14.611377,12.562841,9.65792,7.8998766,7.2887115,6.273875,5.481624,7.7225633,11.053791,9.914458,10.461489,12.838243,11.197151,10.917976,12.702429,16.109108,18.5085,15.07541,5.666483,5.572167,8.13378,9.061845,6.398372,5.2552667,5.511805,7.1378064,9.4127,10.940613,11.465008,11.740409,12.706201,13.287186,10.4049,8.831716,10.272858,9.627739,6.398372,4.6818275,5.093044,6.4474163,7.4282985,7.779153,8.299775,10.069136,13.166461,15.663939,16.120426,13.5663595,13.238141,12.46098,11.208468,9.582467,7.809334,7.3000293,6.8850408,6.3342376,5.4174895,3.904667,2.5880208,2.033445,1.9089483,1.8070874,1.267602,1.6071383,1.2751472,0.94315624,0.8941121,0.995973,0.7922512,0.76207024,0.8601585,0.9620194,0.8601585,0.8262049,0.694163,0.6488915,0.77716076,1.0412445,0.95824677,0.77338815,0.6187105,0.51684964,0.38480774,0.29426476,0.24899325,0.21881226,0.20372175,0.21503963,0.20749438,0.18485862,0.14713238,0.09808825,0.071679875,0.0452715,0.03772625,0.026408374,0.018863125,0.049044125,0.094315626,0.10186087,0.09808825,0.08299775,0.041498873,0.041498873,0.03772625,0.05281675,0.06413463,0.02263575,0.0150905,0.00754525,0.003772625,0.0,0.00754525,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4640329,3.1765501,7.1000805,8.371455,6.25124,3.0860074,0.94315624,0.30181,0.071679875,0.02263575,0.00754525,0.00754525,0.003772625,0.0,0.003772625,0.011317875,0.0150905,0.011317875,0.0,0.00754525,0.011317875,0.011317875,0.011317875,0.030181,0.02263575,0.018863125,0.0150905,0.018863125,0.02263575,0.030181,0.03772625,0.116951376,0.38858038,0.9997456,2.0447628,2.938875,2.8030603,2.1692593,2.9615107,5.511805,7.0170827,7.0812173,5.8664317,4.1197066,3.85185,4.244203,4.2102494,3.6141748,3.2784111,2.6785638,5.081726,5.032682,2.3956168,2.3428001,1.5052774,0.94315624,0.513077,0.21881226,0.23013012,0.30935526,0.40367088,0.47912338,0.60362,0.97333723,2.8181508,3.2255943,4.436607,6.72659,8.443134,6.2663302,3.682082,2.3692086,2.6332922,3.429316,4.52715,5.481624,6.198423,7.141579,9.329701,8.013056,5.4665337,3.338773,2.2183034,1.6637276,1.1619685,0.77338815,0.49044126,0.3169005,0.25276586,0.26408374,0.29426476,0.331991,0.41498876,0.62248313,1.0978339,1.5203679,1.8749946,2.1088974,2.1164427,1.9353566,2.5276587,3.62172,4.640329,4.689373,3.6028569,2.5767028,1.7882242,1.3392819,1.2336484,1.2223305,1.1317875,0.9695646,0.7469798,0.482896,0.30935526,0.21503963,0.16976812,0.1659955,0.20372175,0.41121614,0.422534,0.44894236,0.5394854,0.59607476,0.6187105,0.694163,0.754525,0.7469798,0.6451189,0.52062225,0.39989826,0.34330887,0.38103512,0.48666862,0.4376245,0.4074435,0.38858038,0.3772625,0.35462674,0.18485862,0.05281675,0.06790725,0.07922512,0.033953626,0.0,0.030181,0.060362,0.0452715,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041498873,0.1961765,0.5772116,0.76584285,1.0902886,1.2713746,1.6788181,3.3350005,3.0407357,1.5807298,1.1091517,2.6295197,5.9494295,3.5085413,1.3505998,0.91674787,2.2598023,4.08198,2.505023,2.425798,2.6408374,2.4182527,1.5128226,0.59607476,0.19240387,0.05281675,0.011317875,0.0,0.018863125,0.041498873,0.03772625,0.0150905,0.0452715,0.05281675,0.049044125,0.06413463,0.071679875,0.011317875,0.026408374,0.056589376,0.094315626,0.1056335,0.026408374,0.003772625,0.00754525,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.060362,0.10186087,0.060362,0.030181,0.00754525,0.030181,0.10186087,0.18485862,0.150905,0.3169005,0.43007925,0.5281675,0.9280658,1.448688,1.720317,1.8938577,1.7580433,0.73188925,0.6488915,0.6073926,0.8941121,1.5920477,2.584248,3.7575345,4.8138695,4.749735,4.074435,4.7648253,5.413717,8.937348,13.094781,16.890041,20.557034,20.025093,15.603577,10.891568,7.9338303,7.201941,5.4967146,5.0213637,5.824933,7.201941,7.6923823,5.7683434,4.52715,3.4934506,2.3578906,0.98465514,0.56212115,0.98842776,1.5580941,1.901403,1.9655377,1.9127209,1.9730829,2.335255,3.2067313,4.7912335,5.3684454,5.349582,4.2328854,2.806833,3.1539145,2.8558772,2.052308,1.3317367,1.1242423,1.6863633,1.8259505,1.5882751,1.4335974,1.5203679,1.7165444,1.2638294,1.0827434,1.1732863,1.6071383,2.5238862,2.0258996,1.3732355,1.0148361,1.0336993,1.1695137,1.2902378,1.3204187,1.5580941,1.8485862,1.5958204,1.4826416,2.5276587,3.6443558,4.564876,5.836251,6.375736,5.945657,4.9157305,3.7160356,2.8143783,2.6144292,2.6182017,2.897376,3.308592,3.4934506,2.5314314,2.2183034,1.9429018,1.599593,1.5731846,4.538468,5.583485,4.2328854,2.173032,3.2557755,4.236658,3.8858037,3.6707642,4.055572,4.52715,3.3915899,3.150142,3.5877664,5.13077,8.846806,11.853588,10.336992,7.232122,5.010046,5.692891,6.507778,6.94163,8.001738,9.039209,7.786698,5.80607,5.2137675,5.191132,5.674028,7.3679366,7.3000293,7.069899,6.1342883,5.1647234,6.0550632,7.3905725,7.020855,5.243949,3.1124156,2.4522061,5.05909,7.069899,8.473316,9.0807085,8.518587,7.7376537,8.571404,9.1976595,9.039209,8.737399,6.7869525,7.3377557,7.9413757,7.6923823,7.213259,6.0701537,6.907676,6.7831798,4.961002,2.9464202,2.5917933,2.233394,1.9730829,2.1692593,3.4142256,3.5500402,3.3878171,2.9124665,2.3465726,2.1692593,3.8065786,3.482133,2.3805263,1.4562333,1.4637785,1.4713237,3.0633714,5.43258,6.8359966,4.5799665,2.6031113,2.4559789,3.108643,3.904667,4.564876,6.2851934,11.940358,22.70743,33.31228,32.05977,30.946842,33.410366,36.40583,36.27379,28.732311,24.699375,23.903353,22.7942,20.734346,20.036411,23.250689,23.631723,23.75622,24.242887,23.775084,20.304268,23.171463,25.125683,23.19787,18.715992,16.11288,15.679029,13.792717,10.751981,10.770844,11.0613365,10.140816,7.5263867,5.451443,8.831716,14.883006,13.81158,13.404137,15.286676,14.913187,12.351574,12.917468,18.58395,24.665422,19.84778,9.97482,8.360137,8.91094,9.133525,10.121953,9.929549,10.269085,12.128989,15.516807,19.47429,18.946123,18.742401,17.169216,14.468017,12.804289,14.490653,15.071637,12.811834,8.771353,6.7944975,5.6363015,7.4396167,9.163706,9.495697,8.83926,12.076173,15.271586,17.255987,17.014538,13.679539,15.218769,15.992157,15.509261,13.58145,10.325675,9.397609,9.231613,8.892077,7.7301087,5.406172,3.5651307,3.1916409,3.5085413,3.7348988,3.0897799,3.6368105,2.7691069,1.7052265,1.1883769,1.4826416,1.2713746,1.3166461,1.5165952,1.6486372,1.4147344,1.6033657,1.599593,1.6939086,2.022127,2.5427492,2.2107582,1.9429018,1.6712729,1.3807807,1.0940613,0.694163,0.52439487,0.44894236,0.39989826,0.38480774,0.49044126,0.55080324,0.49044126,0.33953625,0.23767537,0.14335975,0.094315626,0.06413463,0.056589376,0.090543,0.18863125,0.23390275,0.30935526,0.36971724,0.23013012,0.241448,0.271629,0.26031113,0.19240387,0.11317875,0.08299775,0.06790725,0.05281675,0.0452715,0.05281675,0.06413463,0.071679875,0.0754525,0.06790725,0.033953626,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.5885295,2.3956168,4.745962,5.6853456,3.953711,2.3428001,1.146878,0.452715,0.13204187,0.056589376,0.026408374,0.018863125,0.011317875,0.003772625,0.011317875,0.011317875,0.011317875,0.011317875,0.0,0.0,0.00754525,0.0150905,0.018863125,0.026408374,0.026408374,0.018863125,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.041498873,0.090543,0.22258487,0.38858038,0.633801,0.87902164,1.3317367,2.516341,5.9305663,8.409182,8.729855,7.1868505,5.5985756,5.1345425,4.6856003,4.247976,4.0103,4.353609,3.1614597,3.097325,2.5767028,1.8976303,3.2670932,1.4147344,0.51684964,0.19240387,0.14713238,0.150905,0.23390275,0.36971724,0.49044126,0.7507524,1.5580941,3.6896272,3.62172,4.4177437,6.307829,6.700182,6.9491754,5.904158,4.2781568,3.2821836,4.6214657,6.1305156,7.2962565,9.914458,14.407655,19.798737,15.667711,9.291975,4.6290107,2.7879698,2.0070364,1.4373702,0.91674787,0.55457586,0.3470815,0.20372175,0.20749438,0.21881226,0.27540162,0.47535074,0.9695646,1.5354583,1.8599042,2.04099,2.1390784,2.1881225,2.082489,2.7238352,4.044254,5.6551647,6.8359966,5.9532022,4.508287,3.0746894,1.9994912,1.4109617,1.146878,1.0902886,1.1053791,1.0827434,0.9393836,0.6790725,0.49421388,0.38858038,0.35839936,0.38480774,0.60362,0.513077,0.4640329,0.55080324,0.5998474,0.7130261,0.91674787,1.086516,1.1544232,1.0940613,0.87902164,0.67152727,0.55080324,0.5470306,0.6451189,0.6149379,0.5772116,0.573439,0.59607476,0.58475685,0.19994913,0.06413463,0.094315626,0.094315626,0.02263575,0.0,0.011317875,0.08677038,0.08677038,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.211267,0.94315624,2.7011995,2.0787163,1.8863125,3.0897799,6.2399216,11.487643,4.847823,1.9542197,0.8526133,0.77338815,2.0900342,0.9808825,0.39989826,0.8262049,2.1503963,3.6783094,0.965792,0.29803738,0.3470815,0.3772625,0.24522063,0.14713238,0.06790725,0.018863125,0.0,0.0,0.0,0.018863125,0.03772625,0.08299775,0.23013012,0.120724,0.10186087,0.094315626,0.071679875,0.060362,0.03772625,0.02263575,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.018863125,0.041498873,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.09808825,0.24522063,0.1358145,0.041498873,0.10940613,0.27917424,0.3055826,0.392353,0.7582976,0.7469798,0.41498876,0.55080324,0.9016574,1.0450171,0.845068,0.452715,0.3055826,0.27917424,0.7130261,1.3166461,1.7052265,1.388326,1.6939086,3.3727267,4.776143,5.191132,4.8365054,8.243186,14.86037,21.326649,25.253952,25.269043,20.115637,13.426772,8.013056,5.1534057,4.5761943,4.45547,5.5683947,5.824933,5.13077,5.3873086,4.3121104,3.7877154,2.8332415,1.3656902,0.16976812,0.15467763,0.6752999,1.5543215,2.3088465,2.1353056,2.2107582,2.0447628,1.8674494,1.9844007,2.776652,3.410453,3.5990841,3.2444575,2.6521554,2.516341,2.2484846,1.9089483,1.6863633,1.5279131,1.1129243,1.4071891,2.2484846,3.0181,3.218049,2.4710693,1.4335974,1.237421,1.3807807,1.780679,2.7917426,2.595566,1.5580941,1.0525624,1.3392819,1.5731846,1.1431054,0.58098423,0.2263575,0.14335975,0.1056335,0.5583485,3.5274043,5.7909794,6.1908774,5.6287565,6.7643166,5.934339,3.7462165,1.5807298,1.5580941,1.4939595,1.8825399,2.7615614,3.5689032,3.127506,1.1996948,0.7167987,1.418507,2.2673476,1.448688,1.4373702,1.3694628,1.4298248,1.8146327,2.7313805,3.1350515,2.6031113,2.1315331,2.3277097,3.4029078,3.6971724,4.859141,6.432326,8.213005,10.238904,10.616167,7.726336,5.040227,4.6554193,7.277394,6.571913,5.3609,5.66271,6.6360474,4.561104,4.085753,4.214022,4.878004,6.3417826,9.186342,10.650121,11.419736,10.521852,8.409182,6.9567204,7.3377557,7.5490227,7.1793056,6.458734,6.2851934,7.4094353,9.393836,11.548005,12.940104,12.3893,11.608367,12.777881,12.887287,11.117926,8.835487,7.2472124,6.017337,5.1269975,4.61392,4.5761943,3.5877664,1.9051756,0.8563859,0.6752999,0.5055317,0.8941121,1.8976303,2.214531,2.3654358,4.6856003,3.5990841,3.270866,2.867195,2.1088974,1.267602,1.4864142,2.5389767,2.6106565,1.5128226,0.67152727,0.7092535,2.4031622,4.4403796,5.3609,3.5538127,2.6521554,2.5087957,2.1315331,1.720317,2.686109,7.3717093,14.8339615,26.231062,38.771267,45.72799,46.76546,43.958626,43.068287,42.355263,32.57662,28.42673,25.163408,24.925734,27.34776,29.569836,20.88148,12.97783,12.887287,19.146072,21.820864,17.120173,17.071129,14.335975,8.537451,6.2399216,7.5226145,6.19465,6.40969,10.038955,16.693865,18.731083,22.7942,16.592005,5.987156,14.984866,20.88148,17.591751,13.656902,12.947649,14.694374,15.660167,14.535924,13.140053,11.672502,8.729855,12.6345215,11.54046,7.9225125,5.7909794,10.695392,18.18028,14.622695,13.124963,18.02183,24.857826,26.578144,23.48459,17.252214,11.706455,12.815607,11.34051,11.317875,11.819634,11.638548,9.307066,9.382519,9.646602,8.846806,7.605612,8.424272,16.795727,19.074392,17.350302,14.792462,15.611122,18.221779,19.425245,19.01403,16.950403,13.35132,10.9594755,10.005001,9.661693,8.993938,6.94163,5.3080835,4.9723196,6.2889657,7.8961043,6.7152724,6.187105,4.5120597,2.9728284,2.142851,1.8599042,1.4335974,1.3543724,1.50905,1.7542707,1.9391292,3.5236318,4.1310244,4.346064,4.6290107,5.3269467,4.7006907,4.4931965,4.112161,3.4594972,2.897376,1.5920477,1.1016065,0.8941121,0.7130261,0.58098423,1.116697,1.4147344,1.3241913,0.935611,0.58098423,0.35839936,0.20372175,0.124496624,0.116951376,0.150905,0.33576363,0.45648763,0.77338815,1.086516,0.73188925,0.87902164,1.0148361,0.784706,0.331991,0.32067314,0.271629,0.24899325,0.23013012,0.211267,0.19994913,0.26031113,0.29426476,0.31312788,0.29049212,0.1659955,0.094315626,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.056589376,0.18863125,0.362172,0.47157812,0.362172,0.2263575,0.15845025,0.15467763,0.1056335,0.08299775,0.049044125,0.02263575,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.026408374,0.05281675,0.0754525,0.124496624,0.17354076,0.362172,0.6149379,0.62625575,1.1393328,1.5241405,1.8033148,2.2673476,3.4632697,5.342037,5.5004873,4.6554193,3.904667,4.745962,2.3390274,1.237421,1.1581959,1.6071383,1.8787673,1.3392819,0.6451189,0.20749438,0.1056335,0.090543,0.1056335,0.181086,0.26031113,0.3470815,0.52062225,3.5085413,3.863168,3.9612563,4.859141,6.2851934,6.7379084,7.986647,6.741681,4.2328854,6.2097406,8.627994,10.020092,15.475307,24.182526,29.41893,21.55678,10.846297,3.953711,2.2296214,1.7391801,1.3241913,0.83752275,0.482896,0.31312788,0.23013012,0.15467763,0.17354076,0.5093044,1.4222796,3.2029586,4.266839,4.274384,3.4217708,2.3465726,2.1503963,1.871222,2.2748928,3.289729,4.7836885,6.590776,7.54525,6.9755836,5.5495315,3.8141239,2.2258487,1.3958713,0.98842776,0.965792,1.1732863,1.3430545,1.2562841,1.0336993,0.8337501,0.69039035,0.52062225,0.44516975,0.4640329,0.513077,0.56212115,0.6111652,0.7432071,0.91674787,1.1355602,1.3732355,1.5580941,1.4713237,1.1921495,0.90543,0.7167987,0.65643674,0.6073926,0.58475685,0.663982,0.84129536,1.0374719,0.06413463,0.026408374,0.05281675,0.049044125,0.09808825,0.4640329,0.7507524,0.55080324,0.452715,0.49044126,0.14713238,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.011317875,0.094315626,0.73188925,2.7238352,3.6368105,3.5349495,2.7992878,2.41448,3.9725742,1.8523588,0.7582976,0.84129536,2.1164427,4.459243,3.8065786,2.7615614,2.5993385,2.9237845,1.6750455,0.56589377,0.26408374,0.25276586,0.24899325,0.18485862,0.1056335,0.0452715,0.011317875,0.0,0.0,0.0,0.049044125,0.08677038,0.094315626,0.094315626,0.19994913,0.30181,0.2565385,0.10940613,0.09808825,0.071679875,0.041498873,0.02263575,0.026408374,0.06413463,0.011317875,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.32821837,0.18485862,0.02263575,0.0,0.0,0.0,0.00754525,0.011317875,0.02263575,0.060362,0.03772625,0.15845025,0.211267,0.17731337,0.21881226,0.33576363,0.55080324,0.51684964,0.3169005,0.452715,0.6488915,0.8262049,0.7809334,0.66775465,0.9997456,0.41876137,0.52439487,1.2826926,2.425798,3.4255435,3.3123648,3.9348478,4.6290107,4.6629643,3.2255943,7.665974,12.868423,17.784155,20.46649,18.0671,13.743673,9.695646,6.760544,4.9760923,3.5538127,2.6597006,3.470815,4.3121104,4.432834,3.99521,3.7990334,4.0517993,3.1199608,1.177059,0.21503963,1.0035182,1.2864652,1.6561824,2.1692593,2.3201644,3.1048703,3.440634,2.9501927,2.033445,1.8485862,2.082489,2.0296721,1.8485862,1.6712729,1.6260014,1.1619685,0.9393836,0.95824677,1.1016065,1.1242423,1.6524098,1.7354075,1.8787673,1.9240388,1.0299267,0.9205205,0.8639311,0.7507524,0.69039035,1.0110635,1.3128735,0.97710985,0.7922512,0.9507015,1.0450171,0.5319401,0.21503963,0.071679875,0.049044125,0.071679875,1.9768555,5.198677,6.2625575,5.4438977,6.7643166,7.001992,5.3948536,3.3878171,2.5993385,4.8402777,6.587003,5.2364035,3.399135,2.2899833,1.7127718,1.3958713,4.353609,9.371201,12.898605,9.0543,4.2291126,4.1197066,5.511805,6.126743,4.659192,4.3800178,4.1612053,3.6254926,3.0633714,3.4142256,6.1305156,7.745199,7.3377557,5.824933,5.9682927,5.3571277,4.0895257,3.7613072,4.9987283,7.435844,6.319147,6.0739264,7.7187905,9.80128,8.420499,4.183841,3.0860074,3.5990841,4.6516466,5.6098933,6.156924,8.050782,9.567377,9.963503,9.495697,7.454707,7.6320205,8.126234,7.877241,6.700182,6.515323,7.1981683,7.9262853,8.469543,9.178797,9.982366,11.016065,11.812089,12.128989,11.98563,10.710483,8.575176,6.930312,6.349328,6.6662283,6.1531515,3.9310753,1.8372684,0.814887,0.91674787,1.1921495,1.3920987,1.4977322,1.8334957,3.059599,2.6597006,2.0636258,1.5958204,1.3656902,1.2525115,1.8636768,1.9768555,1.5731846,0.9997456,0.9393836,0.5470306,1.2034674,2.203213,2.8407867,2.4182527,2.335255,2.0975795,1.5845025,1.2902378,2.3428001,7.960239,17.569115,29.913143,41.75164,47.878384,40.997116,35.345722,32.0824,29.939552,25.227543,26.321604,23.816582,25.744392,33.995125,44.29062,41.36306,30.320587,20.455173,16.177015,17.022083,24.989868,30.158363,27.328896,18.678267,13.747445,19.1008,21.23988,19.108345,14.43029,11.6875925,23.601542,18.983849,10.657665,7.7225633,15.558306,19.538425,19.127209,17.942604,17.655886,18.014284,18.316093,20.175999,18.65563,14.2944765,13.109872,14.690601,12.366665,10.133271,10.680302,15.369675,14.418973,10.34831,10.257768,14.626467,17.312576,16.15438,16.06761,14.984866,12.366665,9.193887,8.778898,9.699419,9.442881,8.062099,8.171506,11.321648,10.963248,11.472552,14.019074,16.565596,15.641303,17.33144,18.523588,18.417955,18.500954,20.138271,23.016785,23.831673,21.998177,19.636513,16.026112,15.086727,15.143317,14.713238,12.494934,10.733118,8.710991,7.745199,8.028146,8.631766,8.360137,7.462252,6.0324273,4.6214657,4.2404304,3.832987,3.3651814,3.31991,3.6669915,3.8292143,4.5196047,5.20245,6.6813188,8.578949,9.352338,8.322411,7.224577,6.368191,5.802297,5.3269467,4.266839,3.470815,2.886058,2.6219745,2.9351022,2.9766011,2.8785129,2.7615614,2.6144292,2.3013012,1.9542197,1.1016065,0.4640329,0.27540162,0.26408374,0.3169005,1.0638802,1.720317,1.9957186,2.11267,2.2484846,2.2447119,1.9957186,1.6033657,1.3468271,0.995973,0.7582976,0.573439,0.422534,0.331991,0.3169005,0.3734899,0.47157812,0.5470306,0.5357128,0.44139713,0.36594462,0.30181,0.25276586,0.23013012,0.19240387,0.094315626,0.041498873,0.0452715,0.03772625,0.018863125,0.003772625,0.0,0.0,0.0,0.07922512,0.27917424,0.392353,0.3734899,0.35839936,0.35839936,0.35085413,0.30935526,0.21881226,0.071679875,0.0452715,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.011317875,0.003772625,0.0,0.0,0.003772625,0.011317875,0.030181,0.05281675,0.071679875,0.094315626,0.071679875,0.0452715,0.03772625,0.0452715,0.0452715,0.041498873,0.026408374,0.018863125,0.0150905,0.0150905,0.003772625,0.0,0.003772625,0.011317875,0.011317875,0.011317875,0.0150905,0.011317875,0.003772625,0.0150905,0.026408374,0.018863125,0.011317875,0.003772625,0.003772625,0.003772625,0.011317875,0.026408374,0.0452715,0.05281675,0.060362,0.10940613,0.18485862,0.27917424,0.36971724,0.44139713,0.6451189,0.8224323,1.0751982,1.7429527,2.3918443,2.3390274,2.0673985,1.9202662,2.1088974,2.505023,1.4147344,1.3430545,2.2296214,1.4260522,1.8825399,1.1996948,0.44139713,0.09808825,0.06790725,0.060362,0.07922512,0.10186087,0.13204187,0.2263575,1.3317367,1.9542197,2.354118,2.7653341,3.380272,4.466788,7.0472636,9.122208,10.393582,12.253486,13.536179,15.196134,19.410156,25.110592,27.95515,17.086218,7.7602897,2.584248,1.3543724,1.0789708,0.7922512,0.52062225,0.32067314,0.211267,0.15467763,0.181086,0.7582976,2.5276587,5.353355,8.307321,8.469543,7.0887623,4.8138695,2.4823873,1.1280149,0.8639311,1.0110635,1.690136,2.8332415,4.1989317,5.3948536,6.1116524,6.168242,5.7079816,5.2062225,3.983892,2.535204,1.448688,0.9620194,0.9280658,0.98842776,0.90543,0.76207024,0.633801,0.58098423,0.58475685,0.5998474,0.60362,0.60362,0.633801,0.72811663,0.8262049,1.0487897,1.4147344,1.81086,1.8825399,1.9881734,2.0485353,2.04099,1.9994912,1.9693103,1.7542707,1.5505489,1.4147344,1.2562841,0.120724,0.0452715,0.033953626,0.03772625,0.150905,0.6451189,0.62625575,0.44516975,0.41876137,0.48666862,0.18485862,0.05281675,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.018863125,0.030181,0.060362,0.0,0.011317875,0.003772625,0.2565385,1.1921495,3.380272,4.7120085,3.99521,2.463524,1.3204187,1.7165444,0.62248313,0.19994913,0.6187105,2.1277604,5.0515447,4.285702,3.218049,3.0181,3.0256453,0.76207024,0.32444575,0.18485862,0.16976812,0.16222288,0.11317875,0.060362,0.056589376,0.056589376,0.049044125,0.056589376,0.011317875,0.060362,0.094315626,0.08299775,0.071679875,0.63002837,0.98465514,0.7469798,0.18485862,0.20749438,0.2263575,0.181086,0.09808825,0.026408374,0.041498873,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.16976812,0.094315626,0.011317875,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.00754525,0.00754525,0.09808825,0.13958712,0.14335975,0.27917424,0.32821837,0.6073926,0.94692886,1.1808317,1.1581959,0.8941121,0.7054809,0.52062225,0.4678055,0.845068,0.6451189,0.5772116,0.965792,1.7957695,2.7011995,2.8558772,3.640583,4.538468,4.52715,2.071171,6.428553,10.929295,13.687083,13.754991,11.148107,9.378746,7.809334,6.458734,5.0854983,3.1954134,2.1541688,2.505023,3.2859564,3.9273026,4.2328854,4.5196047,4.644101,3.9159849,2.4899325,1.3468271,2.5767028,2.3390274,2.0673985,2.082489,1.5958204,2.2296214,2.8936033,2.8181508,2.0636258,1.5354583,1.9542197,1.8599042,1.6712729,1.5618668,1.4600059,0.91674787,0.7432071,0.84129536,1.1016065,1.4034165,1.4034165,1.0827434,1.0299267,1.1846043,0.83752275,0.67152727,0.56212115,0.47912338,0.49421388,0.76584285,1.2223305,1.0336993,0.7922512,0.73188925,0.7130261,0.49044126,0.241448,0.12826926,0.24899325,0.6375736,2.7917426,4.5120597,4.4705606,3.5236318,4.696918,5.3759904,4.4177437,3.2218218,3.0181,4.8629136,5.2250857,3.572676,2.8219235,3.4330888,3.399135,1.4562333,3.3840446,7.835742,11.348056,8.36391,3.7763977,5.1269975,7.515069,7.5112963,3.1652324,2.8521044,3.097325,3.5764484,4.2027044,5.119452,5.9494295,6.2851934,5.7909794,4.640329,3.5424948,3.2444575,2.7313805,2.746471,3.5236318,4.768598,4.496969,5.0062733,6.673774,8.518587,8.201687,5.7872066,4.5988297,3.7575345,3.0407357,2.848332,2.9652832,4.2592936,5.7079816,6.72659,7.175533,7.183078,7.4396167,7.5792036,7.115171,5.43258,5.0515447,5.7117543,6.5832305,7.432071,8.597813,8.635539,9.258021,10.329447,11.517824,12.294985,10.86516,8.786444,6.8925858,5.670255,5.27413,4.7572803,3.2029586,1.5618668,0.543258,0.6187105,0.79602385,0.94692886,1.0638802,1.3166461,2.052308,2.5578396,2.142851,1.6976813,1.5316857,1.3694628,1.4109617,1.3845534,1.2298758,0.95447415,0.60362,0.55080324,1.0751982,1.3996439,1.3091009,1.146878,1.2562841,1.116697,0.8563859,0.84129536,1.6825907,6.300284,16.233604,28.65686,39.129665,41.615826,30.275316,24.861599,24.148573,25.61235,25.404858,26.491373,23.635496,24.427748,30.592216,37.98656,43.34369,38.854263,31.105293,23.941078,18.459454,23.352549,27.094994,25.186045,18.746174,14.524607,20.06282,19.953413,17.36162,15.675257,18.493408,25.065321,19.447882,15.098045,17.40312,23.65813,21.002203,21.179516,21.986858,22.137764,21.27006,21.304014,22.82438,21.78691,18.293459,16.558052,14.973549,14.188843,13.072145,12.6345215,16.026112,15.301767,12.955194,12.442118,14.679284,18.018057,16.392056,14.977322,14.369928,13.943622,11.819634,10.265312,10.457717,10.042727,9.567377,12.494934,12.434572,12.67602,14.584969,17.84829,20.46649,17.916197,19.296976,21.790682,23.605314,23.978804,23.356321,23.676994,23.145054,21.488873,19.972277,17.87847,17.120173,16.667458,16.592005,18.059555,20.673985,17.595524,14.147344,12.981603,14.0983,12.857106,11.299012,10.076681,9.193887,8.013056,7.352846,6.651138,6.8774953,8.103599,9.484379,10.884023,11.902632,13.490907,15.181043,15.113135,13.340002,12.038446,11.551778,11.947904,13.019329,12.702429,11.691365,10.499215,9.382519,8.360137,7.194396,6.379509,5.7570257,5.194905,4.5912848,4.327201,3.350091,2.2786655,1.5203679,1.2600567,1.5128226,2.3088465,2.9615107,3.3010468,3.663219,3.983892,4.2592936,4.504514,4.557331,4.055572,3.4217708,2.9351022,2.4710693,2.0598533,1.8863125,1.7089992,1.6637276,1.6410918,1.5543215,1.3317367,1.0789708,0.87902164,0.84129536,0.91297525,0.875249,0.7394345,0.62625575,0.6451189,0.7130261,0.56589377,0.32444575,0.21503963,0.2678564,0.44894236,0.66775465,0.91297525,1.1695137,1.2449663,1.1091517,0.9016574,0.6526641,0.47535074,0.35085413,0.24899325,0.15467763,0.120724,0.08677038,0.06790725,0.060362,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.033953626,0.056589376,0.06413463,0.041498873,0.049044125,0.041498873,0.030181,0.0150905,0.00754525,0.00754525,0.011317875,0.011317875,0.00754525,0.00754525,0.00754525,0.003772625,0.02263575,0.0452715,0.02263575,0.02263575,0.011317875,0.011317875,0.0150905,0.00754525,0.0,0.0,0.003772625,0.00754525,0.0150905,0.0150905,0.0150905,0.011317875,0.011317875,0.0150905,0.018863125,0.018863125,0.011317875,0.00754525,0.0,0.00754525,0.011317875,0.018863125,0.030181,0.03772625,0.10940613,0.1358145,0.13204187,0.13958712,0.20372175,0.21881226,0.30935526,0.43385187,0.7922512,1.8334957,1.3845534,4.0782075,4.395108,2.0560806,2.0447628,1.8599042,1.0902886,0.8865669,1.1921495,0.7167987,0.97710985,0.72811663,0.45648763,0.33953625,0.24522063,0.17354076,0.14713238,0.116951376,0.090543,0.1358145,0.36594462,0.69793564,0.9922004,1.8485862,4.5761943,3.6707642,5.6363015,8.631766,11.555551,14.037937,16.188334,18.21046,21.09652,23.518545,21.839725,11.959221,5.0741806,1.6146835,0.7997965,0.63002837,0.47157812,0.32821837,0.21881226,0.14335975,0.10940613,0.43007925,2.3918443,4.719554,7.149124,10.423763,9.857869,7.3679366,4.587512,2.3578906,0.724344,0.47535074,0.4376245,0.70170826,1.2713746,2.0900342,3.1425967,4.002755,4.6327834,5.2099953,6.1418333,6.217286,5.5457587,4.2894745,2.8521044,1.8485862,1.418507,1.1355602,0.90920264,0.7167987,0.60362,0.6375736,0.663982,0.7205714,0.8186596,0.9507015,1.0751982,1.1280149,1.2147852,1.3807807,1.6109109,1.7655885,1.961765,2.0749438,2.082489,2.0673985,2.0975795,1.9655377,1.8184053,1.6939086,1.5580941,0.10940613,0.03772625,0.10186087,0.23013012,0.5583485,1.4373702,0.845068,0.38858038,0.23767537,0.2867195,0.13958712,0.05281675,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.094315626,0.00754525,0.03772625,0.026408374,0.094315626,0.181086,0.049044125,0.13204187,0.543258,1.0789708,2.1315331,4.7120085,5.583485,3.9574835,2.2220762,1.478869,1.5241405,0.39989826,0.20372175,0.8941121,2.4597516,4.9232755,3.8254418,2.7992878,2.655928,2.6521554,0.47535074,0.23390275,0.14335975,0.116951376,0.094315626,0.05281675,0.060362,0.06790725,0.06413463,0.056589376,0.071679875,0.0150905,0.0754525,0.15845025,0.241448,0.392353,0.935611,1.1996948,0.84884065,0.19240387,0.18485862,0.26031113,0.26408374,0.19240387,0.09808825,0.071679875,0.090543,0.041498873,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.003772625,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.00754525,0.02263575,0.0452715,0.10186087,0.2565385,0.241448,0.66020936,1.2713746,1.6637276,1.2638294,0.79602385,0.55457586,0.44894236,0.5017591,0.8563859,0.83752275,0.633801,0.6111652,0.90920264,1.448688,1.8221779,3.2557755,4.376245,4.183841,2.0598533,5.100589,8.428044,10.054046,9.374973,7.1679873,6.741681,6.0550632,5.3910813,4.6818275,3.4896781,2.4522061,2.3956168,3.0105548,3.8782585,4.5007415,4.847823,5.0251365,4.504514,3.4029078,2.493705,3.5462675,2.8407867,2.1692593,1.9466745,1.1921495,1.4713237,2.0560806,2.252257,1.9051756,1.4147344,1.7240896,1.7316349,1.8033148,2.0183544,2.142851,1.3694628,1.0336993,1.1921495,1.6373192,1.8787673,1.3053282,0.8262049,0.724344,0.88279426,0.8111144,0.55080324,0.55080324,0.59607476,0.6375736,0.77338815,1.0374719,0.9242931,0.7507524,0.67152727,0.69039035,0.56212115,0.331991,0.271629,0.5394854,1.2110126,2.5012503,2.7351532,2.3314822,1.9579924,2.5314314,3.5764484,3.4594972,2.8143783,2.3692086,2.9426475,2.5238862,1.6410918,1.9504471,3.2821836,3.6330378,1.5807298,2.1202152,4.406426,6.349328,4.640329,2.6634734,4.847823,7.1264887,7.0359454,3.7273536,4.025391,4.5460134,4.878004,5.194905,6.270103,5.3646727,5.100589,5.149633,4.9232755,3.5689032,2.8898308,2.686109,2.6597006,2.6710186,2.71629,3.1199608,4.115934,5.4476705,6.63982,6.971811,6.541732,5.7192993,4.6629643,3.7198083,3.440634,3.5575855,3.8858037,4.357382,4.8440504,5.1835866,6.296511,6.5832305,6.647365,6.2399216,4.2291126,3.8254418,4.349837,6.092789,8.68081,11.087745,9.665465,8.401636,8.537451,9.865415,10.759526,9.039209,7.062354,5.6551647,5.0213637,4.7120085,3.4217708,2.1051247,1.0638802,0.5017591,0.5017591,0.56589377,0.724344,0.814887,0.90920264,1.3015556,2.0372176,1.871222,1.5430037,1.3392819,1.1204696,0.8601585,0.97333723,1.0035182,0.7582976,0.3055826,0.5093044,0.90920264,0.9242931,0.55457586,0.3772625,0.43385187,0.3772625,0.331991,0.47535074,1.0638802,4.346064,13.845533,26.215971,35.877663,35.059006,21.68505,16.094019,17.384256,22.322622,25.32186,25.850027,23.533634,22.473528,24.122164,27.268534,34.72324,37.043404,35.12691,29.569836,20.68153,22.960196,26.378195,26.02734,20.63626,12.555296,14.392565,12.872196,12.015811,14.392565,21.088974,20.274086,16.984358,17.757746,23.246916,28.245644,24.657877,25.431265,27.476028,28.819082,28.611588,28.015512,26.729048,23.854307,20.040184,17.512526,15.347038,14.818871,13.728582,12.717519,15.301767,16.365646,15.62244,15.290449,16.459963,19.08571,18.202915,17.101309,16.70141,16.471281,14.43029,13.973803,13.607859,14.109617,15.863888,18.866898,14.211478,13.664448,15.614895,18.757492,22.054766,21.447372,22.115128,23.322369,24.7786,26.638506,26.219744,25.042685,23.914669,23.069601,22.183035,22.356575,21.87368,21.4851,22.258488,25.574625,28.377686,26.302742,22.515026,19.591242,19.53088,16.77309,14.641558,15.124454,16.935314,15.509261,14.498198,13.532406,14.898096,18.255732,20.628714,22.167944,23.420456,24.620152,25.072866,23.160145,20.43631,19.500698,19.346022,19.68933,20.975796,21.119154,20.583443,19.957186,19.15739,17.421982,15.154634,13.479589,12.117672,10.895341,9.7296,9.016574,8.096053,7.0284004,5.9305663,4.98741,4.67051,4.908185,5.1760416,5.300538,5.4665337,5.515578,5.87775,6.6058664,7.360391,7.405663,6.752999,6.1116524,5.492942,4.9723196,4.6818275,4.38379,4.0706625,3.7386713,3.3576362,2.8936033,2.425798,2.0183544,1.8900851,2.0145817,2.1277604,2.3692086,2.5804756,2.6446102,2.5087957,2.1805773,1.7240896,1.4335974,1.3505998,1.4675511,1.7052265,1.9881734,2.1541688,2.082489,1.7957695,1.4373702,0.9620194,0.7167987,0.59607476,0.5093044,0.36971724,0.3734899,0.28294688,0.21881226,0.2263575,0.31312788,0.1961765,0.10940613,0.06413463,0.0452715,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.026408374,0.033953626,0.060362,0.08677038,0.1056335,0.090543,0.15845025,0.14335975,0.11317875,0.09808825,0.071679875,0.033953626,0.0150905,0.00754525,0.011317875,0.0150905,0.011317875,0.00754525,0.03772625,0.0754525,0.026408374,0.02263575,0.0150905,0.0150905,0.011317875,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.00754525,0.0150905,0.018863125,0.02263575,0.018863125,0.00754525,0.018863125,0.018863125,0.0150905,0.02263575,0.041498873,0.13204187,0.13958712,0.116951376,0.10940613,0.13204187,0.14713238,0.1961765,0.27917424,0.573439,1.448688,1.3128735,4.61392,5.0025005,2.2560298,2.2598023,1.3392819,0.845068,0.573439,0.41121614,0.32821837,0.271629,0.29803738,0.43007925,0.59230214,0.63002837,0.47157812,0.35085413,0.23013012,0.14713238,0.1961765,0.20749438,0.38858038,0.95824677,2.1390784,4.1574326,2.4710693,3.199186,5.1081343,7.3377557,9.4013815,11.680047,13.434318,15.079182,15.573396,12.434572,6.405917,2.6597006,0.8903395,0.44516975,0.32821837,0.25276586,0.19240387,0.13958712,0.10186087,0.09808825,1.3732355,4.085753,6.952948,9.514561,12.132762,9.752235,6.2323766,3.5877664,2.282438,1.2110126,0.56212115,0.29049212,0.2565385,0.40367088,0.7469798,1.4335974,2.082489,2.7540162,3.6330378,5.0213637,6.33801,7.2283497,7.194396,6.2399216,4.8402777,3.5990841,2.6710186,1.9391292,1.3505998,0.9280658,0.8186596,0.77716076,0.8526133,1.0035182,1.1280149,1.2298758,1.2864652,1.327964,1.3770081,1.4600059,1.5241405,1.6448646,1.7769064,1.9089483,2.0447628,2.033445,1.931584,1.8334957,1.7580433,1.6373192,0.271629,0.120724,0.36971724,0.76207024,1.2713746,2.0862615,1.2110126,0.43007925,0.0754525,0.094315626,0.060362,0.033953626,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16976812,0.3470815,0.049044125,0.011317875,0.018863125,0.15467763,0.33953625,0.32821837,0.41121614,1.2298758,2.11267,3.1652324,5.2779026,5.3458095,3.3274553,1.841041,1.6184561,1.4826416,0.67152727,0.56212115,1.539231,3.4142256,5.4703064,3.7273536,2.4861598,2.0258996,1.7995421,0.41121614,0.22258487,0.14335975,0.09808825,0.05281675,0.018863125,0.0754525,0.060362,0.026408374,0.018863125,0.041498873,0.00754525,0.120724,0.3055826,0.6526641,1.4109617,1.1317875,0.814887,0.44894236,0.124496624,0.049044125,0.14335975,0.211267,0.2263575,0.1961765,0.14713238,0.14335975,0.06413463,0.0150905,0.018863125,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.018863125,0.00754525,0.003772625,0.011317875,0.026408374,0.0150905,0.003772625,0.0,0.00754525,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.003772625,0.0,0.0,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.05281675,0.0754525,0.0150905,0.003772625,0.0,0.0,0.00754525,0.03772625,0.018863125,0.011317875,0.011317875,0.0452715,0.1659955,0.23013012,0.7092535,1.2487389,1.3958713,0.63002837,0.32821837,0.36594462,0.5583485,0.8526133,1.3166461,0.9695646,0.663982,0.44894236,0.43007925,0.7507524,1.1393328,3.0709167,4.2291126,3.8103511,2.5012503,3.6707642,5.560849,7.3981175,8.069645,6.092789,5.1458607,3.9914372,3.470815,3.6896272,4.0103,2.9766011,2.7804246,3.3953626,4.3121104,4.5460134,4.7308717,5.089271,4.67051,3.6066296,3.127506,3.3764994,2.444661,1.7693611,1.6825907,1.418507,1.2562841,1.4637785,1.6335466,1.5731846,1.3128735,1.1921495,1.2411937,1.750498,2.546522,2.9916916,2.1805773,1.7127718,1.9391292,2.505023,2.372981,1.5052774,1.0450171,0.845068,0.7432071,0.56212115,0.49421388,0.70170826,0.8111144,0.7092535,0.56589377,0.52439487,0.5583485,0.69039035,0.83752275,0.7997965,0.56589377,0.47535074,0.76584285,1.3958713,2.0447628,1.7089992,1.3694628,1.5505489,2.0975795,2.173032,2.5616124,2.5578396,1.9844007,1.2525115,1.3392819,1.8334957,1.6939086,1.4939595,1.5128226,1.750498,1.841041,2.4484336,3.1576872,3.2972744,1.9391292,2.305074,3.99521,5.3269467,6.0814714,7.5075235,8.865668,8.654402,7.1868505,5.696664,6.326692,5.6061206,5.6853456,5.9607477,5.9003854,5.05909,3.4217708,3.4179983,3.5651307,3.2255943,2.595566,2.8936033,3.7914882,4.708236,5.3080835,5.485397,5.3269467,4.9760923,5.070408,5.6476197,6.1606965,6.541732,6.3342376,6.1041074,5.975838,5.6363015,5.6551647,5.9796104,6.628502,6.7567716,4.647874,3.5877664,3.591539,6.0022464,10.280403,14.007756,11.864905,8.412953,6.8925858,7.6810646,8.280911,6.828451,4.881777,4.002755,4.398881,4.927048,3.059599,1.6184561,0.8941121,0.77338815,0.73188925,0.70170826,0.69039035,0.6451189,0.5998474,0.67152727,0.97710985,0.94315624,0.7696155,0.60362,0.55080324,0.5394854,0.7167987,0.6413463,0.32444575,0.23013012,0.36971724,0.43385187,0.40367088,0.29803738,0.19994913,0.19240387,0.15467763,0.1358145,0.25276586,0.68661773,3.2218218,11.864905,23.676994,32.75393,30.248907,17.278622,10.925522,11.883769,17.621931,22.394302,24.054256,22.926243,20.36463,18.444365,19.987368,23.563816,28.294687,30.750666,28.841719,21.839725,24.152346,29.056757,30.535627,25.114365,11.883769,8.197914,6.8171334,7.7187905,10.499215,14.354838,10.789707,9.9257765,13.355092,19.447882,23.34123,24.650331,26.781864,29.766012,32.984062,35.149548,33.938534,30.026323,24.73333,19.708193,16.931541,16.878725,15.207452,13.257004,12.608112,15.064092,17.123945,17.497435,18.048239,18.489635,16.395828,16.724047,17.991648,19.081938,18.485863,14.302021,17.410664,17.625704,18.810308,21.454918,22.696112,17.77661,15.961976,16.143063,17.82188,21.088974,23.639269,23.511,22.4773,22.673477,26.585688,27.483574,26.71773,26.55928,27.268534,27.110083,28.951124,29.185026,29.626425,31.131702,33.595226,32.7577,32.644524,30.546946,26.71773,24.393793,20.315586,18.259504,20.741892,25.589716,25.95566,25.253952,23.763765,25.461447,29.939552,32.36535,33.863083,35.247635,36.56428,36.76046,33.693314,29.773556,28.86058,28.347504,27.476028,27.332668,27.645796,28.1551,29.007713,29.600016,28.596497,25.850027,23.61286,21.598278,19.598787,17.508753,15.716756,14.713238,14.083209,13.35132,12.004493,10.70671,10.133271,9.740918,9.265567,8.714764,8.035691,7.8696957,8.356364,9.344792,10.378491,10.197406,9.831461,9.416472,9.005256,8.597813,8.156415,7.492433,6.79827,6.149379,5.5193505,4.8742313,4.2894745,3.8178966,3.5689032,3.712263,4.398881,4.9685473,4.9949555,4.5309224,4.06689,3.6443558,3.2369123,2.9237845,2.746471,2.727608,2.8143783,2.7728794,2.5314314,2.1353056,1.7844516,1.3015556,1.0638802,1.0638802,1.1280149,0.875249,0.87902164,0.66775465,0.4979865,0.4979865,0.68661773,0.4979865,0.35085413,0.2565385,0.18485862,0.06413463,0.056589376,0.03772625,0.026408374,0.018863125,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.0452715,0.056589376,0.06790725,0.08677038,0.120724,0.18485862,0.32821837,0.30935526,0.271629,0.25276586,0.211267,0.14335975,0.090543,0.05281675,0.026408374,0.018863125,0.003772625,0.00754525,0.049044125,0.094315626,0.071679875,0.0452715,0.033953626,0.026408374,0.0150905,0.00754525,0.00754525,0.011317875,0.011317875,0.003772625,0.011317875,0.0150905,0.0150905,0.0150905,0.011317875,0.003772625,0.011317875,0.02263575,0.026408374,0.026408374,0.0150905,0.033953626,0.041498873,0.041498873,0.041498873,0.071679875,0.094315626,0.090543,0.09808825,0.120724,0.1358145,0.120724,0.16222288,0.18863125,0.20749438,0.30935526,1.2261031,2.4220252,2.5578396,1.7919968,1.780679,1.1317875,0.8299775,0.66775465,0.5470306,0.482896,0.33953625,0.3470815,0.5017591,0.77716076,1.0940613,0.91674787,0.6451189,0.38480774,0.241448,0.30181,0.38103512,0.62248313,1.539231,2.4182527,1.3166461,0.754525,0.6073926,0.7507524,1.1393328,1.7844516,2.8709676,3.7575345,4.436607,4.5422406,3.3463185,1.9693103,1.1846043,0.7582976,0.47912338,0.1659955,0.11317875,0.08677038,0.0754525,0.0754525,0.11317875,2.2371666,4.8138695,8.269594,11.808316,13.415455,9.0807085,4.9723196,2.7917426,2.4672968,2.1503963,1.0148361,0.42630664,0.19240387,0.15845025,0.211267,0.49044126,0.9318384,1.4298248,2.0070364,2.8181508,4.4101987,6.436098,8.265821,9.280658,8.873214,7.405663,5.8702044,4.485651,3.308592,2.2598023,1.6222287,1.2713746,1.1695137,1.1846043,1.1242423,1.1129243,1.2034674,1.327964,1.4260522,1.4411428,1.3656902,1.388326,1.5618668,1.8561316,2.142851,1.991946,1.8033148,1.7052265,1.6712729,1.5316857,1.358145,0.5998474,0.995973,1.7240896,1.8146327,0.16976812,0.094315626,0.056589376,0.033953626,0.011317875,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.38858038,0.7922512,0.18485862,0.03772625,0.018863125,0.14713238,0.48666862,1.1431054,0.7432071,0.7130261,2.1013522,3.712263,2.1503963,1.9089483,1.2223305,0.73566186,0.69039035,0.94692886,1.177059,0.91674787,1.5618668,3.9688015,8.424272,5.1873593,3.199186,1.5618668,0.27917424,0.23013012,0.15467763,0.12826926,0.09808825,0.056589376,0.030181,0.030181,0.011317875,0.00754525,0.0150905,0.0150905,0.003772625,0.23013012,0.52062225,1.3015556,3.5839937,1.7429527,0.5319401,0.03772625,0.049044125,0.060362,0.03772625,0.041498873,0.10186087,0.16976812,0.120724,0.060362,0.018863125,0.018863125,0.049044125,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.090543,0.030181,0.0150905,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.00754525,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.09808825,0.2678564,0.36971724,0.0754525,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.026408374,0.033953626,0.071679875,0.29049212,0.7432071,1.0638802,1.1619685,0.9620194,0.41121614,0.26408374,0.23767537,0.47157812,0.9997456,1.7693611,1.0978339,0.8224323,0.6790725,0.56589377,0.52062225,1.1431054,2.8898308,4.4177437,4.357382,1.3430545,1.5279131,3.31991,5.7079816,7.066127,5.1873593,3.4783602,2.4672968,2.233394,2.7653341,3.9386206,3.0709167,3.2029586,4.025391,5.0213637,5.462761,5.7079816,5.1647234,4.719554,4.3724723,3.2482302,2.2975287,1.4826416,1.1053791,1.2223305,1.6637276,0.55080324,0.5319401,0.9393836,1.3015556,1.3128735,1.2525115,0.9242931,1.418507,2.4786146,2.5012503,2.795515,2.867195,3.0633714,3.2029586,2.5804756,1.6637276,1.3505998,0.91674787,0.35462674,0.36594462,0.52439487,0.5470306,0.4979865,0.45648763,0.5017591,0.5017591,0.5394854,0.9808825,1.3958713,0.58098423,0.63002837,0.9620194,2.2748928,3.983892,4.2404304,2.1315331,2.1503963,3.6481283,5.138315,4.3347464,2.565385,1.3241913,0.8111144,1.327964,3.2821836,4.719554,3.470815,1.931584,1.1883769,0.9922004,2.1881225,3.8254418,4.636556,4.2328854,3.097325,2.987919,3.5085413,4.376245,6.3719635,11.351829,13.841762,10.574668,6.930312,5.583485,6.485142,6.937857,6.4436436,5.956975,5.7570257,5.462761,4.496969,4.8138695,4.927048,4.3385186,3.5689032,3.2029586,2.8747404,2.8822856,2.9464202,2.214531,2.2598023,2.4371157,3.187868,4.52715,6.0286546,6.651138,6.549277,6.719045,7.2962565,7.5527954,7.2094865,7.8395147,8.986393,9.6051035,8.039464,5.040227,4.9760923,6.8473144,9.5032425,11.627231,10.725573,8.29223,6.217286,5.3873086,5.692891,6.092789,4.8025517,2.8521044,1.3505998,1.4939595,1.4826416,1.3430545,1.1242423,0.8903395,0.73188925,0.7809334,0.65643674,0.44894236,0.2678564,0.24522063,0.40367088,0.3772625,0.2867195,0.22258487,0.26031113,0.392353,0.34330887,0.211267,0.094315626,0.1056335,0.21503963,0.21503963,0.20372175,0.19994913,0.150905,0.1659955,0.1659955,0.150905,0.211267,0.56589377,3.2255943,10.182315,19.451654,26.283878,23.133736,14.0983,9.544742,9.714509,13.664448,19.255478,23.503454,21.73032,17.527617,14.298248,15.214996,18.119919,20.960705,24.17121,26.234835,23.695858,16.848543,18.746174,21.93027,21.809546,16.633503,9.733373,4.889322,2.8822856,3.2105038,4.0895257,2.625747,2.1315331,3.5047686,6.1531515,7.997965,9.865415,13.343775,17.889788,22.748928,26.94786,26.642279,24.718239,22.892288,21.266287,18.312323,19.859098,19.413929,16.965494,14.588741,16.418465,21.058792,23.69963,23.620405,19.53088,9.582467,11.329193,11.830952,14.400109,17.003222,12.253486,17.429527,19.47429,17.99542,15.663939,18.202915,23.880716,24.74842,21.884998,17.546478,15.165953,21.477554,21.794455,21.805773,24.352295,29.41893,26.280106,24.254206,24.940825,27.502436,28.626678,30.799711,32.95388,33.88572,34.398796,37.292397,38.378914,37.57157,36.6171,35.25518,31.20338,26.834682,25.110592,26.04243,29.554745,35.477764,37.099995,34.549698,32.014496,31.5731,33.17269,37.431984,39.1938,42.45335,46.6221,46.52401,40.982025,38.031834,36.077614,34.45161,33.40282,34.327114,35.61358,36.88873,37.850746,38.254417,35.896526,34.108303,31.886227,28.849264,25.238861,22.269806,20.817345,20.730574,21.368149,21.575642,20.69662,19.791191,18.734856,17.41821,15.746937,14.50197,12.955194,11.581959,11.000975,11.978085,12.966512,13.864397,14.219024,13.996439,13.58145,12.725064,11.796998,10.963248,10.231359,9.476834,8.778898,8.258276,7.122716,5.59103,4.881777,4.7120085,4.8138695,4.768598,4.447925,4.044254,4.115934,3.9989824,3.7952607,3.5575855,3.2670932,2.9124665,2.6295197,2.2899833,1.931584,1.7844516,1.6146835,1.1581959,1.3241913,1.961765,1.8749946,1.6448646,1.3015556,1.0110635,0.8337501,0.7469798,0.6375736,0.65643674,0.6187105,0.47912338,0.32067314,0.28294688,0.19240387,0.1056335,0.05281675,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.0452715,0.094315626,0.07922512,0.07922512,0.15845025,0.36594462,0.5017591,0.52439487,0.5017591,0.4678055,0.44139713,0.392353,0.3169005,0.2263575,0.12826926,0.030181,0.00754525,0.00754525,0.041498873,0.09808825,0.18485862,0.09808825,0.049044125,0.030181,0.030181,0.030181,0.030181,0.02263575,0.0150905,0.011317875,0.0,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.003772625,0.00754525,0.0150905,0.0150905,0.0150905,0.06413463,0.13204187,0.14335975,0.10940613,0.120724,0.071679875,0.071679875,0.08299775,0.10940613,0.18485862,0.2678564,0.24522063,0.17731337,0.124496624,0.1358145,0.23390275,0.5885295,1.0223814,1.2713746,0.97710985,0.694163,0.73566186,0.875249,0.995973,1.0676528,0.69039035,0.66775465,0.77338815,0.9620194,1.388326,1.4260522,0.98465514,0.5470306,0.32821837,0.29049212,0.33953625,0.2867195,0.23390275,0.20372175,0.16976812,0.14335975,0.1358145,0.13204187,0.150905,0.26031113,0.41876137,0.59607476,0.76584285,0.7922512,0.42630664,1.5015048,2.1088974,2.071171,1.388326,0.23013012,0.094315626,0.041498873,0.030181,0.05281675,0.1358145,0.9922004,3.4859054,6.8435416,10.008774,11.657412,8.397863,5.0477724,3.2784111,3.006782,2.3956168,1.7354075,0.8224323,0.241448,0.11317875,0.0754525,0.10186087,0.29049212,0.6375736,1.0827434,1.50905,2.293756,3.6783094,5.9984736,8.8618965,11.170743,11.536687,10.484125,9.114662,7.7037,5.6778007,3.8065786,2.6898816,2.0183544,1.5882751,1.297783,1.0902886,1.2034674,1.3845534,1.4411428,1.2223305,1.2940104,1.358145,1.4449154,1.5430037,1.6184561,1.3619176,1.1959221,1.2562841,1.4826416,1.6184561,0.392353,0.14335975,0.19994913,0.34330887,0.362172,0.033953626,0.018863125,0.011317875,0.00754525,0.003772625,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06790725,0.27540162,0.44516975,0.14713238,0.030181,0.20749438,0.6111652,0.91297525,0.5470306,0.32821837,0.33953625,0.8601585,1.5354583,1.358145,1.0374719,2.1503963,2.7011995,2.2107582,1.7165444,1.3920987,2.7691069,3.7273536,3.85185,4.432834,3.5500402,2.082489,0.8262049,0.26408374,0.5470306,0.55080324,0.2867195,0.08677038,0.049044125,0.041498873,0.02263575,0.071679875,0.18863125,0.30935526,0.30935526,0.150905,0.11317875,0.13958712,0.36971724,1.1091517,0.42630664,0.12826926,0.060362,0.1056335,0.1961765,0.150905,0.08299775,0.0754525,0.11317875,0.08677038,0.033953626,0.02263575,0.018863125,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.00754525,0.0150905,0.018863125,0.00754525,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.011317875,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.00754525,0.0,0.0,0.0,0.003772625,0.0150905,0.011317875,0.003772625,0.00754525,0.011317875,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.06413463,0.16976812,0.241448,0.124496624,0.0754525,0.08299775,0.06790725,0.018863125,0.0,0.0,0.003772625,0.011317875,0.08677038,0.3734899,1.0336993,1.4524606,1.750498,1.961765,2.0485353,1.5580941,1.0601076,0.77338815,1.0336993,2.282438,1.7467253,1.1317875,0.90920264,1.2525115,2.0447628,2.3654358,3.150142,4.1536603,4.304565,1.7089992,1.4034165,3.2369123,5.409944,6.2663302,4.3083377,4.425289,4.395108,3.640583,2.6597006,3.0218725,3.187868,4.217795,4.640329,4.315883,4.4139714,4.715781,4.429062,4.4139714,4.3800178,2.897376,1.3204187,1.6675003,1.6260014,0.8639311,1.0299267,0.9808825,1.358145,1.4977322,1.3920987,1.6675003,1.5845025,1.086516,1.0487897,1.4637785,1.4411428,1.6373192,1.9768555,2.1579416,2.1164427,2.04099,1.5052774,1.6863633,1.3845534,0.55080324,0.27917424,0.32067314,0.6073926,1.0450171,1.388326,1.2223305,0.7469798,0.59607476,1.3807807,2.4295704,1.7769064,0.7394345,0.5394854,0.814887,1.177059,1.177059,0.72811663,1.7429527,3.6368105,4.9949555,3.5651307,1.4826416,0.7582976,0.80356914,1.3543724,2.4861598,2.7087448,1.9504471,1.2751472,1.146878,1.4298248,1.629774,1.8184053,1.7957695,1.6712729,1.8636768,2.8596497,3.2972744,3.6556737,4.7421894,7.7037,8.152642,6.115425,4.142342,3.4481792,3.92353,3.8443048,3.289729,2.6898816,2.4899325,3.1425967,3.7613072,4.5196047,4.919503,4.768598,4.1574326,4.104616,3.8820312,3.9801195,4.217795,3.7499893,3.9273026,3.6971724,3.078462,2.4899325,2.7313805,4.0480266,5.4174895,6.6322746,7.073672,5.7117543,5.0741806,5.6098933,6.730363,7.914967,8.677037,8.846806,8.688355,8.858124,9.442881,9.955957,9.665465,8.382772,6.417235,4.666737,4.640329,5.523123,5.1345425,4.142342,3.3123648,3.5085413,2.5012503,1.8787673,1.5505489,1.4411428,1.478869,1.0072908,0.66020936,0.44139713,0.32444575,0.23013012,0.35085413,0.3169005,0.24899325,0.27917424,0.5394854,0.6451189,0.83752275,1.5543215,2.3201644,1.7542707,0.56589377,0.17354076,0.11317875,0.14713238,0.26408374,0.392353,0.2565385,0.14335975,0.422534,1.5279131,4.727099,8.733627,14.4114275,19.293203,17.591751,11.378237,8.122461,7.2170315,8.458225,12.019584,14.392565,13.324911,11.314102,10.646348,13.419228,15.573396,18.49718,21.541689,22.862108,19.425245,14.675511,13.000465,12.468526,11.815862,10.469034,6.296511,3.3764994,2.0749438,1.9278114,1.6222287,1.9655377,2.3126192,2.3993895,2.3654358,2.7351532,3.783943,5.3344917,8.443134,12.540206,15.448899,17.946377,19.195116,18.632996,17.836971,20.557034,18.542452,17.191853,16.203424,15.690348,16.173243,19.074392,19.57615,18.904623,18.61036,20.557034,15.124454,15.573396,17.708702,18.440592,15.792209,13.487134,14.169979,17.369165,21.45869,23.646814,18.991394,19.610106,21.639776,21.605824,16.42601,14.396337,17.63325,23.560043,27.238352,21.38701,26.725275,30.02255,30.241362,28.287142,27.038403,31.271288,35.41363,38.51473,40.589672,42.600483,50.3985,55.0011,55.529266,52.08109,45.754395,41.06125,36.021023,34.56479,37.330124,41.627144,46.25993,47.15404,44.320797,39.699333,37.175446,36.95286,39.75592,44.43398,49.330845,52.262173,52.46967,49.960873,45.71667,41.64978,40.589672,41.038616,41.48001,42.58162,43.89072,43.845448,39.389977,37.258446,35.45513,32.904835,29.44911,27.547709,26.174473,25.529354,25.729303,26.838455,27.657114,28.185282,28.332415,27.69484,25.574625,23.107328,20.304268,17.780382,16.0827,15.652621,15.497944,15.596032,15.992157,16.497688,16.716501,16.995676,16.437326,15.660167,14.966003,14.347293,13.4644985,12.510024,10.751981,8.627994,7.7150183,6.888813,6.198423,5.6287565,5.138315,4.678055,4.508287,4.349837,4.112161,3.7348988,3.180323,2.6974268,2.335255,2.0070364,1.7089992,1.4939595,1.3996439,1.3392819,1.4034165,1.5543215,1.5958204,1.6373192,1.750498,1.7165444,1.5430037,1.4675511,1.3392819,1.3241913,1.4260522,1.5128226,1.297783,0.84884065,0.5696664,0.41498876,0.33953625,0.28294688,0.5772116,0.35462674,0.1961765,0.271629,0.32821837,0.23013012,0.21503963,0.30935526,0.4376245,0.41121614,0.31312788,0.28294688,0.36594462,0.5357128,0.6828451,0.70170826,0.68661773,0.7469798,0.87147635,0.95447415,0.965792,0.7696155,0.6375736,0.59230214,0.44516975,0.26408374,0.15467763,0.10940613,0.13204187,0.2565385,0.2867195,0.1961765,0.090543,0.030181,0.030181,0.030181,0.02263575,0.0150905,0.0452715,0.16976812,0.271629,0.15845025,0.049044125,0.06790725,0.22258487,0.08299775,0.03772625,0.02263575,0.026408374,0.06413463,0.55080324,0.88279426,0.7130261,0.23013012,0.1358145,0.08677038,0.06790725,0.0754525,0.25276586,0.8903395,1.3392819,1.1544232,0.69793564,0.29049212,0.22258487,0.25276586,0.6111652,1.0186088,1.3317367,1.539231,1.1695137,1.1129243,1.0978339,1.0299267,0.995973,0.94692886,1.2147852,1.4147344,1.4335974,1.3996439,1.0072908,0.8111144,0.7092535,0.6526641,0.6451189,0.5357128,0.4376245,0.32067314,0.1961765,0.120724,0.0754525,0.056589376,0.0452715,0.0452715,0.0754525,0.10940613,0.1659955,0.482896,0.935611,1.0374719,0.694163,0.56212115,0.68661773,0.88279426,0.72811663,0.22258487,0.06413463,0.03772625,0.041498873,0.0754525,0.32444575,1.1732863,2.372981,3.5538127,4.236658,3.289729,2.372981,2.071171,2.1503963,1.5279131,0.8224323,0.41876137,0.1961765,0.07922512,0.05281675,0.0452715,0.09808825,0.241448,0.4979865,0.875249,1.3241913,2.123988,3.4368613,5.300538,7.61693,9.495697,10.374719,10.948157,11.404645,11.449917,10.948157,8.907167,6.3153744,4.044254,2.8332415,2.1088974,1.5958204,1.3128735,1.1921495,1.0487897,0.995973,1.0148361,1.0148361,0.9695646,0.8978847,0.8639311,0.8224323,0.79602385,0.7884786,0.7884786,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.12826926,0.2263575,0.2263575,0.071679875,0.0150905,0.22258487,0.58475685,1.0751982,1.780679,3.7386713,3.0256453,1.6561824,0.9507015,1.5165952,2.3767538,3.0520537,3.0143273,2.3767538,1.8900851,2.2598023,3.8895764,4.115934,2.8256962,2.425798,2.1843498,1.3204187,1.2562841,1.7354075,0.83752275,1.1242423,1.4034165,1.0487897,0.271629,0.14713238,1.0978339,1.8900851,2.0598533,1.841041,2.1956677,1.4335974,0.58475685,0.094315626,0.05281675,0.1961765,0.0452715,0.03772625,0.0754525,0.15845025,0.35839936,0.6073926,0.35085413,0.116951376,0.09808825,0.13958712,0.1659955,0.090543,0.026408374,0.00754525,0.0,0.02263575,0.049044125,0.03772625,0.003772625,0.026408374,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.0150905,0.0,0.0,0.00754525,0.00754525,0.0150905,0.018863125,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.030181,0.026408374,0.011317875,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.003772625,0.003772625,0.0,0.0,0.00754525,0.00754525,0.041498873,0.041498873,0.011317875,0.0150905,0.0150905,0.011317875,0.00754525,0.00754525,0.00754525,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0452715,0.18485862,0.47535074,0.7167987,0.331991,0.12826926,0.25276586,0.211267,0.2565385,0.31312788,0.44516975,0.5394854,0.30181,0.11317875,0.12826926,0.17354076,0.18863125,0.24899325,0.7884786,1.3053282,1.7467253,2.052308,2.173032,2.757789,2.1956677,1.388326,1.0299267,1.6146835,1.9693103,1.6750455,1.4034165,1.4864142,1.9240388,2.3503454,2.727608,3.1765501,3.2444575,1.9089483,2.4786146,2.9011486,3.4066803,3.663219,2.7728794,4.7346444,5.5759397,4.557331,2.8558772,3.5424948,3.1124156,3.6896272,4.217795,4.429062,4.8365054,4.6327834,4.4630156,4.636556,4.4215164,2.0485353,1.1657411,2.2673476,2.3654358,1.3091009,1.7957695,2.2786655,2.282438,1.8674494,1.388326,1.478869,1.5203679,1.1280149,0.87902164,0.9242931,0.9922004,1.4637785,1.9844007,2.2484846,2.2484846,2.3013012,2.052308,1.6825907,1.1808317,0.70170826,0.58098423,0.65643674,1.0299267,1.2940104,1.2487389,0.88279426,0.6149379,0.47912338,0.9620194,1.7316349,1.6373192,0.73188925,0.44139713,0.40367088,0.5093044,0.91674787,1.9466745,2.5578396,2.7917426,2.565385,1.6524098,0.62625575,0.392353,1.2185578,2.4295704,2.3880715,1.6976813,1.5618668,1.6750455,1.8259505,1.9089483,2.1277604,2.9992368,3.863168,3.9763467,2.4710693,3.3161373,4.4139714,5.8702044,7.1340337,7.001992,5.715527,4.640329,4.146115,4.044254,3.5839937,2.7389257,2.2371666,2.2673476,2.7540162,3.350091,3.7763977,4.191386,4.659192,4.919503,4.3686996,3.5047686,3.059599,3.1576872,3.5387223,3.5689032,4.3083377,4.715781,4.719554,4.4516973,4.2328854,4.636556,5.2779026,6.375736,7.4207535,7.1793056,6.8473144,6.541732,6.3342376,6.3455553,6.7643166,7.2472124,7.115171,6.7643166,6.4021444,6.047518,6.1418333,6.1531515,5.515578,4.406426,3.7462165,4.168751,3.802806,3.169005,2.757789,3.0143273,2.5276587,1.9579924,1.6071383,1.5316857,1.5354583,1.1280149,0.8111144,0.6073926,0.5055317,0.48666862,0.6375736,0.66775465,0.58475685,0.48666862,0.5470306,0.452715,0.5055317,0.90543,1.388326,1.2147852,0.5055317,0.17731337,0.071679875,0.1056335,0.24522063,0.3734899,0.2678564,0.29426476,0.935611,2.7879698,6.851087,9.424017,11.61214,13.015556,11.710228,8.371455,5.904158,4.5912848,4.696918,6.4738245,8.544995,8.926031,7.8319697,6.7567716,8.439363,9.480607,10.668983,12.683565,14.483108,13.302276,10.412445,8.243186,6.8661776,5.983383,4.927048,2.9728284,1.8976303,1.448688,1.3091009,1.1091517,1.6373192,1.9391292,2.3126192,2.7502437,2.957738,3.5123138,5.7381625,8.771353,11.487643,12.498707,15.509261,15.169725,14.588741,15.184815,16.716501,19.938324,23.05074,24.503199,25.140774,28.215462,23.1526,19.040438,17.105082,17.927513,21.4436,16.588232,14.222796,13.698401,13.615403,11.834724,13.358865,15.445127,17.429527,19.681786,23.62795,19.149845,21.847271,23.661903,21.122927,15.347038,13.966258,21.752956,29.467974,30.071594,18.776354,24.050484,26.959179,28.294687,28.517273,27.747658,32.199356,36.469967,39.09194,39.601246,38.548683,44.1963,52.66207,55.84617,52.91861,50.326817,55.065235,54.276756,52.14522,51.83964,55.49909,58.34742,58.60396,54.420116,47.25213,41.849728,45.01119,47.014454,48.768723,51.43597,56.434696,59.222668,60.07528,60.45254,60.169598,57.392944,55.2765,54.65779,54.171124,52.424397,47.98779,44.13594,41.928955,39.989826,37.435757,33.881947,32.0824,31.456148,31.218472,31.41842,32.931244,35.16464,36.2172,36.28888,35.406086,33.41414,30.780848,27.66466,24.646559,22.22076,20.772074,20.002459,19.595015,19.534653,19.753464,20.138271,20.458946,20.081682,19.440336,18.844261,18.493408,18.033148,16.856089,14.690601,12.057309,10.272858,9.208978,8.360137,7.7716074,7.4207535,7.2094865,7.0510364,6.651138,6.115425,5.462761,4.640329,3.8367596,3.2972744,2.9049213,2.595566,2.335255,2.1956677,2.161714,2.173032,2.1994405,2.2220762,2.2711203,2.384299,2.41448,2.354118,2.323937,2.2484846,2.1956677,2.1654868,2.082489,1.8146327,1.418507,1.1242423,0.90543,0.7432071,0.6149379,0.7696155,0.77716076,0.8111144,0.9620194,1.2261031,1.3166461,1.3770081,1.4562333,1.5618668,1.6561824,1.9127209,2.0070364,2.0447628,2.0900342,2.173032,2.1692593,2.093807,2.1805773,2.4182527,2.565385,2.4069347,2.0145817,1.6410918,1.3355093,0.935611,0.76584285,0.68661773,0.6451189,0.6149379,0.60362,0.7469798,0.66775465,0.45648763,0.2263575,0.120724,0.10186087,0.10186087,0.17731337,0.30935526,0.41498876,0.52062225,0.41498876,0.35085413,0.3772625,0.33953625,0.094315626,0.026408374,0.018863125,0.026408374,0.06790725,0.3734899,0.58098423,0.47535074,0.16976812,0.10186087,0.08677038,0.08677038,0.1056335,0.23013012,0.6488915,1.1921495,1.2902378,1.0412445,0.6451189,0.392353,0.32067314,0.47912338,0.6451189,0.7997965,1.1280149,1.6109109,1.841041,1.5920477,1.146878,1.297783,1.2751472,1.297783,1.2864652,1.2185578,1.1280149,0.965792,0.97710985,0.9997456,1.0035182,1.0601076,0.95824677,0.8337501,0.6187105,0.35839936,0.20749438,0.11317875,0.060362,0.030181,0.0150905,0.011317875,0.011317875,0.030181,0.17731337,0.41498876,0.5394854,0.29803738,0.14713238,0.181086,0.34330887,0.44139713,0.181086,0.211267,0.19240387,0.06413463,0.041498873,0.124496624,0.3772625,0.694163,0.9808825,1.1280149,0.9507015,0.80734175,0.83752275,0.90920264,0.6149379,0.34330887,0.331991,0.271629,0.10940613,0.06413463,0.0452715,0.041498873,0.08299775,0.19240387,0.4074435,0.8526133,1.478869,2.2560298,3.270866,4.7233267,6.2361493,7.360391,8.314865,9.246704,10.246449,12.468526,12.83447,11.487643,9.0807085,6.760544,4.927048,3.2633207,2.093807,1.4411428,1.026154,0.8903395,0.76584285,0.6790725,0.6187105,0.55080324,0.55457586,0.58098423,0.5696664,0.5093044,0.44139713,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.094315626,0.13204187,0.1056335,0.08677038,0.1358145,0.2867195,0.58475685,1.4335974,3.5839937,5.1571784,3.5953116,1.6410918,0.875249,1.7429527,2.704972,2.6785638,2.3578906,2.1466236,2.1579416,2.6408374,3.399135,3.2331395,2.2296214,1.7542707,1.780679,1.5165952,1.8221779,2.2560298,1.0940613,1.7655885,2.3277097,2.5540671,2.293756,1.4411428,2.5917933,3.3651814,2.9351022,1.8636768,2.1013522,1.4034165,0.5772116,0.094315626,0.018863125,0.02263575,0.12826926,0.9922004,1.0412445,0.29049212,0.32067314,0.7167987,0.48666862,0.21503963,0.14713238,0.16976812,0.20372175,0.12826926,0.049044125,0.02263575,0.02263575,0.0452715,0.08299775,0.0754525,0.030181,0.056589376,0.02263575,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.011317875,0.05281675,0.05281675,0.026408374,0.003772625,0.003772625,0.02263575,0.03772625,0.041498873,0.033953626,0.018863125,0.0150905,0.00754525,0.011317875,0.011317875,0.011317875,0.026408374,0.041498873,0.0452715,0.030181,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.003772625,0.003772625,0.003772625,0.00754525,0.0150905,0.0150905,0.05281675,0.05281675,0.0150905,0.0150905,0.026408374,0.026408374,0.02263575,0.011317875,0.0150905,0.02263575,0.011317875,0.003772625,0.003772625,0.0,0.003772625,0.00754525,0.0754525,0.27917424,0.663982,0.83752275,0.35462674,0.06790725,0.211267,0.362172,0.45648763,0.5055317,0.6149379,0.7130261,0.5093044,0.663982,1.0525624,1.026154,0.6073926,0.482896,0.80734175,1.2185578,1.4977322,1.5656394,1.4901869,2.5276587,2.2447119,1.4901869,0.87147635,0.7582976,1.4034165,1.5015048,1.388326,1.2751472,1.2713746,1.9466745,2.6068838,2.9313297,2.806833,2.3126192,2.9803739,2.6295197,2.493705,2.7653341,2.5880208,4.4743333,5.624984,5.0477724,3.62172,4.074435,3.5236318,3.1954134,3.6028569,4.6026025,5.409944,4.9647746,4.564876,4.429062,3.893349,1.4071891,1.1204696,2.5389767,2.8181508,1.8938577,2.4672968,2.7351532,2.3993895,1.7919968,1.2600567,1.1695137,1.1996948,0.9507015,0.754525,0.8111144,1.20724,2.0145817,2.3805263,2.41448,2.3126192,2.3805263,2.0862615,1.5279131,1.146878,1.0978339,1.2449663,1.0902886,1.1996948,1.146878,0.8601585,0.5998474,0.59607476,0.49421388,0.58098423,0.8337501,0.9205205,0.52062225,0.38858038,0.44894236,0.7432071,1.4600059,2.4823873,2.3163917,1.5580941,0.76584285,0.5017591,0.47535074,0.98842776,2.6823363,4.244203,2.4031622,1.3355093,1.3505998,1.720317,2.1579416,2.7879698,3.8103511,5.2175403,6.013564,5.4476705,3.0256453,3.519859,4.749735,6.5040054,7.6810646,6.273875,4.8666863,4.4403796,4.3686996,4.1083884,3.218049,2.263575,2.1353056,2.7917426,3.7198083,3.9122121,3.470815,3.3689542,3.6896272,4.1083884,3.9084394,3.138824,2.7917426,2.9464202,3.429316,3.7990334,5.1760416,5.9494295,6.138061,5.904158,5.5268955,5.3080835,5.1873593,6.1041074,7.696155,8.311093,7.858378,7.986647,7.6207023,6.7454534,6.387054,6.379509,5.8890676,5.0854983,4.2027044,3.5387223,3.5123138,3.783943,3.8971217,3.640583,3.0709167,2.8030603,2.214531,1.6939086,1.4901869,1.7089992,1.7278622,1.3845534,1.1129243,1.0450171,1.0223814,0.8299775,0.663982,0.59230214,0.6149379,0.663982,0.7884786,0.814887,0.69039035,0.47912338,0.362172,0.2263575,0.18485862,0.271629,0.43385187,0.5017591,0.36971724,0.17731337,0.06413463,0.08677038,0.20749438,0.362172,0.3961256,0.7394345,2.0485353,5.221313,8.646856,9.691874,9.480607,8.661947,7.3868,5.7117543,4.025391,3.0369632,2.9916916,3.6594462,4.949684,5.907931,5.3684454,3.8858037,3.7160356,3.7952607,3.7990334,4.7346444,6.3417826,7.0887623,6.3719635,5.3986263,4.7308717,4.3649273,3.7160356,3.180323,2.9841464,2.727608,2.3201644,1.9806281,1.8297231,2.04099,2.5691576,3.1916409,3.500996,3.783943,5.7381625,8.59404,11.16697,11.872451,14.102073,12.1101265,11.336739,13.015556,14.169979,18.16519,23.48459,26.879953,28.679495,32.746384,27.977787,23.718493,21.734093,22.069857,23.005466,20.093,15.856343,14.464244,15.388537,13.389046,11.438599,13.619176,16.180788,17.89356,20.051502,19.395065,22.307531,22.371666,18.02183,12.513797,13.853079,23.186554,30.135729,29.260479,20.085455,19.104572,20.059048,22.039675,24.250433,26.016022,29.32084,31.656096,33.006695,33.474503,33.278324,33.991352,40.89903,45.603493,46.43724,48.45937,57.00059,59.93569,61.056164,63.20656,68.284515,70.333046,68.70705,62.825523,54.431435,47.584118,51.16434,51.503876,51.232246,53.009155,59.539566,62.37281,63.93845,66.764145,69.638885,67.61298,65.903984,66.32275,65.96435,62.817978,55.751854,52.03959,49.75338,47.75766,45.11682,41.095203,39.46166,38.593952,37.963924,37.91111,39.62765,41.99686,43.109787,42.95888,41.755413,39.944553,37.145267,34.051712,31.071339,28.64177,27.223263,26.94786,26.44233,25.763256,25.084183,24.695602,24.8201,25.216225,25.204908,24.480564,23.118647,22.797974,21.417192,19.379974,17.108854,15.067864,13.792717,12.853333,12.438345,12.438345,12.468526,11.989402,10.910432,9.793735,8.801534,7.7187905,6.6624556,5.775889,5.1458607,4.7535076,4.4516973,4.2404304,4.0970707,4.032936,4.002755,3.942393,3.8858037,3.8556228,3.8254418,3.783943,3.7273536,3.6594462,3.5349495,3.3538637,3.108643,2.8030603,2.4559789,2.1013522,1.7580433,1.4901869,1.3807807,1.9278114,2.7502437,3.7499893,4.817642,5.828706,5.8588867,5.6778007,5.3873086,5.081726,4.8365054,4.617693,4.38379,4.172523,4.014073,3.9310753,3.7047176,3.4029078,3.2444575,3.3048196,3.531177,3.4972234,3.2029586,2.7313805,2.2560298,2.0183544,1.9429018,1.9881734,1.7014539,1.1317875,0.8299775,1.1431054,1.4411428,1.3468271,0.90543,0.56589377,0.36594462,0.29049212,0.33953625,0.46026024,0.52062225,0.5583485,0.55457586,0.58098423,0.5885295,0.392353,0.1056335,0.026408374,0.02263575,0.030181,0.049044125,0.120724,0.19994913,0.19994913,0.124496624,0.08677038,0.090543,0.094315626,0.10940613,0.1659955,0.31312788,0.7922512,1.1506506,1.2110126,0.98465514,0.6828451,0.46026024,0.36971724,0.331991,0.3772625,0.6526641,1.4260522,1.690136,1.4637785,1.1808317,1.6863633,1.841041,1.5505489,1.237421,1.1280149,1.2638294,1.3732355,1.327964,1.2449663,1.267602,1.5505489,1.6146835,1.2600567,0.8526133,0.56589377,0.38480774,0.20749438,0.10940613,0.05281675,0.02263575,0.011317875,0.003772625,0.003772625,0.011317875,0.026408374,0.06413463,0.10186087,0.07922512,0.049044125,0.041498873,0.1056335,0.094315626,0.29803738,0.362172,0.21503963,0.041498873,0.08677038,0.21881226,0.41876137,0.55457586,0.362172,0.211267,0.15845025,0.21503963,0.392353,0.7205714,0.58475685,0.965792,0.9318384,0.41498876,0.19994913,0.18485862,0.17731337,0.150905,0.116951376,0.1358145,0.5093044,1.1619685,1.8334957,2.474842,3.240685,3.942393,4.5724216,5.1760416,5.847569,6.719045,9.318384,11.385782,12.004493,11.144334,9.654147,8.024373,5.9984736,4.2027044,2.8332415,1.6712729,1.20724,0.845068,0.63002837,0.5470306,0.48666862,0.43007925,0.4074435,0.3772625,0.32821837,0.271629,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.003772625,0.02263575,0.08299775,0.19994913,0.49044126,0.58098423,0.76207024,1.7127718,4.4931965,3.2218218,1.4524606,0.55457586,0.86770374,1.6939086,1.5618668,1.4713237,1.7580433,2.4031622,3.0633714,2.5201135,1.9202662,1.8863125,2.1692593,1.6675003,2.082489,2.1503963,1.9089483,1.5279131,1.3091009,2.2183034,2.5804756,3.4896781,4.4177437,3.218049,3.663219,3.410453,2.0975795,0.43385187,0.1659955,0.124496624,0.07922512,0.094315626,0.19994913,0.4074435,1.5165952,2.7011995,2.1654868,0.392353,0.15845025,0.41498876,0.41498876,0.33576363,0.2565385,0.1659955,0.124496624,0.09808825,0.06413463,0.033953626,0.056589376,0.056589376,0.07922512,0.08299775,0.06413463,0.0754525,0.041498873,0.030181,0.018863125,0.00754525,0.0,0.02263575,0.030181,0.0452715,0.071679875,0.120724,0.06413463,0.03772625,0.03772625,0.056589376,0.10186087,0.10940613,0.094315626,0.06413463,0.030181,0.018863125,0.02263575,0.05281675,0.049044125,0.02263575,0.041498873,0.049044125,0.03772625,0.018863125,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.011317875,0.011317875,0.011317875,0.018863125,0.0150905,0.0150905,0.02263575,0.026408374,0.018863125,0.0150905,0.033953626,0.041498873,0.03772625,0.026408374,0.0150905,0.0150905,0.00754525,0.003772625,0.011317875,0.0,0.011317875,0.049044125,0.120724,0.22258487,0.38103512,0.241448,0.08299775,0.0,0.08299775,0.422534,0.5394854,0.573439,0.56212115,0.59230214,0.80734175,1.2789198,1.991946,1.8448136,1.0186088,0.95447415,1.0638802,1.1544232,1.0751982,0.8601585,0.7054809,1.3317367,1.4637785,1.1695137,0.6790725,0.35839936,0.543258,0.7469798,0.8865669,0.91674787,0.8299775,1.7014539,2.8936033,3.3953626,3.0860074,2.6936543,2.4295704,2.354118,2.8143783,3.5349495,3.6179473,3.832987,4.5837393,4.889322,4.5007415,3.904667,4.255521,3.4557245,3.4444065,4.5497856,5.462761,5.119452,4.346064,3.6896272,2.9841464,1.3317367,1.1846043,2.2975287,2.6785638,2.1768045,2.4823873,2.1843498,1.780679,1.3807807,1.0827434,0.9695646,0.8299775,0.663982,0.62248313,0.8563859,1.5241405,2.4107075,2.4861598,2.2183034,1.9994912,2.1277604,1.6976813,1.5807298,1.5920477,1.6448646,1.7655885,1.2261031,0.94692886,0.754525,0.633801,0.724344,0.724344,0.6111652,0.5055317,0.452715,0.38858038,0.43007925,0.5357128,0.73566186,1.056335,1.539231,1.4600059,0.91297525,0.55457586,0.5583485,0.6375736,0.90543,2.04099,4.032936,5.168496,2.0070364,1.1996948,1.0110635,1.3392819,2.1881225,3.663219,5.240176,6.0512905,5.59103,4.1800685,2.9539654,3.0822346,3.5538127,4.244203,4.696918,4.1008434,3.8895764,3.9499383,3.6368105,2.9049213,2.293756,2.0070364,2.4182527,3.169005,3.7462165,3.5160866,2.674791,2.4710693,2.6295197,2.9086938,3.108643,3.5424948,3.772625,3.9612563,4.1574326,4.304565,6.0362,6.888813,6.8359966,6.228604,5.7872066,5.2062225,5.0025005,5.9984736,7.673519,8.186596,7.201941,8.812852,9.710737,8.99771,8.179051,7.635793,6.25124,4.8365054,3.8178966,3.218049,2.727608,2.3163917,2.2069857,2.3503454,2.4559789,1.7316349,1.0902886,0.70170826,0.59607476,0.66775465,0.663982,0.4979865,0.35839936,0.30935526,0.32067314,0.28294688,0.27540162,0.38480774,0.56589377,0.62625575,0.663982,0.6111652,0.45648763,0.2565385,0.150905,0.14335975,0.18485862,0.35462674,0.5394854,0.452715,0.33576363,0.18485862,0.07922512,0.0754525,0.1961765,0.44139713,0.65643674,1.3694628,3.3048196,7.375482,9.118435,8.695901,7.5716586,6.439871,5.2137675,3.832987,2.9124665,2.565385,2.6672459,2.8709676,2.7540162,3.1840954,3.150142,2.323937,1.0374719,0.6073926,0.58475685,0.875249,1.4675511,2.4522061,3.519859,4.006528,4.38379,4.9044123,5.594803,5.6400743,5.6778007,5.2892203,4.4101987,3.31991,2.4295704,2.6219745,2.7087448,2.4861598,2.7087448,2.886058,3.097325,4.825187,7.6395655,9.201432,10.299266,9.14107,8.718536,10.370946,13.777626,14.245432,17.05981,19.930779,21.990631,23.7864,26.495146,25.751938,25.287905,25.627441,24.061802,23.099783,20.142044,20.270313,22.956423,22.035902,10.457717,9.454198,13.389046,16.995676,15.380992,17.80679,18.48209,17.01831,13.600313,8.967529,11.004747,17.701157,22.654613,23.48459,21.805773,14.305794,14.332202,15.565851,16.603323,20.95316,22.522572,22.266033,22.873425,25.087955,27.721249,24.910643,26.989359,31.524054,36.756687,41.615826,46.20334,50.02501,56.114025,64.41757,71.79683,75.727905,73.87554,68.44674,61.618282,55.570766,54.91433,53.15629,51.9,53.111015,59.090626,61.391926,60.992027,62.278492,65.41732,66.36047,67.94498,71.38561,73.4681,72.4344,67.97138,63.91204,60.973164,58.875587,56.68746,52.80166,51.89623,50.096687,48.13115,47.086132,48.41787,49.69679,50.417362,50.02501,48.557457,46.678688,43.453094,40.401043,37.99788,36.541645,36.1757,36.658596,36.08516,34.79115,33.21042,31.897545,32.30876,33.761223,34.598743,33.78763,30.924208,29.686787,28.26828,27.32135,26.64605,25.186045,23.348776,21.62846,20.621168,20.277859,19.87796,18.791445,16.923996,15.226315,13.966258,12.73261,11.593277,10.336992,9.2844305,8.52236,7.8961043,7.54525,7.2472124,7.0246277,6.851087,6.6662283,6.458734,6.300284,6.145606,5.983383,5.8136153,5.66271,5.455216,5.2099953,4.930821,4.61392,4.2328854,4.036709,4.093298,4.4101987,4.9534564,6.2399216,7.537705,9.152389,10.940613,12.321393,11.989402,11.385782,10.608622,9.688101,8.59404,7.2962565,6.417235,5.873977,5.541986,5.2854476,4.708236,4.1536603,3.6669915,3.429316,3.7462165,4.1612053,4.1762958,3.802806,3.4557245,3.9612563,4.014073,3.7877154,2.8332415,1.4977322,0.935611,1.4524606,2.305074,2.5691576,2.093807,1.478869,1.0487897,0.7167987,0.5470306,0.5319401,0.573439,0.48666862,0.543258,0.60362,0.5696664,0.36971724,0.150905,0.0754525,0.05281675,0.049044125,0.0452715,0.071679875,0.17731337,0.21881226,0.16976812,0.11317875,0.10186087,0.08677038,0.08299775,0.10940613,0.19994913,0.5696664,0.98465514,1.2110126,1.1846043,0.9922004,0.65643674,0.362172,0.23013012,0.28294688,0.44516975,0.72811663,0.76207024,0.7582976,0.9620194,1.6524098,2.161714,1.9579924,1.5731846,1.4373702,1.8976303,2.1051247,1.7014539,1.3128735,1.3128735,1.8334957,2.0862615,1.4826416,0.91674787,0.7054809,0.543258,0.30181,0.16222288,0.08677038,0.05281675,0.03772625,0.011317875,0.003772625,0.003772625,0.003772625,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0150905,0.041498873,0.23390275,0.4074435,0.40367088,0.08299775,0.06413463,0.17354076,0.482896,0.7582976,0.4640329,0.30935526,0.26408374,0.3055826,0.573439,1.3543724,1.086516,1.7165444,1.750498,0.98842776,0.51684964,0.47535074,0.46026024,0.34330887,0.14335975,0.0452715,0.1961765,0.80356914,1.539231,2.2673476,3.0218725,3.3425457,3.470815,3.6179473,3.832987,3.983892,4.5120597,6.0739264,7.594294,8.612903,9.273112,9.250477,8.084735,6.470052,4.7535076,2.9501927,2.0258996,1.3468271,0.91674787,0.68661773,0.543258,0.41876137,0.29049212,0.19994913,0.15467763,0.13958712,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.0452715,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.02263575,0.0150905,0.071679875,0.18485862,0.32067314,1.1393328,1.2600567,0.9016574,0.91674787,2.806833,1.0487897,0.55457586,0.72811663,1.1431054,1.5731846,1.2525115,1.5882751,2.595566,3.953711,5.0062733,3.0256453,1.599593,1.1959221,1.4826416,1.3128735,1.8749946,1.5845025,1.327964,1.3958713,1.478869,2.0787163,2.384299,2.0372176,1.6825907,2.9766011,3.2935016,1.9429018,0.7922512,0.4376245,0.23013012,0.20372175,0.1358145,0.27917424,0.8111144,1.7995421,6.3644185,3.8443048,0.91674787,0.1961765,0.24522063,0.2565385,0.34330887,0.40367088,0.3734899,0.23013012,0.1056335,0.041498873,0.0150905,0.018863125,0.030181,0.030181,0.049044125,0.060362,0.06413463,0.0754525,0.10186087,0.08677038,0.06413463,0.03772625,0.0,0.10940613,0.120724,0.18485862,0.27917424,0.1659955,0.08299775,0.07922512,0.14713238,0.23390275,0.26031113,0.26031113,0.20372175,0.120724,0.041498873,0.030181,0.056589376,0.16222288,0.150905,0.026408374,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.026408374,0.0150905,0.0150905,0.02263575,0.03772625,0.041498873,0.0150905,0.0150905,0.02263575,0.02263575,0.0150905,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.19240387,0.26408374,0.150905,0.0150905,0.003772625,0.0,0.0,0.00754525,0.030181,0.32444575,0.543258,0.7507524,1.1242423,1.9542197,0.8563859,0.72811663,0.66020936,0.5017591,0.87147635,0.724344,0.45648763,0.29426476,0.32821837,0.5357128,1.4260522,1.7769064,1.4600059,0.8224323,0.70170826,0.7394345,0.6187105,0.7092535,0.97710985,0.97710985,1.8674494,2.8143783,3.0709167,2.6332922,2.2447119,1.6448646,1.6335466,1.8900851,2.4220252,3.5689032,3.1199608,2.9049213,3.5538127,4.3083377,3.0520537,4.3083377,4.3196554,4.2064767,4.4630156,4.9760923,4.436607,3.7462165,3.1765501,2.674791,1.8297231,2.0749438,1.9240388,1.8297231,1.9579924,2.2107582,1.991946,1.4713237,1.1091517,1.0186088,0.94692886,0.6790725,0.58475685,0.5394854,0.56212115,0.7922512,1.1732863,1.448688,1.7014539,1.9579924,2.2107582,2.2598023,2.372981,2.2748928,1.8523588,1.1431054,0.72811663,0.5696664,0.52062225,0.56589377,0.80734175,0.56589377,0.44894236,0.422534,0.5093044,0.77716076,1.1808317,1.4750963,1.418507,1.0374719,0.6111652,0.4640329,0.392353,0.56589377,0.9318384,1.1732863,1.1996948,1.7731338,2.3390274,2.252257,0.76207024,0.77338815,0.91674787,1.7995421,3.0633714,3.3576362,3.440634,2.7879698,2.1202152,2.0372176,2.9916916,2.0636258,1.4298248,0.95824677,0.6488915,0.6111652,1.0148361,1.7165444,2.1881225,2.233394,2.0145817,2.4786146,3.1161883,3.0897799,2.3692086,1.7089992,2.1353056,2.8030603,3.180323,3.1350515,2.916239,4.0480266,5.0213637,4.8855495,3.731126,2.6710186,4.146115,6.0626082,7.779153,8.714764,8.360137,5.7607985,5.406172,6.2663302,7.541477,8.650629,7.7225633,9.4127,11.00852,11.046246,9.337247,7.654656,5.0439997,3.5236318,3.350091,3.0218725,2.323937,1.6373192,1.3505998,1.4562333,1.5430037,0.79602385,0.4640329,0.40367088,0.4376245,0.35085413,0.27917424,0.17731337,0.1056335,0.0754525,0.0754525,0.124496624,0.23013012,0.32067314,0.38103512,0.44139713,0.47912338,0.36971724,0.24899325,0.17731337,0.150905,0.150905,0.30935526,0.5394854,0.73188925,0.73188925,0.452715,0.24522063,0.10940613,0.071679875,0.18485862,0.5357128,0.87147635,1.8259505,3.4934506,5.4476705,7.2283497,7.3377557,6.598321,5.553304,4.45547,2.9803739,2.2899833,1.9655377,1.7731338,1.6637276,1.2713746,1.1921495,1.3505998,1.3656902,0.55080324,0.15845025,0.08677038,0.30935526,0.6790725,0.9620194,1.4750963,2.214531,2.8558772,3.4330888,4.349837,4.38379,5.5193505,6.1418333,5.5306683,3.8443048,3.0030096,2.6634734,2.4823873,2.354118,2.425798,2.6823363,2.1503963,1.5845025,1.4637785,1.9994912,2.463524,5.040227,5.836251,5.621211,9.857869,16.120426,14.452927,11.815862,10.714255,9.186342,9.895596,7.7942433,9.216523,13.196642,11.476325,16.13929,18.327412,19.519562,21.805773,27.906107,21.4851,14.169979,10.574668,11.242422,12.6345215,15.47908,14.524607,11.68382,8.514814,6.19465,5.6476197,7.798016,10.604849,13.698401,18.387774,13.660675,14.796235,14.124708,11.747954,15.535669,15.814844,15.354584,16.524097,18.161417,15.55076,12.974057,15.150862,19.017803,23.43932,29.177483,33.229282,38.563774,44.686745,51.326565,58.441734,64.568474,67.137634,68.62028,69.40121,67.778984,65.715355,61.320248,55.167095,49.776012,49.606247,54.076805,54.559704,55.76694,58.585094,60.07528,62.57653,68.50333,73.40396,76.61447,81.25102,79.470345,74.411255,71.30261,70.978165,69.85393,70.21987,69.03904,66.26238,63.199013,62.531258,62.57653,62.03327,60.516678,58.23801,55.966892,52.575302,49.59493,48.43296,49.07808,50.077824,49.3233,47.83311,45.91662,44.24912,43.883175,45.652534,47.05595,47.995335,47.980244,46.109024,42.264717,41.423424,43.064514,45.180958,44.26421,41.189518,37.00568,33.074604,29.962187,27.434528,26.140518,24.28816,22.586706,21.300241,20.26277,19.11589,17.840744,16.263786,14.441608,12.6345215,11.902632,11.32542,10.834979,10.401127,10.008774,9.6201935,9.303293,9.020347,8.744945,8.439363,8.182823,7.914967,7.635793,7.3377557,7.0170827,6.8246784,7.7716074,9.952185,12.925014,15.731846,16.758,16.207197,15.4074,14.800008,13.947394,13.347548,12.830698,12.174261,11.072655,9.156161,7.9338303,6.9982195,6.3455553,5.956975,5.798525,5.1647234,4.749735,4.4630156,4.38379,4.7610526,5.455216,5.455216,5.149633,5.243949,6.7454534,6.952948,5.119452,3.078462,1.7882242,1.3128735,1.9579924,2.8634224,3.5047686,3.5424948,2.8219235,2.4823873,1.6260014,1.0299267,0.91674787,0.97710985,0.73188925,0.55080324,0.47157812,0.41876137,0.19994913,0.23390275,0.19994913,0.124496624,0.071679875,0.1056335,0.19240387,0.4074435,0.44139713,0.271629,0.1358145,0.124496624,0.11317875,0.094315626,0.0754525,0.0754525,0.41876137,0.7582976,1.0450171,1.1883769,1.0525624,0.88279426,0.4640329,0.21881226,0.23767537,0.27540162,0.32444575,0.47157812,0.45648763,0.32444575,0.45648763,1.0940613,1.8372684,2.0258996,1.8863125,2.5314314,2.8256962,1.9089483,1.1091517,0.9922004,1.358145,1.5543215,1.2185578,0.87147635,0.69039035,0.52062225,0.33576363,0.18863125,0.10940613,0.08677038,0.060362,0.02263575,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.03772625,0.17731337,0.35085413,0.1659955,0.08299775,0.07922512,0.150905,0.27917424,0.42630664,0.87902164,0.9808825,0.6828451,0.29426476,0.48666862,0.66020936,0.95824677,1.3732355,1.6033657,1.0525624,0.845068,0.7469798,0.47157812,0.094315626,0.0452715,0.071679875,0.241448,0.72811663,1.6410918,3.0218725,3.7047176,3.8480775,3.8593953,3.85185,3.6330378,3.1312788,3.0256453,3.2633207,3.7914882,4.5460134,5.8173876,6.300284,6.0739264,5.3080835,4.255521,3.2444575,2.2484846,1.4260522,0.84884065,0.52062225,0.38480774,0.2678564,0.17731337,0.116951376,0.090543,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.049044125,0.030181,0.02263575,0.16976812,0.4678055,0.7809334,0.31312788,0.5357128,0.88279426,1.0487897,0.965792,1.3732355,2.425798,2.3314822,1.2826926,1.478869,2.9916916,2.4710693,1.3732355,0.7884786,1.448688,1.5316857,1.6788181,2.3126192,2.8332415,1.6373192,1.3166461,1.2487389,1.5618668,1.9127209,1.50905,2.7917426,3.2972744,3.6669915,4.0103,3.9197574,3.3878171,3.3123648,2.4484336,1.4864142,3.0746894,1.5656394,0.90920264,0.56589377,0.3169005,0.26408374,0.49421388,2.0975795,3.8065786,3.9310753,0.35839936,1.3015556,0.90920264,0.44894236,0.3734899,0.3055826,0.18863125,0.23013012,0.29049212,0.29049212,0.20372175,0.10186087,0.0452715,0.033953626,0.041498873,0.041498873,0.041498873,0.05281675,0.06413463,0.0754525,0.0754525,0.10940613,0.071679875,0.060362,0.07922512,0.011317875,0.033953626,0.03772625,0.049044125,0.0754525,0.08299775,0.14335975,0.33953625,0.4640329,0.43385187,0.271629,0.19240387,0.20749438,0.21881226,0.20749438,0.2263575,0.29803738,0.2565385,0.150905,0.0452715,0.0150905,0.0150905,0.0150905,0.018863125,0.026408374,0.026408374,0.03772625,0.033953626,0.026408374,0.026408374,0.026408374,0.026408374,0.030181,0.030181,0.026408374,0.0150905,0.026408374,0.03772625,0.03772625,0.033953626,0.041498873,0.030181,0.030181,0.02263575,0.011317875,0.003772625,0.011317875,0.0150905,0.011317875,0.011317875,0.011317875,0.003772625,0.05281675,0.10186087,0.11317875,0.0754525,0.124496624,0.19240387,0.17354076,0.071679875,0.018863125,0.4678055,0.754525,0.79602385,0.80356914,1.2826926,0.9242931,1.1431054,1.6637276,1.9542197,1.237421,0.69793564,0.4376245,0.5093044,0.76207024,0.8639311,0.6413463,1.1091517,1.4071891,1.3128735,1.2525115,0.8865669,0.7054809,0.76207024,0.9620194,1.0487897,1.8938577,2.5201135,2.1843498,1.2110126,0.98465514,0.845068,1.1996948,1.8749946,2.6483827,3.229367,3.5500402,3.1539145,3.1765501,3.7688525,4.1008434,5.983383,5.938112,5.6589375,5.798525,5.9984736,4.0480266,2.8822856,2.2371666,1.8033148,1.2336484,1.0072908,1.0336993,1.1996948,1.4449154,1.7618159,1.659955,1.2034674,0.84884065,0.73188925,0.69039035,0.6375736,0.8299775,1.1921495,1.4260522,1.0148361,1.3430545,1.6976813,2.0296721,2.2183034,2.0673985,1.9278114,2.0560806,1.9806281,1.5807298,1.0601076,0.6526641,0.47535074,0.4376245,0.46026024,0.47912338,0.5281675,0.44139713,0.392353,0.4376245,0.52062225,0.5357128,0.5772116,0.55080324,0.44516975,0.32821837,0.44516975,0.6828451,0.8563859,0.9242931,0.94315624,0.84884065,0.7884786,0.8526133,1.0601076,1.3355093,2.637065,5.715527,5.798525,2.9501927,2.0636258,2.7841973,2.5502944,1.8259505,1.1431054,1.0978339,0.8563859,1.146878,1.901403,2.4597516,1.5618668,1.7882242,1.8334957,1.7693611,1.6373192,1.4637785,1.6260014,1.7618159,1.7844516,1.7542707,1.9164935,2.8407867,3.5424948,3.8065786,3.4783602,2.4861598,2.305074,2.191895,2.1843498,2.4220252,3.1463692,4.52715,5.481624,6.224831,7.356619,9.861642,7.7225633,7.3490734,7.541477,7.748972,8.088508,6.439871,6.4474163,6.255012,5.1798143,3.7235808,2.7992878,2.161714,2.0447628,2.4786146,3.3010468,2.9766011,1.9353566,1.1846043,1.1016065,1.4298248,0.9695646,0.60362,0.52062225,0.6149379,0.5093044,0.543258,0.38103512,0.26031113,0.2678564,0.34330887,0.34330887,0.392353,0.44894236,0.49044126,0.5017591,0.36594462,0.32821837,0.241448,0.094315626,0.030181,0.049044125,0.094315626,0.18863125,0.3055826,0.35462674,0.181086,0.071679875,0.02263575,0.030181,0.10940613,0.211267,0.34330887,0.68661773,1.3015556,2.1503963,3.561358,4.961002,6.205968,6.964266,6.7152724,4.847823,4.285702,4.666737,5.20245,4.7044635,2.8747404,2.0636258,1.7165444,1.418507,0.9016574,0.55080324,0.32444575,0.2678564,0.34330887,0.39989826,1.9957186,2.6785638,2.5616124,2.2183034,2.6634734,2.8181508,3.0143273,3.9612563,5.1269975,4.7610526,2.7351532,2.323937,2.4031622,2.3692086,2.1202152,1.7995421,1.3807807,1.0336993,1.0450171,1.8297231,2.282438,2.5276587,2.3956168,2.3088465,3.3010468,7.3679366,5.553304,3.5387223,3.2444575,2.8634224,3.3576362,3.3463185,3.821669,4.5007415,3.8443048,5.696664,10.03141,11.981857,10.642575,9.099571,10.321902,9.763554,10.065364,11.940358,14.173752,15.260268,10.884023,7.2358947,6.1078796,4.90064,5.093044,5.753253,6.741681,9.073163,14.93205,13.664448,12.653384,10.397354,7.424526,6.319147,6.0814714,6.802043,8.6732645,11.559323,15.011275,16.576914,16.754227,16.392056,16.218515,16.859861,20.100546,23.488363,26.612097,29.596243,33.089695,38.495865,45.807213,51.715145,55.310455,58.113514,60.305412,59.807423,57.513668,55.25009,55.782032,60.271458,63.22165,65.26264,65.85871,63.297104,64.02145,67.38663,71.159256,74.97337,80.32673,84.86143,89.64134,92.1275,90.618454,84.26913,80.82849,80.232414,78.19143,74.23772,71.721375,69.57475,68.575005,66.662285,62.983974,57.872066,57.819252,59.467888,61.75787,63.489506,63.297104,62.47467,60.712852,59.532024,59.95833,62.512398,66.292564,68.288284,68.19397,66.764145,65.82476,63.512142,60.72417,59.58484,59.852695,58.935947,55.382133,50.941757,47.523758,45.32809,42.85325,39.069305,34.783604,31.093975,28.562544,27.21949,25.56708,24.141027,22.714975,21.1682,19.519562,17.935059,16.531643,15.535669,14.7736,13.660675,13.023102,12.419481,11.883769,11.442371,11.087745,10.812344,10.540714,10.269085,9.989911,9.691874,9.359882,13.015556,18.719765,23.726038,24.484337,21.319103,17.833199,14.818871,12.702429,11.555551,11.785681,11.608367,11.400873,11.0613365,10.020092,9.514561,9.035437,8.560086,8.16396,7.9941926,7.605612,7.3679366,7.515069,8.141325,9.190115,9.205205,8.975075,8.4544525,8.27714,9.759781,9.691874,8.854351,7.5565677,5.956975,4.032936,4.3007927,4.67051,4.5497856,3.8443048,2.969056,2.746471,2.0673985,1.6524098,1.6222287,1.478869,1.026154,0.7394345,0.58475685,0.52439487,0.47912338,0.271629,0.422534,0.45648763,0.30935526,0.32821837,0.15845025,0.17731337,0.24899325,0.26408374,0.150905,0.116951376,0.116951376,0.1056335,0.08677038,0.08677038,0.5772116,0.845068,0.98465514,1.0336993,0.965792,0.7884786,0.513077,0.331991,0.34330887,0.55457586,0.83752275,0.6149379,0.33576363,0.2263575,0.26408374,0.8563859,1.8485862,2.493705,2.6710186,2.886058,2.6634734,2.1579416,1.720317,1.5505489,1.7127718,1.5467763,1.2902378,0.94692886,0.6149379,0.482896,0.3169005,0.24899325,0.21881226,0.17731337,0.08677038,0.049044125,0.026408374,0.0150905,0.0150905,0.011317875,0.011317875,0.003772625,0.011317875,0.02263575,0.0150905,0.018863125,0.10186087,0.211267,0.25276586,0.071679875,0.090543,0.07922512,0.07922512,0.1056335,0.14713238,0.392353,0.52439487,0.422534,0.26408374,0.5357128,0.6187105,1.4826416,1.629774,0.95447415,0.73566186,0.38103512,0.24899325,0.16222288,0.07922512,0.056589376,0.38480774,0.36971724,0.44139713,0.9997456,2.3993895,3.3953626,4.496969,4.9723196,4.7950063,4.6327834,4.2102494,3.610402,3.338773,3.4557245,3.5575855,4.036709,4.5497856,4.825187,4.587512,3.5387223,2.6106565,2.1277604,1.6675003,1.1393328,0.7997965,0.52062225,0.31312788,0.18485862,0.116951376,0.090543,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.06413463,0.27917424,0.35085413,0.181086,0.120724,0.25276586,0.40367088,0.33576363,1.4071891,1.9957186,1.6033657,0.8903395,1.2713746,2.1277604,2.7200627,2.6446102,1.841041,2.2748928,1.7165444,1.20724,1.6675003,3.8895764,3.0256453,2.1805773,2.0636258,2.335255,1.5807298,1.7731338,1.7127718,2.1768045,2.8634224,2.372981,2.384299,2.8709676,2.9841464,2.6823363,2.7087448,2.2069857,2.123988,1.991946,1.8297231,2.1277604,0.8639311,0.633801,1.0412445,1.9504471,3.5047686,2.4220252,2.2296214,2.3918443,2.052308,0.026408374,0.10186087,0.23013012,0.3470815,0.3734899,0.23767537,0.19994913,0.2565385,0.29803738,0.2867195,0.24522063,0.15467763,0.094315626,0.06413463,0.06790725,0.08299775,0.0754525,0.06413463,0.060362,0.06790725,0.1056335,0.090543,0.0452715,0.049044125,0.090543,0.1056335,0.08299775,0.05281675,0.033953626,0.033953626,0.033953626,0.10186087,0.271629,0.5093044,0.6752999,0.5394854,0.33953625,0.271629,0.27917424,0.362172,0.5772116,0.8601585,0.69793564,0.36971724,0.090543,0.033953626,0.011317875,0.02263575,0.041498873,0.05281675,0.0754525,0.05281675,0.03772625,0.033953626,0.041498873,0.049044125,0.041498873,0.033953626,0.026408374,0.018863125,0.0150905,0.026408374,0.041498873,0.049044125,0.05281675,0.026408374,0.030181,0.026408374,0.018863125,0.0150905,0.00754525,0.0150905,0.0150905,0.0150905,0.018863125,0.02263575,0.041498873,0.12826926,0.32444575,0.55457586,0.66020936,0.6451189,0.6187105,0.62625575,0.7809334,1.2525115,1.8863125,1.4750963,0.94315624,0.72811663,0.76584285,0.63002837,0.68661773,0.8903395,1.0223814,0.68661773,0.4979865,0.543258,0.7469798,0.9507015,0.8903395,0.3772625,0.513077,0.8865669,1.2826926,1.6825907,1.5543215,1.2034674,1.0751982,1.388326,2.1466236,2.4069347,2.848332,2.6031113,1.720317,1.1921495,1.2185578,1.6146835,2.173032,2.674791,2.897376,3.2935016,2.8709676,3.1312788,4.5761943,6.7341356,6.40969,6.221059,6.858632,7.3981175,5.2967653,2.7691069,2.0183544,1.780679,1.4260522,0.94692886,0.7582976,0.6790725,0.88279426,1.2713746,1.4826416,1.327964,1.0827434,0.95447415,0.9318384,0.80734175,0.77338815,0.84884065,1.0676528,1.2751472,1.0940613,1.3166461,1.5505489,1.7014539,1.6712729,1.3694628,1.2525115,1.2713746,1.2298758,1.086516,0.95447415,0.91674787,0.94315624,0.77716076,0.482896,0.422534,0.4640329,0.44894236,0.41876137,0.4074435,0.422534,0.39989826,0.3470815,0.29426476,0.271629,0.2867195,0.5055317,0.7054809,0.8903395,1.116697,1.4901869,1.6976813,1.0789708,0.65643674,0.91674787,1.8184053,4.395108,6.8737226,6.224831,2.9841464,1.237421,1.7354075,1.6863633,1.388326,1.1431054,1.2751472,1.0412445,1.0072908,1.3091009,1.6373192,1.2223305,1.0789708,1.0336993,1.0789708,1.1431054,1.1091517,0.9808825,1.1431054,1.5580941,2.0372176,2.233394,2.6182017,2.8936033,2.9313297,2.897376,3.259548,2.8181508,1.9466745,1.5920477,2.1390784,3.410453,5.142088,6.903904,7.7829256,8.039464,9.14107,8.899622,9.940866,10.699164,10.182315,7.9791017,6.3531003,6.247467,6.047518,4.889322,2.686109,1.8561316,1.6561824,1.7014539,1.9202662,2.546522,2.2786655,1.6863633,1.2147852,1.1355602,1.5316857,1.3770081,1.0072908,0.814887,0.845068,0.77716076,0.633801,0.48666862,0.42630664,0.43007925,0.36594462,0.35462674,0.35462674,0.36971724,0.44516975,0.663982,0.67152727,0.58098423,0.35462674,0.090543,0.00754525,0.011317875,0.0150905,0.0452715,0.08677038,0.1056335,0.0452715,0.011317875,0.0,0.00754525,0.03772625,0.05281675,0.090543,0.181086,0.35085413,0.63002837,1.2600567,2.2598023,3.9084394,6.0701537,8.201687,7.284939,6.398372,6.3342376,6.9152217,6.983129,5.172269,4.06689,3.519859,3.1652324,2.4182527,1.6524098,1.1016065,0.7432071,0.55080324,0.51684964,1.146878,1.3468271,1.1959221,1.0525624,1.5203679,1.6448646,1.539231,2.1994405,3.4029078,3.6896272,2.0372176,1.599593,1.6033657,1.6071383,1.5128226,1.2261031,0.98465514,0.87147635,0.965792,1.3543724,1.6675003,1.7240896,1.7240896,1.7240896,1.6373192,2.8747404,2.0862615,1.4977322,2.11267,3.6971724,5.9117036,7.0472636,6.3229194,4.5120597,3.9612563,3.99521,5.7494807,6.477597,5.6061206,4.749735,6.820906,7.586749,11.151879,16.935314,19.681786,21.032385,16.840998,12.083718,9.201432,8.073418,6.006019,4.4403796,4.1008434,5.7570257,10.231359,10.812344,9.793735,7.9715567,5.8437963,3.6368105,3.199186,3.8593953,5.3080835,7.6395655,11.363147,14.019074,14.807553,14.037937,12.287439,10.401127,11.608367,14.652876,17.429527,19.670467,22.941332,27.951378,33.45564,37.835655,41.163113,45.23,47.919884,50.326817,52.058453,53.299644,54.82756,60.316727,66.017166,69.83129,71.00835,70.12556,71.01589,72.95125,75.11674,77.746254,82.13382,86.14035,91.52011,94.98338,95.18333,92.746216,90.24873,90.448685,90.43737,89.18485,87.570175,83.80886,80.92658,74.77343,66.56797,62.86325,61.25611,61.980457,64.681656,68.0657,69.89165,69.823746,68.978676,68.95604,70.74426,74.73947,82.6733,87.36268,87.234406,83.17883,78.54605,75.59209,71.61197,68.16379,65.99075,64.99478,64.08181,61.765415,60.294094,59.20003,55.2765,51.168114,46.512695,42.174175,38.824085,36.926453,34.46293,32.621887,30.860073,29.034122,27.39303,26.563053,24.27307,22.401848,21.447372,20.504217,19.764782,18.568861,17.08999,15.62244,14.603831,14.245432,13.913441,13.626721,13.407909,13.290957,13.445636,16.893814,21.654867,25.325632,25.069094,22.066084,19.353567,16.954176,14.954685,13.502225,13.045737,12.792972,12.785426,12.808062,12.362892,12.113899,11.661184,11.276376,11.076427,11.042474,10.650121,10.740664,11.174516,11.725319,12.102581,12.58925,12.706201,12.626976,12.913695,14.524607,15.049001,14.739646,13.728582,11.970539,9.265567,8.484633,7.986647,7.462252,6.360646,3.893349,3.742444,3.5839937,3.2784111,2.7313805,1.9240388,1.5241405,1.1959221,0.97333723,1.0412445,1.720317,1.6410918,1.1808317,0.76584285,0.55457586,0.4376245,0.2867195,0.20372175,0.16976812,0.150905,0.116951376,0.10186087,0.1056335,0.1056335,0.15467763,0.41121614,0.6526641,0.8337501,0.935611,0.9507015,0.90920264,0.7130261,0.47535074,0.30935526,0.27917424,0.3961256,0.6375736,0.55080324,0.3470815,0.18863125,0.1961765,0.5093044,0.8865669,1.4373702,2.1164427,2.7011995,3.7235808,4.3611546,4.4139714,3.5689032,1.3807807,1.056335,0.90543,0.8639311,0.95447415,1.2789198,1.4071891,1.388326,1.0336993,0.47535074,0.18485862,0.15467763,0.11317875,0.06413463,0.02263575,0.0150905,0.00754525,0.003772625,0.018863125,0.0452715,0.033953626,0.056589376,0.11317875,0.17354076,0.24522063,0.3734899,0.8941121,0.77338815,0.4376245,0.17354076,0.150905,0.2867195,0.35839936,0.34330887,0.49421388,1.3355093,0.8186596,0.95824677,0.9205205,0.55457586,0.39989826,0.16222288,0.07922512,0.056589376,0.049044125,0.05281675,0.271629,0.35839936,0.8865669,2.052308,3.6971724,4.617693,6.326692,7.7829256,8.639311,9.231613,8.299775,6.187105,4.3385186,3.3425457,2.9464202,3.3576362,6.5228686,11.091517,12.811834,4.557331,2.516341,1.720317,1.3732355,1.116697,1.026154,0.7809334,0.5093044,0.3055826,0.19994913,0.1358145,0.00754525,0.0,0.011317875,0.011317875,0.00754525,0.03772625,0.120724,0.124496624,0.06790725,0.003772625,0.0150905,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.049044125,0.041498873,0.0754525,0.29803738,0.5998474,0.6526641,0.3961256,0.060362,0.16976812,0.543258,1.8184053,2.5012503,2.1956677,1.6109109,1.8485862,2.1541688,2.6785638,3.4632697,4.459243,3.4481792,1.931584,1.478869,2.505023,4.2706113,3.3425457,2.3767538,1.9881734,2.0900342,1.8749946,2.0070364,1.8561316,2.3201644,2.9916916,2.1315331,1.3430545,1.5354583,1.4260522,0.8941121,0.98842776,0.8903395,1.327964,1.8485862,1.9881734,1.2525115,1.1053791,1.9579924,2.4333432,2.5880208,3.9386206,2.7615614,1.7089992,0.9393836,0.52439487,0.41876137,0.2678564,0.29426476,0.32821837,0.2867195,0.15845025,0.24522063,0.28294688,0.27917424,0.25276586,0.24522063,0.17731337,0.124496624,0.09808825,0.1056335,0.13204187,0.120724,0.090543,0.06413463,0.060362,0.08677038,0.056589376,0.030181,0.033953626,0.0754525,0.150905,0.17731337,0.16222288,0.14713238,0.13204187,0.094315626,0.13958712,0.19994913,0.36971724,0.59230214,0.69793564,0.5017591,0.41121614,0.4074435,0.482896,0.6488915,0.845068,0.724344,0.44894236,0.18485862,0.11317875,0.033953626,0.026408374,0.060362,0.124496624,0.23013012,0.150905,0.0754525,0.041498873,0.049044125,0.060362,0.049044125,0.0452715,0.041498873,0.03772625,0.026408374,0.030181,0.033953626,0.041498873,0.0452715,0.02263575,0.033953626,0.026408374,0.02263575,0.026408374,0.02263575,0.02263575,0.02263575,0.02263575,0.02263575,0.030181,0.049044125,0.13204187,0.35085413,0.69039035,1.0638802,1.0940613,1.0072908,1.0186088,1.2638294,1.7769064,1.9391292,1.2864652,0.754525,0.6526641,0.65643674,0.4376245,0.3055826,0.24522063,0.241448,0.29426476,0.5394854,0.65643674,0.73188925,0.7922512,0.8299775,0.47157812,0.38480774,0.56589377,1.0110635,1.7052265,2.3503454,1.9655377,1.5203679,1.6448646,2.6446102,2.354118,2.886058,3.078462,2.595566,1.9391292,1.6033657,1.8184053,2.1315331,2.3880715,2.7426984,3.3651814,3.3312278,3.6028569,4.738417,6.862405,5.251494,5.0251365,6.039973,6.696409,3.9273026,1.9164935,1.7957695,1.8485862,1.4637785,1.1431054,0.935611,0.66020936,0.79602385,1.3166461,1.6863633,1.5958204,1.4298248,1.2940104,1.1883769,1.0148361,1.0676528,1.2638294,1.4637785,1.5656394,1.5052774,1.3317367,1.3355093,1.327964,1.1921495,0.91297525,0.845068,0.784706,0.7432071,0.7394345,0.80734175,1.0789708,1.1959221,0.9507015,0.5319401,0.51684964,0.4979865,0.49044126,0.44894236,0.40367088,0.4640329,0.5017591,0.39989826,0.28294688,0.23013012,0.3055826,0.73566186,0.8563859,0.8865669,1.0110635,1.3732355,1.6109109,1.1280149,0.7884786,0.9997456,1.7089992,3.6443558,4.5724216,3.863168,2.0258996,0.69793564,1.1091517,1.116697,1.0676528,1.146878,1.3543724,1.1242423,0.83752275,0.6413463,0.5696664,0.5696664,0.331991,0.3470815,0.5357128,0.76584285,0.8563859,0.59230214,0.7809334,1.2713746,1.8070874,2.0145817,2.1692593,2.3616633,2.354118,2.4899325,3.6934,2.969056,2.1503963,1.690136,1.901403,2.9728284,5.3269467,7.84706,9.574923,10.0465,9.310839,9.027891,9.997457,11.551778,12.2119875,9.699419,7.484888,6.8171334,6.405917,5.402399,3.3689542,3.127506,3.5274043,3.4368613,2.7426984,2.3578906,1.8070874,1.3505998,1.1129243,1.1808317,1.5882751,1.5467763,1.2298758,1.0751982,1.1883769,1.327964,1.0940613,0.9808825,0.90920264,0.7884786,0.52062225,0.38480774,0.35462674,0.40367088,0.5394854,0.7922512,0.8111144,0.6752999,0.41121614,0.13958712,0.06413463,0.026408374,0.00754525,0.011317875,0.02263575,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.02263575,0.056589376,0.1056335,0.21503963,0.56212115,1.6637276,3.742444,6.7341356,7.673519,6.934085,6.2814207,6.368191,6.7454534,5.9305663,5.383536,5.240176,5.191132,4.5120597,3.7009451,2.8294687,2.022127,1.3807807,0.9808825,0.66775465,0.45648763,0.35839936,0.43385187,0.77338815,0.9242931,0.86770374,1.116697,1.6863633,2.0862615,1.3091009,0.90543,0.76584285,0.77716076,0.8186596,0.76584285,0.77338815,0.9016574,1.0374719,0.8978847,1.2487389,1.7165444,2.071171,2.1654868,1.9391292,1.6109109,1.4939595,1.6071383,2.2560298,4.0216184,6.2436943,6.9755836,6.043745,4.4441524,4.315883,3.6594462,3.2972744,3.3915899,3.9801195,4.9534564,6.304056,6.7944975,12.140307,20.975796,24.854053,24.903097,21.232334,17.120173,14.162435,12.257258,8.228095,5.3080835,4.074435,4.5497856,6.1795597,6.802043,6.2021956,5.1647234,4.0404816,2.7653341,2.4069347,2.704972,3.4029078,4.538468,6.4134626,8.182823,9.405154,9.49947,8.428044,6.7077274,6.5266414,8.582722,10.955703,13.490907,17.814335,22.782883,26.280106,29.015259,31.848501,35.783348,39.2353,43.30219,47.025772,50.236275,53.55241,59.23776,65.91153,70.80085,73.52846,76.10894,79.164764,81.79051,83.82018,85.71781,88.57369,90.803314,93.070656,94.42126,94.81738,95.149376,94.07418,94.06286,94.930565,95.9454,95.83599,93.18761,90.158195,83.00907,73.72841,70.00483,68.84286,68.00534,68.26188,69.61248,71.30639,72.60417,74.6942,76.863464,79.24022,82.79025,90.803314,96.63202,98.61265,96.39812,90.9844,86.11017,81.277435,76.65219,72.89466,71.13662,71.31016,70.842354,70.63109,69.69925,65.18342,61.32402,56.91005,52.828068,49.64397,47.565254,44.792377,42.59671,40.506676,38.37514,36.35679,35.877663,33.66313,31.59196,30.377176,29.56229,28.479546,27.140265,25.514263,23.722265,21.990631,20.670212,19.47429,18.48209,17.73511,17.206944,17.372938,19.025349,21.647322,23.92976,23.793945,22.36412,21.032385,19.791191,18.572634,17.25976,16.324148,15.905387,15.863888,15.946886,15.803526,15.569623,15.116908,14.837734,14.803781,14.766054,14.385019,14.807553,15.426264,15.818617,15.758255,16.644821,17.25976,18.127462,19.383747,20.802254,20.994658,20.270313,18.738628,16.542961,13.830443,13.649357,12.81938,12.291212,11.532914,8.514814,8.224322,7.9489207,6.9680386,5.300538,3.6934,3.1727777,2.7389257,2.625747,2.886058,3.3878171,2.9464202,1.9655377,1.1431054,0.73188925,0.56589377,0.41498876,0.34330887,0.28294688,0.211267,0.16976812,0.1358145,0.10940613,0.10940613,0.22258487,0.5998474,0.5772116,0.694163,0.80356914,0.8224323,0.7394345,0.573439,0.36594462,0.2263575,0.1961765,0.24522063,0.38480774,0.4074435,0.331991,0.2263575,0.21881226,0.23013012,0.17354076,0.41876137,1.0110635,1.6825907,3.138824,4.293247,4.6516466,3.863168,1.7165444,0.9922004,0.7884786,0.9507015,1.4034165,2.1503963,2.263575,2.04099,1.4524606,0.7469798,0.45648763,0.51684964,0.3961256,0.23767537,0.11317875,0.05281675,0.030181,0.03772625,0.06413463,0.08299775,0.0452715,0.08677038,0.1358145,0.181086,0.27540162,0.5281675,1.1053791,1.0751982,0.76584285,0.4979865,0.56589377,0.46026024,0.33953625,0.29426476,0.5394854,1.4222796,0.90920264,0.724344,0.60362,0.44516975,0.30935526,0.14335975,0.06413463,0.08299775,0.16976812,0.241448,0.362172,0.8526133,2.2862108,4.398881,6.085244,7.0284004,8.9788475,11.170743,13.083464,14.437836,12.902377,9.0543,5.7683434,4.1197066,3.410453,4.4516973,10.303039,16.87118,18.263277,6.779407,2.7653341,1.2751472,0.87147635,0.754525,0.7696155,0.66775465,0.5017591,0.3470815,0.23390275,0.17354076,0.07922512,0.018863125,0.026408374,0.026408374,0.018863125,0.071679875,0.24899325,0.26031113,0.14335975,0.003772625,0.011317875,0.018863125,0.00754525,0.00754525,0.041498873,0.13958712,0.07922512,0.026408374,0.003772625,0.011317875,0.03772625,0.1358145,0.23767537,0.18863125,0.0452715,0.09808825,0.77716076,1.9730829,1.6373192,0.16976812,0.39989826,0.9280658,1.81086,2.5616124,2.9992368,3.259548,2.8030603,2.6031113,2.546522,3.6481283,8.035691,7.594294,4.217795,2.2748928,2.5314314,2.1541688,2.2899833,2.3126192,2.233394,2.0485353,1.7165444,1.5882751,1.5015048,1.8825399,2.2447119,1.1808317,0.6073926,0.45648763,0.60362,1.0714256,2.04099,1.327964,1.6373192,2.2409391,2.565385,2.1994405,1.8749946,3.4745877,3.519859,1.7542707,1.1657411,1.2034674,1.1280149,0.97710985,0.83752275,0.87902164,0.44894236,0.331991,0.27917424,0.18485862,0.10940613,0.241448,0.23390275,0.1961765,0.18485862,0.20372175,0.1659955,0.13204187,0.12826926,0.14713238,0.1659955,0.1659955,0.13204187,0.090543,0.06413463,0.03772625,0.03772625,0.033953626,0.041498873,0.06413463,0.120724,0.23013012,0.29803738,0.31312788,0.2867195,0.2263575,0.26031113,0.2565385,0.23390275,0.28294688,0.5885295,0.5394854,0.58475685,0.66020936,0.6752999,0.5017591,0.32444575,0.3772625,0.422534,0.36971724,0.26408374,0.1056335,0.049044125,0.07922512,0.18863125,0.3734899,0.3055826,0.1659955,0.0754525,0.060362,0.06413463,0.06413463,0.06413463,0.07922512,0.090543,0.06790725,0.060362,0.0452715,0.03772625,0.03772625,0.05281675,0.060362,0.060362,0.06413463,0.06790725,0.0452715,0.041498873,0.041498873,0.03772625,0.03772625,0.033953626,0.02263575,0.030181,0.124496624,0.41498876,1.0110635,1.1506506,1.0940613,1.0638802,1.1053791,1.0789708,0.5319401,0.32444575,0.33953625,0.49421388,0.7432071,0.40367088,0.26031113,0.2867195,0.38858038,0.41876137,0.7884786,0.68661773,0.5357128,0.55080324,0.7432071,0.6790725,0.66775465,0.6413463,0.7507524,1.3505998,2.8294687,2.7691069,2.123988,1.7316349,2.293756,1.871222,2.5125682,3.0746894,3.0256453,2.4559789,1.5882751,1.6373192,1.9127209,2.2786655,3.1840954,4.2102494,4.5007415,4.146115,3.7386713,4.38379,4.0291634,3.7198083,3.9386206,4.2404304,3.2520027,2.142851,2.2899833,2.3163917,1.901403,1.7693611,1.3656902,0.875249,0.8526133,1.3770081,2.04099,2.1051247,1.8863125,1.5807298,1.3204187,1.1996948,1.4298248,1.931584,2.233394,2.1579416,1.8146327,1.3015556,1.1695137,1.1091517,0.98465514,0.80356914,0.814887,0.8224323,0.7884786,0.73188925,0.7394345,1.0374719,1.0525624,0.8337501,0.56212115,0.5885295,0.5583485,0.5093044,0.44516975,0.42630664,0.55080324,0.5885295,0.44894236,0.271629,0.20372175,0.36971724,0.98842776,1.0676528,0.8526133,0.59607476,0.56212115,0.58098423,0.845068,1.177059,1.4147344,1.4147344,1.2826926,1.1921495,0.9318384,0.56589377,0.44516975,1.0450171,1.0487897,0.90920264,0.80734175,0.67152727,0.62625575,0.56212115,0.44139713,0.29803738,0.25276586,0.21503963,0.241448,0.46026024,0.79602385,0.9695646,0.6526641,0.7205714,0.94692886,1.2411937,1.6222287,1.9240388,2.2748928,2.384299,2.463524,3.2482302,2.1956677,1.9240388,1.6976813,1.5618668,2.323937,5.191132,7.6923823,10.0276375,11.449917,10.246449,8.13378,7.6207023,9.718282,12.921241,13.192869,9.405154,7.1000805,5.6815734,4.7535076,4.08198,4.7006907,5.764571,5.587258,4.1272516,2.9728284,2.1994405,1.4939595,1.177059,1.2638294,1.4524606,1.4750963,1.4335974,1.4600059,1.629774,1.9391292,2.11267,2.1315331,1.8448136,1.3053282,0.7696155,0.452715,0.39989826,0.5319401,0.7167987,0.79602385,0.633801,0.51684964,0.3734899,0.21881226,0.14713238,0.06790725,0.018863125,0.0150905,0.030181,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.0150905,0.0150905,0.018863125,0.0150905,0.026408374,0.09808825,0.3961256,1.1959221,2.897376,5.194905,5.1835866,4.5120597,4.123479,4.274384,4.7308717,5.2967653,5.8173876,6.085244,5.8588867,5.523123,4.6214657,3.531177,2.4710693,1.50905,0.9318384,0.56212115,0.38103512,0.34330887,0.34330887,0.5470306,0.6187105,0.6375736,0.7054809,0.94315624,0.79602385,0.48666862,0.28294688,0.25276586,0.26408374,0.36971724,0.5998474,0.84884065,0.9280658,0.5696664,1.0638802,1.6486372,2.0862615,2.2862108,2.3126192,2.082489,1.8749946,1.6637276,1.5656394,1.8297231,2.1956677,1.8297231,1.629774,1.9202662,2.4371157,1.9844007,1.6712729,2.4899325,4.1989317,5.342037,7.0284004,7.4282985,12.1101265,20.602304,26.389511,23.548725,20.274086,18.62545,17.96524,14.939595,10.502988,7.443389,5.8211603,5.0968165,4.1272516,4.2781568,3.8669407,3.0860074,2.323937,2.191895,1.8900851,1.8259505,1.8976303,2.082489,2.3993895,2.8521044,3.500996,4.1310244,4.508287,4.357382,4.1197066,4.678055,6.039973,8.616675,13.211733,17.72002,20.885252,23.507227,26.189562,29.335932,33.504684,37.89979,41.993088,45.93171,50.54563,55.336864,61.0788,66.45479,71.468605,77.4369,83.28447,88.10211,91.52766,93.662964,95.07015,97.24318,97.858116,97.06587,95.53418,94.4288,92.22936,90.48641,90.856125,92.97257,94.4288,94.29676,92.60663,88.66801,83.17129,78.198975,80.6625,80.47009,78.44797,76.02971,75.241234,77.23318,81.8471,85.472595,87.12123,88.437874,92.01432,96.88478,102.45318,106.5427,105.44109,99.12949,93.55356,88.37751,83.661736,79.86647,78.17256,77.859436,77.56517,76.120255,72.52872,69.133354,65.17964,61.86728,59.44148,57.17036,54.691746,52.70357,50.95307,49.145985,46.920135,45.976982,44.747105,43.30219,41.92141,41.083885,39.718197,38.477,37.22449,35.65508,33.319824,30.607307,28.249416,26.012249,23.914669,22.235851,21.156881,20.48158,21.288923,23.046967,23.62795,23.793945,23.390276,22.892288,22.394302,21.579414,20.828663,20.274086,19.945868,19.779873,19.621422,19.591242,19.43279,19.406384,19.481836,19.334703,19.1423,19.662922,20.29295,20.734346,20.99843,21.956678,23.028103,24.755966,26.834682,28.087193,26.680004,24.872917,22.616886,20.209951,18.312323,19.651604,19.153618,18.648085,18.240643,16.316603,16.060064,15.131999,12.887287,9.767326,7.3113475,6.432326,5.704209,5.613666,5.7909794,5.0138187,3.663219,2.5201135,1.5543215,0.87147635,0.73188925,0.4979865,0.47535074,0.49044126,0.44139713,0.29426476,0.21881226,0.12826926,0.11317875,0.2263575,0.48666862,0.41876137,0.5281675,0.65643674,0.6752999,0.5055317,0.39989826,0.25276586,0.15845025,0.16222288,0.241448,0.33576363,0.29803738,0.271629,0.27917424,0.25276586,0.13204187,0.08299775,0.056589376,0.090543,0.34330887,0.94692886,1.7618159,2.1805773,2.1994405,2.4107075,1.3732355,1.0450171,1.2034674,1.7693611,2.7841973,2.6898816,1.9994912,1.2864652,0.87902164,0.8639311,0.94315624,0.73188925,0.5017591,0.33953625,0.15845025,0.10186087,0.10940613,0.12826926,0.120724,0.060362,0.11317875,0.19240387,0.271629,0.35085413,0.45648763,0.66775465,0.8903395,0.95447415,0.9393836,1.1393328,0.80734175,0.47157812,0.30181,0.392353,0.7469798,0.97710985,1.1091517,0.9280658,0.543258,0.38858038,0.211267,0.08677038,0.13204187,0.32821837,0.513077,0.6752999,1.5958204,3.8782585,6.9189944,8.880759,10.0276375,11.846043,14.158662,16.51278,18.153872,15.7657995,10.838752,7.1604424,5.783434,5.0025005,6.5040054,12.664702,17.169216,16.109108,7.9791017,2.806833,0.91674787,0.43007925,0.27917424,0.20372175,0.23013012,0.27540162,0.2678564,0.21503963,0.19240387,0.33576363,0.07922512,0.0150905,0.0150905,0.011317875,0.0,0.049044125,0.041498873,0.018863125,0.0,0.0,0.02263575,0.011317875,0.03772625,0.21503963,0.70170826,0.3961256,0.12826926,0.011317875,0.049044125,0.120724,0.32821837,0.694163,0.5583485,0.049044125,0.060362,1.2562841,5.036454,4.5912848,0.44894236,0.47157812,1.0223814,2.3126192,3.3953626,4.002755,4.5761943,2.4899325,1.8674494,2.3993895,4.5196047,9.4127,12.332711,7.1378064,2.5314314,1.4939595,1.3128735,1.8976303,2.7879698,2.957738,2.4710693,2.4710693,2.033445,1.4298248,1.3807807,1.8523588,2.0598533,1.388326,0.7432071,1.6222287,4.5912848,9.291975,4.9345937,1.9693103,2.4522061,5.5080323,7.3377557,2.444661,1.5316857,1.6222287,1.237421,0.3961256,0.33576363,0.49421388,0.63002837,0.62248313,0.48666862,0.4376245,0.34330887,0.21503963,0.09808825,0.060362,0.08677038,0.10186087,0.13204187,0.181086,0.23013012,0.19240387,0.1659955,0.15845025,0.1659955,0.1659955,0.21503963,0.19240387,0.14335975,0.09808825,0.060362,0.060362,0.08677038,0.11317875,0.120724,0.120724,0.18485862,0.3169005,0.3772625,0.33576363,0.27540162,0.29803738,0.3961256,0.3961256,0.29426476,0.26031113,0.35839936,0.70170826,1.0601076,1.1619685,0.68661773,0.331991,0.5017591,0.7092535,0.7054809,0.47157812,0.26408374,0.15845025,0.116951376,0.12826926,0.21503963,0.35839936,0.31312788,0.19994913,0.10186087,0.0754525,0.124496624,0.10940613,0.12826926,0.17731337,0.150905,0.1659955,0.150905,0.124496624,0.11317875,0.1358145,0.124496624,0.15845025,0.18485862,0.1659955,0.1056335,0.08299775,0.0754525,0.071679875,0.056589376,0.0452715,0.0452715,0.0452715,0.120724,0.31312788,0.65643674,0.6790725,0.62248313,0.52062225,0.35839936,0.090543,0.13958712,0.271629,0.33953625,0.32821837,0.36594462,0.18485862,0.1358145,0.26031113,0.49044126,0.68661773,0.784706,0.56212115,0.6111652,0.8526133,0.5357128,0.66775465,0.8563859,0.8526133,0.7432071,0.9620194,2.4861598,3.3161373,3.059599,2.2296214,2.2447119,2.2786655,2.4069347,2.7502437,2.9464202,2.1503963,1.5279131,1.7844516,2.4861598,3.4783602,4.881777,5.7004366,5.0553174,3.6443558,2.5389767,3.1727777,6.1041074,5.1798143,3.7990334,3.6934,4.9119577,3.4255435,2.9954643,2.9124665,2.7841973,2.5616124,2.11267,1.3317367,0.94692886,1.1506506,1.6033657,1.5769572,1.4260522,1.3505998,1.3958713,1.418507,1.7014539,1.9353566,1.8146327,1.3128735,0.70170826,0.83752275,0.9507015,0.8299775,0.5470306,0.47157812,0.77716076,1.1016065,1.1921495,1.0676528,1.0072908,1.0299267,0.935611,0.77716076,0.5998474,0.44139713,0.392353,0.392353,0.41498876,0.45648763,0.5017591,0.44139713,0.29803738,0.18485862,0.23390275,0.62625575,0.88279426,0.8262049,0.58475685,0.35462674,0.42630664,0.7205714,1.5731846,2.6219745,3.1840954,2.2447119,1.4864142,1.3053282,1.0789708,0.7130261,0.6413463,0.995973,0.9922004,0.72811663,0.35462674,0.060362,0.08677038,0.19240387,0.35839936,0.52062225,0.59607476,0.59607476,0.63002837,1.0902886,1.7995421,2.0447628,1.4826416,1.5241405,1.7882242,2.0862615,2.4408884,2.0372176,1.780679,1.8297231,2.123988,2.3805263,2.0145817,1.6486372,1.4713237,1.7731338,2.9464202,5.617439,7.696155,8.880759,9.110889,8.575176,6.549277,6.1908774,8.631766,13.106099,16.950403,11.204697,6.990674,4.5497856,3.7877154,4.2894745,4.459243,4.3196554,3.8782585,3.3764994,3.2670932,3.1539145,2.7691069,2.3126192,1.8070874,1.0978339,1.599593,2.3654358,2.505023,2.0636258,2.0145817,3.5160866,3.983892,3.2029586,1.6863633,0.67152727,0.35462674,0.27540162,0.38480774,0.56589377,0.62625575,0.44139713,0.3772625,0.3470815,0.29426476,0.18485862,0.08677038,0.02263575,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.041498873,0.056589376,0.041498873,0.0150905,0.0150905,0.00754525,0.00754525,0.026408374,0.0754525,0.8337501,1.4260522,1.7429527,1.8297231,1.8938577,2.9539654,4.1612053,4.6629643,4.45547,4.395108,4.52715,4.315883,3.8141239,3.0256453,1.8749946,0.935611,0.52062225,0.33576363,0.23390275,0.19994913,0.23390275,0.23390275,0.35085413,0.5885295,0.80734175,0.56589377,0.422534,0.2565385,0.090543,0.090543,0.13958712,0.3169005,0.3169005,0.181086,0.29049212,0.5583485,0.7432071,0.8563859,1.0940613,1.8599042,2.3126192,1.9693103,1.358145,0.87902164,0.7922512,0.7696155,0.965792,1.0638802,0.98465514,0.9016574,0.9242931,1.0676528,2.9124665,5.8513412,7.111398,10.174769,10.38981,10.880251,14.132254,22.01704,18.221779,17.546478,18.274595,18.187824,14.588741,10.461489,7.598067,6.273875,5.8702044,4.881777,6.809588,6.779407,5.6513925,4.304565,3.6330378,2.7653341,2.0447628,1.7089992,1.7655885,1.9844007,2.727608,2.886058,3.0935526,3.4670424,3.6028569,4.1762958,5.2062225,6.571913,8.254503,10.329447,12.404391,14.298248,15.762027,16.946632,18.387774,18.523588,22.024584,27.891016,33.80649,36.164383,40.204865,44.886692,52.016953,61.422108,70.97062,77.40295,83.707,88.21152,90.3355,90.59204,94.76834,99.97456,101.611885,99.2389,96.60184,88.97359,84.16349,84.62375,89.25654,93.42906,92.41799,89.89411,88.18888,87.55885,86.18185,90.9429,94.3458,96.081215,96.29625,95.624725,95.34555,96.36416,96.51129,95.11165,93.002754,92.96503,97.36013,105.53164,114.66894,119.79594,115.15561,108.89682,102.155136,95.20974,87.50981,82.84685,80.83604,79.93438,78.88936,76.75028,74.92056,72.29104,69.89919,67.51112,63.629093,61.444744,60.886395,60.98448,60.90903,59.980965,58.98122,58.483234,57.751343,56.830822,56.562965,55.929165,53.92213,51.454834,48.83663,45.76194,42.890972,40.87262,37.786613,33.67445,30.562035,26.532871,23.7864,22.877197,23.446865,24.21648,26.166927,27.159128,27.39303,27.083675,26.47251,25.800982,25.001186,24.118391,23.280869,22.718748,23.744902,24.457928,24.967232,25.269043,25.269043,25.476536,25.544443,25.816072,26.404602,27.23458,28.664404,30.165909,31.659868,33.323597,35.5834,32.41062,29.939552,28.26828,27.359077,27.053493,27.053493,26.962952,25.702894,23.80149,23.360094,24.227798,23.307278,20.281631,15.992157,12.449662,11.2801485,9.940866,9.06939,8.284684,6.2097406,4.134797,2.8181508,1.8448136,1.1091517,0.8526133,0.6111652,0.5017591,0.5357128,0.56212115,0.3055826,0.27917424,0.1659955,0.08677038,0.09808825,0.18485862,0.36594462,0.58475685,0.7092535,0.663982,0.45648763,0.32444575,0.26408374,0.20749438,0.1659955,0.23013012,0.31312788,0.32821837,0.30181,0.25276586,0.1659955,0.241448,0.13958712,0.041498873,0.0150905,0.0150905,0.08677038,0.573439,1.0374719,1.3128735,1.4939595,1.3355093,1.1695137,1.3091009,1.9768555,3.2972744,3.6141748,2.4031622,1.2525115,0.9016574,1.20724,0.875249,0.70170826,0.7130261,0.73188925,0.36594462,0.23013012,0.16222288,0.1358145,0.1358145,0.120724,0.1961765,0.27917424,0.39989826,0.5281675,0.56589377,0.845068,1.1355602,1.2525115,1.2110126,1.237421,1.1883769,0.8639311,0.56589377,0.47912338,0.68661773,1.5430037,1.4335974,1.0450171,0.66775465,0.23013012,0.181086,0.094315626,0.056589376,0.14713238,0.42630664,0.6111652,1.4524606,3.9197574,7.7678347,11.566868,12.762791,14.086982,15.943113,17.99542,19.180025,14.909414,10.487898,8.073418,7.6622014,7.1264887,7.2094865,9.099571,9.993684,8.416726,4.2404304,1.7391801,0.6451189,0.27917424,0.181086,0.1056335,0.08299775,0.13204187,0.19994913,0.241448,0.23013012,0.43385187,0.35462674,0.16976812,0.0452715,0.030181,0.09808825,0.20372175,0.331991,0.23767537,0.071679875,0.36594462,0.62625575,0.39989826,0.1358145,0.090543,0.32444575,0.47912338,0.45648763,0.2867195,0.08677038,0.071679875,0.97333723,1.6863633,2.1654868,1.9391292,0.09808825,0.7582976,3.6028569,4.3422914,2.252257,0.1659955,0.47157812,0.935611,1.7542707,2.5993385,2.5880208,2.2296214,2.674791,2.9803739,3.3350005,5.0553174,5.726845,4.353609,2.4333432,0.97710985,0.482896,1.2638294,1.8184053,2.776652,4.3385186,6.2814207,4.504514,1.9164935,0.5394854,0.8639311,1.8523588,2.1088974,4.6252384,5.511805,4.168751,3.3123648,2.1164427,2.2560298,3.0822346,4.3309736,6.1418333,2.3126192,1.1091517,1.1317875,1.3505998,1.1053791,0.5357128,3.3651814,3.7235808,1.1657411,0.67152727,0.55457586,0.35462674,0.17731337,0.0754525,0.049044125,0.05281675,0.056589376,0.08677038,0.15467763,0.25276586,0.27540162,0.2263575,0.17731337,0.15467763,0.15467763,0.25276586,0.2565385,0.211267,0.15467763,0.10940613,0.10186087,0.08677038,0.09808825,0.11317875,0.071679875,0.08677038,0.14335975,0.18485862,0.18485862,0.150905,0.26408374,0.392353,0.5319401,0.663982,0.724344,0.4678055,0.35462674,0.62625575,0.9997456,0.663982,0.3169005,0.2678564,0.33576363,0.38480774,0.33953625,0.29803738,0.25276586,0.19240387,0.124496624,0.1056335,0.211267,0.30935526,0.30935526,0.23390275,0.211267,0.150905,0.10940613,0.11317875,0.1659955,0.24899325,0.28294688,0.23390275,0.16976812,0.150905,0.22258487,0.29049212,0.3055826,0.271629,0.20749438,0.15467763,0.13958712,0.116951376,0.090543,0.071679875,0.056589376,0.056589376,0.041498873,0.049044125,0.08677038,0.15467763,0.19994913,0.20372175,0.39989826,0.6073926,0.26408374,0.4376245,0.6149379,0.6111652,0.42630664,0.2678564,0.18485862,0.10186087,0.07922512,0.14713238,0.331991,0.32444575,0.2867195,0.49421388,0.8337501,0.7922512,0.6413463,0.724344,0.7696155,0.72811663,0.7432071,1.0374719,1.8221779,2.323937,2.3088465,2.0975795,2.191895,2.1164427,2.1994405,2.6068838,3.3350005,2.916239,2.8822856,3.2029586,4.1272516,6.1644692,6.8058157,5.8211603,4.22534,2.897376,2.5767028,4.3422914,3.6330378,3.0407357,3.6783094,5.1835866,4.2894745,3.783943,3.4444065,3.0746894,2.5012503,2.625747,2.11267,1.4034165,0.9620194,1.297783,1.6712729,1.8184053,1.8033148,1.690136,1.5279131,1.3619176,1.2411937,1.267602,1.3505998,1.237421,1.5505489,1.6146835,1.5543215,1.478869,1.4750963,1.5052774,1.5052774,1.5467763,1.6146835,1.5920477,1.2261031,0.8601585,0.58475685,0.41498876,0.29426476,0.3169005,0.3734899,0.35839936,0.2867195,0.29426476,0.26408374,0.21503963,0.2565385,0.42630664,0.7092535,0.76207024,0.633801,0.452715,0.4074435,0.7432071,0.8526133,1.7240896,2.372981,2.263575,1.3166461,0.9280658,0.7997965,0.7205714,0.6451189,0.69039035,0.7884786,0.7394345,0.66775465,0.5885295,0.40367088,0.55457586,0.9280658,1.2638294,1.4071891,1.3166461,1.267602,1.3770081,1.6788181,2.052308,2.2296214,1.8599042,1.5354583,1.478869,1.7391801,2.161714,1.5618668,1.1619685,1.0601076,1.3505998,2.123988,2.5087957,2.1768045,2.0900342,2.3993895,2.4559789,3.380272,3.85185,4.006528,4.055572,4.2781568,4.587512,5.8211603,7.432071,8.903395,9.752235,10.220041,9.914458,8.069645,5.560849,4.9119577,2.9615107,1.9051756,1.5920477,2.1164427,3.802806,4.991183,4.7648253,3.682082,2.335255,1.3430545,1.8636768,2.0900342,1.991946,1.8297231,2.173032,2.8143783,2.173032,1.3958713,1.0072908,0.8903395,0.7582976,0.76207024,0.97710985,1.1883769,0.90543,0.44139713,0.23013012,0.18863125,0.18485862,0.08677038,0.03772625,0.030181,0.05281675,0.06413463,0.011317875,0.003772625,0.0,0.0,0.003772625,0.011317875,0.003772625,0.02263575,0.033953626,0.026408374,0.003772625,0.02263575,0.011317875,0.0,0.003772625,0.0150905,0.1659955,0.3055826,0.4376245,0.6413463,1.0638802,2.0560806,3.0860074,3.5538127,3.2972744,2.5993385,2.2371666,1.8900851,1.6410918,1.4034165,0.9507015,1.1129243,0.69039035,0.27917424,0.10940613,0.05281675,0.08677038,0.0754525,0.07922512,0.12826926,0.211267,0.21881226,0.18485862,0.120724,0.06790725,0.06790725,0.1659955,0.331991,0.32821837,0.22258487,0.41121614,0.86770374,1.1506506,1.1921495,1.2034674,1.690136,1.9466745,1.4939595,0.875249,0.47157812,0.513077,0.51684964,0.76584285,0.86770374,0.784706,0.8262049,0.724344,0.72811663,1.4750963,3.048281,4.949684,12.47607,16.490145,17.452164,17.240896,19.149845,16.376965,15.0376835,15.399856,15.113135,9.22784,6.881268,5.802297,5.7570257,6.085244,5.7004366,6.0286546,6.3153744,6.0512905,5.243949,4.436607,4.214022,3.2255943,2.6974268,3.0030096,3.6330378,3.5575855,3.361409,3.350091,3.5538127,3.7348988,3.9688015,4.878004,5.6287565,5.9984736,6.375736,7.326438,8.91094,10.612394,12.053536,12.955194,12.355347,13.128735,15.301767,18.361366,21.236107,25.35204,29.196344,33.88572,40.6274,50.730488,58.82277,67.53376,75.16578,80.76813,84.15972,91.52766,95.51155,96.35661,95.67,96.43207,92.59154,88.17379,88.89059,95.707726,104.84125,103.24165,96.76406,91.1353,88.66801,88.25679,89.05281,90.939125,91.93133,91.50124,90.584496,89.5923,92.44063,97.07719,101.11767,101.82692,103.17752,105.78818,110.07388,114.55199,115.842224,113.03916,109.94184,105.40337,99.416214,93.10084,87.47963,83.224106,80.27014,78.47814,77.6293,77.89716,78.2216,78.07825,77.07095,74.90924,72.09863,70.76313,70.74804,71.43843,71.76287,71.33656,70.69899,69.759605,69.11826,70.05387,71.0008,70.755585,69.71811,67.67712,63.851677,58.072018,53.495823,49.704334,46.290108,42.85702,39.978508,36.37942,33.51977,31.939043,31.222244,31.05625,31.44483,31.96168,32.425713,32.919926,33.22551,33.278324,32.59548,31.075111,28.981306,27.332668,26.785637,26.966724,27.574116,28.34373,30.00746,30.98457,31.109066,31.052477,32.301216,33.54618,35.71167,40.891483,46.814503,46.83714,41.19329,37.32258,35.119366,34.240345,34.108303,32.350258,29.286888,26.378195,25.646305,29.660378,33.708405,32.04845,27.683523,22.892288,19.225298,16.25624,13.996439,12.121444,10.227587,7.8206515,6.828451,5.8098426,4.6516466,3.5123138,2.806833,1.9957186,1.2864652,0.8299775,0.5998474,0.392353,0.3169005,0.24899325,0.18485862,0.150905,0.20749438,0.36971724,0.43385187,0.5357128,0.6073926,0.3734899,0.24899325,0.211267,0.1961765,0.1659955,0.13204187,0.1961765,0.211267,0.211267,0.20372175,0.1659955,0.23013012,0.18863125,0.15845025,0.15467763,0.0754525,0.041498873,0.16976812,0.90920264,1.8297231,1.6410918,1.4826416,1.2261031,1.026154,1.0148361,1.3053282,1.5543215,1.358145,1.1204696,1.1091517,1.4600059,1.327964,0.94692886,0.845068,0.995973,0.80734175,0.56212115,0.38480774,0.38103512,0.5017591,0.5357128,0.47535074,0.38103512,0.3772625,0.47535074,0.5885295,0.6828451,0.7167987,0.7130261,0.73188925,0.845068,1.0601076,1.116697,0.965792,0.724344,0.68661773,1.4449154,1.2449663,0.935611,0.7696155,0.4376245,0.23013012,0.120724,0.094315626,0.25276586,0.80734175,0.73566186,1.1846043,2.3163917,4.2706113,7.1604424,10.612394,13.226823,15.437581,17.180534,17.886015,13.996439,10.797253,8.786444,7.4018903,5.040227,6.511551,12.849561,19.772327,21.869907,12.577931,4.889322,1.4713237,0.35462674,0.1659955,0.094315626,0.060362,0.071679875,0.11317875,0.1659955,0.20372175,0.30181,0.83752275,0.4074435,0.02263575,0.02263575,0.094315626,0.5696664,0.8601585,0.6149379,0.16222288,0.513077,0.7922512,0.5357128,0.19240387,0.02263575,0.090543,0.3169005,0.86770374,1.0186088,0.6111652,0.071679875,0.7130261,2.1768045,4.719554,6.168242,1.9202662,1.0450171,4.346064,4.949684,2.5427492,3.3878171,0.935611,0.68661773,1.4600059,2.354118,2.7238352,3.059599,2.8521044,2.425798,2.6898816,5.119452,4.938366,3.7348988,2.6068838,1.8938577,1.1808317,3.7613072,7.7376537,8.6581745,6.2135134,4.221567,3.1199608,1.448688,0.4074435,1.026154,4.172523,4.112161,5.5457587,6.881268,6.7756343,4.1498876,2.8030603,3.0030096,3.3463185,3.2067313,2.7502437,1.9768555,1.418507,1.0487897,0.8299775,0.73188925,0.35085413,3.2520027,3.5877664,1.0336993,0.7997965,0.59230214,0.34330887,0.15467763,0.060362,0.03772625,0.030181,0.026408374,0.05281675,0.124496624,0.241448,0.32821837,0.29803738,0.21881226,0.16976812,0.23390275,0.42630664,0.35462674,0.24522063,0.18485862,0.15845025,0.10940613,0.08299775,0.08299775,0.08299775,0.033953626,0.07922512,0.14335975,0.26408374,0.4074435,0.47912338,0.47535074,0.4376245,0.5357128,0.77338815,0.965792,0.5093044,0.2678564,0.3772625,0.69793564,0.83752275,0.7696155,0.5470306,0.35462674,0.28294688,0.29426476,0.39989826,0.41876137,0.36594462,0.271629,0.17731337,0.1659955,0.19994913,0.21881226,0.2263575,0.27917424,0.1659955,0.09808825,0.08677038,0.12826926,0.211267,0.23390275,0.1961765,0.13958712,0.10940613,0.150905,0.1659955,0.16976812,0.15845025,0.13958712,0.150905,0.14335975,0.12826926,0.11317875,0.1056335,0.07922512,0.06413463,0.041498873,0.030181,0.033953626,0.041498873,0.060362,0.071679875,0.181086,0.32821837,0.31312788,0.6187105,0.86770374,0.8601585,0.58098423,0.23390275,0.35085413,0.2678564,0.150905,0.120724,0.25276586,0.24522063,0.26408374,0.47912338,0.8186596,0.94692886,0.94692886,1.0186088,0.9922004,0.8224323,0.60362,0.6073926,1.4637785,2.0183544,2.0258996,2.161714,2.071171,1.7957695,2.161714,3.187868,4.0706625,4.4139714,3.5839937,2.9841464,3.3764994,4.8629136,5.674028,5.093044,4.293247,3.8593953,3.7914882,4.9949555,3.821669,2.6597006,2.7653341,4.2592936,4.496969,4.9647746,5.323174,5.2099953,4.236658,3.6179473,2.7804246,1.9127209,1.2864652,1.237421,1.81086,2.1692593,2.0900342,1.7089992,1.539231,1.3732355,1.3015556,1.2261031,1.1317875,1.0638802,1.388326,1.3807807,1.358145,1.4373702,1.5580941,1.690136,1.7429527,1.8184053,1.841041,1.5580941,1.056335,0.67152727,0.41876137,0.2678564,0.15845025,0.150905,0.21503963,0.2565385,0.26031113,0.29049212,0.331991,0.30181,0.29803738,0.3734899,0.55080324,0.5772116,0.59230214,0.6451189,0.7582976,0.935611,0.8262049,1.0412445,1.1959221,1.116697,0.8186596,0.91297525,0.935611,0.845068,0.76584285,0.98465514,0.9507015,0.90543,0.87902164,0.80734175,0.51684964,0.7130261,1.20724,1.6448646,1.8787673,1.9730829,1.9164935,1.8900851,1.7655885,1.6033657,1.6524098,1.4147344,1.1544232,1.1695137,1.4864142,1.8523588,1.388326,0.8601585,0.7054809,0.97333723,1.3166461,1.5128226,1.629774,1.9353566,2.263575,2.0598533,2.3805263,2.655928,2.686109,2.5087957,2.4182527,4.349837,6.779407,8.303548,7.8244243,4.5535583,5.409944,6.8850408,7.61693,6.862405,4.508287,2.1843498,1.1695137,1.0223814,1.6033657,3.0935526,5.3269467,4.9647746,3.4670424,2.071171,1.8070874,2.5427492,2.4484336,1.8749946,1.3015556,1.3619176,1.5920477,1.1657411,0.9318384,1.3204187,2.3390274,2.6823363,2.3163917,1.6410918,0.9808825,0.59230214,0.28294688,0.13958712,0.09808825,0.090543,0.041498873,0.0150905,0.0150905,0.030181,0.05281675,0.07922512,0.0150905,0.011317875,0.018863125,0.0150905,0.00754525,0.0,0.00754525,0.011317875,0.011317875,0.0,0.05281675,0.03772625,0.011317875,0.0,0.0,0.0,0.0150905,0.05281675,0.14713238,0.35085413,0.9016574,1.3392819,1.6448646,1.7165444,1.3355093,0.94315624,0.65643674,0.5281675,0.49421388,0.35839936,0.5885295,0.46026024,0.26408374,0.1358145,0.05281675,0.0452715,0.030181,0.0150905,0.003772625,0.02263575,0.06790725,0.06413463,0.041498873,0.030181,0.060362,0.12826926,0.21503963,0.24522063,0.22258487,0.241448,0.7432071,1.1808317,1.3166461,1.2751472,1.5731846,1.4977322,0.935611,0.41121614,0.181086,0.23013012,0.271629,0.41498876,0.452715,0.38480774,0.4074435,0.4678055,0.56589377,0.9620194,1.81086,3.1652324,7.809334,11.408418,13.211733,13.5663595,13.936077,13.890805,15.335721,16.648594,15.705438,9.884277,7.4811153,7.0510364,6.9265394,6.6662283,7.0585814,6.85486,7.273621,7.2962565,6.752999,6.349328,7.0887623,6.6850915,5.617439,4.3913355,3.5575855,3.3953626,3.4632697,3.6481283,3.742444,3.440634,3.572676,4.2819295,4.5837393,4.3083377,4.104616,4.3083377,4.991183,6.300284,8.035691,9.646602,10.834979,11.615912,12.347801,13.728582,16.761772,19.930779,22.10381,24.657877,28.977533,36.443558,44.430206,53.741043,62.16154,68.6165,73.158745,78.66678,80.80962,81.37552,80.77945,78.0707,79.04404,77.81793,77.67081,80.61345,87.35513,87.71353,85.28019,83.88055,84.83502,86.9741,86.14035,87.50981,88.57746,88.48315,87.98893,87.58526,88.41147,89.28671,89.82997,90.47509,94.560844,98.66169,102.864395,106.6672,108.96473,105.03365,102.8078,100.393326,97.64308,96.15289,93.33474,90.68636,88.43033,86.78547,85.95171,86.21203,86.71756,87.32872,87.63431,86.95523,85.966805,85.389595,85.2236,85.219826,84.850105,84.072945,83.01284,81.63206,80.27392,79.670296,79.44394,78.61396,78.3461,78.02543,75.241234,71.93264,69.40875,66.97541,64.2478,61.142933,58.283283,55.13314,51.91132,48.810223,45.965664,44.200073,43.07206,42.174175,41.166885,39.76724,39.480522,40.446312,40.929207,40.20109,38.522274,36.428467,35.187275,34.25921,33.57259,33.534863,34.69683,36.122883,37.307487,38.031834,38.382687,38.378914,40.917892,46.399513,51.930183,51.29261,46.75037,44.117077,42.5288,40.793396,37.41312,33.244373,29.354795,28.74363,33.331142,43.95108,46.614555,40.14073,31.799456,25.714212,22.877197,21.38701,18.946123,16.146835,13.449409,11.200924,10.246449,9.231613,8.213005,7.4169807,7.250985,6.3342376,4.825187,3.0822346,1.659955,1.2713746,0.87902164,0.62248313,0.46026024,0.3772625,0.4074435,0.573439,0.573439,0.56212115,0.5772116,0.56212115,0.5583485,0.33576363,0.1659955,0.12826926,0.1358145,0.1659955,0.181086,0.17354076,0.18485862,0.2678564,0.18863125,0.16976812,0.21881226,0.271629,0.1659955,0.124496624,0.1056335,0.44139713,0.97333723,1.0299267,1.1280149,0.9620194,0.6790725,0.452715,0.48666862,0.66020936,0.8111144,0.90543,1.0450171,1.4335974,1.4939595,1.0751982,0.784706,0.7884786,0.8337501,0.573439,0.40367088,0.41121614,0.5281675,0.55080324,0.34330887,0.26408374,0.29426476,0.36971724,0.35839936,0.42630664,0.44894236,0.4640329,0.52439487,0.7092535,0.95447415,1.1657411,1.1053791,0.7997965,0.5017591,0.8337501,0.73188925,0.68661773,0.8111144,0.8639311,0.5394854,0.38480774,0.44894236,0.6752999,0.90920264,0.80356914,1.0035182,1.4600059,2.6144292,5.3986263,9.582467,11.23865,12.31762,14.403882,18.689585,16.343012,11.710228,7.6508837,5.6400743,5.772116,12.351574,19.53088,23.733583,21.934042,11.634775,5.240176,1.8749946,0.5055317,0.19240387,0.090543,0.056589376,0.0452715,0.06413463,0.10186087,0.1358145,0.150905,0.7394345,0.35462674,0.0,0.00754525,0.0452715,0.47912338,1.2336484,1.2110126,0.51684964,0.42630664,1.1431054,1.026154,0.56589377,0.14335975,0.0,0.13204187,0.91674787,1.5543215,1.50905,0.5017591,0.3772625,1.8749946,4.4818783,6.013564,2.584248,1.6146835,4.085753,4.678055,3.2746384,4.9421387,1.2525115,0.5772116,1.1393328,2.3088465,4.61392,5.138315,3.4179983,2.0145817,2.173032,3.8443048,3.3727267,2.3126192,1.8372684,2.2258487,2.8407867,6.013564,10.970794,11.174516,6.1908774,1.7014539,1.478869,1.3996439,2.0673985,3.500996,5.149633,4.3385186,4.214022,5.1798143,5.9720654,3.663219,2.5578396,2.384299,2.3163917,1.8523588,0.845068,1.5958204,1.3694628,0.8526133,0.49421388,0.49421388,0.4074435,1.8674494,2.003264,0.7092535,0.67152727,0.46026024,0.2678564,0.13204187,0.060362,0.02263575,0.018863125,0.0150905,0.033953626,0.08299775,0.181086,0.30181,0.3169005,0.26031113,0.211267,0.271629,0.41876137,0.33953625,0.24522063,0.211267,0.1961765,0.1358145,0.11317875,0.09808825,0.071679875,0.033953626,0.08677038,0.17731337,0.32444575,0.5017591,0.59607476,0.62625575,0.5998474,0.6526641,0.7997965,0.935611,0.5998474,0.33953625,0.26408374,0.41121614,0.7469798,0.9695646,0.7507524,0.4678055,0.31312788,0.28294688,0.4678055,0.5470306,0.5696664,0.5583485,0.5017591,0.31312788,0.19994913,0.16222288,0.19240387,0.29426476,0.1961765,0.12826926,0.094315626,0.10186087,0.14335975,0.15467763,0.14713238,0.116951376,0.090543,0.090543,0.07922512,0.06790725,0.06790725,0.08299775,0.120724,0.124496624,0.124496624,0.12826926,0.13204187,0.1056335,0.07922512,0.056589376,0.03772625,0.030181,0.033953626,0.030181,0.03772625,0.0452715,0.08299775,0.241448,0.5017591,0.69039035,0.6752999,0.4678055,0.19994913,0.35085413,0.27917424,0.18485862,0.181086,0.27917424,0.241448,0.23013012,0.3772625,0.7205714,1.20724,1.6146835,1.7391801,1.5316857,1.0525624,0.482896,0.5394854,1.1355602,1.4750963,1.5165952,2.0070364,2.2296214,2.0862615,2.3956168,3.2784111,4.1574326,4.7836885,3.9310753,3.029418,2.9086938,3.783943,4.568649,4.1989317,3.8292143,3.893349,4.0895257,4.357382,3.4859054,2.5804756,2.4220252,3.440634,4.9345937,6.2927384,6.790725,6.1833324,4.7006907,3.7348988,2.837014,2.1768045,1.8448136,1.8372684,2.3805263,2.2371666,1.9164935,1.8184053,2.2409391,2.2409391,1.9655377,1.539231,1.1506506,1.0487897,1.3392819,1.3694628,1.4260522,1.539231,1.4939595,1.5543215,1.7127718,1.7429527,1.5430037,1.1280149,0.7205714,0.4678055,0.3169005,0.2263575,0.15845025,0.1961765,0.23013012,0.29803738,0.41876137,0.56589377,0.49421388,0.44139713,0.41121614,0.422534,0.5319401,0.5885295,0.6375736,0.7092535,0.77338815,0.73188925,0.56589377,0.43007925,0.4074435,0.4979865,0.62248313,0.97710985,0.97710985,0.83752275,0.77716076,0.9922004,0.9808825,1.3505998,1.6410918,1.5430037,0.9016574,1.1506506,1.5052774,1.750498,1.8749946,2.0447628,1.9994912,1.8146327,1.4939595,1.1883769,1.1883769,1.0714256,0.9318384,0.95447415,1.1695137,1.4449154,1.478869,1.1619685,0.9620194,0.97710985,0.95824677,1.1204696,1.5241405,1.8787673,2.0183544,1.901403,2.2899833,2.7087448,2.6785638,2.1654868,1.5920477,3.2520027,5.6513925,9.137298,11.151879,6.217286,4.1574326,4.8327327,6.205968,6.5945487,4.6856003,2.746471,1.7693611,1.5467763,1.9240388,2.7879698,5.2250857,4.274384,2.4899325,1.4750963,1.8863125,2.795515,2.4974778,1.6222287,0.784706,0.6111652,0.69793564,0.7092535,0.8639311,1.388326,2.5276587,2.746471,2.1768045,1.2713746,0.47535074,0.21881226,0.11317875,0.06790725,0.0452715,0.030181,0.018863125,0.003772625,0.0,0.003772625,0.02263575,0.08677038,0.02263575,0.0150905,0.026408374,0.030181,0.00754525,0.0,0.00754525,0.011317875,0.011317875,0.00754525,0.049044125,0.03772625,0.02263575,0.018863125,0.011317875,0.003772625,0.003772625,0.011317875,0.0150905,0.0150905,0.16976812,0.21503963,0.33953625,0.52062225,0.482896,0.27917424,0.14335975,0.10186087,0.116951376,0.1056335,0.19994913,0.20749438,0.17354076,0.124496624,0.071679875,0.041498873,0.030181,0.02263575,0.018863125,0.011317875,0.02263575,0.018863125,0.00754525,0.011317875,0.049044125,0.071679875,0.09808825,0.12826926,0.1659955,0.19994913,1.1204696,2.5125682,3.4029078,3.229367,1.8448136,1.0072908,0.43007925,0.124496624,0.049044125,0.07922512,0.181086,0.24522063,0.22258487,0.13958712,0.14335975,0.2867195,0.44894236,0.754525,1.2713746,2.0296721,3.6066296,5.764571,8.360137,10.985884,12.996693,13.619176,14.871688,15.679029,14.796235,10.831206,8.8618965,9.0957985,9.416472,9.220296,9.4013815,9.382519,10.008774,10.103089,9.5032425,9.065618,8.484633,8.073418,7.7338815,7.1076255,5.5797124,4.6290107,4.5950575,5.040227,5.2552667,4.2706113,3.8443048,4.0291634,4.0895257,3.893349,3.8895764,3.5424948,3.5236318,4.142342,5.462761,7.3415284,9.623966,10.967021,11.781908,12.936331,15.758255,17.471025,17.829426,18.931032,21.798227,26.389511,32.89729,40.55949,47.467167,52.850704,57.08736,60.76567,62.327538,63.259377,63.014156,59.003857,61.463608,62.116272,61.6296,61.573013,64.41757,63.930904,64.52321,66.594376,70.16705,74.90547,75.95426,78.17634,80.398415,82.107414,83.44292,84.797295,84.84634,83.54855,81.85087,81.7226,83.175064,86.83828,91.225845,95.11165,97.533676,94.38353,93.221565,92.47081,91.92378,92.73867,92.38027,91.92378,91.618195,91.36543,90.70899,90.380775,90.22233,90.41096,90.81086,90.973076,91.84456,92.274635,92.46704,92.49345,92.26709,90.86745,89.49044,88.02666,86.555336,85.34055,85.291504,85.170784,86.18185,87.687126,87.215546,87.317406,87.166504,85.89513,83.53346,81.03599,79.08554,77.44444,75.475136,72.93993,70.012375,66.28125,63.157516,60.309185,57.396717,54.027763,52.3414,52.122585,51.439743,49.772243,48.01797,46.32029,44.58488,42.80043,41.2612,40.517994,40.26523,40.842438,42.211903,43.67568,43.86054,43.811493,46.17693,49.88542,52.914837,52.330082,50.406044,50.05896,49.78733,47.9727,42.8872,36.515236,32.527573,33.58768,40.12564,50.311726,48.927174,40.710396,32.286125,27.132719,25.551989,26.638506,24.601288,21.507734,18.659403,16.607096,14.977322,13.487134,12.743927,13.038192,14.317112,12.600568,9.903141,6.5643673,3.5990841,2.704972,2.04099,1.4637785,1.0374719,0.7997965,0.7582976,0.87147635,0.80356914,0.70170826,0.69039035,0.90920264,0.9280658,0.6149379,0.32821837,0.21503963,0.1961765,0.17731337,0.17354076,0.17354076,0.19994913,0.27917424,0.16976812,0.17354076,0.25276586,0.32067314,0.27917424,0.38858038,0.32444575,0.271629,0.34330887,0.5998474,0.663982,0.60362,0.4640329,0.32444575,0.31312788,0.4979865,0.62248313,0.663982,0.724344,1.026154,1.1204696,0.8224323,0.52439487,0.41876137,0.52062225,0.422534,0.29049212,0.271629,0.35085413,0.35839936,0.150905,0.11317875,0.17731337,0.24899325,0.211267,0.24899325,0.2867195,0.30935526,0.35462674,0.51684964,0.68661773,0.84884065,0.8903395,0.79602385,0.66775465,0.6375736,0.62248313,0.7997965,1.1355602,1.3770081,0.9922004,0.965792,1.1808317,1.3807807,1.1581959,1.4600059,1.8448136,1.961765,2.5012503,5.2099953,8.541223,8.967529,8.748717,10.480352,17.13149,16.98813,11.389555,6.0626082,4.0178456,5.5683947,12.875969,17.05981,17.037174,13.004238,6.40969,3.3764994,1.4411428,0.48666862,0.20372175,0.09808825,0.060362,0.033953626,0.033953626,0.05281675,0.06790725,0.06413463,0.13958712,0.06413463,0.049044125,0.094315626,0.0,0.018863125,1.0714256,1.4562333,0.84129536,0.26408374,1.4373702,1.5052774,0.965792,0.32444575,0.08677038,0.20749438,0.6111652,1.4449154,2.1843498,1.6410918,0.52439487,1.0186088,1.6184561,1.7052265,1.5580941,1.8976303,2.4408884,3.31991,4.08198,3.6934,1.1581959,0.482896,0.6149379,1.81086,5.6325293,6.043745,3.5047686,1.6825907,1.3996439,0.63002837,0.20372175,0.15467763,0.44516975,1.3920987,3.682082,5.594803,8.382772,8.073418,4.459243,1.1091517,1.6146835,3.0445085,5.349582,6.8058157,3.99521,2.746471,2.1994405,2.0447628,1.7429527,0.5394854,0.76584285,0.8299775,0.724344,0.663982,1.0525624,1.2449663,0.87147635,0.56589377,0.56212115,0.69039035,0.70170826,0.59607476,0.5055317,0.44894236,0.3470815,0.22258487,0.150905,0.10186087,0.060362,0.0150905,0.011317875,0.0150905,0.018863125,0.041498873,0.094315626,0.21503963,0.29049212,0.3055826,0.27540162,0.24899325,0.24899325,0.241448,0.26408374,0.28294688,0.21503963,0.19240387,0.181086,0.14713238,0.10186087,0.06790725,0.090543,0.18485862,0.27917424,0.34330887,0.38480774,0.6149379,0.80734175,0.91297525,0.9242931,0.8903395,0.9318384,0.66775465,0.422534,0.362172,0.482896,0.7884786,0.69039035,0.56212115,0.52062225,0.452715,0.58098423,0.6187105,0.6790725,0.784706,0.8526133,0.573439,0.35839936,0.23767537,0.21881226,0.27540162,0.24899325,0.18863125,0.13204187,0.10186087,0.10940613,0.120724,0.1358145,0.1358145,0.120724,0.1056335,0.12826926,0.10186087,0.08299775,0.090543,0.1056335,0.11317875,0.124496624,0.1358145,0.14335975,0.1358145,0.116951376,0.08677038,0.056589376,0.030181,0.0150905,0.003772625,0.00754525,0.030181,0.06790725,0.14713238,0.2565385,0.30181,0.2678564,0.18863125,0.15845025,0.17731337,0.1358145,0.150905,0.24522063,0.34330887,0.23390275,0.19240387,0.271629,0.6111652,1.4411428,2.1315331,2.335255,2.082489,1.4600059,0.6413463,0.8563859,1.0601076,1.2223305,1.4071891,1.7580433,2.4031622,2.8181508,2.8332415,2.8445592,3.8065786,3.8405323,3.712263,3.4066803,3.1954134,3.6292653,4.0517993,3.5387223,3.0633714,2.9615107,2.957738,2.2484846,2.233394,2.3805263,2.5691576,3.0633714,5.4363527,7.1868505,7.2170315,5.6476197,3.8103511,3.0746894,2.6483827,2.565385,2.8219235,3.3915899,3.5575855,2.4069347,1.7052265,2.1390784,3.3236825,3.5047686,2.848332,2.033445,1.4713237,1.3053282,1.539231,1.6524098,1.7769064,1.8146327,1.4298248,1.2789198,1.3920987,1.2940104,0.935611,0.6790725,0.5357128,0.44894236,0.3772625,0.33576363,0.35839936,0.4678055,0.44894236,0.452715,0.5696664,0.814887,0.56212115,0.48666862,0.5055317,0.5696664,0.66775465,0.724344,0.66775465,0.5696664,0.46026024,0.3470815,0.29049212,0.31312788,0.38480774,0.482896,0.59230214,0.935611,0.73566186,0.55457586,0.59230214,0.694163,0.7997965,1.7618159,2.6106565,2.6672459,1.5505489,1.5882751,1.5920477,1.5015048,1.3807807,1.448688,1.4147344,1.1846043,0.98465514,0.9242931,0.9997456,1.1053791,1.1016065,1.0601076,1.0751982,1.2751472,2.0145817,2.1164427,1.7542707,1.2864652,1.2638294,1.7957695,2.0372176,2.0296721,1.9051756,1.8825399,2.6219745,3.0445085,2.7313805,1.8259505,1.0714256,1.2600567,2.7728794,8.477088,14.781145,11.619685,6.9227667,5.3910813,5.0138187,4.9119577,5.3571277,4.8666863,3.9008942,3.4557245,3.7009451,3.9461658,5.379763,3.731126,1.8221779,1.0487897,1.4147344,2.233394,1.871222,1.1657411,0.6149379,0.3734899,0.4376245,0.6073926,0.7469798,0.875249,1.1657411,0.84884065,0.5017591,0.2565385,0.14713238,0.0754525,0.030181,0.0150905,0.02263575,0.033953626,0.00754525,0.003772625,0.0,0.0,0.003772625,0.02263575,0.018863125,0.00754525,0.0150905,0.033953626,0.011317875,0.003772625,0.0150905,0.026408374,0.026408374,0.0150905,0.0150905,0.0150905,0.026408374,0.03772625,0.02263575,0.003772625,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.00754525,0.011317875,0.011317875,0.011317875,0.003772625,0.00754525,0.026408374,0.0452715,0.06413463,0.150905,0.08299775,0.030181,0.0452715,0.05281675,0.041498873,0.02263575,0.02263575,0.033953626,0.026408374,0.018863125,0.0150905,0.011317875,0.011317875,0.026408374,0.033953626,0.03772625,0.03772625,0.07922512,0.27917424,1.6448646,3.8782585,5.5382137,5.304311,2.0183544,0.55457586,0.11317875,0.05281675,0.0452715,0.060362,0.19994913,0.26408374,0.21503963,0.116951376,0.1358145,0.20749438,0.3470815,0.60362,1.0035182,1.5618668,2.4522061,3.663219,6.4247804,10.70671,15.196134,14.02662,12.264804,11.59705,11.766817,10.555805,9.986138,11.102836,12.472299,12.989148,11.887542,12.792972,14.524607,15.245177,14.385019,12.6345215,9.205205,7.707473,8.424272,9.918231,9.031664,6.7454534,6.1908774,6.790725,7.3981175,6.304056,5.251494,4.8100967,4.6629643,4.6629643,4.8402777,4.1008434,3.832987,3.7952607,4.134797,5.402399,7.0812173,8.45068,9.884277,11.627231,13.815352,14.290704,13.864397,14.596286,17.006994,20.059048,24.60506,29.581152,34.10453,37.907337,41.33288,44.747105,46.788094,48.183968,48.742313,47.365307,47.76898,48.19906,48.399006,48.49332,48.99885,45.04137,44.773514,46.369335,49.334618,54.51443,58.27951,61.456062,64.80992,68.44296,71.78551,74.43012,75.87881,76.80687,77.63685,78.54228,73.98118,74.47162,77.82548,81.49625,82.56767,82.11873,82.39036,82.68839,82.80534,82.98266,82.97511,83.50706,84.77466,86.19694,86.3818,86.11394,85.7744,85.272644,84.87274,85.185875,86.725105,87.76257,88.81514,90.075195,91.410706,90.39964,89.63757,89.07168,88.79627,89.011314,91.10512,93.23288,95.90767,98.82014,100.86113,102.74367,103.28693,102.000465,99.4049,97.00928,95.93408,95.95672,96.27739,96.266075,95.488914,90.48641,85.963036,81.68865,77.44444,73.04934,69.83506,67.01314,63.515915,59.59993,56.845913,55.121822,52.90729,50.817257,49.225212,48.25942,46.769234,45.76194,45.95812,47.120087,48.07079,49.142212,50.839893,52.51494,53.556183,53.412827,53.11856,53.522232,53.699543,52.64698,49.300663,42.894745,39.646515,40.683987,44.486794,46.856003,41.10275,35.34195,31.15811,29.034122,28.35505,30.62617,29.44911,27.14781,25.046457,23.48459,21.636003,19.794964,19.647831,21.277605,23.163918,18.946123,14.883006,10.344538,6.1531515,4.5761943,3.6066296,2.7351532,1.9957186,1.4713237,1.2713746,1.2298758,1.1053791,0.97710985,0.995973,1.3694628,1.2600567,1.0110635,0.7507524,0.5394854,0.34330887,0.241448,0.18863125,0.1961765,0.23013012,0.20372175,0.1961765,0.25276586,0.29049212,0.30181,0.34330887,0.6073926,0.58098423,0.45648763,0.40367088,0.55080324,0.3470815,0.33576363,0.39989826,0.44516975,0.41121614,0.58475685,0.58475685,0.44516975,0.3055826,0.44516975,0.43385187,0.32067314,0.19994913,0.120724,0.11317875,0.21881226,0.1358145,0.08677038,0.124496624,0.13958712,0.06413463,0.03772625,0.06790725,0.13958712,0.21881226,0.20372175,0.241448,0.2263575,0.17354076,0.23013012,0.30935526,0.35085413,0.52062225,0.84129536,1.1996948,1.056335,1.177059,1.5580941,2.0296721,2.2598023,2.203213,2.474842,2.8181508,2.9011486,2.3088465,3.1048703,3.8065786,3.6292653,3.3915899,5.50426,7.4396167,8.028146,7.360391,7.54525,12.706201,14.434063,9.57115,4.8968673,3.2444575,3.5424948,6.398372,6.3342376,4.587512,2.4597516,1.3355093,0.8526133,0.5055317,0.29049212,0.17354076,0.10186087,0.06790725,0.033953626,0.02263575,0.026408374,0.026408374,0.0150905,0.003772625,0.0,0.23767537,0.47535074,0.0,0.0,0.0,0.116951376,0.30181,0.35085413,0.59607476,0.63002837,0.422534,0.19994913,0.44139713,0.88279426,0.41498876,0.43385187,1.5580941,3.6330378,1.4222796,0.41121614,0.20372175,0.422534,0.7167987,1.2902378,1.8448136,2.1654868,2.2899833,2.5314314,1.2864652,1.1317875,0.91297525,0.51684964,0.87147635,0.784706,0.34330887,0.041498873,0.02263575,0.0452715,0.33953625,0.38480774,0.27540162,0.25276586,0.7167987,1.0487897,3.2633207,4.3007927,3.3425457,1.8146327,4.014073,7.5565677,8.831716,6.802043,3.006782,2.2862108,1.9127209,1.3015556,0.5281675,0.32067314,0.62625575,1.0223814,0.9922004,0.68661773,0.9318384,0.90543,0.845068,0.73566186,0.6413463,0.70170826,0.6149379,0.49421388,0.3734899,0.26408374,0.150905,0.1056335,0.08299775,0.06413463,0.041498873,0.0150905,0.003772625,0.00754525,0.0150905,0.02263575,0.0452715,0.1659955,0.29803738,0.3734899,0.35839936,0.27540162,0.27540162,0.27540162,0.3734899,0.45648763,0.21503963,0.26408374,0.26408374,0.23013012,0.1659955,0.090543,0.116951376,0.18485862,0.21503963,0.21503963,0.27540162,0.543258,0.8563859,1.1317875,1.3166461,1.4034165,1.7580433,1.5731846,1.1808317,0.83752275,0.70170826,0.663982,0.56589377,0.724344,1.0751982,1.1581959,0.97710985,0.694163,0.5093044,0.52062225,0.7167987,0.694163,0.55080324,0.41498876,0.33576363,0.27540162,0.2867195,0.21503963,0.150905,0.120724,0.120724,0.120724,0.150905,0.17354076,0.181086,0.1659955,0.181086,0.1659955,0.14713238,0.14335975,0.1659955,0.15467763,0.16222288,0.17354076,0.18485862,0.19994913,0.18485862,0.14713238,0.090543,0.041498873,0.0150905,0.003772625,0.00754525,0.033953626,0.09808825,0.24522063,0.40367088,0.48666862,0.4376245,0.29426476,0.18485862,0.1358145,0.18485862,0.28294688,0.392353,0.5017591,0.38103512,0.3961256,0.5017591,0.7205714,1.1581959,1.4411428,1.7127718,1.991946,2.1051247,1.6788181,2.2748928,2.7540162,2.9803739,2.806833,2.0749438,1.7957695,3.0143273,3.5764484,3.2331395,3.6481283,2.463524,2.4522061,3.048281,3.531177,3.006782,2.969056,2.584248,2.4672968,2.5540671,2.0900342,2.003264,1.5543215,1.3015556,1.5882751,2.5012503,4.798779,6.7152724,7.0887623,5.934339,4.45547,3.1727777,3.4481792,4.1272516,4.859141,6.1041074,5.323174,3.6971724,2.5767028,2.5314314,3.3727267,3.7499893,3.3312278,2.5201135,1.6863633,1.1581959,1.2449663,1.2487389,1.2411937,1.1883769,0.9318384,1.0035182,0.84884065,0.6828451,0.63002837,0.7167987,0.9242931,0.8941121,0.7469798,0.6375736,0.7469798,0.724344,0.6149379,0.4376245,0.29049212,0.35085413,0.31312788,0.241448,0.27917424,0.4376245,0.59607476,0.58475685,0.56212115,0.52439487,0.482896,0.45648763,0.52062225,0.5998474,0.56589377,0.482896,0.58098423,0.87147635,0.5998474,0.32444575,0.32821837,0.6111652,0.73188925,1.6410918,2.8332415,3.380272,1.9542197,0.87902164,0.5470306,0.4678055,0.4376245,0.5357128,0.4979865,0.41498876,0.3169005,0.3055826,0.55080324,1.1091517,1.5882751,1.8448136,1.9353566,2.1051247,3.410453,3.5462675,2.7540162,1.7391801,1.6788181,2.3390274,2.0258996,1.7467253,1.7731338,1.6637276,2.7125173,3.1576872,2.5804756,1.3770081,0.77716076,0.8865669,2.2447119,5.5268955,9.224068,9.627739,7.1981683,4.878004,3.3727267,3.2105038,4.7610526,8.360137,8.29223,7.937603,8.107371,7.0359454,6.092789,4.5120597,2.7691069,1.3317367,0.67152727,0.9393836,0.77716076,0.8941121,1.1431054,0.52062225,0.543258,0.7054809,0.6488915,0.35839936,0.150905,0.17731337,0.3734899,0.48666862,0.4074435,0.19994913,0.06413463,0.011317875,0.056589376,0.120724,0.0452715,0.02263575,0.00754525,0.0,0.0,0.0,0.011317875,0.00754525,0.00754525,0.011317875,0.0,0.0,0.0,0.011317875,0.026408374,0.0150905,0.0150905,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.0150905,0.00754525,0.011317875,0.026408374,0.0150905,0.003772625,0.0,0.0,0.003772625,0.0150905,0.026408374,0.02263575,0.02263575,0.026408374,0.0150905,0.041498873,0.03772625,0.02263575,0.02263575,0.0452715,0.6790725,1.0789708,1.6939086,2.0673985,0.80734175,0.23390275,0.10940613,0.10940613,0.08677038,0.060362,0.120724,0.1358145,0.11317875,0.0754525,0.0754525,0.17354076,0.34330887,0.62625575,1.026154,1.5241405,2.0749438,2.6710186,4.2517486,7.2623034,11.642321,9.175024,8.303548,8.975075,10.544487,11.763044,12.193124,13.65313,14.928277,14.864142,12.37421,15.339493,20.496672,23.563816,22.496162,17.455936,13.732355,10.567122,9.171251,9.201432,8.7751255,6.330465,5.704209,6.379509,7.564113,8.14887,7.865923,7.413208,6.6662283,5.7079816,4.7912335,3.92353,3.5877664,3.270866,3.0709167,3.6934,4.2781568,5.111907,6.462507,8.054554,9.0807085,9.495697,10.982111,12.864652,15.079182,18.142553,21.636003,25.729303,29.867872,33.71595,37.171673,39.88042,41.163113,41.883682,42.276035,41.94782,40.67644,41.283836,42.574074,43.57759,43.581364,39.22021,37.492348,37.216946,37.58289,38.133694,38.937263,40.28409,42.287354,44.735786,47.089905,47.433212,49.21012,52.526257,57.46085,64.089355,60.814716,58.99254,60.67513,64.91556,67.73371,67.06218,67.00559,67.80539,69.333305,71.09135,69.895424,69.87279,70.57827,71.68365,72.955025,74.309395,75.04128,75.071465,74.75079,74.8602,75.8109,77.04077,78.88936,81.35288,84.06163,86.34407,88.41524,90.38832,92.4029,94.65139,97.993935,100.74418,104.07163,107.92725,111.05099,112.420456,112.23182,110.07765,106.384254,102.41545,98.30329,98.5636,101.038445,103.77737,105.07138,102.47204,98.89936,94.658936,89.871475,84.48794,80.23996,76.878555,73.60014,70.197235,67.06218,63.776226,61.127842,58.78127,56.68369,55.023735,53.62032,52.26972,50.99457,50.33059,51.330338,52.345173,53.19024,54.936966,57.18545,58.07579,55.48777,51.515194,48.56123,47.618073,48.26319,47.040863,47.029545,48.787586,50.055187,45.74685,38.065784,34.08944,32.750156,32.516254,31.358059,30.599762,30.675215,30.59599,30.256453,30.44131,30.818573,30.218727,31.512737,33.712177,31.965452,22.688566,17.697384,13.313594,8.91094,6.8963585,5.1156793,4.2027044,3.3727267,2.4672968,1.9542197,1.659955,1.6410918,1.539231,1.4562333,1.9693103,1.6637276,1.4600059,1.3430545,1.1732863,0.68661773,0.41876137,0.2867195,0.2263575,0.20372175,0.23013012,0.29049212,0.4074435,0.38103512,0.23390275,0.19994913,0.29426476,0.4376245,0.5055317,0.45648763,0.32067314,0.271629,0.27917424,0.32821837,0.422534,0.59607476,0.38858038,0.41876137,0.31312788,0.1056335,0.21503963,0.150905,0.10940613,0.07922512,0.05281675,0.0150905,0.0150905,0.0150905,0.026408374,0.041498873,0.030181,0.030181,0.049044125,0.056589376,0.071679875,0.18485862,0.2565385,0.40367088,0.3470815,0.13204187,0.1056335,0.120724,0.1961765,0.52439487,1.0789708,1.6033657,1.5656394,2.2069857,3.0105548,3.6971724,4.2102494,5.50426,6.0776987,6.375736,6.349328,5.4476705,5.9003854,6.149379,5.4665337,4.478106,5.1873593,7.3377557,10.774617,11.276376,9.06939,8.850578,10.646348,7.5603404,4.508287,3.1048703,1.6637276,1.3845534,1.2411937,1.0186088,0.663982,0.27540162,0.19994913,0.14713238,0.116951376,0.10186087,0.0754525,0.05281675,0.03772625,0.02263575,0.0150905,0.0150905,0.041498873,0.116951376,0.05281675,0.049044125,0.094315626,0.0,0.0,0.0,0.02263575,0.060362,0.071679875,0.23767537,1.8825399,1.8070874,0.452715,1.9089483,4.0178456,2.0485353,0.6413463,1.3996439,2.897376,1.599593,1.1280149,0.90920264,0.6752999,0.5093044,1.0450171,1.7014539,1.8599042,1.5354583,1.3619176,1.9730829,1.6561824,0.98842776,0.40367088,0.211267,0.30935526,0.2867195,0.33576363,0.60362,1.20724,2.4371157,3.029418,2.5125682,2.8143783,8.296002,2.7389257,1.7844516,2.0447628,2.04099,2.1956677,2.9766011,4.6629643,4.776143,3.0218725,1.2864652,1.7769064,1.8599042,1.2826926,0.43007925,0.32067314,0.7997965,1.2713746,1.3128735,0.9922004,0.845068,1.1242423,1.0487897,0.7997965,0.55457586,0.5055317,0.47157812,0.38103512,0.271629,0.15845025,0.07922512,0.060362,0.03772625,0.018863125,0.00754525,0.003772625,0.011317875,0.00754525,0.003772625,0.011317875,0.0452715,0.10940613,0.18863125,0.271629,0.34330887,0.38480774,0.3055826,0.23013012,0.18485862,0.17731337,0.17731337,0.26408374,0.35085413,0.3772625,0.3470815,0.31312788,0.3055826,0.25276586,0.22258487,0.26031113,0.35839936,0.47157812,1.1053791,1.5807298,1.720317,1.8448136,1.8448136,1.7618159,1.5279131,1.297783,1.4449154,1.9089483,1.961765,1.8523588,1.7882242,1.9542197,2.6597006,1.931584,1.086516,0.70170826,0.59607476,0.68661773,0.66020936,0.6111652,0.573439,0.543258,0.45648763,0.32067314,0.2263575,0.20372175,0.1961765,0.17731337,0.14713238,0.124496624,0.116951376,0.14335975,0.116951376,0.12826926,0.14713238,0.16222288,0.15467763,0.13204187,0.12826926,0.14713238,0.17354076,0.18485862,0.19240387,0.2263575,0.18485862,0.07922512,0.0150905,0.011317875,0.00754525,0.03772625,0.116951376,0.24522063,0.35462674,0.5583485,0.67152727,0.6073926,0.392353,0.36971724,0.33576363,0.482896,0.69793564,0.55080324,0.39989826,0.35839936,0.38480774,0.47912338,0.694163,0.97710985,1.2261031,1.6373192,2.1994405,2.6785638,2.9049213,2.5616124,2.2786655,2.2673476,2.3088465,3.2557755,4.0593443,4.195159,3.7877154,3.5990841,2.384299,2.4974778,2.5238862,2.0673985,1.7354075,2.071171,1.448688,1.1393328,1.4750963,1.871222,2.1466236,1.7429527,1.6373192,2.1466236,2.916239,4.0216184,5.4212623,5.753253,4.749735,3.2821836,2.8219235,4.5460134,6.187105,6.934085,7.4471617,5.4250345,3.8707132,2.806833,2.335255,2.6408374,2.704972,2.3503454,1.9466745,1.6939086,1.599593,1.5467763,1.20724,0.84129536,0.5772116,0.41876137,0.6073926,0.68661773,0.73566186,0.7696155,0.7167987,0.67152727,0.5394854,0.48666862,0.573439,0.77338815,0.5017591,0.271629,0.120724,0.071679875,0.094315626,0.116951376,0.08677038,0.124496624,0.29049212,0.59607476,0.59230214,0.58098423,0.5696664,0.5357128,0.43385187,0.4376245,0.42630664,0.33953625,0.23390275,0.31312788,0.91674787,0.9242931,1.0789708,1.3392819,0.86770374,0.95824677,0.90920264,0.9242931,0.9393836,0.62248313,0.38858038,0.38103512,0.44894236,0.4678055,0.35085413,0.44139713,0.48666862,0.41121614,0.35462674,0.66020936,1.1129243,1.1053791,1.0714256,1.146878,1.1544232,1.9730829,2.3277097,2.191895,1.7731338,1.50905,1.6788181,1.7429527,1.5618668,1.3091009,1.4939595,2.8822856,3.1237335,2.372981,1.2185578,0.6790725,0.6828451,1.3656902,2.384299,3.3161373,3.6707642,3.5160866,3.2670932,2.776652,2.5238862,3.6141748,6.7341356,6.3908267,5.0968165,4.221567,4.006528,3.338773,2.897376,2.2484846,1.4222796,0.8903395,1.1996948,1.8523588,2.806833,3.270866,1.690136,1.5279131,1.7919968,1.3732355,0.392353,0.1659955,0.29803738,0.5357128,0.70170826,0.65643674,0.331991,0.10940613,0.13958712,0.29426476,0.362172,0.0452715,0.02263575,0.0150905,0.018863125,0.02263575,0.011317875,0.02263575,0.018863125,0.018863125,0.02263575,0.011317875,0.003772625,0.0,0.00754525,0.026408374,0.06413463,0.026408374,0.0150905,0.011317875,0.003772625,0.0,0.011317875,0.018863125,0.0150905,0.003772625,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.00754525,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.011317875,0.003772625,0.003772625,0.018863125,0.026408374,0.030181,0.026408374,0.02263575,0.13958712,0.21503963,0.33953625,0.41498876,0.16222288,0.056589376,0.049044125,0.09808825,0.14335975,0.10940613,0.26031113,0.55080324,0.7809334,0.7582976,0.30935526,0.19240387,0.24899325,0.49044126,0.9393836,1.6373192,2.233394,2.8634224,4.4177437,6.670001,8.262049,7.2887115,7.149124,7.9526935,9.424017,10.899114,12.14408,13.788944,16.248695,18.806536,19.625195,19.693102,20.847527,23.993895,27.600525,27.698612,23.288414,17.37671,13.045737,11.446144,11.7894535,8.993938,6.779407,5.9305663,6.2927384,6.7341356,6.9491754,7.1679873,6.8699503,5.881522,4.3875628,3.3350005,2.6672459,2.335255,2.3201644,2.6295197,3.2935016,3.6556737,4.0593443,4.485651,4.561104,5.7607985,7.696155,9.778644,12.385528,16.886269,21.881226,26.265015,29.875418,32.776566,35.2665,35.534355,35.24009,35.017506,35.15332,35.587173,34.719467,34.772285,34.95337,34.900555,34.704376,30.875162,30.69785,31.799456,32.61057,32.357803,31.599506,31.320333,31.671186,32.648296,34.07812,34.926964,36.149292,39.156075,44.000126,49.37989,52.20936,50.715397,49.244076,49.04035,48.278282,47.53885,49.41007,52.18672,54.71061,56.38188,56.64974,56.676144,57.355217,58.856724,60.62231,62.135136,63.25183,63.968628,64.685425,66.17939,67.95252,69.37857,71.11398,73.51714,76.625786,80.8134,85.42732,89.34708,92.7198,96.95646,99.50298,103.02284,106.04849,108.21775,110.29646,111.205666,111.933784,112.035645,111.341484,109.9607,108.52333,107.938576,107.4255,106.42575,104.59603,102.33623,100.581955,98.72205,96.318886,93.09329,88.23792,83.563644,78.94218,74.64139,71.31016,68.65046,66.205795,64.210075,62.723663,61.652237,60.414818,59.02649,57.87584,57.083588,56.47997,56.087616,56.19702,57.47594,59.309437,59.81874,56.84214,52.160313,48.482002,47.13895,48.082108,49.59493,52.382896,56.744053,60.128098,57.147724,48.30469,40.55949,36.292652,35.258953,34.56856,34.960915,35.07032,34.46293,33.96117,35.62867,35.764484,33.68577,32.95388,33.267006,30.463947,24.17498,21.036158,16.81459,11.193378,7.7640624,6.5266414,5.4665337,4.5309224,3.712263,3.0633714,2.6144292,2.354118,2.1692593,2.0900342,2.2598023,2.093807,1.9655377,1.961765,1.8825399,1.2487389,0.9695646,0.7469798,0.56212115,0.41121614,0.32821837,0.36971724,0.45648763,0.5055317,0.45648763,0.271629,0.26031113,0.28294688,0.3055826,0.30935526,0.28294688,0.25276586,0.30935526,0.32444575,0.29426476,0.33953625,0.2678564,0.22258487,0.23013012,0.271629,0.26408374,0.13204187,0.071679875,0.041498873,0.018863125,0.003772625,0.003772625,0.003772625,0.003772625,0.00754525,0.00754525,0.0150905,0.05281675,0.06790725,0.071679875,0.120724,0.41876137,0.5696664,0.5357128,0.41121614,0.4376245,0.633801,0.66775465,0.6413463,0.663982,0.8563859,1.0638802,1.7580433,2.9011486,4.870459,8.458225,9.910686,9.9257765,10.457717,11.144334,9.291975,6.7077274,6.360646,7.6320205,9.390063,9.971047,12.2270775,14.596286,16.595778,16.21097,9.88805,10.616167,7.1868505,4.4818783,3.874486,3.2255943,1.7618159,1.0902886,0.7394345,0.4640329,0.23767537,0.1358145,0.071679875,0.041498873,0.033953626,0.041498873,0.026408374,0.018863125,0.018863125,0.0150905,0.0150905,0.018863125,0.056589376,0.026408374,0.003772625,0.00754525,0.0,0.00754525,0.003772625,0.003772625,0.02263575,0.071679875,1.7354075,2.1315331,1.3505998,0.39989826,1.2110126,2.384299,1.3166461,0.4074435,0.8337501,2.5314314,1.1280149,0.62248313,0.4376245,0.29803738,0.19240387,0.513077,0.965792,1.0940613,0.83752275,0.5281675,1.0902886,1.871222,1.9542197,1.3996439,1.2449663,1.7655885,2.093807,3.180323,3.942393,1.267602,2.2786655,2.214531,1.9466745,2.727608,6.1908774,2.867195,1.9391292,2.0975795,2.4295704,2.4182527,2.7992878,2.595566,1.9089483,1.4713237,2.6408374,1.2147852,0.8639311,0.62625575,0.24899325,0.19994913,0.45648763,0.95824677,1.2751472,1.2034674,0.7582976,0.80734175,0.68661773,0.48666862,0.31312788,0.29426476,0.32821837,0.2678564,0.17731337,0.094315626,0.041498873,0.02263575,0.011317875,0.003772625,0.0,0.0,0.003772625,0.003772625,0.003772625,0.011317875,0.026408374,0.05281675,0.094315626,0.19240387,0.35462674,0.5319401,0.5281675,0.4376245,0.38480774,0.36971724,0.27917424,0.35462674,0.59230214,0.7922512,0.9318384,1.1732863,0.845068,1.026154,0.86770374,0.4640329,0.86770374,1.1393328,1.7655885,2.003264,1.7919968,1.7429527,1.2336484,1.4637785,1.841041,2.1692593,2.6672459,4.08198,3.6481283,3.1237335,2.9916916,2.4710693,2.6031113,2.3088465,1.9768555,1.7693611,1.6373192,1.3241913,0.97333723,0.76584285,0.73188925,0.72811663,0.5696664,0.39989826,0.29803738,0.2678564,0.23013012,0.19994913,0.17731337,0.16222288,0.14713238,0.120724,0.13204187,0.15467763,0.15845025,0.14713238,0.14335975,0.120724,0.124496624,0.15467763,0.18863125,0.19994913,0.24899325,0.31312788,0.32821837,0.24899325,0.05281675,0.02263575,0.011317875,0.06790725,0.20372175,0.39989826,0.97333723,1.0487897,0.8111144,0.543258,0.6073926,0.63002837,0.5017591,0.56589377,0.784706,0.70170826,0.7054809,0.56589377,0.44139713,0.40367088,0.452715,1.0035182,1.7014539,2.1654868,2.3088465,2.3428001,2.0673985,1.7957695,1.6637276,1.7919968,2.3013012,2.8558772,3.9876647,4.9421387,5.1081343,4.025391,3.470815,3.380272,2.9728284,2.1994405,1.7580433,2.6332922,2.8709676,2.938875,2.8898308,2.354118,3.0897799,2.565385,2.2598023,2.5804756,2.867195,3.4670424,4.5497856,5.1835866,4.870459,3.5575855,3.7047176,5.2062225,6.677546,7.3075747,6.8661776,4.9534564,3.9348478,3.4745877,3.3010468,3.218049,2.4861598,2.0598533,1.7467253,1.5015048,1.4335974,1.2826926,1.0902886,0.88279426,0.73566186,0.7582976,0.7922512,0.7432071,0.754525,0.8563859,0.94692886,0.6451189,0.44139713,0.51684964,0.8639311,1.2826926,0.9507015,0.59230214,0.3470815,0.241448,0.18485862,0.24522063,0.16976812,0.1961765,0.3772625,0.58475685,0.5696664,0.41498876,0.3055826,0.28294688,0.23390275,0.19994913,0.20372175,0.18863125,0.23390275,0.56589377,0.9242931,1.0638802,1.0676528,0.94692886,0.5998474,0.55457586,0.41876137,0.34330887,0.3470815,0.3169005,0.44516975,0.56212115,0.73188925,0.845068,0.6149379,0.35085413,0.27540162,0.36971724,0.52062225,0.52062225,0.5885295,0.55457586,0.52439487,0.56589377,0.7130261,1.4335974,1.6448646,1.5128226,1.2826926,1.3091009,1.5543215,1.7089992,1.5543215,1.2638294,1.3958713,2.1541688,2.1654868,1.6222287,0.9318384,0.72811663,0.6828451,0.80356914,0.95447415,1.1544232,1.569412,2.4522061,2.6182017,2.1881225,1.6222287,1.7354075,3.059599,2.8936033,2.1881225,1.6637276,1.7957695,1.4524606,1.4071891,1.3543724,1.1506506,0.8186596,0.7997965,1.0940613,1.5052774,1.6184561,0.8111144,0.73566186,0.86770374,0.69793564,0.24899325,0.0754525,0.13958712,0.24522063,0.331991,0.331991,0.17354076,0.05281675,1.2223305,2.003264,1.6373192,0.29426476,0.071679875,0.0150905,0.0150905,0.011317875,0.00754525,0.056589376,0.030181,0.00754525,0.0150905,0.02263575,0.003772625,0.0,0.003772625,0.0150905,0.049044125,0.030181,0.018863125,0.011317875,0.00754525,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.00754525,0.0,0.003772625,0.011317875,0.0150905,0.018863125,0.00754525,0.0,0.0,0.011317875,0.033953626,0.056589376,0.05281675,0.05281675,0.08677038,0.13958712,0.1659955,0.3961256,0.8865669,1.7693611,2.2220762,0.43007925,0.23767537,0.2678564,0.5093044,1.0110635,1.8749946,2.837014,3.6481283,4.979865,6.7643166,8.213005,8.367682,8.688355,9.514561,10.812344,12.174261,13.905896,15.033911,16.87118,19.40261,21.300241,20.919205,19.979822,20.564579,22.90738,25.404858,23.069601,18.417955,14.418973,12.706201,13.585222,11.5857315,9.039209,7.3377557,6.677546,6.0776987,5.9418845,5.8136153,5.4438977,4.7572803,3.8858037,3.1312788,2.3654358,1.8221779,1.6109109,1.7240896,1.9844007,2.3692086,2.674791,2.8785129,3.1237335,4.06689,5.873977,7.888559,10.197406,13.649357,15.931795,17.855835,19.73083,21.492645,22.696112,22.956423,23.118647,23.593996,24.435291,25.325632,26.461191,27.29494,27.434528,27.140265,27.30626,27.185535,28.177736,29.03035,29.354795,29.615107,29.581152,30.486582,30.71294,30.256453,30.750666,31.776821,31.97677,32.621887,34.006443,35.45513,37.15658,36.454876,35.47399,34.632698,32.62566,33.289642,35.590942,37.779068,39.197575,40.291634,41.461147,41.902546,41.977997,41.974224,42.11381,43.05697,44.06803,44.818787,45.49031,46.754143,49.2818,51.98677,54.921875,58.20406,62.01441,66.85469,72.8343,78.84409,84.63507,90.80708,95.692635,100.989395,105.44487,108.704414,111.307526,113.53715,115.604546,117.472,118.95841,119.75821,120.39955,120.188286,119.40358,118.162384,116.415665,114.22754,111.91115,109.749435,107.51227,104.45644,99.97079,95.07392,90.11669,85.34055,80.86622,77.13509,73.396416,70.080284,67.38663,65.28528,64.00259,62.83307,61.91632,61.203297,60.49027,60.411045,60.324272,60.660038,61.101433,60.577038,57.845657,55.551903,54.26921,54.020218,54.288074,54.865284,56.619556,58.43796,58.419098,53.88063,47.569027,41.977997,38.175194,36.258698,35.36836,35.25518,35.79844,35.538128,34.549698,34.428974,35.15332,33.06706,31.558008,30.773302,27.63825,24.190071,22.371666,19.025349,13.924759,9.767326,8.29223,6.930312,5.87775,5.1647234,4.6516466,4.134797,3.7952607,3.5802212,3.4557245,3.4330888,3.4444065,3.199186,2.9954643,2.8143783,2.3126192,1.9240388,1.50905,1.1846043,0.94315624,0.633801,0.51684964,0.44516975,0.44894236,0.45648763,0.30935526,0.241448,0.20749438,0.2263575,0.27540162,0.31312788,0.36594462,0.38858038,0.3470815,0.26408374,0.211267,0.29049212,0.271629,0.2867195,0.35839936,0.40367088,0.23390275,0.116951376,0.041498873,0.003772625,0.0,0.02263575,0.026408374,0.0150905,0.0,0.0,0.003772625,0.03772625,0.11317875,0.16976812,0.060362,0.1961765,0.34330887,0.362172,0.31312788,0.4376245,0.6375736,0.65643674,0.6413463,0.6149379,0.46026024,0.7092535,1.3392819,2.3956168,4.3724723,8.201687,10.533169,10.627484,11.042474,11.996947,11.378237,8.83926,9.0957985,11.989402,15.456445,15.497944,13.63804,12.095036,12.713746,13.600313,9.148616,6.888813,4.3913355,7.1566696,12.102581,7.5716586,3.4972234,2.0447628,1.267602,0.47535074,0.211267,0.12826926,0.056589376,0.018863125,0.0150905,0.02263575,0.0150905,0.0150905,0.0150905,0.0150905,0.00754525,0.00754525,0.00754525,0.060362,0.241448,0.36594462,0.00754525,0.03772625,0.10186087,0.14335975,0.14335975,0.10940613,1.7919968,1.7278622,0.9997456,0.44516975,0.66775465,1.629774,0.90543,0.17731337,0.43385187,1.9655377,0.7582976,0.29803738,0.116951376,0.0,0.00754525,0.120724,0.30181,0.38103512,0.29803738,0.10186087,0.241448,2.3767538,3.5953116,3.1652324,2.516341,2.4522061,2.9086938,4.002755,4.5497856,2.0485353,2.7653341,2.5804756,2.4182527,2.546522,2.5729303,1.9391292,2.2183034,2.3767538,2.0636258,1.6410918,1.8070874,1.1242423,0.7130261,1.2600567,3.0369632,0.8262049,0.25276586,0.2263575,0.19994913,0.16976812,0.19994913,0.6111652,1.0035182,1.0714256,0.5998474,0.422534,0.29049212,0.18863125,0.13204187,0.150905,0.19994913,0.16222288,0.094315626,0.0452715,0.018863125,0.003772625,0.0,0.0,0.018863125,0.09808825,0.120724,0.10186087,0.0754525,0.08677038,0.19994913,0.07922512,0.05281675,0.14713238,0.44139713,1.0601076,1.4977322,1.267602,0.935611,0.724344,0.5357128,0.6790725,0.84884065,1.1129243,1.4411428,1.7089992,1.0148361,1.1431054,1.0374719,0.68661773,1.1053791,1.2600567,1.5543215,1.5958204,1.3656902,1.2487389,0.76584285,1.1996948,1.8184053,2.233394,2.4031622,4.2328854,3.682082,3.0746894,3.006782,2.3314822,2.0108092,2.0900342,2.1956677,2.1994405,2.233394,1.9051756,1.4939595,1.1921495,1.056335,1.0148361,0.7809334,0.5093044,0.35085413,0.31312788,0.27540162,0.20749438,0.19240387,0.21503963,0.241448,0.19994913,0.22258487,0.21503963,0.181086,0.13958712,0.14335975,0.14713238,0.1659955,0.17731337,0.18485862,0.19994913,0.28294688,0.3772625,0.4376245,0.38858038,0.120724,0.049044125,0.030181,0.10940613,0.32821837,0.7054809,2.082489,1.8485862,1.056335,0.49421388,0.6790725,0.694163,0.7130261,1.2411937,1.8900851,1.3807807,1.1016065,0.814887,0.6375736,0.62248313,0.7394345,1.2864652,2.123988,2.9237845,3.2859564,2.7389257,2.1994405,2.2560298,2.5389767,2.8256962,3.0331905,3.5877664,4.402653,5.50426,6.2625575,5.3910813,4.979865,4.1197066,3.240685,2.7502437,3.0218725,3.240685,3.8367596,4.5233774,4.6026025,2.9728284,3.4066803,3.1237335,2.8256962,2.7502437,2.6634734,2.7879698,3.802806,4.8138695,5.1760416,4.478106,4.9647746,5.7607985,6.56814,6.7454534,5.3269467,4.0480266,3.572676,3.561358,3.6481283,3.4594972,2.323937,1.871222,1.6863633,1.5467763,1.4109617,1.1883769,1.1619685,1.177059,1.1280149,0.9507015,0.76584285,0.6413463,0.6413463,0.73566186,0.83752275,0.7205714,0.44894236,0.41876137,0.69039035,0.97710985,0.80356914,0.5696664,0.3772625,0.26408374,0.211267,0.24522063,0.181086,0.1961765,0.3169005,0.4074435,0.41498876,0.23767537,0.120724,0.12826926,0.1358145,0.124496624,0.15467763,0.20749438,0.32821837,0.65643674,0.95824677,1.1129243,0.87902164,0.43385187,0.38858038,0.29049212,0.3055826,0.33953625,0.35839936,0.38480774,0.7394345,0.9922004,1.0487897,0.9016574,0.6526641,0.33953625,0.211267,0.29049212,0.42630664,0.28294688,0.26031113,0.35839936,0.5281675,0.68661773,0.7394345,1.1544232,1.20724,1.1053791,1.0186088,1.0902886,1.3166461,1.478869,1.4524606,1.3204187,1.358145,1.448688,1.2864652,0.9695646,0.6828451,0.7092535,0.69039035,0.543258,0.452715,0.5394854,0.87147635,1.690136,1.871222,1.6146835,1.1619685,0.7997965,0.935611,0.9280658,0.8186596,0.7469798,0.9507015,0.8186596,1.0336993,1.0676528,0.79602385,0.49421388,0.30935526,0.25276586,0.19240387,0.09808825,0.018863125,0.030181,0.060362,0.09808825,0.116951376,0.071679875,0.030181,0.060362,0.23390275,0.38858038,0.13204187,0.11317875,1.2789198,1.9768555,1.539231,0.29426476,0.06413463,0.00754525,0.003772625,0.003772625,0.011317875,0.124496624,0.08299775,0.02263575,0.011317875,0.030181,0.011317875,0.011317875,0.011317875,0.00754525,0.018863125,0.018863125,0.0150905,0.018863125,0.018863125,0.00754525,0.011317875,0.026408374,0.030181,0.018863125,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.033953626,0.09808825,0.18863125,0.17354076,0.12826926,0.120724,0.15845025,0.22258487,0.44894236,0.8563859,1.7052265,2.2484846,0.7582976,0.573439,0.6187105,0.9016574,1.4826416,2.4710693,3.8480775,5.2250857,6.7680893,8.601585,10.801025,12.136535,13.060828,13.8719425,14.634012,15.169725,16.116653,16.395828,16.878725,17.753973,18.519815,18.546225,18.297232,17.803017,17.908651,20.26277,20.013775,17.689838,15.199906,13.890805,14.558559,13.962485,12.257258,10.687846,9.691874,8.869441,8.526133,8.039464,7.7225633,7.4735703,6.760544,6.0626082,4.817642,3.5575855,2.6672459,2.3465726,2.1805773,2.6182017,2.9652832,3.138824,3.6707642,4.1536603,4.7874613,5.560849,6.541732,7.914967,8.013056,8.288457,9.224068,10.601076,11.510279,12.268577,13.038192,14.003984,15.16218,16.316603,18.723537,20.75321,21.967995,22.511253,23.118647,24.888006,26.07261,26.827137,27.445847,28.31355,29.120892,30.550716,31.010977,30.656351,31.407103,33.180237,33.881947,33.783855,33.146282,32.218216,31.671186,30.429993,29.739603,29.984823,30.66767,29.607561,30.573353,31.69005,32.07863,31.871136,32.05977,32.003178,31.825865,31.60328,31.327879,31.71646,32.61057,33.489594,34.255436,35.258953,37.69984,40.533085,43.400276,46.275017,49.46666,52.680935,56.759144,61.29384,65.97944,70.63109,75.426094,80.34182,84.80484,88.56615,91.682335,94.949425,97.59404,99.902885,101.96274,103.67928,105.742905,107.161415,108.30074,109.394806,110.53414,110.97931,110.526596,110.07011,109.68907,108.65537,106.45593,103.509514,100.16319,96.42452,91.94642,88.30961,84.50303,80.71531,76.92382,72.890884,70.4915,68.47691,66.68869,65.1985,64.2893,64.18744,63.802635,63.39142,62.946247,62.225677,60.27523,60.11678,60.41859,60.343136,59.554657,60.671356,62.504852,61.448517,56.306427,48.25942,43.95108,41.129158,38.322327,35.673943,34.904327,34.304478,35.34195,35.92671,35.274044,33.897038,33.078377,31.486328,30.33945,29.283115,26.41592,24.393793,22.941332,20.37972,16.414692,12.1101265,10.269085,8.677037,7.5226145,6.820906,6.4021444,6.0550632,5.7872066,5.560849,5.353355,5.1647234,5.100589,4.7308717,4.3083377,3.9159849,3.4670424,2.9200118,2.41448,1.9844007,1.6033657,1.177059,0.84129536,0.58098423,0.452715,0.41876137,0.331991,0.23767537,0.17354076,0.18863125,0.271629,0.36594462,0.42630664,0.482896,0.46026024,0.35085413,0.19994913,0.29803738,0.35462674,0.392353,0.43007925,0.47157812,0.29049212,0.14713238,0.05281675,0.003772625,0.0,0.02263575,0.026408374,0.033953626,0.041498873,0.030181,0.08299775,0.071679875,0.1056335,0.15467763,0.02263575,0.03772625,0.11317875,0.14713238,0.16222288,0.31312788,0.422534,0.46026024,0.5319401,0.573439,0.36971724,0.51684964,0.90920264,1.5845025,2.8521044,5.281675,7.5188417,8.356364,9.4127,11.310329,13.6682205,12.943876,12.204442,13.804035,16.610868,15.9695215,11.691365,8.096053,6.937857,7.3868,6.013564,3.2482302,2.2107582,6.3417826,11.668729,6.8133607,3.2746384,2.1579416,1.4524606,0.58098423,0.392353,0.31312788,0.13204187,0.018863125,0.00754525,0.00754525,0.0150905,0.0150905,0.011317875,0.00754525,0.0,0.24522063,0.2263575,0.27917424,0.5696664,0.77716076,0.08677038,0.090543,0.2565385,0.33576363,0.24522063,0.071679875,0.23767537,1.0789708,1.1732863,0.573439,0.8224323,2.4597516,1.2110126,0.10186087,0.2867195,1.0450171,0.62248313,0.44516975,0.241448,0.011317875,0.03772625,0.026408374,0.026408374,0.033953626,0.0754525,0.20372175,0.271629,2.9200118,4.727099,4.429062,2.9237845,1.9693103,2.4484336,3.0105548,3.289729,3.8971217,3.9989824,4.0103,3.5387223,2.505023,1.1581959,1.0035182,1.9730829,1.901403,0.69039035,0.33576363,0.23013012,0.2565385,0.6828451,1.327964,1.5920477,0.6488915,0.34330887,0.29803738,0.2867195,0.24522063,0.20372175,0.4074435,0.60362,0.62625575,0.36594462,0.1961765,0.13204187,0.1056335,0.094315626,0.09808825,0.10186087,0.071679875,0.03772625,0.018863125,0.026408374,0.041498873,0.02263575,0.003772625,0.05281675,0.2565385,0.26031113,0.211267,0.17354076,0.23390275,0.48666862,0.1961765,0.10186087,0.21503963,0.694163,1.8448136,2.5389767,2.033445,1.3241913,0.9242931,0.8639311,1.1657411,1.3053282,1.6524098,2.1466236,2.3201644,0.9242931,0.56212115,0.66775465,0.8941121,1.0789708,1.0676528,1.1883769,1.4373702,1.7769064,2.1466236,2.0673985,2.252257,2.5767028,2.6521554,1.8297231,2.746471,2.4031622,2.0183544,1.9579924,1.7278622,1.5769572,1.6750455,1.7919968,1.8825399,2.093807,2.1164427,2.1013522,1.9202662,1.6561824,1.569412,1.3166461,0.8186596,0.48666862,0.41876137,0.38858038,0.2867195,0.23767537,0.26408374,0.331991,0.3470815,0.33576363,0.29049212,0.22258487,0.1659955,0.17731337,0.21881226,0.23013012,0.20749438,0.17354076,0.19994913,0.28294688,0.38858038,0.452715,0.4074435,0.18485862,0.10186087,0.08677038,0.20749438,0.5055317,0.995973,2.6785638,2.263575,1.2902378,0.67152727,0.67152727,0.59230214,0.814887,1.8863125,2.9992368,1.9806281,1.3958713,1.0450171,0.9318384,1.0450171,1.3543724,1.5656394,2.1202152,3.2369123,4.266839,3.6783094,3.2369123,3.5047686,4.0404816,4.38379,4.0480266,5.070408,4.957229,5.323174,6.33801,6.7114997,5.9607477,4.459243,3.4066803,3.3915899,4.425289,3.3274553,3.4557245,4.432834,5.0553174,3.2670932,2.867195,3.138824,3.2067313,2.897376,2.704972,2.2220762,3.0445085,4.055572,4.6742826,4.8629136,5.674028,6.0776987,6.2889657,5.915476,3.9574835,3.2784111,3.2369123,3.2821836,3.1652324,2.916239,1.9127209,1.5882751,1.6373192,1.7278622,1.4901869,1.2525115,1.2751472,1.4034165,1.3656902,0.7582976,0.41498876,0.35839936,0.41876137,0.46026024,0.392353,0.69039035,0.3961256,0.14713238,0.11317875,0.03772625,0.07922512,0.116951376,0.10940613,0.0754525,0.08299775,0.060362,0.060362,0.06413463,0.094315626,0.16976812,0.21881226,0.17354076,0.16222288,0.20749438,0.20749438,0.24522063,0.29049212,0.35085413,0.41121614,0.45648763,0.8941121,1.0035182,0.7130261,0.3055826,0.392353,0.38103512,0.5281675,0.5583485,0.44894236,0.43385187,0.8563859,1.1657411,0.9922004,0.49421388,0.3169005,0.3169005,0.271629,0.1961765,0.120724,0.1056335,0.34330887,0.56589377,0.9016574,1.177059,0.9205205,0.8526133,0.87147635,0.9997456,1.1204696,0.9997456,0.98465514,1.1091517,1.2562841,1.3694628,1.4637785,1.297783,1.0223814,0.7432071,0.5583485,0.55080324,0.56212115,0.44139713,0.32067314,0.3055826,0.44516975,0.663982,0.9393836,1.1204696,1.1544232,1.0751982,1.2638294,1.2789198,1.1921495,1.1355602,1.327964,1.6561824,2.0636258,1.750498,0.8262049,0.32067314,0.18485862,0.090543,0.030181,0.00754525,0.0150905,0.030181,0.0452715,0.049044125,0.060362,0.12826926,0.0452715,0.090543,0.41498876,0.724344,0.28294688,0.23767537,0.25276586,0.23390275,0.150905,0.0452715,0.011317875,0.00754525,0.0150905,0.018863125,0.02263575,0.16222288,0.12826926,0.060362,0.033953626,0.041498873,0.026408374,0.026408374,0.02263575,0.011317875,0.0,0.0,0.00754525,0.02263575,0.030181,0.026408374,0.05281675,0.071679875,0.06413463,0.030181,0.00754525,0.0,0.0150905,0.018863125,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.0,0.0,0.011317875,0.0150905,0.011317875,0.003772625,0.0150905,0.018863125,0.02263575,0.07922512,0.20372175,0.40367088,0.38103512,0.30181,0.2867195,0.32821837,0.29426476,0.4074435,0.58475685,0.754525,0.9393836,1.2449663,1.2449663,1.3732355,1.7957695,2.6144292,3.8707132,5.6098933,7.594294,9.563604,11.608367,14.177525,16.493916,18.010511,18.904623,19.168707,18.632996,17.723793,16.965494,16.11288,15.067864,13.8870325,14.347293,16.15438,16.667458,16.01102,17.067356,17.689838,16.84477,15.294222,13.917213,13.721037,14.339747,13.879487,13.151371,12.691111,12.751472,12.540206,12.076173,11.951676,11.868678,10.638803,9.699419,7.8998766,5.983383,4.4743333,3.682082,3.350091,3.6443558,3.7386713,3.6141748,4.044254,4.2819295,3.591539,2.795515,2.2786655,1.9881734,1.9240388,2.2711203,3.2935016,4.8138695,6.1908774,7.1868505,8.126234,8.975075,9.880505,11.16697,13.392818,16.060064,18.523588,20.345766,21.281378,22.296213,23.107328,24.454155,26.280106,27.732567,29.079393,30.214954,31.27506,32.61434,34.80624,37.662117,39.94078,40.906574,40.567036,39.646515,38.48832,36.17193,34.911873,35.97198,39.657833,35.217453,34.13094,34.34975,34.21771,32.42194,30.799711,29.64906,29.57738,30.42622,31.263742,31.207153,31.916407,32.765247,33.54618,34.470474,35.768257,37.096222,38.209145,39.1938,40.491585,40.748123,40.67644,40.793396,41.283836,41.977997,43.777542,46.037342,48.644226,51.402016,54.06549,56.993046,59.147213,60.788307,62.236996,63.878086,66.46611,69.57098,72.92107,76.523926,80.65118,84.6728,88.03043,91.16548,94.14586,96.67729,98.14484,99.08422,99.42376,98.89182,97.0206,95.9869,94.508026,92.357635,89.21881,84.66525,81.24725,77.848114,74.47162,71.483696,69.6087,68.322235,67.18291,66.31143,65.76817,65.58331,64.8401,65.38336,65.23246,63.78,61.78805,64.89292,67.929886,65.54936,57.094906,46.599464,43.01924,41.381924,38.714676,35.251408,34.45161,34.65156,35.390995,36.42092,37.216946,37.001907,33.621635,31.988087,31.1732,30.116865,27.649569,25.457674,23.69963,21.473782,18.421728,14.70192,12.438345,10.61994,9.265567,8.371455,7.865923,7.854605,7.7829256,7.6697464,7.488661,7.164215,6.692637,6.2097406,5.6589375,5.05909,4.5196047,3.8292143,3.3161373,2.8030603,2.2673476,1.8523588,1.3694628,0.965792,0.6790725,0.513077,0.41876137,0.29803738,0.2263575,0.22258487,0.28294688,0.38480774,0.422534,0.59230214,0.66775465,0.5583485,0.29049212,0.27917424,0.4074435,0.52062225,0.5470306,0.49421388,0.29049212,0.150905,0.06413463,0.0150905,0.0,0.0,0.0,0.03772625,0.090543,0.060362,0.16976812,0.1056335,0.060362,0.06413463,0.02263575,0.060362,0.03772625,0.041498873,0.09808825,0.181086,0.19240387,0.26408374,0.35462674,0.41876137,0.39989826,0.43007925,0.5470306,0.7997965,1.2902378,2.1805773,3.9612563,6.2889657,8.756263,11.649866,15.961976,16.392056,12.909923,11.034928,11.623458,10.853842,8.126234,5.6023483,3.591539,2.3503454,2.0862615,1.4600059,1.6976813,2.3578906,2.6597006,1.50905,1.1242423,1.2562841,1.2789198,1.0072908,0.69039035,0.513077,0.21881226,0.041498873,0.018863125,0.00754525,0.011317875,0.011317875,0.00754525,0.0,0.0,1.1581959,1.0751982,0.7884786,0.482896,0.30935526,0.38103512,0.150905,0.29426476,0.27540162,0.03772625,0.0,0.03772625,0.6488915,0.754525,0.331991,0.44139713,0.6375736,0.33953625,0.06413463,0.00754525,0.030181,0.26408374,0.23013012,0.1056335,0.049044125,0.18485862,0.1358145,0.13204187,0.1659955,0.3734899,1.0223814,1.267602,2.3880715,3.1727777,2.9728284,1.7391801,2.191895,2.9992368,5.20245,7.3868,5.692891,3.2633207,1.6033657,0.6790725,0.52062225,1.20724,1.6561824,1.4298248,0.8224323,0.24899325,0.27540162,0.23767537,0.23767537,0.32821837,0.482896,0.58098423,0.543258,0.44139713,0.362172,0.3169005,0.24522063,0.1961765,0.17354076,0.16222288,0.14713238,0.120724,0.09808825,0.19994913,0.2565385,0.1961765,0.060362,0.03772625,0.02263575,0.0150905,0.041498873,0.1358145,0.211267,0.10940613,0.018863125,0.060362,0.3055826,0.071679875,0.02263575,0.1659955,0.40367088,0.55080324,0.35462674,0.2678564,0.543258,1.2449663,2.2598023,1.7316349,0.9808825,0.5583485,0.65643674,1.0827434,1.50905,2.4672968,3.3915899,4.0895257,4.7610526,1.5015048,0.56589377,0.7205714,1.1506506,1.478869,2.3088465,3.361409,4.5007415,5.8702044,7.8734684,7.5188417,6.6624556,6.643593,6.9567204,5.247721,3.3312278,2.4522061,2.04099,1.750498,1.4335974,1.4713237,1.6071383,1.8448136,2.1051247,2.2296214,2.0560806,2.5540671,2.7389257,2.4823873,2.5314314,2.4484336,1.6033657,0.9242931,0.7167987,0.65643674,0.58098423,0.45648763,0.35085413,0.32444575,0.3961256,0.38480774,0.35462674,0.3055826,0.26408374,0.27540162,0.2867195,0.26408374,0.23767537,0.23390275,0.26031113,0.29426476,0.32444575,0.3169005,0.271629,0.19994913,0.16222288,0.23390275,0.47157812,0.7884786,0.94692886,0.9205205,1.0148361,1.1129243,1.0978339,0.8526133,0.6111652,0.4678055,0.5772116,0.8337501,0.87147635,1.3694628,1.3392819,1.2600567,1.3543724,1.5882751,1.5731846,1.9391292,2.3767538,2.674791,2.7011995,2.6031113,2.8822856,3.0218725,3.0331905,3.4481792,3.5349495,3.3538637,3.5877664,4.4177437,5.5382137,5.2590394,4.8855495,4.7572803,4.6554193,3.8141239,3.169005,2.9501927,3.108643,3.3048196,2.916239,2.425798,2.9803739,3.531177,3.6330378,3.4481792,2.6068838,2.3126192,2.2899833,2.493705,3.127506,4.847823,5.553304,5.7306175,5.3873086,4.044254,3.6292653,4.1197066,4.08198,3.2067313,2.305074,1.3996439,1.4298248,1.5769572,1.4034165,0.8563859,0.694163,0.83752275,1.1204696,1.2223305,0.68661773,0.331991,0.19994913,0.23013012,0.29426476,0.18485862,0.2678564,0.1358145,0.041498873,0.071679875,0.120724,0.09808825,0.071679875,0.060362,0.056589376,0.0452715,0.033953626,0.011317875,0.0,0.049044125,0.24522063,0.27917424,0.29803738,0.35462674,0.40367088,0.3055826,0.34330887,0.3961256,0.44516975,0.45648763,0.3961256,0.43385187,0.47157812,0.3961256,0.27917424,0.36594462,0.4640329,0.87147635,1.0487897,0.8111144,0.33576363,0.31312788,0.13204187,0.00754525,0.0,0.0,0.0,0.0,0.0,0.033953626,0.1659955,0.5696664,0.8639311,0.9808825,0.90920264,0.70170826,0.59230214,0.6451189,0.84129536,1.1091517,1.327964,1.2525115,1.1544232,1.2261031,1.5128226,1.8938577,1.8448136,1.4637785,0.97710985,0.55080324,0.3055826,0.23013012,0.20372175,0.21503963,0.2867195,0.45648763,0.58098423,0.7205714,0.8224323,0.97710985,1.4034165,2.2447119,2.384299,2.1088974,1.8297231,2.0598533,3.9989824,4.1008434,3.138824,1.871222,1.0525624,0.7582976,0.38480774,0.120724,0.041498873,0.0754525,0.10186087,0.05281675,0.02263575,0.030181,0.030181,0.00754525,0.0,0.03772625,0.150905,0.38103512,0.10186087,0.02263575,0.02263575,0.033953626,0.0452715,0.02263575,0.041498873,0.06790725,0.060362,0.0,0.011317875,0.02263575,0.060362,0.10186087,0.0754525,0.05281675,0.03772625,0.02263575,0.011317875,0.0,0.0,0.00754525,0.02263575,0.041498873,0.0754525,0.16222288,0.1659955,0.116951376,0.056589376,0.030181,0.00754525,0.0,0.011317875,0.030181,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.026408374,0.056589376,0.16222288,0.36594462,0.67152727,0.66020936,0.6111652,0.7092535,0.80734175,0.42630664,0.36594462,0.5885295,0.65643674,0.7092535,1.4637785,2.1013522,2.4597516,3.2218218,4.678055,6.730363,8.816625,10.582213,12.102581,13.58145,15.350811,17.512526,18.893307,20.14959,21.051247,20.477808,17.976559,15.901614,14.158662,12.691111,11.506506,12.347801,13.875714,14.543469,14.5283785,15.746937,16.271332,15.17727,12.593022,9.703192,8.729855,9.276885,9.058073,8.959985,9.393836,10.284176,9.967276,9.703192,9.276885,8.514814,7.2924843,6.4134626,5.243949,4.1272516,3.2670932,2.71629,2.5804756,2.5578396,1.9844007,1.0902886,0.9922004,1.2600567,1.3091009,1.237421,1.1242423,1.0374719,1.0487897,1.4373702,2.04099,2.7841973,3.663219,4.979865,6.3908267,7.586749,8.627994,9.933322,11.446144,13.143826,15.116908,17.071129,18.342503,19.304522,20.617395,22.522572,25.05023,28.015512,30.931753,34.123394,37.32258,40.555717,44.143486,47.09745,49.100716,49.64397,48.912083,47.791615,47.022,46.516468,46.369335,46.01848,44.234028,42.306217,40.751896,39.49561,38.035606,35.462673,34.632698,33.738586,33.180237,33.229282,34.010216,33.09724,32.9237,32.35403,31.407103,31.233562,30.686531,30.165909,29.566063,29.015259,28.871899,27.758974,25.412401,23.148827,21.764273,21.53037,22.03213,22.315077,23.465727,25.269043,26.185791,27.24967,28.438047,29.581152,30.860073,32.82561,34.632698,37.043404,39.56729,41.955364,44.17744,46.65605,50.002373,53.688225,57.275993,60.411045,64.91556,70.10669,75.51286,80.61345,84.8237,88.69441,91.53897,93.14989,93.75728,94.04022,92.866936,89.95447,86.23089,82.40167,78.94972,75.72413,73.33606,71.82701,71.0008,70.404724,71.18566,71.993004,70.82349,67.58658,64.13085,65.489,65.92662,62.69348,56.034798,49.225212,47.821796,46.73905,43.381416,38.34496,35.417404,38.563774,36.83591,36.481285,39.295662,42.615574,40.85753,37.53762,34.79115,32.859562,30.090458,27.038403,25.314314,23.062057,20.145817,18.142553,14.894323,12.491161,10.616167,9.208978,8.4544525,8.635539,8.884532,9.242931,9.495697,9.14107,8.103599,7.3377557,6.6813188,6.058836,5.5080323,4.738417,4.0517993,3.4368613,2.8898308,2.425798,2.0598533,1.6109109,1.1883769,0.87147635,0.68661773,0.5281675,0.4979865,0.44894236,0.3470815,0.27540162,0.52062225,0.7432071,0.90920264,0.8865669,0.47157812,0.3734899,0.51684964,0.694163,0.77338815,0.70170826,0.35839936,0.17354076,0.0754525,0.02263575,0.0,0.0,0.0,0.02263575,0.049044125,0.0,0.0,0.0,0.1056335,0.21881226,0.060362,0.03772625,0.030181,0.056589376,0.08299775,0.0452715,0.056589376,0.1056335,0.19994913,0.27917424,0.23013012,0.29049212,0.44139713,0.62625575,1.0223814,2.0598533,5.9305663,10.631257,14.147344,15.728074,15.897841,13.275867,7.8131065,4.323428,4.0895257,4.881777,6.2851934,5.8211603,3.9989824,1.901403,1.20724,1.2525115,1.9240388,2.04099,1.3770081,0.65643674,0.4376245,0.9393836,1.8863125,2.3390274,0.70170826,0.24899325,0.10940613,0.09808825,0.090543,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.7809334,0.65643674,0.87147635,0.694163,0.16976812,0.124496624,0.3734899,1.3241913,1.20724,0.16222288,0.24522063,0.14335975,0.21881226,0.23390275,0.3055826,0.8941121,0.8941121,0.36971724,0.15845025,0.5470306,1.2638294,0.31312788,0.116951376,0.1056335,0.15467763,0.56212115,0.6413463,1.1355602,1.2411937,0.9507015,1.0714256,1.0902886,1.8636768,2.4408884,2.6219745,2.9728284,3.1425967,3.4896781,5.983383,8.8618965,6.6549106,2.957738,1.3958713,0.9280658,0.95824677,1.3392819,1.3619176,0.8601585,0.3772625,0.19240387,0.33576363,0.3169005,0.241448,0.23767537,0.31312788,0.3734899,0.40367088,0.36594462,0.32067314,0.2867195,0.23013012,0.15467763,0.094315626,0.07922512,0.1056335,0.15845025,0.1056335,0.0754525,0.071679875,0.071679875,0.02263575,0.06790725,0.056589376,0.026408374,0.02263575,0.10186087,0.23390275,0.17731337,0.124496624,0.26031113,0.7696155,0.5093044,0.2263575,0.1056335,0.38480774,1.3317367,2.6785638,2.7879698,2.987919,3.5047686,3.4557245,2.2560298,1.5618668,0.95824677,0.70170826,1.7052265,5.9230213,7.7414265,7.484888,6.017337,4.7233267,2.957738,3.350091,3.6556737,3.3123648,3.4557245,4.696918,4.678055,4.285702,4.327201,5.5306683,6.4247804,6.0776987,6.2889657,7.3717093,8.141325,6.40969,5.3759904,4.357382,3.0143273,1.3505998,0.98465514,1.1393328,1.4864142,1.7240896,1.5807298,1.2826926,1.5505489,1.7014539,1.7693611,2.5201135,3.5387223,3.4029078,2.9426475,2.5767028,2.2899833,1.5165952,1.0374719,0.72811663,0.543258,0.52062225,0.4678055,0.36971724,0.34330887,0.41498876,0.49421388,0.38858038,0.27540162,0.241448,0.28294688,0.29426476,0.29426476,0.29049212,0.2678564,0.23013012,0.18485862,0.20749438,0.23767537,0.35462674,0.5772116,0.87147635,0.663982,0.6451189,0.87902164,1.2147852,1.2826926,0.88279426,0.6752999,0.5998474,0.6488915,0.88279426,0.97333723,0.8978847,0.95447415,1.2411937,1.6486372,2.11267,2.4559789,2.7125173,2.8747404,2.9200118,2.305074,2.5691576,2.8936033,2.9124665,2.7540162,3.0445085,3.0407357,2.9615107,3.1161883,3.8782585,4.7610526,4.6214657,4.5309224,4.568649,3.8141239,4.496969,4.9760923,5.8702044,6.4134626,4.5007415,3.7084904,3.2972744,3.3048196,3.5839937,3.802806,2.655928,2.033445,1.599593,1.3317367,1.5165952,2.7200627,3.531177,4.093298,4.447925,4.5196047,4.221567,4.1272516,3.3350005,2.022127,1.4600059,1.5845025,1.7240896,1.4637785,0.90920264,0.6828451,0.543258,0.55457586,0.66775465,0.7394345,0.51684964,0.3961256,0.2678564,0.24522063,0.29803738,0.2565385,0.59607476,0.452715,0.20749438,0.094315626,0.16976812,0.1056335,0.060362,0.05281675,0.071679875,0.071679875,0.018863125,0.003772625,0.03772625,0.271629,0.965792,0.33576363,0.18863125,0.17731337,0.1358145,0.09808825,0.0754525,0.08677038,0.124496624,0.19994913,0.33576363,0.39989826,0.4074435,0.29803738,0.1358145,0.120724,0.120724,0.19994913,0.23013012,0.17354076,0.06790725,0.06413463,0.026408374,0.0,0.0,0.0,0.0,0.0,0.011317875,0.056589376,0.181086,0.38858038,0.48666862,0.47912338,0.43007925,0.44516975,0.6790725,0.98465514,1.4562333,1.9542197,2.1315331,2.8407867,2.474842,1.9844007,1.8674494,2.1466236,1.8938577,1.3468271,0.8262049,0.47912338,0.29426476,0.16976812,0.13958712,0.14713238,0.17354076,0.2263575,0.32821837,0.86770374,1.3543724,1.8485862,2.9313297,3.0105548,2.8407867,2.4107075,1.9089483,1.7316349,2.3805263,2.535204,2.3616633,2.11267,2.1164427,1.3920987,0.76207024,0.362172,0.2263575,0.28294688,0.19240387,0.0754525,0.011317875,0.00754525,0.00754525,0.0,0.0,0.011317875,0.041498873,0.08677038,0.033953626,0.0150905,0.02263575,0.041498873,0.08299775,0.1056335,0.19994913,0.181086,0.060362,0.03772625,0.018863125,0.018863125,0.071679875,0.181086,0.28294688,0.14335975,0.1056335,0.06790725,0.011317875,0.0,0.0,0.030181,0.05281675,0.05281675,0.041498873,0.1358145,0.22258487,0.17354076,0.030181,0.00754525,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.003772625,0.003772625,0.0,0.00754525,0.00754525,0.003772625,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.026408374,0.060362,0.116951376,0.26031113,0.543258,1.026154,0.97333723,0.7922512,0.68661773,0.6413463,0.392353,0.3961256,0.4979865,0.5055317,0.5281675,0.965792,2.0673985,2.2296214,2.8256962,4.123479,5.2779026,6.8774953,8.043237,8.843033,9.378746,9.820143,10.801025,11.3820095,12.623203,14.086982,13.826671,12.543978,11.521597,10.661438,9.869187,9.076936,9.556059,10.095545,9.793735,9.14107,10.008774,9.529651,8.167733,6.300284,4.617693,4.13857,3.8367596,3.4934506,3.3538637,3.429316,3.5085413,3.4481792,3.4368613,3.006782,2.293756,2.071171,2.0975795,1.599593,1.1280149,0.87147635,0.6526641,0.5885295,0.6073926,0.5470306,0.41876137,0.43007925,0.63002837,0.7922512,0.94692886,1.0714256,1.1242423,1.2147852,1.3505998,1.629774,2.161714,3.0407357,4.112161,5.3910813,6.820906,8.345046,9.895596,11.529142,13.407909,15.460217,17.346529,18.440592,19.28566,21.31533,24.378702,27.826881,30.528082,33.504684,35.636215,36.97927,37.862064,38.884445,39.39375,39.895508,40.87262,42.347717,43.86054,45.452587,46.76546,47.618073,47.818024,47.127632,45.992073,43.800175,42.230762,40.891483,37.341442,34.39125,32.433258,31.05625,30.116865,29.728285,28.547453,27.457165,26.87618,26.608324,25.850027,24.842735,24.095757,23.231825,22.130219,20.960705,19.711966,18.614132,17.572887,16.724047,16.403374,16.014793,15.69412,15.543215,15.490398,15.282904,15.701665,16.422237,17.599297,19.168707,20.858843,22.997923,25.397312,27.80802,30.067822,32.112583,33.82913,35.390995,36.737823,37.99788,39.47675,41.774277,44.369843,47.05595,50.062733,54.03908,58.03429,61.95782,66.02471,70.182144,74.09435,77.19923,79.21004,80.126785,79.90797,78.47437,77.21432,76.05989,74.92811,74.25658,75.00733,76.29379,75.96935,73.21533,69.24653,67.3074,66.982956,64.45907,59.54711,53.756134,50.323044,51.360516,51.55292,49.417614,45.61858,42.98529,43.566273,42.736298,41.540375,40.578354,40.031322,39.657833,39.186256,38.85049,38.81654,39.159847,35.666397,31.31656,27.14781,23.737356,21.1682,18.19537,15.924251,13.909668,12.132762,11.004747,10.378491,10.223814,10.374719,10.442626,9.8239155,9.118435,8.650629,8.231868,7.654656,6.7039547,5.915476,5.2552667,4.6026025,3.9159849,3.218049,2.746471,2.2862108,1.8523588,1.4713237,1.1506506,0.845068,0.66775465,0.56589377,0.49044126,0.4074435,0.58475685,0.80734175,0.90920264,0.8563859,0.754525,0.65643674,0.51684964,0.44516975,0.44139713,0.4074435,0.29049212,0.18485862,0.10940613,0.06413463,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.03772625,0.08677038,0.10940613,0.049044125,0.033953626,0.030181,0.030181,0.030181,0.033953626,0.056589376,0.090543,0.120724,0.14713238,0.20372175,0.46026024,0.41876137,0.5357128,1.0450171,1.9730829,4.644101,8.122461,10.56335,11.019837,9.442881,7.284939,4.7535076,3.3878171,3.8065786,5.7117543,5.798525,4.38379,2.6106565,1.3355093,1.1091517,1.1846043,1.3807807,1.3505998,1.1544232,1.2525115,0.59607476,0.62248313,0.7696155,0.6752999,0.19994913,0.071679875,0.056589376,0.05281675,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.0,0.35839936,0.30181,0.5017591,0.41876137,0.090543,0.09808825,0.9016574,1.5354583,1.4864142,0.9205205,0.67152727,0.22258487,0.10940613,0.09808825,0.2678564,1.026154,1.026154,0.41121614,0.07922512,0.34330887,0.9016574,0.48666862,0.18485862,0.18485862,0.45648763,0.7582976,0.6828451,1.0525624,1.0751982,0.6828451,0.52439487,0.84129536,1.4071891,1.7052265,1.8485862,2.584248,2.1315331,1.9466745,3.4444065,5.481624,4.353609,1.9844007,2.354118,3.361409,3.6858547,2.7841973,3.180323,3.9461658,3.3576362,1.50905,0.29426476,0.28294688,0.23767537,0.19994913,0.19240387,0.21881226,0.23767537,0.23013012,0.20749438,0.181086,0.14713238,0.090543,0.0452715,0.033953626,0.049044125,0.08677038,0.090543,0.26031113,0.5017591,0.6187105,0.3169005,0.10186087,0.030181,0.05281675,0.17354076,0.45648763,0.48666862,0.3772625,0.27917424,0.35462674,0.80356914,0.87147635,1.750498,3.0633714,4.2064767,4.327201,3.3953626,2.41448,1.8863125,1.9278114,2.2598023,1.7957695,1.6260014,1.7618159,2.9615107,6.722818,10.838752,8.461998,5.402399,4.38379,5.0553174,4.7912335,4.938366,4.0517993,2.354118,1.7278622,2.2484846,2.1202152,1.841041,1.7769064,2.1692593,2.6106565,2.6144292,2.9237845,3.651901,4.2894745,3.8103511,4.255521,5.089271,5.3571277,3.6971724,2.384299,1.8636768,1.720317,1.6863633,1.6373192,1.5656394,1.4675511,1.5015048,1.7240896,2.0975795,2.5276587,2.6974268,2.6634734,2.4182527,1.8787673,1.4600059,1.4750963,1.3732355,1.056335,0.8978847,0.72811663,0.62625575,0.73566186,0.94315624,0.87902164,0.65643674,0.513077,0.43007925,0.39989826,0.3961256,0.44139713,0.39989826,0.35085413,0.32821837,0.32067314,0.49044126,0.56589377,0.6073926,0.6752999,0.845068,0.72811663,0.94315624,1.026154,0.8978847,0.8299775,0.6828451,0.8337501,0.9205205,0.9016574,1.0601076,1.1657411,1.0978339,1.0676528,1.3053282,2.0673985,2.9086938,3.5764484,4.0404816,4.214022,3.9273026,2.727608,2.305074,2.444661,2.7087448,2.4408884,2.987919,2.969056,2.6521554,2.3692086,2.5201135,3.561358,3.9801195,4.1083884,3.9612563,3.2369123,4.3385186,6.043745,6.9982195,6.6360474,5.1835866,5.3194013,4.5497856,3.8782585,3.731126,3.9914372,3.482133,2.655928,2.2258487,2.3503454,2.6144292,2.9728284,2.9841464,3.5575855,4.6554193,5.3269467,4.7572803,4.478106,3.399135,1.7655885,1.1431054,1.4675511,1.4411428,1.0676528,0.62625575,0.68661773,0.7130261,0.7582976,0.7696155,0.7054809,0.49044126,0.4678055,0.3055826,0.20372175,0.2263575,0.32067314,0.47535074,0.30935526,0.116951376,0.03772625,0.071679875,0.0452715,0.03772625,0.056589376,0.0754525,0.041498873,0.00754525,0.0,0.049044125,0.1961765,0.49421388,0.14713238,0.06413463,0.05281675,0.026408374,0.018863125,0.003772625,0.003772625,0.02263575,0.0754525,0.19240387,0.19240387,0.17354076,0.11317875,0.03772625,0.02263575,0.0150905,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.06790725,0.18485862,0.2678564,0.27540162,0.3169005,0.43007925,0.59230214,0.7922512,1.0299267,1.2789198,1.5052774,1.6863633,2.2862108,2.5314314,2.372981,2.003264,1.8636768,1.2751472,0.80734175,0.55457586,0.4640329,0.34330887,0.150905,0.08677038,0.07922512,0.090543,0.120724,0.211267,0.66020936,1.4335974,2.5201135,3.9348478,4.0291634,4.323428,4.2592936,3.7914882,3.3764994,2.9841464,2.5993385,2.2975287,2.293756,2.9464202,2.3654358,1.5505489,0.9808825,0.7205714,0.4074435,0.16222288,0.0452715,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.02263575,0.018863125,0.0150905,0.026408374,0.08299775,0.11317875,0.15467763,0.13204187,0.0754525,0.1358145,0.060362,0.02263575,0.05281675,0.181086,0.4074435,0.1358145,0.10186087,0.10186087,0.0754525,0.090543,0.041498873,0.03772625,0.03772625,0.030181,0.011317875,0.071679875,0.18863125,0.16976812,0.03772625,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.02263575,0.056589376,0.16222288,0.35085413,0.5998474,0.8299775,0.694163,0.5319401,0.45648763,0.46026024,0.39989826,0.49044126,0.70170826,0.7469798,0.6526641,0.7582976,1.3619176,1.5015048,1.8448136,2.5691576,3.3651814,4.376245,5.2665844,5.881522,6.1795597,6.221059,6.628502,6.983129,7.575431,8.258276,8.473316,7.911195,7.4509344,7.0359454,6.537959,5.775889,5.583485,5.372218,5.1081343,4.8063245,4.5460134,4.5196047,4.1008434,3.0709167,1.9164935,1.8184053,1.2713746,1.1581959,1.1393328,1.0223814,0.7922512,0.8639311,0.875249,0.6752999,0.38858038,0.43385187,0.543258,0.41876137,0.3055826,0.26031113,0.15467763,0.07922512,0.0754525,0.1056335,0.15845025,0.25276586,0.5772116,0.90543,1.1242423,1.20724,1.2185578,1.3053282,1.388326,1.5769572,1.9844007,2.7389257,3.6330378,4.6931453,5.9720654,7.4282985,8.899622,10.186088,11.793225,13.532406,15.094273,16.063837,16.818363,18.689585,21.55678,24.76351,27.166672,28.694586,29.69056,29.924461,29.622652,29.47552,30.22627,31.686277,33.93099,36.730278,39.555973,41.306473,42.68348,43.736042,44.2378,43.668133,43.01924,41.679962,40.800938,40.26523,38.642998,35.847485,32.474754,29.822601,28.502182,28.419184,25.774574,24.39002,23.763765,23.401592,22.813063,22.398075,22.17549,21.503962,20.315586,19.093256,17.591751,16.648594,15.845025,15.052773,14.452927,13.717264,13.158916,12.679792,12.325166,12.283667,11.966766,12.045992,12.411936,13.004238,13.792717,14.754736,16.018566,17.346529,18.69713,20.209951,21.934042,23.548725,25.080412,26.532871,27.887243,29.464201,31.237335,32.88597,34.693058,37.533848,39.9521,42.5288,45.520493,48.855495,52.126358,55.340637,58.022972,60.39218,62.519943,64.345894,66.17939,67.45076,68.52973,70.28023,74.105675,77.34636,76.93514,74.034,70.891396,70.84612,70.89894,67.71484,62.104954,56.163067,53.299644,53.92213,53.869312,52.763935,50.90403,49.27048,49.01017,49.081852,47.829338,45.24509,42.951336,41.612053,42.483532,43.702087,44.12085,43.339916,40.01623,35.855026,31.72023,28.215462,25.680258,23.318596,21.477554,19.613878,17.761518,16.539188,15.343266,14.366156,13.804035,13.370183,12.283667,11.2801485,10.604849,10.057818,9.405154,8.386545,7.7829256,7.115171,6.432326,5.726845,4.9119577,4.085753,3.4444065,2.8822856,2.3805263,1.9994912,1.6410918,1.267602,0.995973,0.83752275,0.6790725,0.68661773,0.7997965,0.87902164,0.8865669,0.87147635,0.83752275,0.59607476,0.3734899,0.26031113,0.20749438,0.16976812,0.116951376,0.06790725,0.030181,0.0,0.0,0.0150905,0.0150905,0.0,0.0,0.0,0.018863125,0.033953626,0.033953626,0.018863125,0.0150905,0.011317875,0.02263575,0.041498873,0.041498873,0.049044125,0.06790725,0.071679875,0.071679875,0.09808825,0.21881226,0.2565385,0.32444575,0.5319401,0.97333723,2.0673985,3.6028569,4.7233267,4.979865,4.357382,4.2517486,4.2328854,4.9044123,7.062354,11.680047,9.024119,4.8629136,1.901403,0.9318384,0.83752275,0.80356914,0.814887,0.845068,0.845068,0.72811663,0.3470815,0.27917424,0.27917424,0.241448,0.21503963,0.150905,0.08299775,0.033953626,0.003772625,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.08299775,0.5470306,0.95447415,0.8111144,0.2678564,0.09808825,1.1053791,1.1091517,0.95824677,0.8978847,0.58475685,0.16976812,0.24522063,0.62625575,0.9393836,0.633801,0.65643674,0.2678564,0.0150905,0.08299775,0.32444575,0.51684964,0.26031113,0.17731337,0.38480774,0.49421388,0.49044126,0.58098423,0.5055317,0.26408374,0.12826926,0.513077,1.0374719,1.1431054,1.0902886,1.9579924,2.384299,1.9730829,1.9164935,2.2786655,2.003264,1.2411937,3.4745877,5.0175915,4.564876,3.199186,3.772625,4.436607,3.99521,2.2862108,0.19994913,0.21503963,0.1961765,0.14335975,0.090543,0.09808825,0.09808825,0.1056335,0.09808825,0.0754525,0.056589376,0.35462674,0.30181,0.13958712,0.026408374,0.02263575,0.3772625,0.56589377,0.694163,0.7394345,0.55080324,0.25276586,0.14335975,0.18863125,0.36594462,0.67152727,0.724344,0.6149379,0.935611,1.478869,1.2487389,1.1695137,2.191895,3.6179473,4.6818275,4.564876,2.655928,1.388326,1.1921495,2.4710693,5.587258,4.5007415,3.380272,2.938875,3.9650288,7.322665,9.322156,6.307829,3.8065786,3.9310753,5.3910813,4.9157305,4.1008434,2.6446102,0.995973,0.33576363,0.181086,0.13958712,0.29049212,0.5583485,0.7469798,0.3169005,0.31312788,0.52439487,0.76207024,0.8639311,1.3694628,2.3880715,3.802806,5.0741806,5.2552667,4.7912335,3.451952,2.142851,1.3996439,1.3807807,1.5430037,1.4524606,1.4335974,1.5052774,1.3694628,1.3053282,1.4600059,1.6033657,1.5656394,1.2110126,1.20724,1.4750963,1.448688,1.1280149,1.0789708,0.73188925,0.633801,0.76207024,0.9280658,0.7507524,0.59230214,0.5470306,0.47912338,0.3961256,0.42630664,0.5319401,0.51684964,0.4640329,0.41876137,0.38858038,0.5017591,0.55080324,0.56212115,0.6375736,0.9242931,0.7205714,1.0940613,1.2562841,0.995973,0.694163,0.5772116,0.91297525,1.1921495,1.2034674,1.0299267,1.0374719,0.9016574,0.7696155,0.87902164,1.5279131,2.3088465,3.229367,3.9914372,4.323428,3.983892,3.4330888,2.9916916,3.0445085,3.2670932,2.5804756,3.0935526,3.289729,2.969056,2.354118,2.0673985,3.0558262,3.8254418,4.0706625,3.731126,2.987919,3.7990334,5.715527,6.5568223,6.1041074,6.092789,6.579458,5.96452,5.406172,5.2854476,5.2137675,5.1571784,4.2819295,3.9159849,4.2027044,4.115934,4.478106,4.074435,4.0404816,4.67051,5.4212623,4.4894238,4.0291634,3.1048703,1.7014539,0.7394345,0.90543,0.90920264,0.754525,0.59230214,0.69793564,0.6828451,0.7507524,0.754525,0.6526641,0.4979865,0.5772116,0.40367088,0.21881226,0.1659955,0.30181,0.27540162,0.124496624,0.0150905,0.0,0.0,0.0,0.0150905,0.03772625,0.0452715,0.00754525,0.0,0.0,0.030181,0.071679875,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.018863125,0.06413463,0.033953626,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0452715,0.116951376,0.15845025,0.18863125,0.30935526,0.4979865,0.6149379,0.68661773,0.7432071,0.7696155,0.8337501,1.1091517,1.5052774,1.8221779,1.7429527,1.327964,1.0412445,0.573439,0.41876137,0.5055317,0.67152727,0.6790725,0.7696155,0.7167987,0.55457586,0.4376245,0.67152727,0.88279426,1.0223814,1.418507,2.1994405,3.2746384,3.8480775,4.8138695,5.4250345,5.4363527,5.1043615,4.5007415,3.7084904,3.0746894,2.8256962,3.0709167,2.637065,1.9504471,1.3732355,0.9507015,0.4074435,0.116951376,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.011317875,0.003772625,0.00754525,0.0452715,0.06413463,0.06413463,0.05281675,0.056589376,0.1358145,0.06790725,0.026408374,0.060362,0.21881226,0.55457586,0.16976812,0.071679875,0.07922512,0.1358145,0.32444575,0.15467763,0.090543,0.08299775,0.0754525,0.00754525,0.03772625,0.13204187,0.150905,0.0754525,0.018863125,0.003772625,0.0,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.003772625,0.0150905,0.03772625,0.120724,0.26031113,0.39989826,0.422534,0.3055826,0.23390275,0.23013012,0.271629,0.29426476,0.36594462,0.56212115,0.633801,0.5696664,0.573439,0.633801,0.7205714,0.91674787,1.2261031,1.5731846,2.0900342,2.7125173,3.2444575,3.5424948,3.4896781,3.6066296,3.8254418,3.9612563,4.0593443,4.4177437,4.1272516,4.0706625,3.9386206,3.5839937,3.029418,2.565385,2.2220762,2.2069857,2.173032,1.2034674,1.5203679,1.6788181,1.297783,0.65643674,0.70170826,0.32444575,0.33576363,0.39989826,0.32821837,0.10186087,0.17731337,0.18485862,0.18485862,0.20372175,0.23013012,0.20372175,0.20372175,0.23767537,0.271629,0.23013012,0.120724,0.11317875,0.17354076,0.35085413,0.7469798,1.1619685,1.267602,1.20724,1.0940613,1.0336993,1.20724,1.448688,1.7580433,2.1881225,2.8521044,3.4594972,4.357382,5.3948536,6.4738245,7.5565677,8.507269,9.756008,11.0613365,12.174261,12.864652,13.343775,14.852824,17.033401,19.334703,21.043703,21.164427,21.511507,21.93027,22.537663,23.737356,26.08393,28.649315,31.478783,34.459156,37.27731,38.86558,40.023777,40.98957,41.604507,41.329105,41.381924,40.993343,40.793396,40.834892,40.5859,37.484802,33.504684,30.407358,28.905853,28.660633,25.544443,24.141027,23.307278,22.49239,21.75673,21.605824,21.605824,21.224789,20.341993,19.251705,17.867151,17.01831,16.331694,15.799753,15.777118,14.724555,14.022847,13.611631,13.389046,13.230596,13.000465,12.536433,12.151625,11.996947,12.079946,12.264804,12.66093,13.091009,13.5663595,14.302021,15.667711,16.81459,18.221779,19.734602,20.575897,21.337967,22.628204,23.895807,25.125683,26.827137,28.347504,30.230043,32.474754,34.83642,36.828365,39.03535,40.970707,42.8872,45.05646,47.74634,50.753124,53.024246,55.20105,58.76995,66.0813,69.842606,69.57852,67.797844,66.847145,68.89945,69.84638,67.53753,62.957565,57.951294,55.219913,55.257637,55.208595,54.405025,52.61303,50.02878,49.447796,50.077824,50.436222,49.776012,48.063244,46.70887,46.78432,46.886185,46.06375,43.811493,40.389725,37.111313,33.72727,30.735577,29.366114,27.8382,26.464964,24.929506,23.446865,22.77911,21.394556,19.836462,18.640541,17.708702,16.275105,14.84528,13.807808,12.925014,12.004493,10.899114,9.952185,9.175024,8.495952,7.816879,6.9869013,5.907931,5.0741806,4.3347464,3.6745367,3.187868,2.7841973,2.3126192,1.8938577,1.5618668,1.267602,1.177059,1.2336484,1.2600567,1.1996948,1.1393328,1.0336993,0.724344,0.41498876,0.211267,0.120724,0.094315626,0.056589376,0.02263575,0.0,0.0,0.0,0.0150905,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.0452715,0.056589376,0.06790725,0.026408374,0.026408374,0.033953626,0.033953626,0.026408374,0.018863125,0.026408374,0.09808825,0.124496624,0.120724,0.211267,0.73188925,1.3505998,1.4864142,1.2562841,1.4826416,2.6219745,3.8178966,6.092789,9.771099,14.475562,11.050018,5.6363015,1.8599042,0.73188925,0.6526641,0.55457586,0.47912338,0.4979865,0.513077,0.2565385,0.24522063,0.23013012,0.20372175,0.18863125,0.23013012,0.16976812,0.07922512,0.0150905,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,1.0035182,1.7278622,1.4600059,0.5017591,0.14713238,1.0676528,0.94315624,0.482896,0.1659955,0.24899325,0.181086,0.633801,1.5279131,1.9466745,0.150905,0.090543,0.1659955,0.1659955,0.0754525,0.1056335,0.32444575,0.21881226,0.06413463,0.0,0.00754525,0.271629,0.23767537,0.13958712,0.1056335,0.15467763,0.29049212,0.84884065,0.90920264,0.80734175,2.1164427,3.5877664,3.5085413,2.4559789,1.3128735,1.2940104,0.95824677,3.429316,4.217795,2.6898816,2.0372176,2.3201644,1.720317,1.7618159,2.0296721,0.18485862,0.17354076,0.19994913,0.18485862,0.11317875,0.018863125,0.018863125,0.033953626,0.030181,0.0150905,0.02263575,0.6488915,0.62625575,0.4640329,0.35462674,0.150905,0.72811663,0.7582976,0.5583485,0.41121614,0.56589377,0.4376245,0.362172,0.3772625,0.47157812,0.59607476,0.77716076,0.7394345,1.780679,3.0897799,1.7316349,1.3053282,1.6184561,2.071171,2.4182527,2.7691069,2.5691576,2.3390274,3.3953626,6.4247804,11.449917,8.088508,5.587258,4.266839,4.0593443,4.478106,4.2819295,4.093298,4.274384,4.719554,4.847823,3.2105038,1.8863125,1.3920987,1.599593,1.7618159,0.41876137,0.071679875,0.2867195,0.7205714,1.1091517,0.34330887,0.150905,0.16976812,0.20749438,0.24522063,0.8903395,1.1921495,1.4147344,2.1390784,4.2630663,5.6891184,4.2781568,2.354118,1.2562841,1.3317367,1.5128226,1.5656394,1.4600059,1.2562841,1.0978339,1.1581959,1.116697,1.1317875,1.2261031,1.2826926,1.3091009,1.3958713,1.2298758,0.9242931,1.026154,0.62248313,0.49044126,0.46026024,0.40367088,0.2565385,0.29049212,0.40367088,0.41876137,0.3470815,0.41498876,0.51684964,0.5319401,0.48666862,0.41876137,0.40367088,0.28294688,0.20749438,0.26408374,0.55457586,1.1581959,0.6149379,0.8601585,1.3166461,1.5015048,1.0223814,0.6828451,0.8865669,1.2298758,1.3355093,0.875249,0.59607476,0.35085413,0.19240387,0.1659955,0.3055826,0.9016574,1.8599042,2.7200627,3.1840954,3.1237335,4.172523,4.3385186,4.398881,4.2894745,3.097325,3.1916409,3.7198083,3.7084904,3.0746894,2.6182017,3.4368613,4.074435,4.266839,3.9310753,3.150142,3.6066296,4.5988297,5.2628117,5.670255,6.7944975,6.9982195,6.907676,7.1000805,7.3905725,6.858632,6.790725,5.9984736,5.4967146,5.3194013,4.5422406,5.2665844,5.05909,4.3875628,3.9461658,4.647874,3.4330888,2.6936543,2.0862615,1.3317367,0.20372175,0.181086,0.392353,0.55080324,0.56589377,0.5470306,0.3470815,0.38858038,0.44516975,0.44139713,0.46026024,0.6451189,0.5093044,0.29049212,0.150905,0.21503963,0.15845025,0.056589376,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.071679875,0.15845025,0.2867195,0.40367088,0.39989826,0.40367088,0.35462674,0.3772625,0.56212115,0.9393836,1.2562841,1.0336993,0.6488915,0.36971724,0.362172,0.35462674,0.67152727,1.026154,1.2789198,1.4298248,2.5201135,2.5729303,1.9693103,1.3430545,1.5845025,1.8749946,1.6524098,1.2713746,1.0940613,1.4939595,2.5502944,3.942393,5.1534057,5.836251,5.836251,5.6589375,4.9534564,4.236658,3.6254926,2.837014,2.3126192,1.9089483,1.4562333,0.9205205,0.44516975,0.22258487,0.120724,0.06413463,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.011317875,0.011317875,0.00754525,0.00754525,0.03772625,0.030181,0.033953626,0.094315626,0.271629,0.6111652,0.24522063,0.06790725,0.030181,0.15467763,0.543258,0.29426476,0.19994913,0.20749438,0.20749438,0.0452715,0.041498873,0.094315626,0.13204187,0.124496624,0.05281675,0.011317875,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.003772625,0.0,0.003772625,0.011317875,0.0150905,0.011317875,0.0150905,0.011317875,0.011317875,0.003772625,0.003772625,0.011317875,0.011317875,0.026408374,0.05281675,0.0754525,0.0754525,0.06413463,0.0754525,0.094315626,0.1056335,0.09808825,0.07922512,0.09808825,0.15467763,0.241448,0.32067314,0.19240387,0.17731337,0.32821837,0.5017591,0.34330887,0.55080324,0.8299775,1.2110126,1.50905,1.3015556,1.2751472,1.3241913,1.4373702,1.5920477,1.7655885,1.4977322,1.7278622,1.8070874,1.5807298,1.3845534,1.0978339,1.0299267,1.0902886,0.97710985,0.181086,0.2867195,0.29803738,0.23767537,0.16222288,0.1659955,0.13204187,0.06790725,0.150905,0.28294688,0.120724,0.10186087,0.1358145,0.19994913,0.2565385,0.24522063,0.18485862,0.1659955,0.21503963,0.30935526,0.35839936,0.26408374,0.2678564,0.38103512,0.6828451,1.327964,1.6222287,1.3128735,0.9242931,0.7092535,0.65643674,0.9205205,1.3241913,1.780679,2.293756,2.9351022,3.3689542,4.2291126,5.0741806,5.7192993,6.277648,7.0548086,8.009283,8.959985,9.718282,10.106862,10.182315,11.23865,12.600568,13.804035,14.622695,14.245432,14.456699,15.603577,17.852062,21.187061,24.722012,27.408121,29.841463,32.240852,34.428974,36.485058,37.967697,39.129665,40.15959,41.14802,42.600483,43.61532,44.39248,44.860283,44.649017,41.185745,37.605526,34.870373,33.165146,31.916407,29.852781,28.626678,27.509981,26.182018,24.718239,23.824127,23.035648,22.518799,22.009495,20.8098,19.870417,19.368656,19.029121,19.006485,19.885506,18.75372,18.018057,17.697384,17.440845,16.531643,16.825907,15.924251,15.060319,14.690601,14.471789,14.618922,14.803781,14.886778,14.856597,14.856597,15.433809,15.377219,15.690348,16.290195,15.99593,15.716756,16.320375,17.157898,17.976559,18.89708,20.440083,22.503708,24.910643,27.23458,28.807764,30.456402,31.867363,32.919926,33.81781,35.100502,37.009453,38.484547,40.14073,43.754906,52.28481,54.186214,53.81272,53.669365,55.223686,58.905766,60.199776,59.256622,57.125088,54.884148,53.64673,54.604973,55.84617,54.97092,51.29261,45.82985,44.58488,45.554447,48.89322,52.590393,52.473442,51.956593,50.17591,47.735023,45.162094,42.890972,39.66538,36.869865,33.998898,31.74664,32.010723,31.539145,30.490355,29.151073,28.113602,28.256962,26.781864,25.03514,23.533634,22.311304,20.904116,19.349794,17.987877,16.716501,15.475307,14.25675,12.543978,11.434827,10.63503,9.88805,8.971302,7.828197,6.8963585,6.0362,5.221313,4.561104,4.074435,3.6368105,3.1727777,2.6785638,2.214531,2.0749438,2.11267,2.0560806,1.8485862,1.6637276,1.3619176,0.9620194,0.58475685,0.31312788,0.17354076,0.120724,0.06790725,0.03772625,0.026408374,0.0,0.0,0.018863125,0.030181,0.030181,0.02263575,0.018863125,0.00754525,0.0,0.0,0.0,0.07922512,0.10186087,0.11317875,0.10186087,0.0,0.02263575,0.02263575,0.00754525,0.0,0.0,0.018863125,0.018863125,0.011317875,0.018863125,0.03772625,0.7922512,1.5165952,1.3128735,0.49044126,0.5772116,1.4524606,2.4823873,5.149633,8.899622,11.159425,9.325929,5.406172,2.1541688,0.7092535,0.5998474,0.5470306,0.422534,0.32444575,0.30935526,0.3772625,0.7167987,0.62248313,0.35085413,0.116951376,0.1056335,0.06413463,0.02263575,0.00754525,0.011317875,0.00754525,0.00754525,0.00754525,0.00754525,0.003772625,0.0150905,0.0,0.3772625,0.5281675,0.392353,0.20749438,0.48666862,1.6222287,2.6672459,1.9466745,0.26408374,0.8865669,0.7394345,1.3694628,1.9240388,1.7957695,0.62625575,0.331991,0.754525,0.7582976,0.23013012,0.0452715,0.00754525,0.0,0.0,0.00754525,0.030181,0.2263575,0.32821837,0.35839936,0.362172,0.41121614,0.5583485,1.0072908,1.116697,1.4449154,3.7386713,1.9202662,2.8294687,2.848332,1.6863633,2.3805263,0.7092535,0.56589377,0.58475685,0.3772625,0.55080324,0.5357128,0.8186596,1.3920987,1.6712729,0.48666862,0.1961765,0.44139713,0.6451189,0.5055317,0.030181,0.030181,0.030181,0.02263575,0.033953626,0.1056335,0.02263575,0.26408374,1.0035182,1.6146835,0.68661773,0.35839936,0.5394854,0.73566186,0.70170826,0.45648763,0.3470815,0.40367088,0.40367088,0.35085413,0.47157812,0.5583485,0.55080324,1.7354075,2.9652832,0.67152727,1.0751982,2.5767028,4.4743333,5.8098426,5.372218,7.201941,8.280911,9.522105,10.401127,8.971302,3.832987,3.5387223,5.3269467,7.405663,8.956212,8.469543,5.772116,3.289729,2.11267,2.0145817,1.5015048,1.6373192,3.4745877,6.156924,6.911449,1.6260014,0.120724,0.0,0.0,0.0,0.011317875,0.02263575,0.02263575,0.011317875,0.0,0.14713238,0.19994913,0.1961765,0.22258487,0.44139713,0.9318384,1.4449154,1.9844007,2.625747,3.5387223,3.429316,2.7691069,2.191895,2.1013522,2.686109,2.7351532,2.535204,2.4522061,2.4786146,2.2598023,2.052308,2.2560298,2.1013522,1.5128226,1.0978339,1.086516,0.8903395,0.6111652,0.3772625,0.36594462,0.4376245,0.55080324,0.6111652,0.5998474,0.55080324,0.513077,0.392353,0.28294688,0.3055826,0.6111652,0.40367088,0.26031113,0.48666862,1.0450171,1.5731846,0.76584285,0.56589377,1.0223814,1.5467763,0.9016574,0.66775465,0.7394345,1.0072908,1.2525115,1.1431054,0.76584285,0.5696664,0.41876137,0.27917424,0.24522063,1.5128226,2.4069347,2.9200118,3.1237335,3.1576872,4.9044123,4.881777,4.5535583,4.3686996,3.7688525,3.218049,3.5387223,4.1197066,4.376245,3.7537618,3.6934,3.6783094,3.7952607,3.772625,2.9916916,4.112161,4.3385186,4.4931965,4.878004,5.2967653,6.247467,6.8963585,7.213259,7.1264887,6.515323,6.515323,5.873977,4.8968673,3.904667,3.2331395,2.516341,2.2899833,2.3578906,2.7426984,3.7084904,2.3767538,1.4411428,0.7922512,0.35085413,0.0452715,0.02263575,0.116951376,0.12826926,0.0452715,0.0452715,0.02263575,0.07922512,0.1659955,0.25276586,0.35085413,0.48666862,0.42630664,0.29803738,0.18863125,0.150905,0.06790725,0.018863125,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.03772625,0.060362,0.10940613,0.120724,0.1056335,0.1056335,0.23013012,0.30181,0.35839936,0.55080324,0.86770374,1.0978339,1.1581959,1.0299267,0.83752275,0.80356914,1.20724,1.1581959,1.9391292,2.4522061,2.4672968,2.625747,5.7872066,6.0626082,4.5799665,2.6446102,1.7542707,1.5958204,1.0336993,0.5470306,0.43007925,0.80734175,1.750498,2.9803739,4.172523,5.028909,5.311856,5.2137675,5.1043615,4.738417,4.1083884,3.4481792,2.6672459,2.1164427,1.6448646,1.2147852,0.8865669,0.69039035,0.48666862,0.28294688,0.11317875,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.02263575,0.041498873,0.08677038,0.16976812,0.24522063,0.23013012,0.12826926,0.056589376,0.116951376,0.3961256,0.32444575,0.331991,0.36971724,0.35085413,0.1659955,0.056589376,0.06790725,0.116951376,0.1358145,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.018863125,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.00754525,0.011317875,0.0,0.011317875,0.0150905,0.00754525,0.003772625,0.0150905,0.05281675,0.05281675,0.026408374,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.033953626,0.06413463,0.0754525,0.026408374,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.05281675,0.33953625,0.6073926,0.1056335,0.1056335,0.16976812,0.3470815,0.58098423,0.70170826,0.59230214,0.72811663,0.8563859,0.8111144,0.52062225,0.19994913,0.0754525,0.041498873,0.033953626,0.0452715,0.0452715,0.03772625,0.02263575,0.018863125,0.030181,0.19994913,0.16222288,0.34330887,0.6073926,0.23013012,0.094315626,0.09808825,0.12826926,0.14713238,0.18485862,0.23013012,0.21503963,0.24899325,0.35839936,0.52062225,0.5319401,0.48666862,0.4640329,0.48666862,0.5357128,0.33953625,0.29049212,0.32067314,0.39989826,0.5357128,0.58475685,0.7054809,0.97333723,1.4109617,1.9844007,2.9728284,3.953711,4.647874,5.0213637,5.2628117,5.873977,6.5040054,7.2924843,8.130007,8.66572,8.495952,8.601585,8.858124,9.21275,9.688101,9.910686,10.0276375,10.412445,11.351829,13.045737,15.135772,17.048492,18.995167,21.09652,23.394047,26.604551,29.128437,31.410875,34.029076,37.703613,41.759186,46.671143,50.394726,52.18295,52.59794,52.22822,49.289345,46.399513,44.426434,42.509937,41.91009,41.257427,40.12187,38.367596,36.13043,33.508453,30.543173,28.819082,28.132465,26.532871,25.800982,25.518036,25.548216,25.695349,25.695349,25.657623,25.291677,24.933279,24.393793,22.963968,22.537663,21.021067,19.519562,18.549997,18.03692,17.644567,17.640795,17.527617,17.210714,16.969267,17.320122,17.244669,17.033401,16.72782,16.127972,15.920478,15.961976,15.931795,15.8676605,16.173243,16.761772,17.244669,18.044466,19.236614,20.55326,22.213217,23.782627,25.231316,26.61587,28.090965,28.947351,29.728285,31.169428,33.617863,37.05095,35.67017,34.783604,35.462673,37.933743,41.596962,42.11004,41.687508,42.034588,43.80772,46.614555,50.681446,54.82756,54.748333,49.613792,42.083633,39.314526,40.96316,47.157814,54.03531,53.741043,51.360516,49.45534,47.338898,45.188503,44.05294,43.30596,40.567036,37.26599,34.987324,35.477764,36.40583,35.45513,33.68954,32.248398,32.331398,30.135729,28.260735,26.695095,25.468992,24.627695,23.601542,21.990631,20.432537,19.18757,18.127462,16.199652,14.369928,12.958967,11.84227,10.435081,9.25425,8.371455,7.5527954,6.700182,5.8437963,5.2590394,4.8553686,4.496969,4.0593443,3.4481792,3.0331905,2.9011486,2.8596497,2.7238352,2.335255,1.9429018,1.4713237,1.0148361,0.6375736,0.38103512,0.26031113,0.21881226,0.1961765,0.1358145,0.0,0.0,0.090543,0.15845025,0.15845025,0.120724,0.09808825,0.03772625,0.0,0.0,0.0,0.0,0.06413463,0.14335975,0.15845025,0.0,0.120724,0.1056335,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.1358145,0.2565385,0.32067314,0.32067314,0.4074435,0.5998474,1.2562841,2.4823873,4.164978,3.6783094,3.218049,2.1164427,0.7432071,0.48666862,0.573439,0.47535074,0.38480774,0.48666862,0.97710985,2.0372176,1.4335974,0.56212115,0.1056335,0.030181,0.030181,0.02263575,0.033953626,0.056589376,0.030181,0.030181,0.041498873,0.033953626,0.026408374,0.0754525,0.0,0.14335975,0.19994913,0.1358145,0.0754525,0.2678564,1.7278622,2.6295197,1.9051756,0.29803738,0.38480774,0.9808825,1.327964,1.4147344,1.5241405,2.2371666,2.1013522,0.97710985,0.18485862,0.071679875,0.0452715,0.030181,0.011317875,0.0,0.0150905,0.07922512,0.44894236,0.5696664,0.5696664,0.5357128,0.4979865,0.38858038,0.5055317,0.56212115,0.7092535,1.5279131,0.5583485,0.8526133,1.1317875,0.9997456,0.965792,0.30935526,0.2565385,0.31312788,0.2867195,0.29426476,0.8262049,1.50905,1.5807298,0.95447415,0.21881226,0.211267,0.2565385,0.271629,0.21503963,0.07922512,0.041498873,0.02263575,0.05281675,0.23013012,0.754525,0.73566186,0.7054809,0.84129536,0.94692886,0.41876137,0.21503963,0.1659955,0.27540162,0.8299775,2.4107075,2.0183544,1.297783,0.724344,0.51684964,0.66775465,0.9997456,1.0450171,1.5354583,2.1768045,1.659955,2.2598023,3.0256453,3.1312788,2.6182017,2.4031622,3.9612563,4.9232755,5.0968165,4.6327834,4.0178456,3.240685,3.289729,3.9159849,4.5120597,4.0970707,3.218049,2.1843498,1.6448646,1.8938577,2.8822856,3.7047176,4.889322,5.9532022,6.0022464,3.7009451,0.9242931,0.120724,0.049044125,0.03772625,0.0,0.02263575,0.03772625,0.026408374,0.011317875,0.03772625,0.0754525,0.090543,0.1056335,0.16222288,0.28294688,0.28294688,0.422534,0.69793564,1.0336993,1.2449663,1.1732863,1.0601076,1.0714256,1.3166461,1.8448136,1.9806281,2.0598533,2.3201644,2.686109,2.757789,2.463524,2.916239,3.289729,3.2029586,2.7087448,2.71629,1.6486372,0.6752999,0.2678564,0.20749438,0.17354076,0.18485862,0.1961765,0.1961765,0.1961765,0.3055826,0.41498876,0.47535074,0.5357128,0.73188925,0.935611,0.87902164,1.0601076,1.4977322,1.7165444,1.4675511,1.3317367,1.3166461,1.3241913,1.1581959,0.845068,0.7884786,0.8941121,1.1053791,1.3770081,1.1921495,1.0450171,0.7997965,0.482896,0.27917424,1.2562841,2.04099,2.6483827,3.1840954,3.8556228,4.447925,5.032682,5.4288073,5.541986,5.342037,5.349582,5.6061206,5.4288073,4.561104,3.1539145,2.7540162,3.6028569,4.2027044,4.1008434,3.893349,3.8443048,3.6254926,3.663219,4.3724723,6.1229706,7.360391,7.54525,7.4697976,7.2887115,6.541732,5.904158,5.7419353,5.553304,5.2137675,4.991183,4.115934,2.848332,1.8749946,1.4449154,1.3656902,0.845068,0.5281675,0.3055826,0.12826926,0.00754525,0.003772625,0.02263575,0.026408374,0.00754525,0.00754525,0.003772625,0.02263575,0.0452715,0.06790725,0.1056335,0.19240387,0.21881226,0.18863125,0.13204187,0.1056335,0.08677038,0.06413463,0.033953626,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.00754525,0.03772625,0.07922512,0.08677038,0.06413463,0.08299775,0.13958712,0.22258487,0.31312788,0.35839936,0.6187105,0.80734175,0.80734175,0.6451189,0.80734175,1.0487897,1.3091009,1.5354583,1.6939086,1.9957186,2.305074,2.5767028,2.516341,1.5505489,2.0183544,1.9504471,1.4600059,0.8337501,0.5470306,0.56212115,0.38103512,0.27917424,0.4074435,0.784706,1.3732355,2.252257,3.1916409,4.002755,4.5761943,4.930821,5.1269975,5.1232247,4.9119577,4.485651,4.055572,3.6141748,3.1048703,2.5691576,2.142851,1.7240896,1.3355093,0.97333723,0.65643674,0.43007925,0.241448,0.08677038,0.011317875,0.018863125,0.03772625,0.018863125,0.018863125,0.030181,0.033953626,0.00754525,0.011317875,0.011317875,0.00754525,0.003772625,0.011317875,0.06413463,0.05281675,0.06790725,0.124496624,0.15845025,0.08677038,0.033953626,0.030181,0.08677038,0.19994913,0.31312788,0.4640329,0.55457586,0.55457586,0.5093044,0.29049212,0.18863125,0.14713238,0.12826926,0.08677038,0.026408374,0.003772625,0.0,0.0,0.0,0.011317875,0.03772625,0.03772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.00754525,0.003772625,0.011317875,0.003772625,0.003772625,0.00754525,0.0150905,0.026408374,0.06413463,0.08677038,0.0754525,0.0452715,0.02263575,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.00754525,0.0,0.0,0.003772625,0.003772625,0.011317875,0.041498873,0.10186087,0.090543,0.03772625,0.003772625,0.003772625,0.003772625,0.003772625,0.033953626,0.27540162,0.56212115,0.3734899,0.13958712,0.060362,0.07922512,0.19240387,0.422534,0.241448,0.31312788,0.43007925,0.48666862,0.45648763,0.40367088,0.5281675,0.392353,0.0452715,0.00754525,0.00754525,0.00754525,0.003772625,0.003772625,0.00754525,0.041498873,0.12826926,0.2565385,0.30935526,0.056589376,0.030181,0.02263575,0.026408374,0.033953626,0.060362,0.07922512,0.07922512,0.10940613,0.18863125,0.29803738,0.38103512,0.392353,0.36971724,0.35462674,0.362172,0.29426476,0.2867195,0.2565385,0.21881226,0.26408374,0.24522063,0.29049212,0.49421388,0.87902164,1.4222796,2.0296721,2.6068838,3.1161883,3.4859054,3.591539,3.772625,4.0970707,4.561104,5.089271,5.5193505,5.8173876,5.824933,5.7419353,5.8136153,6.307829,6.692637,7.0246277,7.3188925,7.7150183,8.443134,10.035183,12.095036,14.2944765,16.471281,18.617905,20.69662,22.122673,23.333685,24.703148,26.55928,28.483318,31.350513,34.202618,36.66237,38.914627,41.057476,42.034588,42.67216,42.90229,41.76673,39.733288,39.17494,39.22021,39.171165,38.48832,37.45462,36.398285,35.70035,35.432495,35.334404,33.440548,32.289898,31.497646,30.905344,30.55449,29.969732,29.064302,28.339958,27.547709,25.71044,24.412657,23.32614,23.375185,24.680513,26.532871,22.820608,20.394812,19.221525,18.961214,18.980076,19.395065,18.814081,17.999193,17.323895,16.776863,16.509007,15.946886,15.486626,15.358356,15.611122,15.70921,15.845025,16.324148,17.214487,18.357594,18.8254,19.87796,21.092747,22.382984,23.967487,25.163408,26.446102,28.434275,31.007204,33.31228,31.320333,29.351023,28.479546,28.928488,30.071594,29.61888,29.264252,30.52431,33.58768,37.303715,40.05773,41.54792,40.736805,37.733795,33.795174,33.670677,37.71116,43.985035,49.278027,49.089397,47.003136,45.392223,42.879654,39.684242,37.620617,35.39854,31.565554,27.747658,25.585943,26.747911,32.248398,35.647533,38.05447,40.401043,43.464413,44.95083,45.237545,44.328342,42.22322,38.922173,34.704376,30.954388,27.657114,24.76351,22.167944,19.57615,17.222033,15.720529,14.886778,13.743673,12.355347,11.065109,9.812597,8.616675,7.5792036,6.719045,6.115425,5.670255,5.2892203,4.8629136,4.244203,3.7688525,3.361409,2.9992368,2.7238352,2.4823873,2.1051247,1.6939086,1.297783,0.90543,0.5998474,0.38103512,0.29803738,0.29049212,0.1961765,0.03772625,0.018863125,0.030181,0.041498873,0.071679875,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.041498873,0.08299775,0.07922512,0.0,0.071679875,0.09808825,0.07922512,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.05281675,0.06413463,0.06413463,0.120724,0.20749438,0.3961256,0.875249,1.9579924,5.1873593,4.8063245,2.776652,0.80734175,0.35462674,0.331991,0.2678564,0.26408374,0.52062225,1.3317367,1.7957695,1.0940613,0.45648763,0.36971724,0.58098423,0.3055826,0.38858038,0.7130261,0.94315624,0.52062225,0.2565385,0.15467763,0.120724,0.10186087,0.10186087,0.0,0.033953626,0.0452715,0.049044125,0.14713238,0.543258,1.0186088,1.569412,1.6712729,1.146878,0.1659955,0.5772116,0.76584285,0.7092535,0.7167987,1.4298248,1.6863633,0.87902164,0.32444575,0.32821837,0.19240387,0.11317875,0.049044125,0.011317875,0.00754525,0.03772625,0.20372175,0.32444575,0.32444575,0.23767537,0.20749438,0.13958712,0.150905,0.16976812,0.211267,0.392353,0.094315626,0.15845025,0.3169005,0.3961256,0.29803738,0.10940613,0.10186087,0.13958712,0.14713238,0.120724,0.5696664,0.80356914,0.724344,0.43007925,0.18863125,0.22258487,0.19994913,0.16976812,0.14335975,0.10186087,0.060362,0.033953626,0.033953626,0.120724,0.41121614,0.40367088,0.35839936,0.3470815,0.35085413,0.23013012,0.4640329,1.1431054,3.3727267,5.9117036,5.198677,3.9574835,2.867195,2.6521554,3.4066803,4.5912848,3.0105548,2.6823363,2.9992368,3.338773,3.059599,3.1576872,3.2633207,3.2029586,3.3764994,4.7572803,7.0284004,6.590776,5.4401255,4.8138695,5.1760416,4.2027044,2.8785129,2.0673985,2.003264,2.2786655,2.7841973,2.7841973,2.2673476,1.6825907,1.9429018,2.372981,2.6634734,2.7804246,2.4484336,1.177059,0.3055826,0.049044125,0.02263575,0.018863125,0.0,0.011317875,0.0150905,0.011317875,0.00754525,0.0452715,0.030181,0.02263575,0.033953626,0.06413463,0.116951376,0.0754525,0.09808825,0.19240387,0.3055826,0.35085413,0.3470815,0.32821837,0.44516975,0.7582976,1.2562841,1.3732355,1.4109617,1.5656394,1.8523588,2.123988,1.8938577,2.082489,2.4371157,2.897376,3.5689032,4.146115,2.4597516,1.1091517,0.91297525,0.935611,0.7582976,0.44516975,0.20749438,0.11317875,0.08677038,0.2565385,0.3772625,0.4678055,0.52062225,0.5055317,0.58475685,0.6828451,0.9393836,1.2638294,1.3053282,1.6939086,1.7165444,1.629774,1.6033657,1.7240896,1.5052774,0.9808825,0.70170826,0.784706,0.8941121,0.7092535,0.6451189,0.5885295,0.482896,0.32821837,0.7167987,1.539231,2.1088974,2.505023,3.5689032,4.3309736,5.3609,6.156924,6.537959,6.643593,6.5266414,6.6058664,6.458734,5.7494807,4.22534,3.5160866,3.832987,4.3007927,4.7535076,5.692891,5.292993,4.859141,4.123479,3.6745367,4.949684,5.9984736,7.586749,8.461998,8.492179,8.669493,6.9680386,5.885295,5.372218,5.2364035,5.1571784,4.425289,2.9049213,1.5241405,0.7205714,0.43007925,0.42630664,0.3055826,0.23767537,0.21881226,0.071679875,0.06413463,0.07922512,0.071679875,0.041498873,0.018863125,0.026408374,0.03772625,0.030181,0.0150905,0.018863125,0.049044125,0.071679875,0.120724,0.16222288,0.10940613,0.05281675,0.030181,0.018863125,0.003772625,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.003772625,0.0,0.00754525,0.00754525,0.003772625,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.003772625,0.02263575,0.049044125,0.056589376,0.033953626,0.120724,0.18863125,0.181086,0.14335975,0.1961765,0.44516975,0.59230214,0.5281675,0.32444575,0.43385187,0.65643674,0.845068,0.98465514,1.1846043,1.6109109,1.720317,1.6260014,1.2902378,0.5583485,0.46026024,0.39989826,0.31312788,0.2263575,0.24522063,0.33576363,0.28294688,0.26031113,0.362172,0.63002837,0.94315624,1.5769572,2.3767538,3.1840954,3.8556228,4.353609,4.659192,4.817642,4.881777,4.8742313,4.7308717,4.659192,4.3611546,3.7877154,3.1614597,2.6710186,2.252257,1.8523588,1.4675511,1.1280149,0.7507524,0.45648763,0.28294688,0.20749438,0.1659955,0.124496624,0.10940613,0.08677038,0.060362,0.03772625,0.041498873,0.030181,0.018863125,0.011317875,0.0150905,0.0452715,0.056589376,0.120724,0.18863125,0.071679875,0.02263575,0.011317875,0.030181,0.06790725,0.08677038,0.181086,0.31312788,0.44139713,0.55457586,0.66775465,0.38858038,0.18485862,0.11317875,0.16222288,0.26408374,0.271629,0.15845025,0.056589376,0.0150905,0.0,0.003772625,0.03772625,0.041498873,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.0150905,0.00754525,0.0,0.0,0.00754525,0.018863125,0.041498873,0.0452715,0.060362,0.06790725,0.056589376,0.030181,0.0150905,0.00754525,0.003772625,0.0,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0150905,0.06413463,0.181086,0.1961765,0.094315626,0.018863125,0.00754525,0.00754525,0.0,0.03772625,0.24522063,0.49044126,0.3961256,0.14713238,0.041498873,0.018863125,0.05281675,0.150905,0.06413463,0.12826926,0.20749438,0.23390275,0.20372175,0.3470815,0.56212115,0.4678055,0.124496624,0.00754525,0.0452715,0.049044125,0.030181,0.00754525,0.0,0.0,0.049044125,0.094315626,0.094315626,0.00754525,0.0150905,0.018863125,0.026408374,0.0452715,0.0754525,0.06790725,0.041498873,0.049044125,0.1056335,0.181086,0.241448,0.29049212,0.29803738,0.271629,0.2565385,0.1961765,0.20749438,0.16976812,0.08677038,0.09808825,0.0754525,0.090543,0.18863125,0.41121614,0.7884786,1.1846043,1.569412,1.9768555,2.3465726,2.516341,2.6672459,2.7653341,2.837014,2.9464202,3.2105038,3.5877664,3.6745367,3.6292653,3.6443558,3.9348478,4.244203,4.4818783,4.659192,4.851596,5.1798143,6.0211096,7.326438,8.993938,10.955703,13.170234,15.294222,16.961721,18.289686,19.455427,20.69662,21.722775,22.628204,23.514772,24.650331,26.464964,28.256962,30.192318,32.45212,34.768513,36.443558,36.63596,37.371624,37.662117,37.435757,37.541393,36.832138,36.481285,36.209656,35.87389,35.458904,34.093212,33.380184,32.844475,32.297443,31.807001,30.652578,29.784874,29.139755,28.32487,26.61587,24.80501,24.348522,24.85028,25.8538,26.853544,24.107073,20.945614,19.010258,18.674494,19.081938,18.851807,18.30855,17.923742,17.784155,17.57666,16.739138,16.105335,15.720529,15.588487,15.656394,15.62244,15.712983,16.01102,16.539188,17.248442,17.682293,18.429274,19.43279,20.60985,21.862362,23.137508,24.593742,26.495146,28.521046,29.769783,28.015512,25.453901,23.48459,22.590479,22.322622,21.817091,22.035902,23.329912,25.502945,27.804247,28.807764,28.747402,28.079647,27.426983,27.604298,29.600016,34.04794,38.72222,41.525284,40.495358,38.582638,38.21669,37.57157,36.156837,34.828873,31.788137,26.208426,20.62494,17.022083,16.867407,22.07363,25.808527,28.675722,31.652325,36.107796,40.72926,44.71315,47.9727,50.206093,50.881393,49.232758,45.769485,41.185745,36.164383,31.361832,27.359077,23.020557,19.595015,17.440845,16.01102,14.671739,13.290957,12.027128,10.982111,10.216269,9.208978,8.228095,7.3415284,6.6134114,6.096562,5.4703064,4.8327327,4.327201,3.8669407,3.1237335,2.8219235,2.4672968,2.1541688,1.8674494,1.4675511,0.9808825,0.6488915,0.44516975,0.32821837,0.23390275,0.0452715,0.0,0.0,0.003772625,0.02263575,0.003772625,0.0,0.0,0.011317875,0.06413463,0.071679875,0.116951376,0.09808825,0.033953626,0.056589376,0.07922512,0.09808825,0.08677038,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.041498873,0.071679875,0.2565385,0.9016574,4.346064,5.349582,4.0178456,1.6448646,0.7054809,0.51684964,0.28294688,0.1659955,0.41498876,1.3656902,2.1051247,2.1164427,1.7240896,1.1544232,0.5357128,0.23767537,0.3470815,0.84129536,1.4675511,1.7391801,0.94692886,0.56589377,0.41876137,0.3772625,0.38103512,0.0,0.0,0.0,0.018863125,0.12826926,0.45648763,0.3169005,0.5281675,0.9318384,1.0525624,0.08677038,0.55457586,0.5998474,0.362172,0.13958712,0.38103512,0.66775465,0.47157812,0.3169005,0.3169005,0.17354076,0.10186087,0.0452715,0.018863125,0.018863125,0.02263575,0.030181,0.094315626,0.08677038,0.0150905,0.00754525,0.011317875,0.00754525,0.003772625,0.011317875,0.060362,0.2263575,0.18485862,0.17731337,0.20749438,0.07922512,0.033953626,0.033953626,0.049044125,0.05281675,0.033953626,0.22258487,0.14713238,0.09808825,0.15467763,0.17731337,0.19240387,0.17731337,0.14713238,0.11317875,0.08299775,0.056589376,0.033953626,0.05281675,0.24522063,0.8526133,0.7507524,0.35462674,0.120724,0.35085413,1.177059,3.1727777,3.9763467,6.0626082,8.571404,7.3151197,5.5382137,3.99521,3.4934506,4.3083377,6.1908774,5.4250345,5.753253,6.247467,6.349328,5.855114,5.100589,4.4441524,4.323428,5.4438977,8.778898,8.6732645,6.375736,4.5724216,4.2404304,4.6516466,3.531177,2.293756,1.3619176,0.98465514,1.237421,2.0749438,2.3088465,1.8184053,0.9922004,0.7432071,0.68661773,0.38858038,0.150905,0.06413463,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.0452715,0.02263575,0.0150905,0.011317875,0.0150905,0.02263575,0.030181,0.03772625,0.0452715,0.060362,0.094315626,0.116951376,0.08677038,0.16222288,0.43385187,0.9280658,1.0525624,1.0299267,1.0072908,1.116697,1.4713237,1.2864652,1.1808317,1.2940104,1.8599042,3.2520027,4.768598,3.6028569,2.2975287,2.123988,3.0746894,2.8747404,1.9429018,1.1242423,0.7130261,0.43007925,0.49044126,0.45648763,0.44516975,0.452715,0.35462674,0.31312788,0.44516975,0.6149379,0.724344,0.69039035,1.237421,1.4373702,1.4524606,1.5128226,1.8938577,2.1843498,1.8033148,1.3656902,1.0902886,0.784706,0.422534,0.32067314,0.362172,0.43007925,0.41121614,0.48666862,1.3053282,1.81086,1.9881734,2.8634224,4.214022,5.251494,6.058836,6.934085,8.390318,8.465771,7.8432875,7.2962565,6.8737226,5.885295,5.8437963,5.855114,5.50426,5.040227,5.372218,5.0779533,4.5422406,3.591539,2.704972,3.0030096,3.7499893,5.824933,7.575431,8.507269,9.303293,7.699928,6.2399216,5.311856,4.90064,4.5724216,3.9159849,2.6182017,1.388326,0.65643674,0.5394854,0.7167987,0.6413463,0.5998474,0.5772116,0.27917424,0.2867195,0.241448,0.15845025,0.07922512,0.03772625,0.1056335,0.24899325,0.23767537,0.07922512,0.0,0.003772625,0.0150905,0.06790725,0.12826926,0.07922512,0.0150905,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.0452715,0.03772625,0.018863125,0.00754525,0.00754525,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.02263575,0.094315626,0.15467763,0.17731337,0.15845025,0.12826926,0.06790725,0.124496624,0.14713238,0.094315626,0.0150905,0.06790725,0.24899325,0.38480774,0.43385187,0.48666862,0.9393836,0.77338815,0.62248313,0.7922512,1.2449663,1.569412,1.3732355,0.8903395,0.36971724,0.0754525,0.041498873,0.03772625,0.05281675,0.090543,0.18485862,0.29803738,0.29426476,0.2565385,0.26408374,0.38858038,0.56212115,1.1129243,1.9051756,2.704972,3.187868,3.7763977,4.195159,4.346064,4.4101987,4.817642,5.089271,5.2326307,5.0553174,4.5233774,3.7914882,3.5047686,3.2029586,2.9426475,2.686109,2.3201644,1.7693611,1.8146327,1.8976303,1.6184561,0.73188925,0.724344,0.7054809,0.62625575,0.49421388,0.392353,0.33576363,0.23390275,0.16976812,0.1659955,0.17354076,0.18485862,0.1659955,0.21881226,0.28294688,0.10940613,0.056589376,0.05281675,0.05281675,0.041498873,0.041498873,0.12826926,0.1659955,0.2263575,0.35462674,0.56589377,0.41121614,0.23390275,0.17354076,0.27540162,0.5017591,0.513077,0.35085413,0.18485862,0.094315626,0.056589376,0.018863125,0.0452715,0.05281675,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0,0.0,0.0,0.00754525,0.018863125,0.033953626,0.026408374,0.033953626,0.041498873,0.0452715,0.02263575,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.090543,0.24899325,0.3169005,0.2263575,0.13204187,0.07922512,0.02263575,0.003772625,0.026408374,0.13958712,0.27917424,0.2678564,0.1358145,0.071679875,0.041498873,0.03772625,0.06413463,0.026408374,0.071679875,0.14335975,0.17354076,0.1056335,0.362172,0.62248313,0.59230214,0.29803738,0.08299775,0.2565385,0.3734899,0.331991,0.15845025,0.02263575,0.003772625,0.0,0.0,0.003772625,0.011317875,0.06413463,0.090543,0.1056335,0.120724,0.1358145,0.124496624,0.08677038,0.07922512,0.10940613,0.13204187,0.15467763,0.19240387,0.20749438,0.19240387,0.1659955,0.10186087,0.1056335,0.08299775,0.02263575,0.018863125,0.011317875,0.0150905,0.041498873,0.11317875,0.27917424,0.49044126,0.7130261,0.965792,1.2223305,1.4147344,1.599593,1.6373192,1.6071383,1.6184561,1.8184053,2.1390784,2.354118,2.4899325,2.6106565,2.7804246,2.9916916,3.1539145,3.270866,3.3689542,3.5047686,3.7575345,4.236658,5.2552667,6.677546,7.9262853,10.001229,11.84227,13.449409,14.913187,16.41092,17.799244,18.617905,19.232841,19.934551,20.934296,21.55678,22.639523,24.386248,26.75923,29.467974,31.584417,33.195328,33.847992,34.244118,36.239838,35.191048,34.802467,34.195072,33.25946,32.65584,31.71646,30.935526,29.871645,28.521046,27.30626,26.510237,26.087702,25.650078,24.95214,23.865625,22.933788,23.16769,23.609087,23.744902,23.488363,21.835953,19.398838,17.957695,18.044466,18.934805,18.097282,17.074902,16.667458,16.950403,17.255987,16.350557,15.943113,15.79598,15.75071,15.746937,15.871433,16.143063,16.433554,16.693865,16.97304,17.569115,18.248188,19.047983,19.972277,21.013521,22.209444,23.401592,24.60506,25.43881,25.133228,23.631723,21.34174,19.568605,18.734856,18.372684,18.632996,19.568605,20.485353,21.092747,21.507734,21.617142,20.870161,20.175999,20.424992,22.4773,24.578651,27.60807,30.203636,31.33165,30.301723,29.569836,30.618624,32.17672,33.202873,32.863335,28.31355,21.83218,15.660167,11.378237,9.910686,13.419228,15.569623,16.897587,18.485863,21.964222,26.600779,31.512737,36.503918,41.140476,44.799923,47.286083,47.01068,44.58111,40.778305,36.586918,32.935017,28.566317,24.672968,21.722775,19.451654,17.338985,15.633758,14.1926155,13.04951,12.419481,11.514051,10.446399,9.461743,8.605357,7.7225633,6.8699503,5.994701,5.2779026,4.617693,3.6368105,3.2067313,2.8332415,2.6219745,2.463524,2.0598533,1.4826416,1.1053791,0.76207024,0.4376245,0.30181,0.15845025,0.090543,0.060362,0.049044125,0.041498873,0.0754525,0.071679875,0.03772625,0.011317875,0.06413463,0.071679875,0.1961765,0.1659955,0.011317875,0.056589376,0.07922512,0.09808825,0.094315626,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.003772625,0.003772625,0.06790725,0.34330887,2.1768045,3.6066296,3.482133,2.1390784,1.4147344,1.4071891,0.784706,0.2565385,0.26031113,0.9922004,1.7957695,2.3163917,2.3314822,1.8372684,1.0450171,0.52062225,0.3734899,0.6413463,1.2336484,1.9542197,1.6260014,1.20724,0.845068,0.69793564,0.9318384,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.018863125,0.041498873,0.06413463,0.056589376,0.84884065,0.7997965,0.513077,0.2678564,0.011317875,0.003772625,0.00754525,0.0150905,0.011317875,0.0,0.060362,0.16222288,0.19994913,0.15467763,0.094315626,0.116951376,0.14335975,0.14335975,0.1056335,0.033953626,0.094315626,0.10186087,0.060362,0.030181,0.15845025,0.6488915,0.9280658,0.8526133,0.47535074,0.06413463,0.026408374,0.018863125,0.02263575,0.026408374,0.0150905,0.026408374,0.03772625,0.060362,0.08677038,0.120724,0.1358145,0.13958712,0.10940613,0.06413463,0.041498873,0.033953626,0.018863125,0.21503963,0.7432071,1.6561824,1.6675003,0.94692886,0.91297525,1.961765,3.4934506,6.9680386,7.1604424,6.8058157,7.039718,7.413208,5.9909286,4.466788,3.3123648,3.097325,4.485651,6.6020937,8.20546,8.816625,8.582722,8.307321,7.1566696,5.613666,4.8063245,5.80607,9.612649,5.8890676,2.8709676,1.4977322,1.4562333,1.1921495,1.1695137,1.5920477,1.7089992,1.2223305,0.2565385,0.14713238,0.120724,0.124496624,0.120724,0.08299775,0.03772625,0.011317875,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0,0.00754525,0.018863125,0.02263575,0.03772625,0.03772625,0.030181,0.02263575,0.02263575,0.011317875,0.0150905,0.0150905,0.0150905,0.018863125,0.026408374,0.026408374,0.018863125,0.06790725,0.25276586,0.66020936,0.83752275,0.9280658,0.90920264,0.9016574,1.1732863,0.9997456,0.814887,0.7092535,0.9393836,1.9730829,4.187614,4.459243,3.5802212,2.9539654,4.5950575,4.745962,3.6368105,2.5125682,1.7882242,1.0714256,0.9997456,0.87147635,0.7054809,0.55457586,0.5357128,0.45648763,0.4678055,0.41876137,0.2867195,0.19994913,0.45648763,0.754525,1.0789708,1.4826416,2.1051247,2.565385,2.5993385,2.203213,1.5467763,0.9922004,0.5093044,0.32821837,0.30935526,0.36594462,0.43007925,0.52439487,1.2562841,1.7769064,1.9278114,2.2711203,4.146115,5.062863,5.6778007,6.8246784,9.522105,9.933322,8.548768,7.3151197,6.8850408,6.6360474,7.488661,7.696155,6.511551,4.45547,3.338773,3.3764994,3.0746894,2.7841973,2.5201135,1.9655377,2.2484846,3.1350515,4.7572803,6.6586833,7.8017883,7.5188417,6.5455046,5.462761,4.5460134,3.7914882,3.0746894,2.1503963,1.3732355,0.98842776,1.1355602,1.2638294,1.1393328,0.98465514,0.80734175,0.41876137,0.44516975,0.32821837,0.18863125,0.090543,0.041498873,0.181086,0.46026024,0.45648763,0.15845025,0.0,0.0150905,0.030181,0.03772625,0.030181,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.071679875,0.05281675,0.026408374,0.00754525,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.033953626,0.056589376,0.20372175,0.32821837,0.362172,0.3055826,0.22258487,0.11317875,0.06413463,0.0452715,0.041498873,0.0452715,0.08299775,0.30181,0.513077,0.7167987,1.1242423,1.9844007,1.4147344,1.0110635,1.4335974,2.372981,2.0372176,1.3543724,0.663982,0.19994913,0.06790725,0.02263575,0.0150905,0.018863125,0.03772625,0.07922512,0.18863125,0.22258487,0.1961765,0.150905,0.16222288,0.35462674,1.20724,2.2296214,2.9351022,2.8407867,3.3425457,3.7575345,3.8178966,3.8556228,4.8100967,5.7872066,5.6098933,5.20245,4.8742313,4.3309736,4.2102494,4.085753,3.9499383,3.7613072,3.4594972,2.8521044,3.338773,3.7613072,3.338773,1.6939086,1.7580433,1.6976813,1.5015048,1.2223305,0.97710985,0.845068,0.6488915,0.56589377,0.6111652,0.6488915,0.5583485,0.422534,0.3772625,0.3961256,0.29049212,0.20749438,0.16976812,0.10940613,0.03772625,0.033953626,0.14713238,0.1056335,0.05281675,0.10186087,0.34330887,0.42630664,0.38858038,0.32444575,0.35462674,0.63002837,0.694163,0.58098423,0.41121614,0.26031113,0.1659955,0.056589376,0.05281675,0.06413463,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.02263575,0.026408374,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.1056335,0.29803738,0.43007925,0.3734899,0.3055826,0.24522063,0.056589376,0.011317875,0.0,0.0,0.018863125,0.10186087,0.10186087,0.10940613,0.10186087,0.094315626,0.150905,0.09808825,0.1056335,0.18485862,0.271629,0.26408374,0.5055317,0.73566186,0.73188925,0.5093044,0.31312788,0.62248313,0.8941121,0.8224323,0.43385187,0.071679875,0.02263575,0.00754525,0.003772625,0.011317875,0.05281675,0.16222288,0.211267,0.241448,0.26408374,0.27540162,0.26031113,0.1961765,0.15845025,0.15845025,0.1358145,0.15845025,0.17354076,0.181086,0.1659955,0.1056335,0.05281675,0.033953626,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.05281675,0.10940613,0.1659955,0.23767537,0.34330887,0.4640329,0.55080324,0.66775465,0.8337501,1.0412445,1.2713746,1.5316857,1.7957695,2.0372176,2.2711203,2.505023,2.746471,2.9200118,3.0105548,3.0709167,3.0860074,3.1237335,3.6481283,4.3422914,4.115934,5.5797124,6.9227667,8.431817,10.148361,11.879996,13.958713,16.188334,18.519815,20.583443,21.707684,21.82841,21.790682,22.164171,23.163918,24.650331,26.578144,27.906107,28.98885,30.724258,34.56479,33.591454,33.02556,32.05977,30.890253,30.705395,29.928234,28.675722,26.197107,22.839472,20.040184,20.017548,19.938324,19.568605,18.97253,18.534906,19.11589,19.840235,20.213724,20.130728,19.893051,18.0671,16.939087,16.822134,17.614386,18.806536,17.931286,16.331694,15.343266,15.358356,15.79598,15.445127,15.354584,15.335721,15.335721,15.422491,15.773345,16.248695,16.603323,16.780636,16.946632,17.655886,18.406637,19.047983,19.696875,20.783392,21.820864,22.443346,22.699884,22.29244,20.568352,19.108345,17.795471,17.28994,17.57666,17.99542,19.168707,20.428764,20.794708,20.175999,19.353567,19.54597,18.7839,17.908651,17.80679,19.429018,19.859098,20.606077,21.553007,22.31885,22.239624,23.246916,26.321604,30.29795,33.07083,31.625916,24.378702,17.80679,12.577931,8.990166,6.9567204,8.846806,9.325929,9.092027,9.012801,10.1294985,12.098808,14.871688,17.946377,21.051247,24.1448,28.788902,32.19181,33.964943,34.161118,33.27455,31.950361,30.101774,28.034376,25.800982,23.171463,20.232588,18.104828,16.309057,14.758509,13.773854,12.992921,12.121444,11.3820095,10.642575,9.431562,8.284684,7.2396674,6.2135134,5.221313,4.3686996,3.7688525,3.338773,3.1161883,2.957738,2.5314314,1.9693103,1.5882751,1.146878,0.6752999,0.4640329,0.36971724,0.26408374,0.181086,0.1358145,0.116951376,0.18485862,0.17354076,0.09808825,0.018863125,0.0150905,0.011317875,0.1961765,0.18863125,0.003772625,0.02263575,0.05281675,0.09808825,0.10186087,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.00754525,0.003772625,0.011317875,0.1358145,0.70170826,1.297783,1.6976813,1.8749946,2.2748928,1.3543724,0.42630664,0.124496624,0.4074435,0.83752275,1.2638294,1.629774,1.8599042,1.8372684,1.0940613,0.6111652,0.4640329,0.7696155,1.6712729,1.9127209,1.5882751,1.1657411,1.0412445,1.5543215,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.02263575,0.00754525,0.018863125,0.030181,0.2867195,0.3961256,0.8903395,1.267602,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.3055826,0.8111144,0.9280658,0.58098423,0.23013012,0.29049212,0.48666862,0.58475685,0.46026024,0.1056335,0.362172,0.42630664,0.2565385,0.03772625,0.18485862,1.0751982,2.927557,2.8521044,0.90543,0.0754525,0.041498873,0.030181,0.02263575,0.0150905,0.0150905,0.0150905,0.033953626,0.06413463,0.094315626,0.1056335,0.094315626,0.08299775,0.056589376,0.030181,0.030181,0.030181,0.011317875,0.663982,1.3770081,0.23013012,1.20724,1.5052774,3.62172,6.7152724,6.6058664,7.0359454,7.2057137,6.4964604,5.1534057,4.2894745,4.398881,4.9647746,4.957229,4.2404304,3.5689032,4.436607,5.670255,5.6589375,4.889322,5.9494295,6.156924,3.7009451,1.6448646,1.0940613,1.1921495,0.38480774,0.19994913,0.23767537,0.241448,0.1056335,0.19240387,0.88279426,1.3505998,1.146878,0.18485862,0.18485862,0.211267,0.19994913,0.13204187,0.0452715,0.02263575,0.0150905,0.00754525,0.003772625,0.0150905,0.003772625,0.0,0.0,0.003772625,0.0150905,0.003772625,0.00754525,0.026408374,0.03772625,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.011317875,0.0150905,0.02263575,0.026408374,0.0150905,0.003772625,0.0,0.00754525,0.02263575,0.060362,0.21881226,0.7092535,0.97710985,0.91674787,0.8563859,0.8186596,0.73566186,0.63002837,0.55457586,0.58098423,2.2296214,3.5462675,3.2520027,1.7165444,0.94692886,2.1315331,2.8558772,3.0143273,2.5616124,1.50905,1.6335466,1.901403,1.6448646,1.0450171,1.1431054,0.7054809,0.5772116,0.51684964,0.38480774,0.150905,0.26408374,0.47157812,1.5958204,3.2670932,3.9348478,2.4710693,1.5580941,0.8903395,0.41876137,0.32067314,0.211267,0.19240387,0.20372175,0.19994913,0.1358145,0.16222288,0.8262049,1.5430037,2.0258996,2.3201644,4.564876,6.1342883,6.7643166,6.79827,7.201941,6.72659,5.873977,5.160951,4.768598,4.561104,4.085753,3.904667,3.3161373,2.6936543,3.4481792,3.92353,4.7572803,5.406172,5.323174,3.9688015,3.1840954,2.4597516,2.5314314,3.832987,6.470052,7.250985,6.356873,5.040227,3.9386206,3.0822346,2.3880715,1.6712729,1.2034674,1.1242423,1.4637785,1.5618668,1.1393328,0.58475685,0.16222288,0.0150905,0.003772625,0.0452715,0.08299775,0.0754525,0.0150905,0.08677038,0.16222288,0.150905,0.060362,0.0,0.02263575,0.056589376,0.056589376,0.033953626,0.0452715,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.090543,0.1056335,0.08299775,0.041498873,0.0150905,0.003772625,0.0,0.030181,0.094315626,0.1659955,0.20372175,0.7167987,1.1317875,1.3656902,1.8297231,1.9881734,1.6448646,1.539231,2.214531,3.9989824,1.7769064,0.67152727,0.23013012,0.1056335,0.030181,0.00754525,0.00754525,0.0150905,0.018863125,0.030181,0.07922512,0.12826926,0.14713238,0.1358145,0.1358145,0.4678055,2.4182527,4.1083884,4.478106,3.2821836,3.048281,2.9086938,2.9200118,3.5387223,5.613666,7.7150183,6.3531003,5.194905,5.379763,5.5382137,4.7950063,4.727099,4.2894745,3.4594972,3.2520027,2.8596497,2.6974268,2.5767028,2.4861598,2.6106565,2.7426984,2.4295704,1.9844007,1.599593,1.3430545,1.2223305,1.1544232,1.267602,1.5052774,1.6033657,1.1016065,0.8111144,0.66020936,0.58475685,0.5357128,0.5093044,0.38480774,0.23767537,0.120724,0.0452715,0.02263575,0.00754525,0.00754525,0.08677038,0.38103512,0.5017591,0.5696664,0.392353,0.15467763,0.41121614,0.9242931,0.9620194,0.76584285,0.5055317,0.27540162,0.07922512,0.030181,0.056589376,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.1056335,0.3961256,0.52062225,0.392353,0.41876137,0.52062225,0.1659955,0.033953626,0.0,0.0,0.003772625,0.0150905,0.0150905,0.08677038,0.19994913,0.271629,0.19994913,0.23390275,0.24522063,0.2565385,0.32444575,0.52062225,0.55457586,0.5017591,0.48666862,0.59230214,0.8224323,1.0072908,1.2261031,1.116697,0.6451189,0.120724,0.071679875,0.041498873,0.02263575,0.041498873,0.1358145,0.24899325,0.31312788,0.4074435,0.543258,0.6413463,0.56589377,0.35839936,0.19994913,0.15845025,0.18485862,0.3055826,0.38103512,0.392353,0.32444575,0.150905,0.090543,0.049044125,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.026408374,0.056589376,0.10186087,0.150905,0.19994913,0.271629,0.362172,0.4979865,0.7092535,1.0374719,1.478869,1.9164935,2.3201644,2.655928,2.897376,3.0218725,3.0897799,3.150142,3.2255943,3.3123648,3.9348478,4.327201,5.323174,6.692637,7.1566696,8.36391,10.955703,14.769827,18.934805,21.866135,23.05074,23.593996,24.506971,25.846254,26.68755,26.664913,26.676231,27.102537,28.08342,29.509472,30.59599,30.46772,30.777075,31.595734,31.38824,31.999405,31.886227,28.770039,23.118647,18.112373,17.30503,16.637276,15.954432,15.237633,14.603831,14.724555,15.422491,16.11288,16.878725,18.478317,16.573141,15.852571,16.0412,16.765545,17.546478,17.523844,17.16167,16.335466,15.260268,14.464244,14.524607,14.596286,14.407655,14.117163,14.313339,14.592513,14.966003,15.23386,15.516807,16.252468,17.497435,18.23687,18.840488,19.58747,20.658894,21.51528,21.62846,21.394556,20.862616,19.715738,18.470772,18.150099,18.678267,19.73083,20.704166,21.696367,22.179262,21.843498,20.85507,19.866644,19.987368,19.791191,19.63274,20.002459,21.53037,20.455173,19.821371,20.194862,21.175745,21.409647,22.688566,30.094229,38.37137,41.706367,33.738586,22.945105,15.562078,11.076427,8.446907,6.1041074,5.9192486,6.205968,6.6247296,6.9567204,7.066127,7.1981683,8.412953,9.49947,10.27663,11.581959,13.50977,15.762027,18.044466,20.040184,21.409647,22.311304,23.288414,23.752447,23.58645,23.148827,21.97554,20.1345,18.35382,16.739138,14.784918,13.5663595,12.709973,11.861133,10.921749,10.054046,9.250477,8.616675,7.61693,6.319147,5.4174895,4.52715,3.953711,3.4594972,2.969056,2.5804756,2.1277604,1.6750455,1.2713746,0.9393836,0.67152727,0.5357128,0.422534,0.3055826,0.19994913,0.150905,0.150905,0.150905,0.12826926,0.08677038,0.0754525,0.06413463,0.02263575,0.0,0.02263575,0.1056335,0.02263575,0.10940613,0.10940613,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.030181,0.0,0.0,0.0,0.071679875,0.10186087,0.10186087,0.27540162,1.0072908,1.3996439,0.8639311,0.271629,0.030181,0.090543,0.33576363,0.29426476,0.3772625,0.7130261,1.1883769,1.1280149,0.875249,0.814887,1.5015048,3.663219,1.539231,0.814887,0.9997456,1.539231,1.8448136,0.011317875,0.02263575,0.011317875,0.0,0.0,0.0,0.011317875,0.018863125,0.12826926,0.34330887,0.58098423,0.55457586,0.36594462,0.59230214,0.9997456,0.55080324,0.14713238,0.071679875,0.42630664,0.8262049,0.40367088,0.16222288,0.36971724,0.42630664,0.20372175,0.0452715,0.20372175,0.23013012,0.18863125,0.13958712,0.1056335,0.12826926,0.1358145,0.094315626,0.06790725,0.1961765,0.452715,0.724344,0.77338815,0.724344,1.0789708,2.3201644,2.0598533,1.1204696,0.23767537,0.05281675,0.033953626,0.02263575,0.0452715,0.071679875,0.033953626,0.030181,0.056589376,0.19994913,0.30935526,0.00754525,0.0150905,0.18863125,0.7054809,1.237421,0.9507015,1.2411937,1.8372684,2.7351532,3.561358,3.5802212,8.156415,8.529905,6.8171334,4.666737,3.2746384,3.0143273,3.3764994,3.6028569,3.2821836,2.3880715,2.323937,3.0105548,3.3425457,3.108643,2.9954643,3.3425457,2.4333432,1.4411428,0.94692886,0.94692886,0.4640329,0.18485862,0.07922512,0.071679875,0.033953626,0.1961765,0.392353,0.55457586,0.6451189,0.66020936,0.7092535,0.42630664,0.15467763,0.03772625,0.02263575,0.00754525,0.003772625,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0,0.00754525,0.018863125,0.018863125,0.0,0.011317875,0.056589376,0.0754525,0.06790725,0.09808825,0.060362,0.030181,0.011317875,0.003772625,0.003772625,0.0,0.0,0.026408374,0.1358145,0.41498876,1.1091517,1.5807298,1.3505998,0.68661773,0.58475685,0.6187105,0.55080324,0.49421388,0.4640329,0.422534,0.8563859,1.4864142,1.9806281,2.2409391,2.4107075,2.6182017,2.293756,2.3578906,2.5880208,1.6448646,1.7467253,2.2975287,2.4899325,2.082489,1.388326,1.7014539,2.0598533,2.5578396,3.3689542,4.779916,4.183841,3.1954134,2.2975287,1.7240896,1.4600059,1.0299267,0.694163,0.41498876,0.35839936,0.8941121,0.76584285,0.43385187,0.20372175,0.1358145,0.06413463,0.060362,0.271629,0.73188925,1.4147344,2.2447119,4.2592936,6.436098,7.0246277,6.462507,7.3717093,7.2472124,6.439871,5.726845,5.402399,5.281675,5.5306683,5.349582,4.779916,4.164978,4.168751,4.1574326,3.5802212,3.9763467,4.719554,3.0030096,2.444661,2.0485353,1.9240388,2.3503454,3.7348988,5.0741806,5.409944,4.9685473,4.1498876,3.5085413,2.6483827,1.841041,1.2638294,0.9695646,0.8903395,0.814887,0.49044126,0.18863125,0.033953626,0.003772625,0.011317875,0.18863125,0.211267,0.10940613,0.28294688,0.44516975,0.21881226,0.030181,0.011317875,0.0,0.02263575,0.041498873,0.07922512,0.13204187,0.19240387,0.071679875,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.026408374,0.049044125,0.08677038,0.1659955,0.30935526,0.3055826,0.24522063,0.33576363,0.55457586,0.65643674,0.60362,0.80356914,1.1393328,1.478869,1.6486372,1.7769064,1.9089483,1.8184053,1.5467763,1.3845534,0.5885295,0.271629,0.15467763,0.08677038,0.041498873,0.026408374,0.018863125,0.018863125,0.0452715,0.116951376,0.08677038,0.23390275,0.5281675,0.814887,0.79602385,0.8224323,1.4373702,2.0900342,2.3163917,1.7542707,1.5920477,1.7957695,2.2899833,3.0331905,4.0517993,4.881777,4.353609,4.1310244,4.5761943,4.745962,6.4134626,5.6815734,4.617693,4.1083884,3.8593953,3.4896781,3.1576872,2.8332415,2.5276587,2.2786655,2.11267,1.8221779,1.4260522,1.0072908,0.73188925,0.6790725,0.6451189,0.6526641,0.6790725,0.6488915,0.5093044,0.392353,0.32067314,0.29803738,0.27917424,0.25276586,0.19240387,0.13204187,0.08299775,0.056589376,0.041498873,0.030181,0.026408374,0.05281675,0.150905,0.271629,0.3470815,0.27540162,0.13958712,0.181086,0.694163,0.7432071,0.6451189,0.51684964,0.27540162,0.090543,0.026408374,0.056589376,0.094315626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.018863125,0.00754525,0.00754525,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.08299775,0.33576363,0.38858038,0.32067314,0.39989826,0.5470306,0.35085413,0.120724,0.030181,0.00754525,0.0,0.003772625,0.003772625,0.018863125,0.049044125,0.10186087,0.17354076,0.181086,0.17731337,0.30181,0.5281675,0.663982,0.67152727,0.55080324,0.46026024,0.4979865,0.69039035,1.3430545,1.3505998,0.8941121,0.32067314,0.14713238,0.116951376,0.090543,0.060362,0.0452715,0.124496624,0.24522063,0.3055826,0.44516975,0.6526641,0.7507524,0.65643674,0.5319401,0.41876137,0.41121614,0.62248313,0.68661773,0.7922512,0.8186596,0.73188925,0.58098423,0.38103512,0.2263575,0.1056335,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.011317875,0.026408374,0.041498873,0.041498873,0.05281675,0.071679875,0.1056335,0.15845025,0.24522063,0.392353,0.58098423,0.814887,1.0789708,1.3732355,1.659955,2.0183544,2.867195,3.6783094,2.9954643,3.4594972,4.0706625,4.689373,5.0968165,4.983638,5.2364035,6.511551,8.75249,11.736636,15.067864,18.459454,21.088974,23.299732,25.148317,26.419693,26.374422,26.110338,25.695349,25.186045,24.639013,24.514517,23.752447,22.960196,22.465982,22.307531,22.99415,23.620405,22.303759,19.217752,16.588232,15.222542,14.460471,13.992666,13.63804,13.343775,13.358865,13.358865,13.555041,13.928532,14.219024,13.924759,14.007756,14.230342,14.577423,15.252723,15.297995,14.883006,14.475562,14.320885,14.464244,14.147344,13.645585,13.268322,13.249459,13.728582,13.615403,13.532406,13.494679,13.65313,14.298248,15.339493,16.263786,17.271078,18.459454,19.806282,20.719257,21.228561,21.594505,21.651094,20.775846,20.175999,20.741892,21.688822,22.515026,23.013012,25.555761,26.713957,25.767029,23.609087,22.748928,23.31105,24.371157,27.517527,32.818066,38.812767,36.51901,31.852272,27.804247,25.468992,24.031622,24.239115,27.875927,31.41842,31.358059,24.21648,16.490145,11.717773,8.993938,7.435844,6.1644692,6.458734,7.0548086,7.2396674,6.8246784,6.1116524,6.296511,6.964266,7.4094353,7.5905213,8.175279,8.6581745,9.646602,10.917976,12.193124,13.12119,14.656648,15.528125,16.150608,16.7995,17.618158,17.599297,17.912424,17.610613,16.588232,15.592259,14.683057,13.641812,12.506252,11.32542,10.167224,9.125979,8.484633,7.7640624,6.832224,5.9305663,5.0477724,4.568649,4.104616,3.5274043,2.9803739,2.6483827,2.203213,1.7089992,1.2411937,0.91674787,0.7432071,0.62248313,0.513077,0.3961256,0.29803738,0.26031113,0.20749438,0.150905,0.10940613,0.0754525,0.08299775,0.08677038,0.1056335,0.14335975,0.181086,0.17354076,0.090543,0.02263575,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.011317875,0.0,0.03772625,0.08677038,0.03772625,0.018863125,0.00754525,0.0,0.0,0.0,0.0150905,0.018863125,0.018863125,0.056589376,0.19994913,0.27917424,0.17354076,0.05281675,0.033953626,0.150905,0.22258487,0.1659955,0.12826926,0.20372175,0.44516975,0.56212115,0.8563859,1.0487897,1.1317875,1.3807807,1.1695137,1.4222796,1.7429527,1.8599042,1.6260014,0.0150905,0.011317875,0.003772625,0.0,0.00754525,0.03772625,0.13204187,0.181086,0.26031113,0.3734899,0.422534,0.29803738,0.15845025,0.46026024,1.1242423,1.539231,0.5772116,0.6111652,1.0299267,1.177059,0.33953625,0.6187105,0.62625575,0.39989826,0.09808825,0.018863125,0.14335975,0.2678564,0.36971724,0.39989826,0.3169005,0.1358145,0.116951376,0.1358145,0.1358145,0.1358145,0.181086,0.19240387,0.29049212,0.5357128,0.9242931,1.3807807,1.2223305,0.724344,0.3470815,0.7394345,0.6488915,0.41498876,0.36594462,0.44139713,0.18863125,0.049044125,0.06790725,0.1961765,0.2678564,0.0,0.003772625,2.1088974,4.4818783,5.4174895,3.3538637,3.9084394,3.4444065,3.3689542,3.9914372,4.5422406,12.200669,9.906913,5.855114,4.006528,4.093298,2.191895,1.7542707,1.8825399,1.8787673,1.2223305,1.0525624,1.4298248,1.7014539,1.6033657,1.2525115,1.388326,1.1619685,0.7997965,0.4979865,0.4074435,0.20372175,0.071679875,0.018863125,0.033953626,0.07922512,0.18863125,0.20749438,0.3169005,0.5470306,0.7507524,0.5055317,0.23767537,0.08677038,0.071679875,0.07922512,0.02263575,0.00754525,0.003772625,0.0,0.0,0.030181,0.0754525,0.094315626,0.071679875,0.03772625,0.0452715,0.094315626,0.09808825,0.049044125,0.0,0.003772625,0.026408374,0.03772625,0.033953626,0.049044125,0.030181,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.02263575,0.13204187,0.43007925,1.2034674,1.5920477,1.3317367,0.72811663,0.6451189,0.6451189,0.5319401,0.482896,0.5281675,0.55457586,0.5583485,0.62625575,0.94315624,1.4335974,1.7693611,2.04099,1.7731338,1.81086,2.2296214,2.3390274,1.5128226,1.659955,2.191895,2.5578396,2.2447119,2.1164427,2.2258487,2.6823363,3.380272,4.002755,3.9159849,3.1916409,2.2296214,1.4335974,1.1959221,0.8865669,0.52062225,0.25276586,0.21503963,0.5055317,0.7092535,0.482896,0.23767537,0.12826926,0.06413463,0.0452715,0.090543,0.32444575,0.7696155,1.3770081,3.0520537,5.0025005,6.145606,6.5568223,7.462252,8.156415,7.8395147,7.254758,6.809588,6.579458,6.722818,6.4549613,5.8928404,5.1647234,4.432834,4.3347464,3.651901,3.410453,3.361409,1.991946,2.9652832,2.6408374,2.052308,1.9844007,2.969056,4.3083377,4.8553686,4.847823,4.429062,3.6443558,2.3465726,1.2449663,0.63002837,0.47157812,0.42630664,0.5017591,0.32067314,0.116951376,0.00754525,0.0,0.026408374,0.1056335,0.17354076,0.19240387,0.1659955,0.21881226,0.094315626,0.0,0.0,0.0,0.011317875,0.0150905,0.03772625,0.071679875,0.10186087,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.02263575,0.0150905,0.00754525,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.10186087,0.15845025,0.20749438,0.26408374,0.35085413,0.482896,0.3961256,0.2565385,0.2867195,0.52439487,0.8224323,0.9205205,1.1732863,1.418507,1.5165952,1.3656902,1.5241405,1.5467763,1.3204187,0.9280658,0.6413463,0.4074435,0.3169005,0.25276586,0.1961765,0.211267,0.32444575,0.35839936,0.32821837,0.27917424,0.28294688,0.241448,0.3055826,0.51684964,0.7696155,0.7884786,0.7092535,0.8224323,1.0186088,1.1732863,1.1355602,1.2525115,1.5580941,1.8976303,2.233394,2.6106565,3.150142,3.451952,4.036709,5.1571784,6.809588,8.009283,6.8661776,5.617439,5.081726,4.6629643,4.3196554,3.9876647,3.572676,3.0709167,2.5917933,2.252257,1.9089483,1.5052774,1.0940613,0.8262049,0.7922512,0.77338815,0.7432071,0.68661773,0.60362,0.5394854,0.47912338,0.43385187,0.41121614,0.4074435,0.40367088,0.362172,0.29803738,0.24522063,0.21503963,0.16222288,0.1358145,0.12826926,0.124496624,0.1358145,0.23767537,0.31312788,0.30181,0.21881226,0.18485862,0.41876137,0.52062225,0.60362,0.6413463,0.4376245,0.16222288,0.056589376,0.0452715,0.056589376,0.018863125,0.011317875,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.02263575,0.02263575,0.018863125,0.018863125,0.026408374,0.018863125,0.011317875,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.03772625,0.1659955,0.26031113,0.27540162,0.482896,0.7922512,0.73566186,0.30935526,0.11317875,0.030181,0.0,0.0,0.00754525,0.018863125,0.030181,0.056589376,0.1659955,0.21881226,0.20749438,0.31312788,0.5470306,0.76584285,0.7092535,0.5885295,0.56212115,0.6451189,0.7205714,0.90920264,1.0676528,1.2261031,1.2487389,0.8111144,0.4376245,0.21881226,0.11317875,0.09808825,0.18485862,0.2565385,0.27540162,0.3470815,0.47912338,0.58475685,0.67152727,0.6375736,0.55457586,0.58098423,0.9695646,0.9318384,0.98842776,1.0450171,1.026154,0.8865669,0.5696664,0.35085413,0.181086,0.05281675,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.00754525,0.018863125,0.049044125,0.09808825,0.17354076,0.27917424,0.41498876,0.6073926,0.8903395,1.5316857,2.305074,2.5012503,2.6521554,3.0822346,3.6368105,4.0480266,3.9461658,3.832987,4.2819295,5.2854476,6.8397694,8.944894,12.053536,15.47908,18.829172,21.55678,22.975286,24.008986,24.808783,25.363358,25.435038,24.556017,23.443092,22.058538,20.500444,19.221525,19.010258,20.096773,20.836208,19.813826,17.240896,14.958458,13.766309,13.400364,13.215506,12.928786,12.608112,12.581704,12.193124,11.955449,11.996947,12.053536,12.004493,12.15917,12.449662,12.823153,13.241914,13.604086,13.936077,14.32843,14.618922,14.381247,13.573905,13.106099,12.879742,12.842015,12.966512,12.845788,12.917468,12.917468,12.90615,13.249459,13.800262,14.66042,15.697892,16.931541,18.531134,19.979822,21.164427,21.949133,22.232079,21.97554,22.062311,23.401592,25.363358,27.253443,28.306005,31.210926,31.780594,29.852781,26.898817,26.031113,27.155355,29.98105,35.12691,41.642235,46.999363,43.826584,38.031834,33.331142,30.992115,29.822601,27.41944,25.555761,23.646814,20.719257,15.418718,11.419736,9.329701,7.8696957,6.8774953,7.3075747,7.8244243,8.258276,8.179051,7.4773426,6.3417826,5.6513925,5.715527,5.96452,6.1795597,6.5002327,6.72659,7.1566696,7.7338815,8.356364,8.888305,9.88805,10.525623,11.080199,11.69891,12.408164,12.66093,13.245687,13.536179,13.536179,13.8719425,13.713491,13.011784,12.147853,11.276376,10.321902,9.484379,8.888305,7.967784,6.749226,5.836251,5.089271,4.568649,4.1008434,3.640583,3.2369123,2.9615107,2.625747,2.2296214,1.81086,1.4147344,1.1581959,0.995973,0.8186596,0.62625575,0.5093044,0.4376245,0.3734899,0.30935526,0.25276586,0.18485862,0.17731337,0.19994913,0.25276586,0.32821837,0.42630664,0.46026024,0.27540162,0.08677038,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.10940613,0.124496624,0.090543,0.041498873,0.018863125,0.003772625,0.06413463,0.06413463,0.0,0.0,0.071679875,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.06790725,0.11317875,0.09808825,0.056589376,0.03772625,0.1056335,0.1961765,0.4376245,0.65643674,0.73566186,0.6073926,0.7884786,1.0827434,1.3317367,1.4562333,1.4600059,0.06413463,0.124496624,0.090543,0.10940613,0.30181,0.724344,0.3734899,0.31312788,0.42630664,0.5772116,0.6375736,0.30181,0.38480774,0.73188925,1.4373702,2.8558772,0.9808825,0.9016574,1.0714256,0.7884786,0.18485862,0.73188925,0.69039035,0.38480774,0.11317875,0.16976812,0.16222288,0.23390275,0.38103512,0.56212115,0.6828451,0.2867195,0.181086,0.181086,0.23390275,0.422534,0.23767537,0.331991,0.39989826,0.3772625,0.44894236,0.29803738,0.29426476,0.30181,0.3772625,0.7582976,0.7054809,0.8262049,1.0223814,1.0223814,0.38480774,0.31312788,0.3961256,0.41121614,0.2867195,0.10940613,0.03772625,4.8666863,7.594294,6.092789,3.1350515,5.402399,3.9008942,3.029418,4.093298,5.2779026,12.717519,9.201432,4.3422914,2.6898816,3.7273536,1.8259505,0.8978847,0.67152727,0.7205714,0.43385187,0.44139713,0.69039035,0.875249,0.91674787,0.94692886,0.8865669,0.694163,0.5017591,0.33576363,0.120724,0.02263575,0.02263575,0.041498873,0.09808825,0.27917424,0.16222288,0.12826926,0.22258487,0.422534,0.63002837,0.3169005,0.14713238,0.0754525,0.06413463,0.071679875,0.02263575,0.00754525,0.00754525,0.00754525,0.018863125,0.05281675,0.10186087,0.116951376,0.08677038,0.049044125,0.05281675,0.090543,0.094315626,0.0452715,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.090543,0.27917424,0.79602385,1.1016065,1.0412445,0.7432071,0.633801,0.5583485,0.4376245,0.41121614,0.49421388,0.6111652,0.62625575,0.573439,0.6149379,0.7394345,0.7696155,1.026154,0.9620194,0.97333723,1.2411937,1.7467253,0.9922004,1.0978339,1.7429527,2.5616124,3.1048703,2.9351022,3.3350005,3.6858547,3.561358,2.7691069,2.5578396,2.1164427,1.5731846,1.2638294,1.7316349,1.7014539,1.1619685,0.59607476,0.27540162,0.24899325,0.573439,0.49421388,0.3470815,0.3734899,0.694163,0.5017591,0.39989826,0.41498876,0.5696664,0.875249,1.8976303,3.410453,4.938366,6.368191,7.956466,9.190115,9.001483,8.560086,8.337502,8.118689,7.745199,7.3490734,6.7567716,5.938112,5.0175915,4.5233774,3.92353,3.127506,2.1843498,1.2902378,2.7540162,2.5917933,2.293756,2.6672459,3.8254418,4.7874613,4.557331,3.9008942,3.2557755,2.7238352,1.9542197,1.1506506,0.573439,0.30181,0.21503963,0.31312788,0.2263575,0.094315626,0.0150905,0.03772625,0.03772625,0.026408374,0.07922512,0.14335975,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.018863125,0.00754525,0.003772625,0.0150905,0.030181,0.0452715,0.060362,0.06790725,0.05281675,0.0150905,0.011317875,0.003772625,0.0,0.0,0.00754525,0.011317875,0.018863125,0.03772625,0.07922512,0.15467763,0.19240387,0.21503963,0.23767537,0.28294688,0.35839936,0.29049212,0.17731337,0.19994913,0.46026024,0.965792,0.98465514,1.237421,1.4373702,1.4109617,1.0789708,1.1280149,1.0374719,0.8865669,0.754525,0.70170826,0.5998474,0.5470306,0.5055317,0.5357128,0.77716076,1.0751982,1.1129243,0.9997456,0.84884065,0.76584285,0.6790725,0.5696664,0.56212115,0.6526641,0.72811663,0.8111144,0.90920264,0.88279426,0.784706,0.86770374,1.1204696,1.3732355,1.5505489,1.6825907,1.931584,2.5616124,3.3915899,4.4139714,5.753253,7.6584287,8.050782,7.2623034,6.4474163,6.0286546,5.670255,5.402399,5.0741806,4.5950575,4.002755,3.4632697,3.1199608,2.7879698,2.4031622,1.9881734,1.6448646,1.5656394,1.5241405,1.4675511,1.3656902,1.237421,1.1355602,1.0487897,0.965792,0.8865669,0.83752275,0.8224323,0.7582976,0.663982,0.5696664,0.4979865,0.3772625,0.3055826,0.2678564,0.25276586,0.24899325,0.30935526,0.35839936,0.36971724,0.33576363,0.271629,0.271629,0.3734899,0.5093044,0.5885295,0.49421388,0.19240387,0.071679875,0.030181,0.018863125,0.02263575,0.011317875,0.00754525,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.018863125,0.018863125,0.018863125,0.041498873,0.03772625,0.018863125,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.150905,0.30181,0.5394854,0.8601585,1.20724,0.9016574,0.6073926,0.30935526,0.06790725,0.00754525,0.0150905,0.049044125,0.06790725,0.0754525,0.13204187,0.181086,0.15845025,0.23013012,0.47912338,0.875249,0.8903395,0.7809334,0.7696155,0.8526133,0.7922512,0.543258,0.62625575,1.0035182,1.3807807,1.2336484,0.7507524,0.33576363,0.11317875,0.1056335,0.25276586,0.2565385,0.23013012,0.25276586,0.34330887,0.4640329,0.62625575,0.69793564,0.68661773,0.72811663,1.056335,1.267602,1.4147344,1.3845534,1.2110126,1.0940613,0.72811663,0.47157812,0.26031113,0.094315626,0.041498873,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.0754525,0.20372175,0.49421388,1.0601076,2.033445,2.0560806,2.1805773,2.444661,2.7502437,2.848332,2.8030603,2.8898308,3.1576872,3.6896272,4.610148,6.692637,9.665465,13.008011,15.988385,17.663431,19.081938,20.768301,22.326395,23.450638,23.922215,23.707176,22.522572,20.941841,19.640285,19.38752,19.711966,19.749691,18.62545,16.4826,14.50197,13.513543,13.075918,12.683565,12.234623,12.019584,12.2270775,12.200669,12.042219,11.879996,11.883769,11.59705,11.7026825,12.012038,12.359119,12.593022,13.000465,13.792717,14.713238,15.403628,15.403628,14.426518,13.65313,13.158916,12.902377,12.728837,12.774108,12.981603,13.113645,13.275867,13.932304,13.6833105,14.188843,15.135772,16.335466,17.723793,19.391293,21.066338,22.183035,22.726294,23.258234,24.378702,26.608324,29.396294,32.067314,33.82913,35.29668,34.88169,33.161373,31.425966,31.67496,34.22148,37.8847,42.200584,45.68649,45.86003,42.687252,39.38243,38.397778,39.389977,39.20512,34.587425,28.573862,22.039675,15.912932,11.170743,9.6051035,8.431817,7.3151197,6.7756343,8.179051,9.25425,9.748463,9.544742,8.695901,7.4282985,6.258785,6.009792,6.1908774,6.470052,6.6662283,6.900131,7.326438,7.6697464,7.805561,7.7716074,7.8923316,8.103599,8.367682,8.661947,8.941121,9.190115,9.5032425,9.846551,10.299266,11.031156,11.438599,11.52537,11.355601,10.872705,9.899368,9.2995205,8.76758,7.884786,6.7114997,5.802297,5.1232247,4.6516466,4.2102494,3.7801702,3.5123138,3.2746384,3.006782,2.7238352,2.4069347,2.0070364,1.7127718,1.4562333,1.1921495,0.9393836,0.77716076,0.663982,0.59607476,0.55080324,0.5055317,0.46026024,0.3961256,0.43007925,0.5055317,0.6187105,0.7997965,0.8337501,0.6111652,0.3470815,0.16222288,0.07922512,0.0150905,0.0,0.0,0.0,0.0,0.29803738,0.32444575,0.18863125,0.030181,0.0,0.0,0.06413463,0.06413463,0.0,0.0,0.071679875,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.08299775,0.06790725,0.02263575,0.02263575,0.060362,0.12826926,0.241448,0.35839936,0.36971724,0.56589377,0.7469798,0.8526133,0.9280658,1.0940613,0.11317875,0.24899325,0.1961765,0.27540162,0.7054809,1.5769572,0.7394345,0.543258,0.87147635,1.3920987,1.5467763,0.7809334,0.91674787,1.116697,1.5580941,3.451952,1.1846043,0.77338815,0.543258,0.05281675,0.116951376,0.34330887,0.3470815,0.21881226,0.13958712,0.36594462,0.211267,0.06790725,0.10186087,0.36971724,0.8224323,0.35839936,0.18485862,0.14335975,0.26408374,0.7394345,0.35462674,0.41876137,0.41876137,0.2263575,0.11317875,0.150905,0.27917424,0.3961256,0.38103512,0.1056335,0.15467763,0.97710985,1.5656394,1.4260522,0.5696664,1.0072908,0.9922004,0.72811663,0.513077,0.72811663,0.5998474,6.6247296,7.8734684,3.1840954,1.1581959,5.80607,3.6292653,1.8259505,2.9351022,4.8666863,9.457971,7.1566696,3.6707642,2.0070364,2.4484336,1.629774,0.7696155,0.271629,0.1659955,0.120724,0.29049212,0.4640329,0.62248313,0.845068,1.3355093,1.1619685,0.8601585,0.6111652,0.42630664,0.1358145,0.026408374,0.056589376,0.10940613,0.211267,0.513077,0.20372175,0.120724,0.12826926,0.1961765,0.40367088,0.35462674,0.27917424,0.150905,0.02263575,0.0,0.011317875,0.018863125,0.018863125,0.033953626,0.071679875,0.19240387,0.27917424,0.4074435,0.47912338,0.21881226,0.06413463,0.011317875,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.0150905,0.02263575,0.003772625,0.0,0.0,0.003772625,0.0,0.0,0.018863125,0.06790725,0.150905,0.24899325,0.38103512,0.6413463,0.7884786,0.7205714,0.45648763,0.3169005,0.25276586,0.26031113,0.34330887,0.5055317,0.66775465,0.7922512,0.7922512,0.6413463,0.35839936,0.36594462,0.271629,0.17731337,0.15467763,0.24522063,0.5885295,1.0940613,1.629774,2.263575,3.2520027,3.7009451,4.617693,4.7648253,3.8556228,2.5502944,1.659955,1.1883769,0.86770374,0.8941121,1.8863125,2.516341,1.9504471,1.116697,0.60362,0.66020936,1.2751472,1.0110635,0.6375736,0.6752999,1.3958713,1.0638802,0.8601585,0.7809334,0.80734175,0.91674787,1.146878,2.263575,3.682082,5.383536,7.91874,9.171251,8.692128,8.511042,9.103344,9.416472,8.465771,8.160188,7.7942433,7.0963078,6.2663302,5.0515447,4.3611546,3.4368613,2.3654358,2.0598533,2.493705,2.505023,3.0445085,4.1800685,5.1081343,5.1873593,3.8593953,2.3013012,1.3543724,1.5543215,1.8523588,1.6222287,1.0525624,0.47535074,0.362172,0.2867195,0.1358145,0.041498873,0.06790725,0.2263575,0.13958712,0.06413463,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.03772625,0.02263575,0.018863125,0.033953626,0.056589376,0.06413463,0.10186087,0.120724,0.094315626,0.0150905,0.003772625,0.0150905,0.041498873,0.094315626,0.18485862,0.2263575,0.211267,0.18863125,0.181086,0.18863125,0.116951376,0.060362,0.026408374,0.033953626,0.071679875,0.124496624,0.14713238,0.26408374,0.5583485,1.0902886,0.8601585,0.8941121,1.0412445,1.1053791,0.84884065,0.7469798,0.73566186,0.8299775,0.94315624,0.9016574,0.84129536,0.8299775,0.8299775,0.94315624,1.4147344,1.8146327,1.8184053,1.6675003,1.5128226,1.4562333,1.2789198,0.9922004,0.7997965,0.814887,1.0601076,1.3807807,1.5430037,1.3468271,0.9242931,0.76584285,0.9393836,1.2261031,1.4750963,1.6976813,2.0560806,2.546522,3.3538637,4.2781568,5.160951,5.87775,6.1644692,6.2361493,6.224831,6.2135134,6.2135134,6.115425,5.824933,5.3684454,4.8440504,4.3875628,4.1310244,3.8820312,3.5575855,3.1312788,2.637065,2.474842,2.3805263,2.2748928,2.123988,1.9391292,1.7882242,1.6486372,1.4939595,1.3355093,1.1921495,1.1317875,1.0336993,0.91297525,0.7884786,0.6828451,0.5357128,0.41876137,0.35085413,0.33576363,0.34330887,0.36594462,0.38480774,0.40367088,0.40367088,0.32821837,0.271629,0.331991,0.3734899,0.3734899,0.41121614,0.19240387,0.071679875,0.0150905,0.003772625,0.011317875,0.003772625,0.0,0.011317875,0.02263575,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.03772625,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.071679875,0.30935526,0.47535074,0.6790725,1.4147344,1.4147344,1.1053791,0.65643674,0.25276586,0.08299775,0.041498873,0.0754525,0.10186087,0.09808825,0.08677038,0.120724,0.071679875,0.1056335,0.34330887,0.875249,1.0487897,0.9507015,0.9280658,1.0110635,0.90543,0.5394854,0.2867195,0.2867195,0.5998474,1.2298758,0.94315624,0.41121614,0.06413463,0.06413463,0.26408374,0.23390275,0.19240387,0.22258487,0.331991,0.45648763,0.5885295,0.76207024,0.875249,0.9205205,0.98465514,1.6222287,1.9240388,1.7693611,1.3543724,1.2110126,0.88279426,0.59607476,0.33953625,0.14713238,0.07922512,0.06790725,0.05281675,0.030181,0.003772625,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.16222288,0.5470306,1.3996439,1.5165952,1.4675511,1.3430545,1.297783,1.5580941,1.7429527,1.8561316,1.9051756,2.0070364,2.4031622,3.6066296,5.5495315,7.9526935,10.453944,12.596795,14.034165,16.029884,17.795471,19.312067,21.31533,22.97906,22.714975,21.77559,20.945614,20.541943,19.549744,18.599041,17.4333,16.086473,14.890551,13.958713,13.140053,12.419481,11.921495,11.898859,12.381755,12.996693,13.275867,13.226823,13.29473,12.97783,13.091009,13.264549,13.381501,13.562587,13.6682205,14.268067,15.17727,16.177015,17.006994,16.641048,15.633758,14.784918,14.358611,14.071891,14.475562,14.366156,14.25675,14.622695,15.897841,15.347038,15.573396,16.501461,17.70493,18.395319,19.866644,21.866135,23.62795,24.955914,26.219744,27.804247,30.46772,33.489594,36.122883,37.586662,36.65105,35.934254,36.209656,37.74134,40.28786,44.76974,48.312237,49.923145,48.440506,42.521255,40.12564,40.551945,43.430458,46.742825,46.83714,41.985542,34.576107,25.608578,17.056038,11.84227,11.053791,8.89585,7.201941,6.9227667,8.126234,9.786189,10.872705,11.083972,10.416218,9.186342,8.348819,8.122461,8.179051,8.326183,8.518587,8.439363,9.058073,9.522105,9.408927,8.744945,8.160188,7.8432875,7.6810646,7.598067,7.567886,7.8395147,8.069645,8.182823,8.254503,8.488406,8.986393,9.7069645,10.159679,9.989911,9.001483,8.692128,8.145098,7.496206,6.790725,5.9909286,5.3344917,5.0213637,4.6516466,4.191386,3.9801195,3.7009451,3.4444065,3.2557755,3.0369632,2.5691576,2.2975287,1.9768555,1.6561824,1.3732355,1.1242423,0.9280658,0.8299775,0.7922512,0.784706,0.7922512,0.6828451,0.73566186,0.84129536,0.9695646,1.1732863,1.1846043,0.9695646,0.7054809,0.4678055,0.25276586,0.09808825,0.05281675,0.030181,0.003772625,0.018863125,0.3961256,0.39989826,0.23390275,0.06790725,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.03772625,0.05281675,0.033953626,0.003772625,0.011317875,0.018863125,0.00754525,0.003772625,0.00754525,0.0,0.02263575,0.08299775,0.08299775,0.033953626,0.049044125,0.060362,0.11317875,0.11317875,0.09808825,0.21503963,0.4640329,0.62248313,0.6111652,0.5093044,0.543258,0.0150905,0.003772625,0.08299775,0.271629,0.5772116,0.9922004,1.2864652,1.2864652,2.082489,3.2331395,2.7313805,1.388326,0.8978847,0.8186596,0.9507015,1.327964,1.1204696,0.6111652,0.20749438,0.06790725,0.090543,0.1056335,0.060362,0.03772625,0.09808825,0.3055826,0.120724,0.030181,0.0,0.003772625,0.0150905,0.003772625,0.026408374,0.0452715,0.041498873,0.030181,0.00754525,0.0,0.0,0.003772625,0.0150905,0.0150905,0.38103512,0.59607476,0.45648763,0.090543,0.056589376,0.694163,1.1242423,1.0601076,0.83752275,2.3390274,1.4713237,0.56589377,0.875249,2.546522,2.6332922,4.606375,5.379763,4.3686996,3.4783602,9.0807085,5.9230213,2.4371157,2.5616124,5.723072,8.409182,7.394345,5.8928404,5.0213637,3.8141239,1.1431054,0.49044126,0.41121614,0.24522063,0.120724,0.3772625,0.331991,0.30935526,0.44139713,0.68661773,0.271629,0.48666862,0.48666862,0.1358145,0.0150905,0.003772625,0.056589376,0.15845025,0.3055826,0.48666862,0.5017591,0.30181,0.150905,0.120724,0.120724,0.2678564,0.38858038,0.32067314,0.10940613,0.0,0.060362,0.08677038,0.07922512,0.08299775,0.1659955,0.72811663,1.1091517,1.7957695,2.2711203,0.97710985,0.2565385,0.030181,0.0,0.0,0.0,0.011317875,0.041498873,0.03772625,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.056589376,0.23013012,0.5017591,0.7469798,0.6375736,0.8941121,1.0714256,0.90920264,0.33576363,0.1659955,0.15845025,0.19994913,0.27540162,0.45648763,0.58098423,0.6187105,0.62625575,0.6413463,0.70170826,1.0186088,0.84129536,0.5017591,0.27917424,0.42630664,1.026154,1.5241405,1.8334957,1.9353566,1.8599042,2.5314314,2.2598023,1.5354583,0.97710985,1.3430545,1.2336484,1.1581959,1.0148361,0.8111144,0.70170826,1.750498,1.3996439,0.9507015,1.0487897,1.7089992,4.112161,2.9841464,1.2864652,0.47912338,0.5017591,0.6149379,0.694163,0.87902164,1.0148361,0.68661773,0.55080324,1.20724,2.1466236,3.2935016,4.991183,6.013564,5.511805,6.017337,7.997965,9.842778,8.511042,9.020347,9.740918,9.597558,8.073418,6.4964604,5.956975,5.541986,5.3080835,6.270103,5.515578,5.243949,5.7079816,6.145606,4.7912335,3.0331905,1.6146835,1.1619685,1.6750455,2.516341,2.2975287,1.5279131,0.7092535,0.35085413,0.9620194,0.814887,0.31312788,0.056589376,0.26408374,0.76207024,0.5319401,0.23390275,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.041498873,0.090543,0.13958712,0.150905,0.041498873,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.071679875,0.20372175,0.45648763,0.87147635,1.0299267,0.9393836,0.7507524,0.55457586,0.3961256,0.18863125,0.071679875,0.041498873,0.056589376,0.0452715,0.120724,0.30181,0.5394854,0.77338815,0.9318384,0.80734175,0.5319401,0.4376245,0.58098423,0.70170826,0.77338815,0.875249,0.9318384,0.9393836,0.97710985,1.0978339,1.1657411,1.0940613,0.9997456,1.2223305,1.4034165,1.4600059,1.5203679,1.6637276,1.9089483,1.6524098,1.2562841,1.056335,1.2826926,2.0749438,2.2447119,2.0975795,1.7655885,1.3770081,1.0223814,1.1091517,1.871222,2.3654358,2.372981,2.4107075,1.9353566,1.9730829,2.1503963,2.3503454,2.71629,3.1312788,3.5538127,4.0178456,4.504514,4.9421387,5.138315,5.168496,5.0213637,4.7421894,4.425289,4.168751,3.9499383,3.663219,3.2482302,2.686109,2.4522061,2.3126192,2.161714,1.9504471,1.6939086,1.5354583,1.3770081,1.1996948,0.9997456,0.77716076,0.7167987,0.6187105,0.5017591,0.40367088,0.36594462,0.3055826,0.25276586,0.21503963,0.20749438,0.24522063,0.2678564,0.29426476,0.32444575,0.33953625,0.29049212,0.31312788,0.392353,0.38103512,0.31312788,0.41121614,0.29049212,0.11317875,0.00754525,0.0,0.0,0.0,0.00754525,0.026408374,0.0452715,0.0452715,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.00754525,0.056589376,0.21881226,0.48666862,0.77716076,0.59607476,0.422534,0.452715,0.5696664,0.35085413,0.14335975,0.090543,0.08677038,0.08677038,0.1358145,0.29426476,0.20749438,0.07922512,0.1056335,0.47157812,0.6073926,0.55080324,0.73188925,1.1129243,1.1732863,0.6488915,0.30935526,0.32821837,0.7167987,1.327964,1.0714256,0.44894236,0.0452715,0.030181,0.150905,0.21503963,0.19240387,0.21503963,0.31312788,0.3961256,0.663982,0.91674787,1.1431054,1.267602,1.1431054,1.6335466,1.7919968,1.7731338,1.6146835,1.237421,1.0035182,0.69793564,0.39989826,0.17731337,0.090543,0.090543,0.1358145,0.11317875,0.02263575,0.0,0.011317875,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.17731337,0.34330887,0.5017591,0.69039035,1.0072908,1.2147852,1.5958204,1.81086,1.8146327,1.8749946,2.3880715,4.0103,5.9682927,8.069645,10.680302,14.25675,16.690092,17.976559,18.546225,19.240387,20.277859,20.621168,20.43631,19.821371,18.7839,18.663176,17.67852,16.316603,15.022593,14.2077055,13.498452,13.29473,13.434318,13.59654,13.290957,13.411682,13.52486,13.860624,14.539697,15.562078,15.894069,15.829934,15.577168,15.39231,15.562078,15.403628,15.482853,15.984612,16.690092,16.984358,18.470772,19.055529,19.206434,19.063074,18.417955,19.60256,18.485863,17.112627,16.652367,17.410664,18.715992,19.508244,20.613623,21.77559,21.666185,23.107328,25.800982,29.21898,32.433258,34.11962,33.433002,34.68174,37.348988,39.612564,38.32987,36.341698,37.269764,40.944298,46.24484,51.115295,56.62333,60.441227,60.93544,57.679665,51.46615,49.892967,49.82883,47.636936,43.539864,41.612053,39.729515,33.421684,25.404858,18.251959,14.358611,13.88326,10.431308,7.673519,6.930312,7.1868505,8.262049,10.38981,12.189351,12.736382,11.566868,11.3820095,11.2650585,11.076427,11.019837,11.642321,10.665211,11.125471,11.706455,11.634775,10.695392,9.782416,9.103344,8.503497,7.960239,7.567886,7.8961043,8.311093,8.07719,7.4509344,7.6584287,7.8432875,7.8696957,8.00551,8.269594,8.4544525,8.952439,8.126234,7.1264887,6.477597,6.089017,5.6476197,5.3759904,5.13077,4.908185,4.821415,4.2592936,4.063117,4.0895257,3.9499383,3.0218725,2.776652,2.5502944,2.282438,1.9542197,1.5882751,1.2449663,1.0299267,0.935611,0.91297525,0.9016574,0.8526133,0.98465514,1.1431054,1.2562841,1.3430545,1.3543724,1.1581959,0.9242931,0.7167987,0.47157812,0.32821837,0.271629,0.15467763,0.018863125,0.090543,0.018863125,0.0,0.0,0.041498873,0.19994913,0.041498873,0.0,0.0,0.0,0.0,0.1961765,0.26408374,0.1659955,0.011317875,0.060362,0.08677038,0.03772625,0.018863125,0.03772625,0.0,0.011317875,0.033953626,0.041498873,0.02263575,0.0,0.011317875,0.25276586,0.29049212,0.12826926,0.21503963,0.24899325,0.18485862,0.1056335,0.06790725,0.090543,0.003772625,0.0,0.0150905,0.08299775,0.19994913,0.331991,0.7507524,1.0789708,1.6033657,1.9579924,1.0940613,0.72811663,1.0827434,0.9922004,1.0525624,3.5990841,1.2826926,0.3772625,0.13958712,0.1056335,0.07922512,0.071679875,0.05281675,0.05281675,0.11317875,0.27917424,0.30181,0.29049212,0.27540162,0.26031113,0.22258487,0.124496624,0.060362,0.03772625,0.041498873,0.018863125,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.0754525,0.12826926,0.120724,0.06790725,0.44139713,1.0827434,1.0601076,0.5357128,0.754525,1.4750963,2.7389257,2.595566,1.3996439,1.8033148,2.5427492,3.0897799,3.712263,4.7572803,6.63982,8.054554,4.6629643,2.1541688,2.3503454,3.2067313,3.783943,3.8480775,4.3385186,4.859141,3.682082,2.0145817,1.3656902,0.8941121,0.36971724,0.16976812,0.22258487,0.14713238,0.13204187,0.271629,0.56589377,0.3734899,0.5885295,0.543258,0.24522063,0.35839936,0.88279426,0.9205205,0.7507524,0.633801,0.80734175,0.633801,0.35085413,0.150905,0.08677038,0.08677038,0.06413463,0.11317875,0.116951376,0.06413463,0.071679875,0.124496624,0.08677038,0.049044125,0.03772625,0.0452715,0.1659955,0.25276586,0.392353,0.47535074,0.1961765,0.05281675,0.02263575,0.06413463,0.124496624,0.1358145,0.07922512,0.056589376,0.030181,0.00754525,0.03772625,0.056589376,0.0452715,0.026408374,0.011317875,0.0,0.011317875,0.02263575,0.32067314,0.69793564,0.44139713,0.3734899,0.73188925,1.0186088,0.9393836,0.44516975,0.29426476,0.20372175,0.181086,0.23390275,0.4074435,0.65643674,0.95824677,1.146878,1.1393328,0.8978847,0.6790725,0.482896,0.36971724,0.36594462,0.4640329,0.66020936,1.2336484,2.493705,4.06689,4.9119577,3.8480775,2.8558772,2.0447628,1.5958204,1.7467253,1.7240896,2.0975795,2.252257,1.8259505,0.69039035,0.8978847,0.9922004,0.86770374,0.67152727,0.7922512,1.3317367,1.7014539,1.7957695,1.6788181,1.5769572,0.52439487,0.30935526,0.41876137,0.4979865,0.34330887,0.35839936,0.6451189,1.177059,2.022127,3.3161373,4.244203,3.7688525,3.7386713,5.1534057,8.171506,8.548768,8.318638,8.548768,9.0957985,8.631766,9.714509,10.008774,9.14107,7.4999785,6.198423,4.768598,3.6028569,2.7351532,2.214531,2.1164427,1.9994912,2.4861598,2.7389257,2.4031622,1.6146835,1.267602,0.79602385,0.392353,0.21503963,0.3772625,0.35462674,0.22258487,0.14713238,0.24899325,0.60362,0.73188925,0.45648763,0.18863125,0.09808825,0.09808825,0.030181,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.13204187,0.13204187,0.09808825,0.13958712,0.116951376,0.09808825,0.0754525,0.0754525,0.17354076,0.4678055,0.6187105,0.7167987,0.8639311,1.1506506,1.2487389,1.1996948,1.0374719,0.80356914,0.52062225,0.25276586,0.32067314,0.45648763,0.47535074,0.27917424,0.30181,0.6413463,0.875249,0.875249,0.80734175,0.724344,0.814887,1.0148361,1.2034674,1.237421,1.0374719,0.845068,0.7469798,0.7997965,1.0148361,1.1846043,1.2940104,1.1695137,0.9808825,1.20724,1.4109617,1.3619176,1.2902378,1.297783,1.3468271,1.1393328,0.97710985,0.9620194,1.1657411,1.6486372,1.81086,1.7014539,1.5656394,1.7052265,2.463524,3.1614597,3.399135,3.0143273,2.252257,1.750498,1.5580941,1.2713746,1.0374719,0.94315624,1.0072908,1.0902886,1.2034674,1.3845534,1.6222287,1.8561316,1.9240388,1.901403,1.841041,1.7769064,1.7014539,1.6410918,1.5505489,1.4071891,1.2110126,0.9997456,0.90543,0.83752275,0.76584285,0.6828451,0.58475685,0.5319401,0.4640329,0.3961256,0.32821837,0.25276586,0.27917424,0.26408374,0.21881226,0.17731337,0.16976812,0.13958712,0.094315626,0.06790725,0.071679875,0.09808825,0.10186087,0.120724,0.16222288,0.211267,0.241448,0.27540162,0.29803738,0.3055826,0.3055826,0.32821837,0.22258487,0.094315626,0.02263575,0.011317875,0.011317875,0.02263575,0.041498873,0.08299775,0.13204187,0.14335975,0.049044125,0.011317875,0.003772625,0.011317875,0.0,0.011317875,0.00754525,0.00754525,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.026408374,0.18485862,0.39989826,0.39989826,0.1961765,0.1056335,0.12826926,0.20372175,0.21503963,0.25276586,0.482896,0.5998474,0.48666862,0.22258487,0.35085413,0.3961256,0.3169005,0.23013012,0.39989826,0.5357128,0.63002837,0.86770374,1.1280149,1.0035182,0.4678055,0.38858038,0.59230214,0.875249,0.98465514,0.6111652,0.23013012,0.02263575,0.0150905,0.06790725,0.10940613,0.09808825,0.11317875,0.18485862,0.29803738,0.47912338,0.6187105,0.80356914,1.0110635,1.1431054,1.5241405,2.022127,2.2484846,1.9655377,1.0902886,0.90543,0.7884786,0.6413463,0.44894236,0.27540162,0.1659955,0.120724,0.090543,0.0754525,0.10940613,0.181086,0.16976812,0.10940613,0.049044125,0.03772625,0.026408374,0.018863125,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0452715,0.10940613,0.2263575,0.41876137,0.72811663,0.9808825,1.3392819,1.5543215,1.6373192,1.8636768,1.7731338,2.2899833,3.3651814,4.98741,7.1906233,10.114408,13.026875,16.15438,19.379974,22.243397,23.156372,23.077147,22.57916,22.243397,22.639523,22.371666,22.21699,21.651094,20.572124,19.296976,18.433046,17.697384,17.052265,16.358103,15.377219,15.041456,14.7321005,14.535924,14.5132885,14.698147,15.260268,16.158154,16.644821,16.509007,16.063837,15.973294,18.078419,19.123436,18.685812,19.1423,19.998686,20.934296,22.201899,23.55627,24.276842,24.423975,24.48811,24.8201,25.276588,25.22377,24.586197,24.276842,24.597515,25.340723,25.816072,27.366621,29.758467,32.98029,36.39074,38.707134,38.90331,41.28761,45.150776,48.746086,49.293118,48.425415,51.153023,53.631638,54.11076,52.937473,54.348434,55.7179,56.042343,55.699036,56.449787,61.603195,61.64469,57.362762,50.21741,42.343945,33.723495,25.706667,19.911915,16.708956,15.237633,12.702429,10.20495,8.405409,7.6018395,7.7602897,9.684328,10.676529,11.830952,12.925014,12.396846,13.20796,13.902123,14.471789,14.800008,14.667966,13.713491,13.336229,12.936331,12.37421,11.989402,11.876224,11.216014,10.197406,9.073163,8.167733,7.7942433,7.9715567,7.937603,7.6093845,7.564113,7.61693,7.6886096,7.7942433,7.9262853,8.050782,7.964011,8.062099,7.635793,6.760544,6.270103,5.8626595,5.594803,5.4363527,5.3571277,5.311856,4.9345937,4.727099,4.7421894,4.647874,3.742444,3.2029586,2.8898308,2.686109,2.4559789,2.052308,1.9127209,1.8523588,1.629774,1.3053282,1.2525115,1.1091517,1.1431054,1.2261031,1.2940104,1.3807807,1.50905,1.4637785,1.2826926,1.0110635,0.7167987,0.52062225,0.3961256,0.2867195,0.19240387,0.17731337,0.124496624,0.07922512,0.15845025,0.25276586,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.03772625,0.05281675,0.033953626,0.003772625,0.011317875,0.018863125,0.10940613,0.18485862,0.18863125,0.120724,0.0754525,0.13958712,0.16976812,0.120724,0.03772625,0.03772625,0.18863125,0.32444575,0.3169005,0.090543,0.10940613,0.06790725,0.030181,0.0150905,0.030181,0.14713238,0.24899325,0.10940613,0.056589376,0.32821837,1.0940613,0.94315624,1.2940104,1.8297231,2.214531,2.0598533,0.8978847,1.4260522,1.4373702,0.98842776,2.3993895,1.3845534,0.94315624,0.59230214,0.23013012,0.150905,0.094315626,0.06413463,0.049044125,0.05281675,0.10940613,0.13958712,0.181086,0.23013012,0.24522063,0.14713238,0.06790725,0.026408374,0.0150905,0.0150905,0.00754525,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.24522063,0.62248313,0.7130261,0.5772116,0.79602385,2.282438,3.9650288,3.6707642,1.9844007,2.2673476,2.8256962,3.3689542,4.285702,5.798525,7.9715567,7.877241,5.485397,3.6066296,2.9766011,2.2296214,1.4298248,1.5279131,2.2598023,2.9200118,2.3465726,1.9994912,1.5769572,1.0148361,0.4979865,0.44894236,0.24522063,0.08677038,0.19994913,0.59230214,1.0751982,0.4640329,0.452715,0.46026024,0.362172,0.48666862,0.8111144,0.7394345,0.5394854,0.452715,0.7092535,0.49044126,0.331991,0.26408374,0.23390275,0.094315626,0.049044125,0.120724,0.17354076,0.14713238,0.071679875,0.071679875,0.071679875,0.18863125,0.392353,0.52062225,0.44894236,0.46026024,0.41876137,0.2867195,0.10940613,0.21881226,0.32444575,0.4074435,0.41121614,0.241448,0.14713238,0.0754525,0.026408374,0.003772625,0.018863125,0.033953626,0.026408374,0.0150905,0.003772625,0.0,0.003772625,0.00754525,0.211267,0.47912338,0.32067314,0.43385187,0.51684964,0.573439,0.5470306,0.29049212,0.3055826,0.44516975,0.5583485,0.5998474,0.62625575,0.7582976,1.1506506,1.5882751,1.8297231,1.6146835,1.0638802,0.77716076,0.67152727,0.694163,0.8299775,1.1091517,1.6976813,2.41448,3.0520537,3.380272,2.776652,2.3088465,1.9466745,1.6712729,1.4524606,1.8938577,3.059599,3.9084394,3.9914372,3.440634,2.776652,3.0671442,2.776652,1.871222,1.8297231,1.2185578,1.4071891,1.7693611,1.9429018,1.81086,0.7809334,0.32444575,0.30935526,0.5885295,0.9922004,1.0789708,0.9205205,0.90543,1.297783,2.2220762,2.9652832,2.5804756,2.191895,2.6483827,4.5309224,7.2698483,9.156161,10.284176,10.616167,10.020092,10.499215,10.303039,9.144843,7.3075747,5.621211,3.8971217,2.6144292,1.9957186,2.123988,2.9615107,2.776652,2.5540671,2.2069857,1.6750455,0.9016574,0.86770374,0.73566186,0.5017591,0.27917424,0.28294688,0.29426476,0.23013012,0.18485862,0.21503963,0.32821837,0.39989826,0.25276586,0.1056335,0.049044125,0.049044125,0.02263575,0.02263575,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.033953626,0.033953626,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.011317875,0.003772625,0.00754525,0.06790725,0.26408374,0.36594462,0.36594462,0.3055826,0.24522063,0.2565385,0.34330887,0.34330887,0.29803738,0.25276586,0.24899325,0.4640329,0.5772116,0.6488915,0.72811663,0.845068,0.7997965,0.7167987,0.62248313,0.513077,0.3470815,0.30935526,0.49421388,0.5885295,0.49044126,0.29049212,0.3169005,0.6375736,0.875249,0.8903395,0.79602385,0.8337501,1.0223814,1.1431054,1.116697,0.9997456,0.86770374,0.8262049,0.9205205,1.0789708,1.1242423,1.2261031,1.3694628,1.4373702,1.3920987,1.2864652,1.3920987,1.3241913,1.2487389,1.2034674,1.0789708,0.9620194,0.875249,0.7997965,0.79602385,0.97333723,1.1921495,1.6184561,2.282438,2.9766011,3.2444575,2.686109,2.1768045,1.7014539,1.267602,0.90920264,0.7507524,0.5093044,0.32067314,0.23767537,0.23013012,0.23013012,0.24522063,0.29426476,0.36971724,0.452715,0.4678055,0.44516975,0.42630664,0.42630664,0.42630664,0.41498876,0.38858038,0.3470815,0.3055826,0.31312788,0.32067314,0.2678564,0.20372175,0.15845025,0.13958712,0.116951376,0.094315626,0.07922512,0.06413463,0.056589376,0.071679875,0.06790725,0.06413463,0.060362,0.0754525,0.05281675,0.030181,0.018863125,0.0150905,0.033953626,0.033953626,0.056589376,0.094315626,0.1358145,0.19240387,0.23767537,0.25276586,0.23013012,0.19240387,0.21503963,0.150905,0.071679875,0.026408374,0.02263575,0.02263575,0.02263575,0.041498873,0.07922512,0.116951376,0.11317875,0.060362,0.03772625,0.02263575,0.011317875,0.0,0.011317875,0.00754525,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.049044125,0.12826926,0.18863125,0.120724,0.03772625,0.011317875,0.018863125,0.0452715,0.08299775,0.23013012,0.56589377,0.633801,0.3772625,0.1056335,0.20749438,0.4979865,0.66020936,0.5998474,0.4376245,0.52062225,0.7394345,1.0676528,1.2449663,0.7884786,0.36594462,0.52439487,0.8563859,1.0412445,0.8526133,0.5093044,0.2263575,0.056589376,0.00754525,0.0452715,0.08299775,0.071679875,0.060362,0.08299775,0.18485862,0.2678564,0.362172,0.4678055,0.573439,0.6488915,0.9393836,1.2864652,1.4675511,1.4411428,1.3166461,0.88279426,0.94692886,1.0412445,0.94692886,0.6790725,0.59607476,0.40367088,0.241448,0.17354076,0.19240387,0.21881226,0.19994913,0.15467763,0.116951376,0.12826926,0.071679875,0.05281675,0.05281675,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.06413463,0.15467763,0.29049212,0.47157812,0.7394345,0.9507015,1.0940613,1.3015556,1.2110126,1.3430545,1.8448136,2.8256962,4.3686996,6.1229706,8.526133,11.740409,15.69412,20.066593,23.507227,25.32186,25.717985,25.314314,25.133228,24.56356,23.990122,23.778856,23.58268,22.352802,21.107838,20.11941,19.274342,18.323639,16.897587,16.218515,15.313085,14.611377,14.302021,14.351066,14.7170105,15.098045,15.573396,16.146835,16.712729,16.637276,19.421474,21.564325,22.100037,22.631977,23.458181,23.533634,23.816582,24.537153,25.212452,26.287651,27.721249,29.437794,30.924208,31.22979,30.033867,29.056757,28.366367,28.24187,29.143528,32.301216,35.52681,38.756176,41.43097,42.50239,44.226482,47.116314,51.19075,55.163322,56.472424,57.064724,60.354454,62.538803,61.73901,58.011654,56.170612,56.762917,58.241783,60.497814,64.870285,70.21987,70.13687,65.61726,57.125088,44.603745,31.508965,22.990377,19.119663,17.953922,15.513034,12.702429,10.774617,9.450426,8.650629,8.507269,9.654147,10.842525,12.521342,14.132254,14.086982,14.8339615,15.494171,16.203424,16.923996,17.440845,17.301258,16.67123,15.554533,14.279386,13.494679,12.89106,12.151625,11.423509,10.744436,10.038955,9.26934,8.684583,8.224322,7.9036493,7.8206515,8.243186,8.43559,8.333729,8.103599,8.167733,8.186596,8.130007,7.752744,7.201941,7.01331,6.6549106,6.228604,5.87775,5.6513925,5.4967146,5.304311,5.081726,4.878004,4.606375,4.0404816,3.5764484,3.2067313,2.927557,2.686109,2.3578906,2.1768045,2.1051247,1.9881734,1.8372684,1.8184053,1.5807298,1.539231,1.599593,1.6410918,1.4977322,1.6260014,1.6410918,1.5279131,1.3468271,1.20724,0.8601585,0.66020936,0.513077,0.3961256,0.38103512,0.30935526,0.27917424,0.30181,0.29049212,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0150905,0.033953626,0.026408374,0.033953626,0.1659955,0.049044125,0.090543,0.16222288,0.19240387,0.16222288,0.18863125,0.23013012,0.28294688,0.30181,0.211267,0.24899325,0.27540162,0.30181,0.3055826,0.23390275,0.36594462,0.5093044,0.4376245,0.21503963,0.18863125,0.17731337,0.30935526,0.1358145,0.181086,0.73188925,1.8485862,1.146878,1.2789198,1.690136,2.0258996,2.1277604,0.9205205,1.1204696,1.4826416,1.5354583,1.569412,2.1843498,2.0145817,1.3430545,0.6375736,0.52062225,0.3055826,0.3169005,0.24899325,0.071679875,0.03772625,0.02263575,0.06790725,0.116951376,0.124496624,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.27540162,0.47157812,0.6488915,1.1393328,3.218049,3.7386713,2.927557,1.8146327,2.2183034,3.3915899,3.9159849,4.4101987,5.247721,6.56814,6.6247296,5.534441,3.893349,2.2975287,1.358145,0.4678055,0.392353,0.7205714,1.0940613,1.1921495,1.5580941,1.3694628,0.94315624,0.573439,0.5281675,0.21881226,0.07922512,0.24522063,0.6488915,0.9997456,0.3961256,0.36594462,0.41498876,0.35839936,0.32821837,0.5055317,0.5055317,0.44894236,0.5281675,0.98465514,0.55457586,0.392353,0.3772625,0.3470815,0.071679875,0.049044125,0.116951376,0.181086,0.211267,0.2263575,0.422534,1.0299267,1.3694628,1.2562841,1.0148361,0.80734175,0.6451189,0.5319401,0.482896,0.52439487,0.724344,0.7507524,0.663982,0.49044126,0.23390275,0.15467763,0.094315626,0.049044125,0.0150905,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.07922512,0.1961765,0.20372175,0.362172,0.32444575,0.2678564,0.2263575,0.11317875,0.26031113,0.6413463,1.0148361,1.2185578,1.1695137,1.0638802,1.2223305,1.5731846,1.9164935,1.901403,1.4222796,1.1242423,0.9695646,0.935611,1.0072908,1.2034674,1.5731846,1.7957695,1.8976303,2.2786655,2.2598023,2.1315331,1.991946,1.8070874,1.3958713,1.690136,2.848332,4.3347464,5.5306683,5.772116,4.7346444,4.5950575,4.22534,3.4066803,2.8181508,1.8070874,1.5279131,1.7354075,1.931584,1.3807807,0.7054809,0.31312788,0.26408374,0.5281675,0.9808825,1.1280149,0.91297525,0.694163,0.73566186,1.1959221,1.690136,1.7429527,1.5618668,1.4562333,1.8146327,5.6551647,9.64283,11.932813,12.076173,10.982111,10.0465,9.107117,7.99042,6.5832305,4.8402777,3.7499893,3.682082,3.5689032,3.169005,3.0746894,2.4597516,1.8636768,1.4449154,1.2713746,1.3053282,1.8485862,1.8146327,1.2600567,0.6111652,0.6488915,0.58098423,0.31312788,0.15845025,0.17354076,0.181086,0.1659955,0.20372175,0.18485862,0.094315626,0.011317875,0.011317875,0.018863125,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.026408374,0.041498873,0.026408374,0.011317875,0.124496624,0.3470815,0.5357128,0.44516975,0.38103512,0.34330887,0.34330887,0.4074435,0.44139713,0.42630664,0.38858038,0.3470815,0.29803738,0.33953625,0.35839936,0.3961256,0.452715,0.48666862,0.33953625,0.27917424,0.2678564,0.2678564,0.23013012,0.29426476,0.45648763,0.52439487,0.44516975,0.30935526,0.35462674,0.55457586,0.694163,0.7469798,0.8337501,1.026154,1.0902886,1.0186088,0.87902164,0.814887,0.87902164,1.0412445,1.2487389,1.3845534,1.2826926,1.3694628,1.5279131,1.5845025,1.4524606,1.116697,1.1431054,1.1506506,1.1808317,1.2185578,1.1808317,1.116697,0.90920264,0.67152727,0.52062225,0.59607476,0.9922004,1.8448136,2.7804246,3.2444575,2.4672968,1.3128735,0.68661773,0.44139713,0.38480774,0.27917424,0.1659955,0.071679875,0.0150905,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.018863125,0.011317875,0.00754525,0.011317875,0.018863125,0.011317875,0.00754525,0.00754525,0.02263575,0.08299775,0.11317875,0.07922512,0.03772625,0.011317875,0.018863125,0.003772625,0.0,0.011317875,0.033953626,0.041498873,0.00754525,0.003772625,0.011317875,0.030181,0.056589376,0.041498873,0.026408374,0.011317875,0.00754525,0.0150905,0.018863125,0.041498873,0.06790725,0.09808825,0.15467763,0.18863125,0.19994913,0.18485862,0.15845025,0.1659955,0.12826926,0.06413463,0.026408374,0.02263575,0.030181,0.026408374,0.033953626,0.056589376,0.08299775,0.06413463,0.056589376,0.0452715,0.030181,0.011317875,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.056589376,0.03772625,0.0,0.0,0.0,0.003772625,0.026408374,0.08299775,0.18863125,0.3772625,0.36594462,0.150905,0.00754525,0.12826926,0.5885295,0.9318384,0.9242931,0.5772116,0.5998474,0.9280658,1.2298758,1.2147852,0.6149379,0.42630664,0.6488915,0.84129536,0.80356914,0.56212115,0.4376245,0.2678564,0.10940613,0.0150905,0.026408374,0.05281675,0.056589376,0.03772625,0.026408374,0.07922512,0.10186087,0.15845025,0.19994913,0.21503963,0.241448,0.41876137,0.5470306,0.62625575,0.7432071,1.1053791,0.83752275,1.1695137,1.5467763,1.6109109,1.2147852,0.935611,0.633801,0.3961256,0.26031113,0.21503963,0.1961765,0.16976812,0.15845025,0.15845025,0.15845025,0.094315626,0.090543,0.090543,0.06413463,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.026408374,0.10186087,0.23013012,0.362172,0.48666862,0.6187105,0.69039035,0.7696155,0.9922004,1.4600059,2.2598023,3.3878171,4.776143,6.9454026,10.182315,14.547242,19.836462,24.412657,27.634478,29.234072,29.298206,28.049467,26.404602,25.65385,25.68403,24.997414,23.72981,22.590479,21.620914,20.685303,19.455427,18.429274,17.120173,16.097792,15.482853,14.981093,14.811326,14.569878,14.800008,15.728074,17.286167,17.47857,19.251705,21.360603,23.1526,24.571106,25.56708,25.506718,25.15209,25.129456,25.92925,27.740112,30.346996,32.776566,34.36484,34.760967,34.357296,33.553726,32.62566,32.25217,33.512226,37.26222,40.72926,43.362553,44.92442,45.497856,48.07079,50.50036,53.499596,56.559193,57.985245,58.856724,62.180405,65.8474,67.609215,65.09287,60.109234,60.10546,63.67814,69.35971,75.629814,76.36548,74.0604,67.526215,56.5856,42.07986,29.66415,22.398075,19.40261,18.350048,15.475307,13.298503,12.0082655,11.140562,10.359629,9.461743,9.718282,10.906659,13.000465,15.301767,16.429781,16.927769,17.40312,17.91997,18.500954,19.149845,19.934551,19.896824,19.074392,17.738882,16.380737,14.981093,13.551269,12.66093,12.253486,11.664956,10.816116,10.042727,9.378746,8.846806,8.469543,8.809079,9.0543,8.971302,8.76758,9.0957985,9.099571,8.684583,8.031919,7.4735703,7.4811153,7.1793056,6.6813188,6.1833324,5.794752,5.564622,5.4891696,5.3080835,5.0062733,4.6214657,4.2291126,3.8593953,3.4896781,3.1576872,2.867195,2.595566,2.3428001,2.2183034,2.1692593,2.1768045,2.282438,2.1390784,2.0183544,1.9655377,1.9164935,1.7014539,1.81086,1.7769064,1.6675003,1.5580941,1.5430037,1.20724,1.0035182,0.8224323,0.66020936,0.6073926,0.5319401,0.5281675,0.4640329,0.32067314,0.18485862,0.15467763,0.13204187,0.1056335,0.08677038,0.09808825,0.033953626,0.15845025,0.25276586,0.2867195,0.4074435,0.20372175,0.12826926,0.13204187,0.1659955,0.15467763,0.22258487,0.26031113,0.32444575,0.39989826,0.38858038,0.49421388,0.47535074,0.44894236,0.513077,0.72811663,1.177059,1.3619176,1.1695137,0.7432071,0.49421388,0.06413463,0.124496624,0.056589376,0.2867195,0.9507015,1.8749946,1.1544232,0.9620194,0.9808825,0.97333723,0.7696155,0.84129536,0.4979865,0.965792,1.9768555,1.750498,2.8596497,2.6068838,1.8787673,1.3392819,1.4260522,0.88279426,0.8299775,0.73566186,0.5055317,0.4979865,0.47535074,0.35085413,0.18485862,0.056589376,0.030181,0.0150905,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25276586,0.36594462,0.7092535,2.4408884,3.7613072,2.3465726,1.1204696,1.146878,1.6260014,4.429062,4.9723196,4.557331,4.093298,4.115934,4.3724723,4.104616,2.6634734,0.8224323,0.77338815,0.59607476,0.29426476,0.124496624,0.2263575,0.6111652,0.91674787,0.87902164,0.7205714,0.55080324,0.36971724,0.124496624,0.06790725,0.16222288,0.29426476,0.30181,0.211267,0.41876137,0.47535074,0.27917424,0.071679875,0.4376245,0.5885295,0.633801,0.7884786,1.3732355,0.76207024,0.46026024,0.36594462,0.3055826,0.056589376,0.071679875,0.0754525,0.09808825,0.19240387,0.4376245,0.9242931,2.0975795,2.5427492,2.071171,1.7429527,1.7655885,1.2034674,0.7507524,0.7432071,1.146878,1.2185578,0.98842776,0.6451189,0.331991,0.15467763,0.10940613,0.10186087,0.07922512,0.033953626,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.011317875,0.033953626,0.06790725,0.11317875,0.18863125,0.20372175,0.1358145,0.033953626,0.19994913,0.633801,1.1619685,1.569412,1.5882751,1.358145,1.1921495,1.3053282,1.6373192,1.8749946,1.659955,1.4260522,1.2940104,1.2713746,1.2713746,1.0601076,0.95824677,1.086516,1.5769572,2.5917933,2.637065,2.4295704,2.2371666,2.0673985,1.6825907,1.9579924,1.9127209,3.048281,5.2062225,6.5455046,5.587258,4.7535076,4.610148,4.7120085,3.640583,2.7238352,1.9202662,1.750498,1.81086,0.7809334,0.33576363,0.20749438,0.20372175,0.21503963,0.2263575,0.41498876,0.4678055,0.39989826,0.3169005,0.3961256,0.6828451,1.1581959,1.4901869,1.5354583,1.3355093,4.172523,8.480861,11.348056,11.800771,10.774617,9.216523,8.186596,7.4811153,6.571913,4.61392,4.515832,5.6513925,5.5004873,3.7537618,2.2899833,1.4524606,1.8259505,2.1768045,2.2786655,2.9011486,3.399135,3.0256453,2.052308,1.1544232,1.3958713,1.0789708,0.44139713,0.124496624,0.2565385,0.43385187,0.49421388,0.55080324,0.46026024,0.23390275,0.041498873,0.030181,0.08299775,0.08299775,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.049044125,0.049044125,0.0452715,0.10186087,0.392353,0.73566186,0.6149379,0.241448,0.1961765,0.27917424,0.38858038,0.5470306,0.47912338,0.44516975,0.41121614,0.36971724,0.34330887,0.2867195,0.23013012,0.2263575,0.271629,0.32821837,0.211267,0.211267,0.23767537,0.25276586,0.30935526,0.331991,0.35839936,0.41121614,0.452715,0.3961256,0.46026024,0.513077,0.5055317,0.5281675,0.8224323,1.1129243,1.0186088,0.8224323,0.73566186,0.8639311,1.0789708,1.297783,1.3958713,1.3505998,1.2147852,1.3770081,1.5769572,1.5128226,1.2110126,1.0072908,1.0751982,1.1657411,1.2638294,1.3770081,1.5128226,1.4373702,1.0902886,0.724344,0.543258,0.73188925,1.1921495,1.8900851,2.2862108,1.9806281,0.7092535,0.20749438,0.049044125,0.02263575,0.018863125,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.030181,0.06790725,0.06413463,0.011317875,0.00754525,0.033953626,0.06413463,0.09808825,0.08677038,0.041498873,0.0150905,0.0150905,0.011317875,0.02263575,0.033953626,0.05281675,0.08677038,0.13958712,0.14335975,0.13958712,0.16976812,0.21881226,0.19994913,0.15845025,0.08299775,0.02263575,0.00754525,0.030181,0.041498873,0.041498873,0.05281675,0.071679875,0.056589376,0.049044125,0.033953626,0.02263575,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.00754525,0.011317875,0.003772625,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.08677038,0.2678564,0.19240387,0.11317875,0.05281675,0.02263575,0.0,0.13958712,0.58475685,0.94315624,0.995973,0.7167987,0.7469798,1.1695137,1.4071891,1.2185578,0.7205714,0.67152727,0.73566186,0.60362,0.29803738,0.16222288,0.3055826,0.29049212,0.17354076,0.03772625,0.0,0.011317875,0.026408374,0.026408374,0.0150905,0.018863125,0.0150905,0.030181,0.041498873,0.060362,0.116951376,0.17354076,0.20372175,0.21881226,0.271629,0.452715,0.66775465,1.2638294,1.8636768,2.1541688,1.8749946,1.1657411,0.73566186,0.49044126,0.35462674,0.271629,0.19240387,0.1358145,0.124496624,0.13958712,0.10940613,0.07922512,0.09808825,0.094315626,0.05281675,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.003772625,0.0,0.02263575,0.06790725,0.124496624,0.25276586,0.35839936,0.52439487,0.7696155,1.0299267,1.9994912,2.4484336,3.3312278,5.2062225,8.246958,13.396591,19.87419,26.491373,31.995632,35.077866,34.900555,33.263233,31.878681,31.354286,31.207153,30.32436,29.143528,27.970242,26.90636,25.846254,24.046711,22.266033,20.889025,19.794964,18.33873,17.301258,16.59955,16.35433,16.848543,18.523588,19.1008,19.270569,20.225042,22.209444,24.491882,25.676485,26.604551,26.962952,27.215717,28.577635,30.105547,33.002922,35.35704,36.469967,36.851,37.873383,38.25819,38.31478,38.62036,39.98228,42.67216,45.033825,46.456104,47.38417,49.342163,52.118813,53.186466,53.869312,54.816242,56.02348,56.464878,60.06019,66.3982,72.34763,72.05714,63.719635,61.85219,66.18316,74.04908,80.37955,77.184135,73.61146,65.258865,51.764187,36.80573,28.456911,23.446865,20.217497,17.818108,15.8676605,14.3095665,13.705947,13.347548,12.619431,10.989656,10.853842,11.374464,13.060828,15.705438,18.361366,19.229069,20.126955,20.53817,20.440083,20.30804,21.258741,22.107582,22.303759,21.65864,20.349539,18.557543,16.33924,14.769827,13.920986,12.823153,11.989402,11.566868,11.099063,10.431308,9.718282,9.352338,9.352338,9.352338,9.431562,10.114408,10.001229,9.661693,9.035437,8.409182,8.409182,7.7187905,7.01331,6.4021444,5.9494295,5.674028,5.6778007,5.553304,5.3458095,5.032682,4.534695,4.134797,3.7801702,3.440634,3.1124156,2.8181508,2.535204,2.3692086,2.2673476,2.2711203,2.4823873,2.6144292,2.5201135,2.335255,2.1579416,2.052308,2.2296214,2.0485353,1.8523588,1.7618159,1.659955,1.5203679,1.4034165,1.2298758,1.0148361,0.8563859,0.77716076,0.7696155,0.6752999,0.51684964,0.482896,0.44516975,0.38858038,0.30935526,0.24522063,0.2565385,0.07922512,0.27540162,0.513077,0.6187105,0.573439,0.36971724,0.26408374,0.2678564,0.3055826,0.211267,0.17354076,0.211267,0.27540162,0.35085413,0.44516975,0.6111652,0.63002837,0.6790725,0.875249,1.2940104,1.9806281,2.0296721,1.7316349,1.3128735,0.90920264,0.0150905,0.0150905,0.00754525,0.02263575,0.27917424,1.1431054,1.2411937,0.83752275,0.3772625,0.18485862,0.42630664,1.720317,1.0299267,0.22258487,0.10186087,0.38103512,1.0035182,1.0676528,1.3845534,2.1805773,3.097325,2.0485353,1.4298248,1.4411428,1.8749946,2.1202152,2.1579416,1.4524606,0.69039035,0.2263575,0.090543,0.056589376,0.03772625,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026408374,0.041498873,1.1959221,5.8588867,4.395108,1.7957695,0.63002837,1.3204187,2.1503963,6.398372,8.552541,8.341274,6.5341864,4.8968673,3.187868,2.6446102,2.161714,1.7014539,2.2899833,2.0673985,0.98842776,0.21881226,0.071679875,0.0,0.071679875,0.1358145,0.271629,0.4074435,0.32067314,0.11317875,0.02263575,0.0,0.02263575,0.1056335,0.14335975,0.5281675,0.6187105,0.33953625,0.1659955,0.83752275,0.7507524,0.45648763,0.33576363,0.58098423,0.49421388,0.25276586,0.08677038,0.094315626,0.23013012,0.30181,0.24899325,0.1358145,0.09808825,0.3055826,0.5357128,0.5394854,0.72811663,1.5958204,3.7084904,5.149633,3.9688015,2.444661,1.6712729,1.5882751,1.0638802,0.6111652,0.35462674,0.26408374,0.1659955,0.08299775,0.07922512,0.060362,0.0150905,0.0150905,0.003772625,0.00754525,0.00754525,0.003772625,0.0150905,0.003772625,0.0,0.00754525,0.018863125,0.030181,0.06790725,0.06790725,0.06790725,0.071679875,0.0452715,0.14335975,0.331991,0.56589377,0.784706,0.9318384,1.0412445,1.1242423,1.5580941,2.2673476,2.7313805,2.3277097,2.071171,2.1164427,2.4069347,2.7011995,2.0787163,1.3920987,0.995973,0.9922004,1.237421,1.6637276,1.9240388,2.052308,1.9881734,1.5731846,4.429062,2.323937,0.754525,2.3088465,6.6662283,5.583485,4.9534564,5.172269,5.9003854,6.058836,5.1798143,2.8634224,1.4298248,1.2562841,0.7922512,0.41498876,0.28294688,0.241448,0.21503963,0.21503963,0.32444575,0.3772625,0.3734899,0.3961256,0.6413463,0.94692886,0.84884065,1.0676528,1.8259505,2.837014,2.7653341,4.979865,7.2396674,8.541223,9.14107,8.518587,8.790216,8.778898,7.8961043,6.1644692,5.726845,4.817642,3.8292143,3.4142256,4.5007415,3.4745877,5.2250857,5.9796104,5.0741806,4.927048,3.1576872,1.8749946,1.4147344,1.7391801,2.4107075,1.6033657,0.5885295,0.23013012,0.6790725,1.3732355,1.6788181,1.2336484,0.63002837,0.21503963,0.090543,0.12826926,0.41121614,0.422534,0.1358145,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.43007925,0.80356914,0.8941121,0.38103512,0.0754525,0.21881226,0.452715,0.59607476,0.65643674,0.8639311,0.8978847,0.77338815,0.56212115,0.36594462,0.32821837,0.29426476,0.2678564,0.27917424,0.36594462,0.40367088,0.392353,0.29049212,0.22258487,0.5017591,0.724344,0.62248313,0.4640329,0.3961256,0.45648763,0.5319401,0.52062225,0.47912338,0.482896,0.6413463,0.8224323,0.8601585,0.7507524,0.6073926,0.65643674,0.8526133,0.9922004,0.90543,0.63002837,0.3961256,0.63002837,0.9997456,1.3204187,1.5807298,1.9240388,2.214531,2.2069857,2.071171,1.9051756,1.7089992,1.6222287,1.4637785,1.1581959,0.9280658,1.2826926,1.1355602,0.7884786,0.3772625,0.06413463,0.0150905,0.026408374,0.02263575,0.02263575,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.030181,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.018863125,0.03772625,0.041498873,0.0150905,0.003772625,0.00754525,0.0754525,0.16976812,0.18485862,0.120724,0.05281675,0.0150905,0.011317875,0.0,0.0,0.00754525,0.033953626,0.07922512,0.150905,0.116951376,0.116951376,0.15845025,0.22258487,0.26031113,0.211267,0.124496624,0.0452715,0.00754525,0.030181,0.041498873,0.056589376,0.06790725,0.08299775,0.1056335,0.056589376,0.026408374,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.00754525,0.011317875,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.030181,0.18485862,0.6111652,0.27917424,0.1056335,0.041498873,0.02263575,0.0,0.011317875,0.24522063,0.513077,0.6790725,0.65643674,0.8526133,1.3770081,1.7957695,1.8561316,1.4637785,1.0751982,0.8111144,0.52439487,0.23390275,0.1358145,0.271629,0.34330887,0.2678564,0.09808825,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.018863125,0.0150905,0.026408374,0.056589376,0.090543,0.07922512,0.049044125,0.060362,0.120724,0.18485862,0.27917424,0.8262049,1.4600059,2.0598533,2.7313805,1.6675003,0.935611,0.5885295,0.5394854,0.56589377,0.30935526,0.14335975,0.071679875,0.060362,0.060362,0.049044125,0.03772625,0.018863125,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.00754525,0.0150905,0.0150905,0.026408374,0.094315626,0.29049212,0.60362,0.94692886,1.056335,1.3128735,1.8372684,2.8030603,4.425289,8.209232,13.713491,20.813572,29.39252,39.352253,46.467422,48.787586,48.71968,47.931202,47.331352,46.731506,45.852486,44.577335,42.728752,40.06905,36.334152,33.11233,30.773302,29.143528,27.49489,25.174726,23.314823,21.892544,21.258741,22.126446,22.624432,23.1526,23.514772,23.782627,24.307022,25.79721,27.668432,29.641514,31.422194,32.716206,33.482048,34.77606,36.386967,38.220463,40.28409,41.917637,44.39625,46.625874,48.078335,48.79513,50.02878,50.183456,50.549404,52.46967,57.325035,61.086346,60.362,57.86452,56.000847,56.85346,58.622818,63.553642,71.70628,78.746,75.92785,64.074265,57.679665,57.28731,60.814716,63.52346,66.33029,70.42736,68.0242,56.65351,39.186256,31.882454,28.019285,24.118391,19.825144,17.882242,15.954432,15.599804,15.490398,14.920732,13.807808,13.468271,13.226823,13.536179,14.920732,17.961468,20.534397,23.277096,24.257978,23.458181,22.748928,22.081175,22.726294,23.34123,23.48459,23.620405,22.288668,20.704166,19.025349,17.120173,14.558559,13.422999,12.725064,12.336484,12.1252165,11.978085,10.831206,10.012547,9.420244,9.148616,9.491924,10.005001,10.582213,11.329193,12.019584,12.068627,9.699419,7.9451485,6.9152217,6.417235,5.96452,6.138061,5.915476,5.798525,5.7306175,5.0968165,4.606375,4.1762958,3.7952607,3.440634,3.0520537,2.6974268,2.463524,2.335255,2.3126192,2.4107075,2.8143783,3.0520537,3.0331905,2.8332415,2.686109,3.150142,2.704972,2.384299,2.3314822,1.8297231,1.8561316,1.8976303,1.7693611,1.478869,1.237421,1.0789708,0.94692886,0.9695646,1.0789708,1.0072908,0.77338815,0.62625575,0.47912338,0.34330887,0.3055826,0.20749438,0.12826926,0.2867195,0.55080324,0.42630664,0.29426476,0.46026024,0.7469798,0.88279426,0.5017591,0.17354076,0.10940613,0.13958712,0.18863125,0.27540162,0.422534,0.45648763,0.56589377,0.84129536,1.2826926,1.5015048,1.4373702,1.3015556,1.2638294,1.4335974,0.003772625,0.05281675,0.1358145,0.35085413,0.55457586,0.3772625,1.3920987,2.3126192,1.7618159,0.41121614,0.97710985,1.3317367,1.0940613,0.8337501,0.7092535,0.44139713,0.6073926,0.9808825,1.4637785,1.7995421,1.5731846,1.478869,3.6896272,4.429062,2.8936033,1.2525115,1.2600567,1.5958204,1.6033657,1.1883769,0.8111144,0.73566186,0.34330887,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.05281675,0.44139713,1.7354075,1.2562841,0.70170826,0.5281675,0.91674787,1.7844516,5.6513925,8.009283,8.054554,6.598321,6.058836,4.8742313,3.6254926,2.637065,2.6898816,5.0213637,3.0445085,1.2638294,0.55080324,0.6752999,0.27917424,0.090543,0.05281675,0.10940613,0.16976812,0.124496624,0.11317875,0.0452715,0.071679875,0.150905,0.02263575,0.049044125,0.20372175,0.241448,0.14335975,0.120724,0.28294688,0.2565385,0.241448,0.35462674,0.6149379,0.72811663,0.66775465,0.4376245,0.16222288,0.08299775,0.17354076,0.21881226,0.18863125,0.38480774,1.4524606,2.444661,3.2859564,4.825187,6.4210076,5.915476,4.6931453,3.85185,3.4444065,3.2331395,2.7087448,1.3958713,0.5696664,0.211267,0.14713238,0.071679875,0.033953626,0.056589376,0.05281675,0.011317875,0.003772625,0.0,0.0,0.00754525,0.011317875,0.0150905,0.011317875,0.003772625,0.0,0.00754525,0.018863125,0.026408374,0.049044125,0.071679875,0.08677038,0.08299775,0.13204187,0.241448,0.362172,0.47535074,0.5998474,0.60362,0.5583485,0.70170826,1.1355602,1.8033148,2.2107582,2.2899833,2.2107582,2.1088974,2.0787163,1.8070874,1.4637785,1.2336484,1.1619685,1.1619685,1.3656902,3.1840954,3.9348478,2.9841464,1.7316349,2.214531,1.4713237,0.8601585,1.1619685,2.5804756,3.229367,3.651901,4.9685473,6.8133607,7.3151197,5.772116,3.7235808,3.1312788,3.8141239,3.4179983,1.3807807,0.62248313,0.5696664,0.8978847,1.5430037,2.425798,2.4974778,2.071171,1.7089992,2.214531,1.6033657,0.83752275,0.4376245,0.513077,0.77338815,0.91674787,1.4071891,2.674791,4.5497856,6.270103,7.152897,6.930312,6.881268,7.2698483,7.360391,7.752744,5.726845,4.055572,3.6179473,3.4142256,3.6783094,3.8669407,3.9461658,4.006528,4.2819295,4.1800685,2.6332922,1.3166461,0.9318384,1.2034674,0.8865669,0.38480774,0.18863125,0.3470815,0.49421388,0.7507524,0.724344,0.56589377,0.513077,0.8978847,1.7429527,1.3807807,0.69039035,0.19240387,0.049044125,0.03772625,0.02263575,0.00754525,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.08677038,0.2678564,0.43007925,0.4376245,0.29049212,0.1358145,0.116951376,0.15467763,0.2263575,0.29803738,0.35085413,0.41121614,0.3734899,0.27540162,0.18485862,0.18485862,0.392353,0.422534,0.35839936,0.30935526,0.41498876,0.6752999,0.84884065,0.77338815,0.52439487,0.4074435,0.392353,0.47535074,0.47157812,0.35839936,0.27540162,0.33953625,0.362172,0.5017591,0.7469798,0.94692886,0.69793564,0.5772116,0.6073926,0.7205714,0.7432071,0.58475685,0.573439,0.52062225,0.40367088,0.3470815,0.56212115,0.8526133,1.1732863,1.4977322,1.7995421,2.123988,2.354118,2.3578906,2.161714,1.9655377,2.0560806,2.0862615,1.9391292,1.6109109,1.2336484,0.65643674,0.3470815,0.211267,0.1659955,0.124496624,0.15845025,0.1056335,0.0452715,0.018863125,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.018863125,0.026408374,0.018863125,0.0150905,0.0150905,0.011317875,0.011317875,0.0,0.0,0.003772625,0.00754525,0.00754525,0.003772625,0.0,0.00754525,0.03772625,0.08677038,0.14713238,0.17354076,0.116951376,0.0452715,0.003772625,0.011317875,0.030181,0.030181,0.02263575,0.033953626,0.116951376,0.10940613,0.10186087,0.13958712,0.20749438,0.22258487,0.1358145,0.08299775,0.03772625,0.0,0.00754525,0.03772625,0.06413463,0.06790725,0.060362,0.0452715,0.026408374,0.011317875,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0150905,0.071679875,0.1961765,0.10186087,0.041498873,0.018863125,0.0150905,0.0,0.003772625,0.11317875,0.271629,0.40367088,0.4376245,0.4640329,0.7582976,1.2562841,1.720317,1.720317,0.9507015,0.44516975,0.17354076,0.08677038,0.124496624,0.211267,0.20372175,0.124496624,0.030181,0.0,0.0,0.0150905,0.0150905,0.003772625,0.00754525,0.003772625,0.003772625,0.003772625,0.0150905,0.030181,0.03772625,0.026408374,0.033953626,0.071679875,0.1358145,0.20372175,0.543258,0.8865669,1.0902886,1.1581959,0.8865669,0.6526641,0.49421388,0.3961256,0.28294688,0.18485862,0.13958712,0.15467763,0.17731337,0.09808825,0.094315626,0.07922512,0.041498873,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.018863125,0.026408374,0.030181,0.071679875,0.1961765,0.44894236,0.90920264,1.448688,2.0560806,2.3880715,2.5125682,2.886058,4.2592936,6.8397694,10.902886,16.867407,25.314314,36.496376,46.456104,53.352463,55.880123,53.288326,50.54186,47.52753,44.82256,42.66839,40.985798,39.52579,38.307236,37.303715,36.13043,34.051712,32.376667,30.939297,30.090458,29.852781,29.95087,29.660378,29.309525,28.905853,28.592726,28.626678,29.207663,31.199608,34.557243,38.81654,43.090923,42.91361,41.959137,42.14022,43.800175,45.72799,47.31249,49.112034,51.213383,53.49205,55.608494,55.974438,54.054173,51.534058,50.134415,51.601963,54.75588,55.84994,55.84617,56.03857,58.026745,61.15425,65.496544,69.92183,71.97037,67.8733,61.22216,59.467888,61.531513,64.71938,64.69297,69.62002,77.25959,77.470856,66.89619,48.94981,39.499382,33.07083,28.207916,24.269297,21.398329,19.94964,18.75372,17.444618,16.180788,15.663939,16.414692,16.237377,15.992157,16.263786,17.350302,19.183798,22.039675,24.386248,25.533127,25.593489,25.559534,25.442583,25.189817,24.846508,24.55979,23.892035,23.001694,22.043447,20.700394,18.157644,17.365393,15.230087,13.671993,13.211733,12.966512,12.336484,11.98563,11.393328,10.612394,10.26154,10.695392,10.789707,10.880251,11.208468,11.910177,11.680047,11.25374,10.344538,9.016574,7.6886096,7.1566696,6.609639,6.1833324,5.855114,5.4740787,5.6400743,5.481624,4.9647746,4.2706113,3.783943,3.5085413,3.1010978,2.7917426,2.6597006,2.6295197,3.0030096,3.338773,3.451952,3.410453,3.5274043,3.572676,3.500996,3.2935016,2.916239,2.3201644,2.1202152,2.0258996,1.9127209,1.7278622,1.4939595,1.2864652,1.2600567,1.3694628,1.4335974,1.1053791,1.2147852,1.1808317,0.9808825,0.73566186,0.7092535,0.63002837,0.5998474,0.69793564,0.8186596,0.66020936,0.45648763,0.47535074,0.7394345,0.91674787,0.34330887,0.21881226,0.30935526,0.38480774,0.36594462,0.33576363,0.422534,0.56212115,0.7167987,1.026154,1.8184053,2.0673985,2.003264,1.8636768,1.8184053,1.9579924,0.00754525,0.071679875,0.38103512,0.633801,0.62248313,0.211267,1.1242423,2.0673985,1.8146327,0.79602385,1.0789708,2.655928,2.3956168,1.629774,1.0186088,0.55080324,1.0450171,1.1695137,1.086516,1.026154,1.2826926,1.2600567,2.6106565,3.1161883,2.335255,1.6146835,1.4298248,1.6335466,1.4939595,1.0638802,1.1657411,1.3091009,1.0940613,0.6375736,0.16976812,0.056589376,0.033953626,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026408374,0.15467763,0.52062225,0.3734899,0.27540162,0.32067314,0.6828451,1.5731846,5.0251365,6.6813188,6.6549106,5.753253,5.4778514,4.957229,3.7273536,3.229367,3.4557245,2.9615107,1.5165952,0.66775465,0.7092535,1.0638802,0.2867195,0.090543,0.094315626,0.14335975,0.14335975,0.0754525,0.12826926,0.07922512,0.07922512,0.120724,0.00754525,0.056589376,0.16976812,0.241448,0.26408374,0.33576363,0.29049212,0.25276586,0.3470815,0.5583485,0.7167987,0.60362,0.46026024,0.27917424,0.1056335,0.0452715,0.071679875,0.094315626,0.090543,0.4074435,1.7844516,2.6332922,3.440634,4.3196554,4.8553686,4.134797,3.7650797,2.9992368,2.2975287,1.9202662,1.9278114,1.2223305,0.482896,0.094315626,0.06413463,0.026408374,0.011317875,0.02263575,0.02263575,0.011317875,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.0150905,0.011317875,0.003772625,0.0,0.00754525,0.0150905,0.026408374,0.049044125,0.07922512,0.10186087,0.116951376,0.14713238,0.20372175,0.3055826,0.47157812,0.5055317,0.48666862,0.66775465,1.2223305,2.2598023,2.9766011,3.0369632,2.7389257,2.372981,2.1881225,1.9466745,1.6373192,1.418507,1.3392819,1.3355093,1.3355093,2.173032,2.535204,2.1956677,1.9994912,3.5085413,3.2633207,1.9806281,0.7809334,1.1619685,2.4974778,3.6896272,4.636556,5.3646727,6.009792,5.458988,3.874486,2.9992368,3.218049,3.5424948,2.8558772,2.1541688,1.5656394,1.1921495,1.1355602,1.5882751,1.7655885,1.6184561,1.5543215,2.4371157,3.3274553,3.2670932,3.1312788,2.9200118,1.780679,1.5279131,1.7467253,2.384299,3.3350005,4.4743333,6.9454026,8.160188,8.477088,8.160188,7.3490734,7.6886096,6.3455553,4.889322,4.134797,4.123479,4.13857,3.8141239,3.3538637,3.187868,3.983892,4.285702,2.8256962,1.5580941,1.1921495,1.2034674,0.8111144,0.9016574,1.1808317,1.2487389,0.58475685,0.42630664,0.9016574,1.4260522,1.659955,1.4826416,1.6335466,1.2110126,0.7997965,0.69793564,0.9393836,0.452715,0.13958712,0.011317875,0.049044125,0.211267,0.14335975,0.071679875,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.026408374,0.011317875,0.00754525,0.026408374,0.071679875,0.1961765,0.32444575,0.31312788,0.25276586,0.47157812,0.1961765,0.13204187,0.16976812,0.22258487,0.21881226,0.18485862,0.124496624,0.08299775,0.10186087,0.211267,0.41876137,0.482896,0.46026024,0.44894236,0.573439,0.694163,0.6451189,0.49421388,0.32067314,0.2263575,0.24899325,0.3169005,0.3734899,0.39989826,0.43007925,0.43385187,0.45648763,0.55457586,0.724344,0.9016574,0.5281675,0.33953625,0.43385187,0.68661773,0.72811663,0.6488915,0.633801,0.69039035,0.8186596,1.0148361,0.875249,0.84129536,0.814887,0.80356914,0.9280658,1.1846043,1.3996439,1.5769572,1.8297231,2.3692086,2.7011995,2.3993895,1.8674494,1.297783,0.7092535,0.2678564,0.09808825,0.071679875,0.08677038,0.07922512,0.10186087,0.06790725,0.033953626,0.02263575,0.0150905,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.011317875,0.00754525,0.0150905,0.011317875,0.00754525,0.003772625,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.03772625,0.08299775,0.13204187,0.124496624,0.071679875,0.0150905,0.00754525,0.030181,0.026408374,0.011317875,0.011317875,0.060362,0.060362,0.06413463,0.09808825,0.150905,0.150905,0.094315626,0.060362,0.026408374,0.0,0.0,0.0150905,0.03772625,0.041498873,0.030181,0.011317875,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.090543,0.08299775,0.041498873,0.011317875,0.003772625,0.0,0.0,0.03772625,0.120724,0.23767537,0.392353,0.33576363,0.35085413,0.6375736,1.1317875,1.4939595,0.845068,0.30935526,0.041498873,0.018863125,0.049044125,0.07922512,0.06790725,0.033953626,0.003772625,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.011317875,0.0150905,0.0150905,0.02263575,0.049044125,0.13204187,0.27917424,0.40367088,0.4678055,0.47157812,0.49044126,0.482896,0.41498876,0.33953625,0.36971724,0.5055317,0.452715,0.3470815,0.23767537,0.08677038,0.08677038,0.060362,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.02263575,0.030181,0.06790725,0.15467763,0.34330887,0.7092535,1.3694628,2.1881225,2.776652,3.048281,3.199186,3.6066296,4.5007415,6.187105,9.201432,14.290704,22.982832,33.16892,42.86834,50.138187,53.084606,51.83587,48.648,44.99987,41.86859,39.740833,38.85049,37.669662,36.624645,35.738075,34.628925,33.606544,32.316307,31.739094,32.00695,32.399303,31.912636,31.735321,31.739094,31.825865,31.96168,31.874908,32.9237,35.88521,40.00869,43.011696,43.841675,43.355007,42.845703,42.702343,42.374123,42.03836,42.06477,43.09847,44.8716,46.180702,47.636936,48.00288,47.237038,45.799667,44.64147,45.822304,47.09745,48.757404,51.402016,55.955574,60.282776,62.79534,62.999065,60.86753,56.823277,54.793606,56.51015,61.56924,68.133606,72.93239,79.364716,80.63232,74.07549,61.508877,49.24785,44.16235,38.582638,32.984062,28.162645,25.253952,24.148573,22.567842,20.873934,19.40261,18.43682,18.704676,18.327412,18.002966,18.055782,18.406637,19.123436,20.806026,22.914925,24.888006,26.1707,27.015768,27.547709,27.819336,27.770292,27.24967,26.1707,25.227543,24.352295,23.394047,22.141537,21.911406,20.206179,18.221779,16.516552,15.026365,14.019074,13.479589,13.12119,12.947649,13.234368,12.985375,12.694883,12.1252165,11.427281,11.129244,11.902632,12.245941,12.042219,11.404645,10.691619,9.601331,8.20546,7.039718,6.3116016,5.8890676,5.9796104,5.7909794,5.5306683,5.2137675,4.708236,4.3724723,4.115934,3.904667,3.6783094,3.3463185,3.3878171,3.4670424,3.591539,3.783943,4.0782075,4.0517993,3.8895764,3.6368105,3.2859564,2.7879698,3.0218725,2.8106055,2.5767028,2.3503454,1.7655885,1.5543215,1.418507,1.3694628,1.3845534,1.4034165,1.4222796,1.3015556,1.1695137,1.0978339,1.1091517,1.0525624,0.9280658,0.9620194,1.0676528,0.8526133,0.5394854,0.47535074,0.59607476,0.7130261,0.51684964,0.44139713,0.5055317,0.62625575,0.7394345,0.7809334,0.8978847,1.0186088,1.1204696,1.358145,2.052308,2.493705,2.916239,2.8898308,2.4672968,2.1654868,0.00754525,0.049044125,0.482896,1.3053282,1.9127209,1.1091517,1.0940613,1.2600567,1.2110126,0.9922004,1.0827434,2.7691069,3.2105038,2.727608,1.7580433,0.8224323,1.5430037,1.3732355,0.91297525,0.663982,1.0374719,0.8941121,1.0299267,1.1695137,1.3543724,1.9693103,2.2069857,1.8561316,1.3166461,0.9507015,1.0978339,1.3996439,1.4449154,1.0299267,0.43007925,0.40367088,0.30181,0.11317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.06413463,0.2867195,0.20749438,0.13958712,0.95447415,2.3013012,2.6295197,8.145098,9.469289,8.922258,8.224322,8.503497,6.828451,4.357382,3.0860074,2.7351532,0.7394345,0.21881226,0.14713238,0.4640329,0.73566186,0.15845025,0.116951376,0.18485862,0.20372175,0.14335975,0.0754525,0.09808825,0.06790725,0.05281675,0.056589376,0.02263575,0.06413463,0.17354076,0.271629,0.35085413,0.452715,0.35085413,0.3055826,0.39989826,0.5583485,0.55080324,0.35839936,0.24899325,0.1659955,0.116951376,0.16222288,0.15845025,0.13204187,0.11317875,0.34330887,1.3166461,1.7089992,2.4031622,2.7804246,2.8143783,3.059599,3.7801702,2.6823363,1.3807807,0.86770374,1.5241405,1.1544232,0.5055317,0.124496624,0.08677038,0.0150905,0.003772625,0.0,0.00754525,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.00754525,0.0,0.0,0.011317875,0.0150905,0.026408374,0.05281675,0.08677038,0.10186087,0.09808825,0.10940613,0.16976812,0.30935526,0.36594462,0.4074435,0.694163,1.4147344,2.674791,3.5236318,3.4029078,2.9086938,2.5125682,2.5616124,2.535204,2.1843498,1.7995421,1.5543215,1.4901869,1.3958713,1.3392819,1.4071891,1.7655885,2.674791,4.191386,3.712263,2.1805773,0.7507524,0.79602385,1.7542707,2.8332415,3.3915899,3.5953116,4.447925,4.6327834,3.5274043,2.3465726,1.9466745,2.8407867,3.7160356,3.6292653,3.108643,2.6295197,2.6182017,2.293756,1.7995421,1.4335974,1.4939595,2.263575,3.7877154,4.515832,4.772371,4.4931965,3.2067313,2.5389767,2.3126192,2.203213,2.2296214,2.7653341,6.2399216,8.68081,9.563604,8.944894,7.488661,7.4509344,6.360646,5.1571784,4.587512,5.2137675,4.5497856,3.7499893,2.9652832,2.5917933,3.2520027,3.3236825,2.3993895,1.6335466,1.3958713,1.2826926,1.1959221,1.4562333,1.8485862,1.9957186,1.3543724,1.1431054,1.5769572,1.9730829,2.0145817,1.7467253,1.5618668,1.2864652,1.1280149,1.1506506,1.2525115,0.56212115,0.17354076,0.030181,0.08299775,0.271629,0.181086,0.09808825,0.03772625,0.00754525,0.0,0.0,0.0,0.011317875,0.0452715,0.09808825,0.0452715,0.0150905,0.030181,0.094315626,0.16222288,0.21503963,0.29426476,0.30181,0.38858038,0.94692886,0.422534,0.2263575,0.18863125,0.1961765,0.18485862,0.1056335,0.090543,0.13958712,0.23013012,0.331991,0.4979865,0.5998474,0.60362,0.5696664,0.633801,0.5885295,0.392353,0.2263575,0.150905,0.13958712,0.17354076,0.23767537,0.331991,0.41876137,0.44139713,0.41876137,0.41498876,0.422534,0.47912338,0.63002837,0.41876137,0.2867195,0.35462674,0.5583485,0.6451189,0.6828451,0.663982,0.7432071,0.9205205,1.026154,0.7809334,0.8111144,0.7997965,0.6375736,0.44516975,0.69039035,1.0336993,1.2789198,1.5769572,2.4220252,2.3201644,1.7278622,1.0940613,0.6111652,0.2263575,0.06413463,0.033953626,0.0452715,0.041498873,0.018863125,0.026408374,0.0150905,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0150905,0.018863125,0.018863125,0.0150905,0.018863125,0.0150905,0.011317875,0.003772625,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.026408374,0.06790725,0.120724,0.150905,0.124496624,0.00754525,0.02263575,0.02263575,0.0150905,0.011317875,0.02263575,0.033953626,0.049044125,0.0754525,0.094315626,0.0754525,0.060362,0.03772625,0.0150905,0.0,0.0,0.0,0.0150905,0.018863125,0.00754525,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.056589376,0.05281675,0.026408374,0.018863125,0.090543,0.13204187,0.090543,0.03772625,0.003772625,0.0,0.0,0.003772625,0.033953626,0.120724,0.31312788,0.29803738,0.17354076,0.20749438,0.49044126,0.9205205,0.55457586,0.19994913,0.0150905,0.018863125,0.071679875,0.0150905,0.0,0.0,0.0,0.00754525,0.0,0.0,0.003772625,0.0150905,0.018863125,0.00754525,0.00754525,0.003772625,0.0,0.00754525,0.00754525,0.011317875,0.00754525,0.0,0.00754525,0.07922512,0.12826926,0.1659955,0.21881226,0.32444575,0.40367088,0.41498876,0.38103512,0.4376245,0.83752275,1.1016065,0.86770374,0.5055317,0.23013012,0.10186087,0.0754525,0.033953626,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.060362,0.120724,0.23767537,0.4640329,1.0525624,1.8599042,2.5880208,3.0860074,3.3274553,3.500996,3.7462165,4.236658,5.311856,7.466025,12.004493,19.059301,28.02683,37.71116,46.33538,50.70408,51.085114,48.598957,44.532066,40.35577,38.424187,36.598236,35.119366,34.168663,33.866856,33.451866,32.286125,31.493874,31.376923,31.399557,31.063795,31.222244,31.358059,31.452375,31.99186,32.13522,32.81052,34.9081,37.937515,40.02755,41.668644,42.143993,41.298927,39.42016,37.22449,36.156837,36.066296,37.00568,38.277054,38.458138,40.186,42.966427,45.12814,45.810986,44.96969,45.060234,46.056206,48.168877,51.59442,56.517696,60.77699,62.757618,62.259632,59.58861,55.555676,52.620575,52.67339,55.570766,60.89394,67.96007,72.90221,69.05413,60.0451,50.383408,45.448814,44.8301,41.77805,37.14904,32.289898,29.041668,27.49489,25.917934,24.567333,23.443092,22.311304,21.55678,20.8513,20.52308,20.526854,20.424992,20.274086,20.85507,22.043447,23.609087,25.19359,26.581915,27.830654,28.996395,29.958416,30.429993,29.754694,28.845491,27.785383,26.68755,25.672712,25.631214,24.888006,23.345003,21.23988,19.146072,17.467255,16.177015,15.475307,15.331948,15.497944,15.086727,15.135772,14.841507,13.977575,12.868423,12.902377,12.917468,12.898605,12.868423,12.875969,12.162943,10.725573,9.21275,8.016829,7.281166,6.730363,6.40969,6.1908774,5.904158,5.342037,5.142088,5.1873593,5.2779026,5.1571784,4.496969,4.244203,4.06689,4.044254,4.191386,4.432834,4.504514,4.236658,3.9386206,3.7047176,3.4179983,3.4142256,3.2482302,3.2670932,3.2482302,2.4182527,2.173032,1.8599042,1.5618668,1.3958713,1.5430037,1.4901869,1.2789198,1.2525115,1.4335974,1.4939595,1.6524098,1.4260522,1.297783,1.3015556,1.0374719,0.814887,0.6413463,0.5772116,0.60362,0.63002837,0.65643674,0.6413463,0.7054809,0.8563859,0.9695646,1.1506506,1.3015556,1.4335974,1.690136,2.372981,2.916239,3.5689032,3.5990841,2.9426475,2.1805773,0.018863125,0.033953626,0.3734899,1.8221779,3.4896781,2.7917426,2.123988,1.2298758,0.7696155,0.8337501,0.97710985,1.4713237,2.8143783,3.1954134,2.2296214,0.97333723,1.4977322,1.7919968,1.7014539,1.2487389,0.6413463,0.49044126,0.3470815,0.31312788,0.6111652,1.5845025,2.546522,1.9806281,1.3920987,1.3053282,1.2713746,1.1619685,1.1695137,0.95447415,0.63002837,0.72811663,0.56589377,0.21881226,0.00754525,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.14335975,0.05281675,0.08299775,1.9051756,4.745962,5.379763,12.106354,13.777626,13.392818,12.845788,12.940104,8.854351,4.7346444,2.0673985,0.95824677,0.14335975,0.041498873,0.02263575,0.0150905,0.003772625,0.026408374,0.1358145,0.20372175,0.181086,0.094315626,0.06413463,0.03772625,0.026408374,0.03772625,0.060362,0.03772625,0.03772625,0.120724,0.2263575,0.35462674,0.5470306,0.3734899,0.32821837,0.35839936,0.392353,0.30181,0.36971724,0.4074435,0.33576363,0.21881226,0.29049212,0.32821837,0.3055826,0.26031113,0.29426476,0.543258,0.7469798,1.4826416,2.0485353,2.474842,3.5160866,4.06689,2.6597006,1.2411937,0.84884065,1.6109109,1.056335,0.5055317,0.20749438,0.14335975,0.011317875,0.003772625,0.0,0.00754525,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.00754525,0.003772625,0.0,0.011317875,0.011317875,0.0150905,0.02263575,0.05281675,0.08677038,0.094315626,0.07922512,0.060362,0.08677038,0.116951376,0.17731337,0.4678055,1.146878,2.3088465,3.361409,3.2784111,2.757789,2.4182527,2.7879698,3.1010978,2.7841973,2.2560298,1.7957695,1.5618668,1.50905,1.5165952,1.6486372,2.0900342,3.1237335,3.0445085,2.2862108,1.5279131,1.0487897,0.72811663,0.84129536,1.3920987,2.1013522,2.848332,3.6896272,4.014073,3.5085413,2.474842,1.6184561,2.052308,3.3878171,4.0291634,4.2630663,4.5460134,5.534441,4.949684,3.519859,2.4484336,2.1654868,2.3201644,2.7992878,3.7952607,4.395108,4.3875628,4.2517486,4.3309736,3.31991,1.9768555,1.1355602,1.6939086,4.9987283,7.8961043,9.178797,8.952439,8.646856,7.937603,6.541732,5.704209,5.7872066,6.273875,4.949684,3.4783602,2.5087957,2.1956677,2.1881225,1.9278114,1.7731338,1.5467763,1.3053282,1.3053282,1.6561824,1.7278622,1.8976303,2.2258487,2.463524,2.7502437,2.6068838,2.0900342,1.5618668,1.7089992,1.8448136,1.6486372,1.4147344,1.1921495,0.77338815,0.33953625,0.23013012,0.3055826,0.41498876,0.38858038,0.181086,0.12826926,0.120724,0.090543,0.026408374,0.00754525,0.0,0.026408374,0.08677038,0.16222288,0.0452715,0.03772625,0.120724,0.23767537,0.32067314,0.35462674,0.32067314,0.2867195,0.44516975,1.1091517,0.6187105,0.32444575,0.18485862,0.14713238,0.15845025,0.08677038,0.15467763,0.28294688,0.40367088,0.47535074,0.6187105,0.73188925,0.7054809,0.5772116,0.5357128,0.46026024,0.35085413,0.26031113,0.211267,0.1659955,0.14335975,0.23390275,0.32821837,0.34330887,0.2263575,0.22258487,0.181086,0.15467763,0.18485862,0.32821837,0.38103512,0.35462674,0.3470815,0.41121614,0.5470306,0.6111652,0.5470306,0.5394854,0.55457586,0.35839936,0.35085413,0.7696155,1.0789708,1.0223814,0.5998474,0.875249,1.2902378,1.3770081,1.2751472,1.7316349,0.97333723,0.452715,0.16222288,0.05281675,0.011317875,0.02263575,0.06413463,0.08677038,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.0150905,0.018863125,0.026408374,0.030181,0.033953626,0.041498873,0.018863125,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.124496624,0.2867195,0.35085413,0.018863125,0.0150905,0.02263575,0.02263575,0.011317875,0.011317875,0.033953626,0.06413463,0.06790725,0.0452715,0.02263575,0.02263575,0.018863125,0.00754525,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.116951376,0.120724,0.06413463,0.0150905,0.071679875,0.14713238,0.13204187,0.071679875,0.011317875,0.0,0.0,0.0,0.0,0.030181,0.14713238,0.23767537,0.16976812,0.08299775,0.1056335,0.32821837,0.20749438,0.1056335,0.0452715,0.05281675,0.150905,0.033953626,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0150905,0.03772625,0.049044125,0.02263575,0.0150905,0.00754525,0.0,0.0,0.011317875,0.011317875,0.00754525,0.003772625,0.011317875,0.0452715,0.07922512,0.124496624,0.20372175,0.35085413,0.41121614,0.3734899,0.36594462,0.62625575,1.4977322,1.659955,1.1657411,0.5696664,0.19240387,0.124496624,0.06413463,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.02263575,0.0452715,0.0754525,0.13958712,0.27917424,0.7054809,1.327964,1.9429018,2.4371157,2.7540162,2.938875,3.1652324,3.4783602,4.002755,4.930821,6.330465,9.865415,15.814844,24.005213,33.821583,43.96617,50.424904,52.72998,51.002117,45.965664,41.129158,37.51121,34.987324,33.51977,33.16892,33.063286,32.286125,31.259972,30.169682,28.954897,28.551226,28.468227,28.08342,27.702385,28.566317,29.56229,30.686531,32.157856,34.08944,36.47374,38.137466,39.16362,38.548683,36.436012,34.093212,34.300705,36.30397,38.737312,40.389725,40.204865,40.8198,43.54741,46.701324,49.25162,50.817257,52.160313,53.95608,56.110252,58.385143,60.38841,62.882114,65.9304,68.74854,69.74452,66.50383,58.505867,52.79034,49.666607,49.80242,54.22771,53.684452,48.255646,42.743843,39.80874,39.929462,41.00089,40.548172,38.62036,35.64376,32.429485,30.169682,28.732311,27.811792,27.117628,26.389511,24.974777,24.088211,23.680767,23.4695,22.933788,22.56407,22.65084,22.933788,23.39782,24.27307,25.544443,26.740366,28.238098,30.158363,32.357803,33.165146,33.021786,32.327625,31.15811,29.268024,28.528591,28.01174,27.053493,25.56708,24.016531,22.08872,20.213724,18.859352,17.95015,16.856089,16.497688,17.184307,17.784155,17.738882,17.105082,15.860115,15.030138,14.468017,14.154889,14.222796,14.298248,13.751218,12.6345215,11.2801485,10.280403,8.899622,8.20546,7.496206,6.6020937,5.885295,5.8588867,6.0814714,6.4134626,6.519096,5.8626595,5.5268955,5.3194013,5.160951,5.0477724,5.0515447,5.1081343,4.7950063,4.432834,4.172523,3.983892,3.1954134,3.1840954,3.6858547,4.06689,3.3274553,3.0633714,2.6446102,2.2220762,1.8825399,1.6260014,1.7278622,1.4373702,1.4147344,1.7014539,1.750498,2.2560298,2.0485353,1.7240896,1.5241405,1.3468271,1.358145,1.0751982,0.8299775,0.73566186,0.663982,0.7922512,0.72811663,0.68661773,0.7582976,0.91297525,1.0110635,1.1996948,1.418507,1.780679,2.5804756,3.1199608,3.6179473,3.6481283,3.1199608,2.282438,0.090543,0.116951376,0.15845025,0.694163,2.022127,4.255521,5.2099953,3.5047686,1.4600059,0.34330887,0.36594462,1.2826926,1.4939595,1.0148361,0.31312788,0.29049212,0.47157812,3.0897799,4.3196554,3.0445085,0.8865669,0.77338815,0.5017591,0.29803738,0.241448,0.23013012,0.8526133,1.1355602,1.3845534,1.9202662,3.0671442,1.2487389,0.663982,0.58098423,0.4979865,0.16976812,0.13204187,0.049044125,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.030181,0.1056335,0.23013012,0.071679875,0.030181,1.1846043,4.244203,9.567377,7.454707,9.5183325,12.37421,13.060828,9.031664,4.3347464,1.8787673,0.7432071,0.27917424,0.1056335,0.033953626,0.00754525,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.011317875,0.026408374,0.0150905,0.026408374,0.041498873,0.1056335,0.16976812,0.060362,0.011317875,0.08299775,0.23390275,0.5357128,1.1431054,0.72811663,0.56212115,0.5055317,0.52062225,0.65643674,1.1808317,1.1016065,0.7092535,0.29049212,0.1056335,0.20372175,0.27540162,0.27917424,0.2867195,0.45648763,1.2751472,1.901403,2.1956677,2.2598023,2.4408884,1.8674494,1.1921495,0.6187105,0.2565385,0.120724,0.03772625,0.033953626,0.041498873,0.02263575,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.041498873,0.08299775,0.094315626,0.06413463,0.0150905,0.0150905,0.0150905,0.1056335,0.41498876,1.0978339,2.6106565,3.3463185,3.1652324,2.5314314,2.5314314,2.6672459,2.535204,2.2862108,2.003264,1.7089992,1.780679,1.901403,1.9127209,1.8146327,1.7542707,1.7542707,1.9089483,2.123988,2.0447628,1.0676528,1.056335,2.2069857,3.3048196,3.7499893,3.5538127,4.640329,5.243949,4.6856003,3.0181,0.9922004,1.8599042,2.5880208,3.2784111,4.1083884,5.342037,5.87775,5.160951,4.104616,3.270866,2.867195,2.3428001,3.1840954,4.4516973,5.4967146,5.934339,9.7069645,8.892077,5.5797124,2.5616124,3.3425457,4.817642,8.382772,9.42779,8.477088,11.200924,9.050528,8.733627,9.405154,9.7296,7.8734684,5.6891184,3.942393,2.6898816,1.9693103,1.7844516,1.5165952,1.8334957,1.8334957,1.5882751,2.1353056,1.599593,1.750498,2.1013522,2.584248,3.5236318,4.52715,3.8895764,2.7841973,1.9164935,1.5241405,1.3317367,1.0072908,0.7432071,0.5998474,0.5017591,0.392353,0.724344,1.3204187,1.7542707,1.327964,0.5357128,0.4074435,0.48666862,0.45648763,0.1358145,0.041498873,0.00754525,0.011317875,0.026408374,0.0150905,0.0150905,0.16976812,0.32821837,0.38103512,0.26031113,0.331991,0.21503963,0.1961765,0.34330887,0.48666862,0.3169005,0.15467763,0.08677038,0.09808825,0.060362,0.049044125,0.1358145,0.26031113,0.40367088,0.6111652,0.6828451,0.65643674,0.5470306,0.41498876,0.36594462,0.3772625,0.42630664,0.42630664,0.33953625,0.1659955,0.241448,0.23013012,0.1659955,0.090543,0.090543,0.07922512,0.056589376,0.056589376,0.120724,0.29049212,0.32821837,0.271629,0.25276586,0.32821837,0.47157812,0.65643674,0.59230214,0.47157812,0.38103512,0.32067314,0.5281675,0.8903395,1.0072908,0.845068,0.7469798,0.8941121,0.5357128,0.16976812,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.026408374,0.0150905,0.026408374,0.030181,0.030181,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.090543,0.422534,0.663982,0.030181,0.00754525,0.00754525,0.00754525,0.0,0.0,0.011317875,0.060362,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.0754525,0.06413463,0.0,0.0,0.02263575,0.056589376,0.0452715,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.071679875,0.17354076,0.211267,0.19240387,0.23013012,0.27917424,0.21503963,0.13204187,0.06790725,0.030181,0.018863125,0.00754525,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.018863125,0.049044125,0.060362,0.03772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.011317875,0.00754525,0.03772625,0.1056335,0.1659955,0.181086,0.19994913,0.2867195,0.7054809,1.9391292,1.7165444,1.1242423,0.55457586,0.211267,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.011317875,0.033953626,0.06413463,0.120724,0.24522063,0.513077,0.95447415,1.5052774,2.0560806,2.4710693,2.6785638,2.886058,3.2029586,3.953711,5.6778007,5.4438977,6.9227667,9.439108,12.838243,17.486116,25.204908,35.975754,48.127377,57.770206,58.80768,48.58764,39.857784,34.266754,31.79191,30.716713,30.131956,30.331905,30.192318,29.139755,27.159128,25.585943,24.103302,23.201643,23.084692,23.680767,24.95214,26.238607,27.430756,28.487091,29.464201,31.34674,32.88597,33.900806,34.202618,33.62918,35.632442,40.28786,45.18473,48.49332,48.979992,48.79513,47.99156,47.448303,47.938747,50.11178,55.699036,61.316475,65.05892,65.77194,63.048107,62.293583,66.05866,73.241745,80.39464,81.72637,72.21559,62.67839,57.966385,58.634136,60.927895,51.285065,41.2197,34.69683,32.47098,32.105038,32.72752,33.45941,34.5082,35.432495,35.142002,33.60277,31.972998,30.41113,29.185026,28.67195,27.755201,27.23458,26.78941,26.265015,25.680258,25.92548,25.857573,25.66894,25.593489,25.910389,26.348013,26.385738,26.800728,28.158873,30.807257,32.799202,34.64779,36.08516,36.469967,34.83642,32.06354,29.815056,28.007969,26.691322,26.031113,25.129456,24.159891,23.201643,21.967995,19.821371,17.976559,18.157644,18.678267,19.180025,20.643805,20.621168,20.145817,18.964987,17.482344,16.7995,16.248695,16.42601,16.33924,15.762027,15.211224,13.381501,11.623458,9.835234,8.20546,7.2170315,6.741681,6.6662283,6.7152724,6.802043,7.0359454,6.8737226,6.983129,7.043491,6.94163,6.760544,6.319147,5.73439,5.0741806,4.4215164,3.8593953,3.3350005,3.2972744,3.7348988,4.217795,3.874486,3.7914882,3.4557245,3.3312278,3.2029586,2.2107582,2.6634734,2.161714,1.7957695,1.8259505,1.6788181,2.3390274,2.372981,2.0447628,1.750498,2.0296721,2.04099,1.780679,1.3958713,1.056335,0.94692886,0.8978847,0.83752275,0.8526133,0.98465514,1.267602,0.83752275,0.814887,0.97333723,1.2864652,1.9240388,2.5087957,2.9841464,3.1614597,3.0520537,2.867195,1.0940613,1.7316349,1.3204187,0.8111144,0.90920264,2.0485353,2.0447628,2.1654868,1.6939086,0.9016574,1.0601076,0.73566186,0.58475685,0.46026024,0.422534,0.72811663,0.5319401,1.4147344,1.9127209,1.6561824,1.3619176,2.052308,1.3053282,0.51684964,0.24899325,0.23013012,0.90920264,0.814887,0.7394345,1.0601076,1.7014539,0.7884786,1.0487897,1.2940104,1.0487897,0.5357128,0.17354076,0.049044125,0.0150905,0.0,0.003772625,0.003772625,0.090543,0.120724,0.06790725,0.0,0.0,0.094315626,0.5885295,1.2449663,1.2789198,0.36971724,0.0754525,2.5804756,7.322665,10.982111,7.2887115,6.9265394,8.990166,10.902886,8.446907,3.640583,1.2600567,0.3772625,0.20749438,0.094315626,0.030181,0.00754525,0.0,0.0,0.003772625,0.003772625,0.0,0.00754525,0.0150905,0.003772625,0.003772625,0.030181,0.06413463,0.08677038,0.071679875,0.033953626,0.07922512,0.1659955,0.3961256,0.98465514,1.1355602,1.0827434,0.90543,0.73566186,0.754525,1.4449154,1.4449154,1.3694628,1.4147344,1.3392819,0.52062225,0.35462674,0.31312788,0.23390275,0.2867195,0.9205205,1.5656394,1.9466745,1.9881734,1.8184053,1.4713237,1.0487897,0.6187105,0.27540162,0.16976812,0.06413463,0.049044125,0.056589376,0.05281675,0.03772625,0.026408374,0.018863125,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.011317875,0.003772625,0.00754525,0.018863125,0.026408374,0.011317875,0.060362,0.07922512,0.0452715,0.026408374,0.018863125,0.0150905,0.041498873,0.19240387,0.62248313,1.7957695,2.8709676,3.4934506,3.5575855,3.2029586,3.0369632,2.9539654,2.7879698,2.4371157,1.8787673,1.7278622,1.7316349,1.750498,1.7580433,1.8636768,1.991946,1.901403,1.871222,1.8938577,1.6788181,1.5279131,1.4449154,1.5241405,1.8825399,2.6634734,3.31991,3.7763977,3.531177,2.505023,1.0638802,0.965792,1.1393328,1.539231,2.052308,2.4861598,3.2670932,3.8480775,4.1008434,3.9197574,3.2218218,3.1161883,3.62172,3.7198083,3.1463692,2.384299,4.183841,4.1800685,3.1652324,1.9466745,1.3392819,1.7429527,3.470815,4.8025517,6.477597,11.69891,9.484379,8.424272,8.050782,8.028146,8.152642,8.45068,9.469289,8.4544525,5.3873086,3.006782,1.9957186,1.6788181,1.6712729,1.6939086,1.599593,1.3543724,1.4675511,1.720317,2.2899833,3.7575345,5.323174,4.402653,3.2972744,2.7200627,1.780679,1.0902886,1.0148361,1.1996948,1.2789198,0.87147635,0.69039035,1.5316857,2.233394,2.1654868,1.2411937,0.7997965,1.6939086,2.1277604,1.5052774,0.4074435,0.14335975,0.060362,0.041498873,0.026408374,0.003772625,0.003772625,0.06413463,0.14335975,0.181086,0.08677038,0.08299775,0.1056335,0.16976812,0.21881226,0.120724,0.116951376,0.06413463,0.026408374,0.049044125,0.15845025,0.28294688,0.5394854,0.9997456,1.2562841,0.3772625,0.34330887,0.33953625,0.29803738,0.271629,0.42630664,0.47912338,0.5093044,0.5281675,0.513077,0.39989826,0.181086,0.12826926,0.13204187,0.150905,0.18863125,0.090543,0.090543,0.181086,0.35085413,0.5696664,0.5394854,0.39989826,0.34330887,0.3734899,0.32821837,0.2867195,0.2678564,0.26408374,0.29803738,0.44139713,0.45648763,0.3734899,0.26408374,0.17731337,0.150905,0.17731337,0.1056335,0.033953626,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.033953626,0.030181,0.018863125,0.0150905,0.018863125,0.011317875,0.011317875,0.018863125,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08299775,0.25276586,0.35839936,0.1056335,0.018863125,0.0150905,0.02263575,0.011317875,0.0,0.011317875,0.02263575,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.018863125,0.0,0.0,0.003772625,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.0,0.0150905,0.049044125,0.19994913,0.41876137,0.5357128,0.7696155,0.63002837,0.362172,0.13204187,0.018863125,0.00754525,0.0,0.003772625,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.026408374,0.049044125,0.0452715,0.030181,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.0,0.003772625,0.0,0.018863125,0.049044125,0.08299775,0.11317875,0.16976812,0.27540162,0.55457586,1.2298758,1.2751472,0.90543,0.47535074,0.17731337,0.05281675,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.011317875,0.026408374,0.0452715,0.08677038,0.15845025,0.35085413,0.7054809,1.2411937,1.8561316,2.3503454,2.704972,2.9351022,3.169005,3.5349495,4.1612053,4.4403796,5.0439997,6.2889657,8.446907,11.763044,16.822134,23.714722,31.995632,41.20461,50.873848,56.13289,53.899494,47.244583,39.371113,33.621635,30.535627,28.611588,27.211945,26.049976,25.19359,23.36764,21.983086,21.27006,21.273832,21.862362,22.243397,22.696112,23.001694,23.1526,23.337458,24.269297,25.363358,26.366877,27.46471,29.271797,31.54669,34.398796,38.36005,42.408077,43.939762,46.599464,48.76495,50.3985,51.111523,50.17214,52.179176,55.940483,59.464115,61.248566,60.30164,61.237247,65.76817,70.17837,71.7176,68.60519,66.30011,66.88487,71.144165,75.75808,73.31719,57.10245,45.131912,37.386715,33.289642,31.712687,30.256453,29.166164,28.966215,29.716967,31.01475,31.67496,31.554235,31.075111,30.414904,29.501928,28.204145,27.411894,26.90636,26.668686,26.853544,27.498663,28.057013,28.649315,29.252934,29.716967,30.214954,30.422447,30.694077,31.459919,33.21042,34.40257,35.994614,38.41664,40.808483,41.034843,40.736805,39.529564,36.726505,32.64075,28.581408,25.989614,25.238861,23.748674,21.719002,22.126446,20.29295,18.704676,18.429274,19.1008,18.923487,20.36463,21.643549,22.703657,23.126192,22.111355,20.123182,18.94235,17.795471,16.67123,16.346785,16.35433,15.441354,13.8719425,11.966766,10.110635,8.873214,8.235641,7.748972,7.284939,7.0472636,7.0246277,7.164215,7.5301595,7.9941926,8.262049,8.231868,7.786698,6.8963585,5.772116,4.847823,4.4894238,3.9801195,3.6179473,3.610402,4.0706625,4.093298,3.9914372,3.8254418,3.470815,2.625747,2.9615107,2.3654358,1.7995421,1.7882242,2.4220252,2.263575,2.8256962,2.8181508,2.1768045,2.0787163,2.1881225,1.8259505,1.4637785,1.3204187,1.3355093,1.4449154,1.3732355,1.0978339,0.83752275,1.0601076,0.8262049,0.814887,1.1242423,1.6561824,2.1051247,2.535204,2.4974778,2.384299,2.3013012,2.052308,0.65643674,1.5015048,1.3128735,1.2713746,1.5731846,1.4147344,1.1996948,2.5540671,2.9049213,1.9806281,1.841041,1.3807807,1.5316857,2.1315331,2.6446102,2.1579416,1.2789198,1.5052774,1.9730829,2.1994405,2.082489,2.2862108,1.4071891,0.65643674,0.452715,0.422534,0.5394854,0.392353,0.36594462,0.5583485,0.7997965,0.6488915,0.8601585,0.8903395,0.663982,0.5357128,0.38858038,0.24522063,0.12826926,0.049044125,0.026408374,0.033953626,0.21881226,0.29803738,0.211267,0.120724,0.060362,0.69793564,1.1204696,1.0751982,0.965792,1.599593,4.0782075,7.360391,9.544742,7.877241,4.06689,3.3161373,4.6742826,6.3719635,5.847569,2.6898816,1.0978339,0.56212115,0.52439487,0.38480774,0.18485862,0.060362,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.030181,0.041498873,0.05281675,0.06413463,0.0754525,0.12826926,0.17354076,0.1961765,0.29426476,0.69793564,1.0789708,1.2940104,1.4034165,1.4373702,1.3807807,1.7052265,1.7919968,1.8334957,1.8485862,1.6675003,1.3543724,1.3694628,1.4109617,1.5052774,2.0183544,3.3953626,4.195159,4.3800178,4.0517993,3.4670424,2.5276587,1.6033657,0.9620194,0.63002837,0.392353,0.15845025,0.060362,0.030181,0.02263575,0.018863125,0.0150905,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.0150905,0.02263575,0.011317875,0.026408374,0.03772625,0.041498873,0.06790725,0.041498873,0.026408374,0.02263575,0.060362,0.23013012,0.77338815,1.4637785,2.0862615,2.4899325,2.595566,2.7804246,2.969056,2.9426475,2.6219745,2.052308,1.7391801,1.5920477,1.569412,1.6448646,1.780679,1.8523588,1.8033148,1.7995421,1.8674494,1.8938577,1.6976813,1.327964,1.0336993,1.0751982,1.7278622,2.6710186,2.938875,2.8634224,2.6332922,2.282438,2.2484846,1.7882242,1.599593,1.8221779,2.0258996,2.2748928,2.746471,3.3764994,3.9763467,4.2630663,4.715781,5.5382137,5.794752,5.3609,4.8930945,4.168751,3.9650288,4.247976,4.1574326,2.0108092,1.3166461,1.8033148,2.6031113,3.9159849,7.001992,7.726336,8.66572,9.039209,8.710991,8.20546,8.065872,8.179051,7.8244243,6.8359966,5.6363015,3.9574835,3.0105548,2.535204,2.2371666,1.81086,2.214531,2.8294687,3.2784111,3.62172,4.3649273,4.2328854,3.2670932,2.5578396,2.2748928,1.6637276,1.1091517,0.965792,1.1355602,1.3053282,0.94315624,1.4071891,2.5616124,2.8558772,1.9768555,0.845068,0.7394345,1.2411937,1.3807807,0.8941121,0.21503963,0.07922512,0.03772625,0.033953626,0.026408374,0.00754525,0.0,0.018863125,0.049044125,0.06413463,0.03772625,0.041498873,0.08299775,0.124496624,0.11317875,0.02263575,0.041498873,0.041498873,0.1358145,0.45648763,1.116697,1.1355602,0.90920264,0.7469798,0.63002837,0.19994913,0.19240387,0.31312788,0.38480774,0.36594462,0.331991,0.28294688,0.29049212,0.41121614,0.58098423,0.6149379,0.56212115,0.573439,0.543258,0.46026024,0.41498876,0.30935526,0.271629,0.35839936,0.52439487,0.6413463,0.65643674,0.6187105,0.55457586,0.44894236,0.271629,0.211267,0.20372175,0.2565385,0.38103512,0.58475685,0.47912338,0.331991,0.16976812,0.0452715,0.026408374,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.018863125,0.030181,0.030181,0.026408374,0.033953626,0.033953626,0.018863125,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.42630664,1.0751982,1.6675003,0.331991,0.00754525,0.011317875,0.003772625,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.120724,0.23013012,0.14713238,0.14713238,0.2678564,0.34330887,0.49421388,0.46026024,0.3055826,0.11317875,0.02263575,0.011317875,0.003772625,0.00754525,0.0150905,0.00754525,0.0150905,0.011317875,0.00754525,0.00754525,0.018863125,0.018863125,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0150905,0.02263575,0.02263575,0.0452715,0.10186087,0.18863125,0.36594462,0.7432071,1.6410918,1.056335,0.4640329,0.3169005,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.041498873,0.08299775,0.20372175,0.41876137,0.7582976,1.1695137,1.5505489,1.8448136,2.0900342,2.3465726,2.6634734,3.059599,3.610402,4.22534,5.0477724,6.2889657,8.20546,12.189351,18.342503,26.121656,35.236317,45.622353,54.012672,60.154507,62.7463,60.87885,54.03908,46.29388,40.778305,36.300198,32.65584,30.652578,28.81531,27.872154,26.90259,25.736847,24.971004,24.827644,24.60506,24.910643,25.729303,26.381968,26.434784,26.796955,27.90988,29.524563,30.690304,33.116104,35.402313,37.76775,40.182228,42.39676,46.663597,51.156796,55.782032,59.71688,61.39947,61.456062,61.920094,62.297356,62.625576,63.478188,67.35268,70.92912,70.6424,66.06621,59.90174,59.249077,62.003094,66.53779,69.80488,67.33381,57.706074,48.58764,41.744095,37.33767,33.912125,31.124157,29.29066,28.132465,27.69484,28.34373,29.743376,30.59599,30.995888,31.02984,30.780848,30.237589,29.566063,28.943579,28.54368,28.554998,28.464457,28.381458,28.487091,28.634224,28.336185,28.577635,28.788902,29.13221,29.826374,31.169428,32.961426,34.847736,37.78284,41.510193,44.528294,46.40706,47.77275,47.25213,44.588654,40.61608,36.892498,33.78763,30.603535,27.69484,26.457418,24.582424,23.039421,22.239624,21.75673,20.30804,19.855326,20.798481,22.628204,24.178753,23.62795,22.933788,22.209444,20.870161,19.097027,17.840744,17.542706,16.98813,16.233604,15.226315,13.819125,12.559069,11.306557,10.106862,9.06939,8.348819,7.7112455,7.4584794,7.484888,7.7037,8.069645,8.348819,8.190369,7.6093845,6.7341356,5.8098426,5.413717,4.7874613,4.274384,4.06689,4.191386,4.1762958,4.2064767,4.1762958,4.0178456,3.6745367,3.2557755,2.9086938,2.5427492,2.2786655,2.4710693,2.565385,3.108643,3.180323,2.674791,2.3201644,2.3578906,2.161714,1.9240388,1.8033148,1.9089483,1.8297231,1.7542707,1.5241405,1.2110126,1.1242423,1.0601076,1.3619176,1.5618668,1.5882751,1.7580433,2.11267,2.04099,1.931584,1.9051756,1.7919968,0.6149379,1.0072908,0.935611,1.3505998,2.2409391,2.6144292,2.6785638,3.2331395,3.0218725,2.2409391,2.516341,2.293756,2.584248,3.108643,3.2670932,2.1390784,1.7882242,1.9240388,2.071171,2.0183544,1.8448136,1.8146327,1.2185578,0.73566186,0.573439,0.45648763,0.23390275,0.13958712,0.16976812,0.26408374,0.31312788,0.6149379,0.6488915,0.47157812,0.33576363,0.6790725,1.7655885,1.599593,0.9922004,0.42630664,0.0754525,0.049044125,0.19994913,0.46026024,0.7432071,0.91674787,1.0827434,1.5354583,1.3204187,0.76207024,1.4637785,2.584248,6.903904,8.850578,6.8774953,3.470815,1.6184561,1.1883769,1.690136,2.5389767,3.0633714,1.7316349,1.0525624,0.8563859,0.88279426,0.77338815,0.482896,0.25276586,0.10186087,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.041498873,0.049044125,0.071679875,0.1056335,0.20749438,0.2565385,0.29426476,0.3772625,0.5696664,0.77716076,1.0601076,1.4298248,1.7844516,1.9202662,1.9240388,2.0749438,2.1805773,2.1654868,2.0560806,2.3767538,2.41448,2.3314822,2.463524,3.3274553,5.3269467,6.5002327,6.858632,6.360646,4.908185,3.6028569,2.7615614,2.3993895,2.11267,1.0902886,0.59230214,0.29049212,0.271629,0.3734899,0.18863125,0.041498873,0.00754525,0.003772625,0.003772625,0.018863125,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.003772625,0.00754525,0.026408374,0.06790725,0.049044125,0.041498873,0.02263575,0.011317875,0.041498873,0.30181,0.97333723,1.750498,2.3201644,2.3805263,2.5616124,2.7653341,2.757789,2.4823873,2.0636258,1.7580433,1.5467763,1.4901869,1.5882751,1.7769064,1.8221779,1.8070874,1.8485862,1.931584,1.9127209,1.6071383,1.3015556,1.026154,0.86770374,0.9808825,1.750498,2.173032,2.41448,2.5729303,2.674791,2.6408374,2.1277604,1.7957695,1.7919968,1.7467253,1.5656394,2.1692593,2.7238352,3.0746894,3.7575345,4.8327327,6.1606965,6.719045,6.6360474,7.2170315,5.8098426,5.9909286,6.8435416,7.2094865,5.696664,2.837014,1.9655377,1.9429018,2.5314314,4.436607,5.8513412,7.594294,8.601585,8.518587,7.7301087,7.3415284,6.688864,6.4549613,6.719045,6.9680386,6.2851934,4.870459,3.863168,3.5160866,3.1727777,3.62172,3.6707642,3.8858037,4.432834,5.0779533,3.338773,2.3993895,1.9693103,1.8297231,1.8297231,1.5316857,1.2261031,1.1204696,1.1242423,0.8337501,1.5467763,2.5201135,2.5012503,1.4449154,0.5281675,0.7582976,0.8526133,0.694163,0.36594462,0.15467763,0.181086,0.13204187,0.06413463,0.0150905,0.00754525,0.026408374,0.030181,0.018863125,0.0150905,0.030181,0.0452715,0.060362,0.06413463,0.06790725,0.1056335,0.17731337,0.2678564,0.49044126,0.845068,1.2147852,1.0525624,0.66775465,0.29803738,0.1056335,0.1659955,0.17354076,0.32444575,0.48666862,0.543258,0.41876137,0.21881226,0.19240387,0.30181,0.452715,0.48666862,0.59607476,0.6526641,0.6526641,0.6111652,0.55080324,0.49421388,0.43007925,0.41876137,0.46026024,0.47535074,0.5470306,0.59230214,0.55457586,0.43007925,0.26408374,0.28294688,0.41121614,0.6073926,0.70170826,0.4074435,0.30935526,0.241448,0.15467763,0.056589376,0.033953626,0.026408374,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.0754525,0.14335975,0.16976812,0.09808825,0.030181,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.018863125,0.0150905,0.018863125,0.030181,0.041498873,0.049044125,0.0452715,0.03772625,0.018863125,0.003772625,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.38858038,1.267602,2.6710186,0.5357128,0.0,0.0,0.003772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.030181,0.120724,0.23767537,0.20372175,0.181086,0.2867195,0.5772116,0.41498876,0.27540162,0.15845025,0.06413463,0.018863125,0.011317875,0.003772625,0.00754525,0.0150905,0.011317875,0.011317875,0.00754525,0.003772625,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.011317875,0.00754525,0.00754525,0.02263575,0.060362,0.11317875,0.21503963,0.4074435,1.2940104,0.87147635,0.452715,0.38480774,0.041498873,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.003772625,0.00754525,0.003772625,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.026408374,0.08677038,0.1961765,0.362172,0.5772116,0.83752275,1.0374719,1.2638294,1.5165952,1.8259505,2.2447119,2.8181508,3.482133,4.168751,4.90064,5.794752,8.563859,13.551269,20.564579,29.20389,38.839176,47.67089,57.521214,66.511375,72.38535,72.54381,67.48849,60.731716,52.937473,45.652534,41.28761,39.405067,38.394005,37.00568,35.002415,33.134964,32.387985,31.358059,31.226017,32.25217,33.768764,34.43652,35.402313,36.41715,37.164127,37.2509,38.710907,40.272774,41.11784,41.442287,42.449577,45.45636,49.832603,55.450043,61.64469,67.24704,69.92183,70.66504,70.01992,69.333305,70.770676,75.271416,76.04858,71.823235,64.4553,58.93972,58.55114,59.70179,60.98448,61.15048,59.132126,56.55542,51.760414,46.976727,42.74007,37.888474,34.22148,31.71646,29.95087,28.770039,28.302233,29.196344,30.116865,30.920435,31.554235,32.01827,32.184265,32.172947,31.923952,31.47501,30.954388,30.305496,29.773556,29.422703,29.090712,28.404093,28.290915,28.151327,27.98156,27.947605,28.377686,29.988596,31.64478,34.10453,37.514984,41.41588,45.18473,48.681953,51.03607,51.832096,51.103977,49.632656,46.65605,43.07206,39.480522,36.1757,33.31605,31.625916,30.509218,29.332159,27.404348,26.068838,25.397312,25.355812,25.472763,24.831417,25.118137,25.370903,25.084183,23.918442,21.734093,20.353312,19.210207,18.444365,17.927513,17.229578,16.044973,14.618922,13.102326,11.747954,10.899114,9.737145,8.797762,8.065872,7.6395655,7.745199,8.111144,8.096053,7.8017883,7.2585306,6.4511886,5.926794,5.3194013,4.908185,4.7044635,4.4441524,4.3913355,4.4215164,4.436607,4.38379,4.255521,3.7084904,3.6028569,3.451952,3.1765501,3.0935526,3.097325,3.3538637,3.4783602,3.3236825,2.9766011,2.8558772,2.7728794,2.5691576,2.354118,2.5012503,2.2899833,2.2560298,2.2711203,2.1541688,1.6675003,1.6561824,1.9881734,2.0673985,1.9278114,2.252257,2.463524,2.2598023,2.0485353,2.1692593,2.9124665,1.6033657,0.98465514,0.633801,0.8978847,1.9504471,3.7763977,4.538468,3.3840446,2.0900342,1.7127718,2.5729303,2.7917426,2.7841973,2.5238862,2.0258996,1.3392819,1.8749946,1.8787673,1.4034165,0.84129536,0.9016574,1.1091517,0.97710985,0.724344,0.49044126,0.32821837,0.1961765,0.124496624,0.1056335,0.120724,0.14335975,0.543258,0.6073926,0.41876137,0.29426476,0.7922512,2.9615107,2.927557,2.0145817,1.0601076,0.41121614,0.13958712,0.2678564,0.94692886,1.7769064,1.8297231,2.2447119,2.071171,1.4034165,1.1129243,2.867195,3.2821836,6.8925858,6.2399216,1.4750963,0.33576363,1.026154,0.8601585,0.62248313,0.73188925,1.237421,1.0223814,0.9393836,0.9695646,1.056335,1.0902886,0.8903395,0.66020936,0.4074435,0.17354076,0.0452715,0.011317875,0.0,0.0,0.0,0.003772625,0.030181,0.03772625,0.060362,0.10186087,0.13958712,0.22258487,0.2565385,0.41498876,0.6488915,0.68661773,0.47157812,0.5394854,0.9016574,1.4298248,1.8599042,1.8599042,2.1805773,2.5691576,2.8822856,3.0935526,3.3576362,3.1010978,2.8936033,3.097325,3.8556228,5.583485,7.0963078,8.14887,8.00551,5.413717,4.3724723,4.4743333,4.67051,4.074435,1.961765,1.3845534,0.84129536,0.68661773,0.7582976,0.38103512,0.12826926,0.033953626,0.00754525,0.00754525,0.03772625,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.03772625,0.041498873,0.030181,0.018863125,0.030181,0.38858038,1.4637785,2.6823363,3.410453,2.9728284,2.637065,2.5389767,2.4031622,2.1466236,1.8976303,1.7165444,1.5807298,1.5543215,1.659955,1.8599042,1.9391292,1.8976303,1.9089483,1.9579924,1.8221779,1.5015048,1.2487389,1.0374719,0.8186596,0.55080324,0.6828451,1.3656902,1.9089483,2.052308,1.9806281,1.6939086,1.6109109,1.5731846,1.4373702,1.0902886,0.7922512,1.8221779,2.1994405,1.7165444,1.9127209,3.1237335,4.4931965,5.2062225,5.4740787,6.549277,6.156924,7.062354,7.9225125,8.469543,9.507015,5.7381625,3.380272,2.4295704,3.006782,5.3873086,4.7610526,5.3269467,6.319147,7.183078,7.5603404,7.0812173,6.749226,6.398372,6.255012,6.9567204,7.647111,6.2021956,5.0968165,5.089271,5.2288585,5.4174895,3.8443048,3.2444575,4.3385186,5.8437963,3.591539,2.6898816,2.1994405,1.8976303,2.2711203,2.0108092,1.6410918,1.3015556,1.0186088,0.66775465,1.0601076,1.5618668,1.5807298,1.1204696,0.76207024,1.1204696,1.0978339,0.80356914,0.44139713,0.2867195,0.36594462,0.27540162,0.124496624,0.00754525,0.003772625,0.049044125,0.049044125,0.026408374,0.011317875,0.033953626,0.030181,0.030181,0.0754525,0.19240387,0.38103512,0.47535074,0.5696664,0.73566186,0.7997965,0.34330887,0.11317875,0.041498873,0.08299775,0.18485862,0.26031113,0.27540162,0.331991,0.46026024,0.59230214,0.56589377,0.3169005,0.28294688,0.28294688,0.23390275,0.150905,0.271629,0.32821837,0.422534,0.5281675,0.5017591,0.47535074,0.4074435,0.3169005,0.24899325,0.24899325,0.31312788,0.33953625,0.3470815,0.35839936,0.36971724,0.45648763,0.7696155,1.026154,0.8941121,0.02263575,0.003772625,0.0150905,0.030181,0.030181,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0452715,0.15467763,0.28294688,0.34330887,0.1961765,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.018863125,0.033953626,0.03772625,0.033953626,0.02263575,0.030181,0.041498873,0.056589376,0.06413463,0.041498873,0.02263575,0.00754525,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09808825,0.6149379,2.1013522,0.41876137,0.0,0.0,0.011317875,0.049044125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.12826926,0.23013012,0.41498876,0.9507015,0.55080324,0.21881226,0.049044125,0.02263575,0.0,0.0,0.011317875,0.0452715,0.07922512,0.05281675,0.0150905,0.0150905,0.011317875,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.00754525,0.003772625,0.011317875,0.033953626,0.049044125,0.08299775,0.1358145,0.20372175,0.26031113,0.362172,0.42630664,0.36594462,0.10186087,0.041498873,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.011317875,0.0150905,0.018863125,0.011317875,0.003772625,0.0,0.00754525,0.0150905,0.011317875,0.003772625,0.011317875,0.00754525,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.0754525,0.16222288,0.29049212,0.47157812,0.6187105,0.79602385,0.995973,1.2525115,1.6373192,2.093807,2.6483827,3.2746384,3.8820312,4.3121104,5.4212623,7.8998766,12.419481,19.217752,28.075874,37.71116,46.158066,54.846424,64.296844,74.13586,78.02543,74.85642,67.49226,59.162304,53.43546,50.93421,48.96113,47.025772,44.965916,42.909836,41.69128,40.15959,39.212666,39.389977,40.906574,42.819294,45.309227,46.561737,46.373108,46.15052,45.96189,46.391968,46.444786,45.7129,44.373615,44.33966,46.425922,50.587128,56.7516,64.84388,72.31745,76.71633,78.693184,79.60616,81.50379,83.98995,80.994484,74.290535,67.050865,63.847904,63.65173,62.787796,61.16557,58.79636,55.797123,55.453815,53.658047,50.88894,47.21063,42.28358,38.2846,35.089184,32.844475,31.358059,30.094229,29.898052,30.120638,30.746893,31.622143,32.455894,33.044422,33.75745,34.20639,34.134712,33.433002,32.931244,32.501163,32.07863,31.629688,31.165655,30.716713,30.192318,29.36234,28.35505,27.675978,28.060785,28.913399,30.25268,32.116356,34.56479,39.039124,43.079605,46.90882,50.492813,53.522232,56.26493,56.446014,54.687973,51.74155,48.512184,44.716923,42.377895,41.00466,39.99737,38.642998,38.450596,36.583145,33.915897,31.320333,29.671696,29.27557,29.667923,30.392267,30.384722,27.966469,26.197107,24.506971,22.89606,21.553007,20.82489,19.47429,17.938831,16.335466,14.950912,14.237886,12.913695,11.400873,9.955957,9.012801,9.159933,8.695901,8.265821,7.8923316,7.4697976,6.7643166,6.119198,5.4967146,5.1647234,5.040227,4.719554,4.6856003,4.689373,4.6554193,4.52715,4.2706113,4.1989317,4.1612053,4.1083884,4.093298,4.2706113,3.7877154,3.7650797,3.9725742,4.164978,4.0706625,3.8141239,3.7047176,3.4179983,3.0558262,3.1048703,2.9803739,2.9539654,3.108643,3.1916409,2.6219745,2.6106565,2.6295197,2.5917933,2.6710186,3.2972744,3.3840446,2.9426475,2.595566,2.9841464,4.798779,3.0822346,1.3015556,0.48666862,0.32444575,0.5319401,0.8865669,2.886058,2.8030603,2.2447119,1.8297231,1.1431054,2.4371157,1.9278114,1.5316857,2.1202152,3.5236318,2.0975795,1.1996948,0.784706,0.7582976,0.97710985,0.7922512,0.76584285,0.55080324,0.241448,0.35085413,0.32821837,0.24899325,0.181086,0.15467763,0.1659955,0.362172,0.56589377,0.40367088,0.0,0.0,0.29426476,0.8978847,1.3619176,1.5354583,1.5731846,0.5583485,1.1016065,2.4823873,3.2331395,1.1581959,0.97710985,1.4977322,2.1088974,2.595566,3.1576872,4.7950063,5.855114,4.5761943,1.690136,0.3961256,0.63002837,0.45648763,0.36594462,0.5319401,0.8224323,0.8224323,0.7432071,0.77716076,0.965792,1.1732863,1.3468271,1.3317367,1.0638802,0.6073926,0.1659955,0.0452715,0.00754525,0.0,0.003772625,0.0150905,0.05281675,0.071679875,0.13204187,0.18863125,0.090543,0.150905,0.1659955,0.5017591,0.9922004,0.9318384,0.44139713,0.19240387,0.24899325,0.5281675,0.80734175,1.0638802,1.961765,3.2369123,4.447925,4.9760923,4.191386,3.5953116,3.9801195,5.0175915,5.247721,5.2854476,6.5228686,8.424272,9.246704,6.013564,5.6325293,6.7379084,6.5228686,4.429062,2.1202152,2.305074,1.6712729,0.7507524,0.041498873,0.0150905,0.211267,0.11317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.018863125,0.030181,0.29803738,1.20724,2.4597516,3.4972234,3.5085413,2.8521044,2.4823873,2.214531,1.9466745,1.6788181,1.5580941,1.5731846,1.7165444,1.871222,1.7844516,1.7957695,1.8561316,1.8485862,1.750498,1.6033657,1.7957695,1.478869,0.9507015,0.5017591,0.44139713,0.6488915,0.84884065,1.0751982,1.3468271,1.6637276,1.5882751,1.5543215,1.4864142,1.358145,1.1732863,0.62625575,0.8262049,1.1393328,1.2902378,1.388326,1.2411937,1.297783,2.6597006,4.3875628,3.5085413,3.169005,3.029418,3.399135,4.6742826,7.3075747,9.616421,6.300284,4.172523,4.9459114,5.2628117,4.191386,3.9386206,5.1232247,7.4396167,9.673011,6.096562,5.240176,6.092789,7.515069,8.224322,6.5040054,5.8702044,5.66271,5.775889,6.6662283,7.816879,5.198677,3.6368105,4.719554,6.820906,4.8440504,4.0103,3.169005,2.2598023,2.3201644,1.7089992,1.5203679,1.3958713,1.1204696,0.59607476,0.8526133,1.2826926,1.6222287,1.8372684,2.1051247,1.9353566,1.297783,0.7432071,0.43385187,0.150905,0.150905,0.150905,0.10940613,0.041498873,0.0150905,0.003772625,0.018863125,0.030181,0.033953626,0.0452715,0.033953626,0.06790725,0.29426476,0.663982,0.9318384,0.77338815,0.422534,0.12826926,0.0,0.0,0.03772625,0.06413463,0.15467763,0.29426476,0.38103512,0.51684964,0.48666862,0.362172,0.23767537,0.21503963,0.23767537,0.30935526,0.30935526,0.23767537,0.21503963,0.3734899,0.47535074,0.52439487,0.48666862,0.3055826,0.1358145,0.06413463,0.13204187,0.27540162,0.33576363,0.31312788,0.241448,0.26408374,0.44139713,0.7469798,0.784706,1.0223814,0.77716076,0.14713238,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.026408374,0.011317875,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.041498873,0.06413463,0.071679875,0.056589376,0.0452715,0.033953626,0.041498873,0.0452715,0.041498873,0.030181,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.0,0.06413463,0.211267,0.32067314,0.1358145,0.05281675,0.030181,0.018863125,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.071679875,0.120724,0.1659955,0.15467763,0.26408374,0.43385187,0.5017591,0.19994913,0.10186087,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.041498873,0.03772625,0.02263575,0.0150905,0.0150905,0.003772625,0.00754525,0.00754525,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026408374,0.0754525,0.14335975,0.23013012,0.31312788,0.4640329,0.66020936,0.90543,1.237421,1.6637276,2.3465726,3.1576872,3.9084394,4.349837,4.4818783,4.817642,5.8400235,8.175279,12.619431,19.885506,27.468483,34.65156,41.370605,48.21792,55.61604,62.01441,65.19473,64.73824,62.040817,57.498577,53.782543,50.956844,48.89322,47.2559,46.573055,46.03357,45.33941,44.42266,43.456867,44.030308,46.55419,49.821285,52.35272,52.41308,51.75287,51.560467,52.073544,52.41685,50.598446,49.61002,49.545883,51.730232,56.861004,65.00233,71.75156,77.742485,84.00127,90.49018,96.13026,96.87347,90.99949,82.02064,73.21156,67.59789,65.92285,65.16833,63.602684,60.34691,55.34441,54.563477,52.115044,49.88542,48.082108,45.21114,41.87991,38.820312,35.749393,32.889744,30.95816,30.177227,29.61888,29.524563,30.015005,31.052477,32.478527,32.92747,33.48582,34.296932,34.591198,34.67797,34.13094,33.451866,32.89729,32.47098,31.701368,31.64478,31.633461,31.38824,31.022295,30.837437,31.248653,32.06354,32.976517,33.599,35.809757,38.477,41.10275,43.51346,45.867577,49.07808,51.51142,53.209103,54.21262,54.563477,52.74507,50.681446,48.89322,47.908566,48.26319,48.90831,48.878128,47.750114,45.51672,42.585392,40.17091,38.431732,37.216946,36.096478,34.36107,34.5082,34.73833,32.82561,29.151073,26.672459,24.903097,22.062311,19.70442,18.350048,17.471025,16.0412,14.777372,13.392818,12.67602,14.494425,10.993429,9.061845,8.152642,7.677292,7.020855,6.349328,5.5570765,5.1232247,5.0025005,4.6252384,4.587512,4.749735,4.8742313,4.8327327,4.6252384,4.3196554,4.22534,4.255521,4.3913355,4.6856003,4.659192,4.636556,4.825187,5.1835866,5.402399,5.194905,5.0515447,4.708236,4.2027044,3.8593953,3.983892,3.7386713,3.4255435,3.3161373,3.6481283,3.7801702,3.6028569,3.2746384,2.9803739,2.9464202,3.2255943,3.0030096,3.059599,3.821669,5.372218,2.6446102,1.0638802,0.4678055,0.513077,0.7922512,0.8224323,1.0299267,0.9280658,1.1506506,2.2409391,4.6214657,6.1229706,5.1081343,5.2854476,6.9189944,6.820906,5.070408,3.0746894,1.6448646,0.9695646,0.62248313,0.48666862,0.4074435,0.573439,0.90543,1.0336993,0.3961256,0.211267,0.18485862,0.16222288,0.14335975,0.181086,0.5394854,0.46026024,0.033953626,0.16976812,0.38480774,0.49421388,0.63002837,0.7922512,0.8262049,0.48666862,1.0148361,1.4675511,1.3807807,0.7696155,1.7089992,1.539231,1.5958204,2.8596497,5.9418845,4.666737,3.1237335,1.6788181,0.6073926,0.116951376,0.13204187,0.150905,0.1659955,0.241448,0.49421388,0.33953625,0.32821837,0.47912338,0.73566186,0.94315624,1.1544232,1.3694628,1.4373702,1.2525115,0.76584285,0.35085413,0.14335975,0.049044125,0.0150905,0.026408374,0.241448,0.19994913,0.13204187,0.13958712,0.18863125,0.32821837,0.43007925,0.573439,0.7054809,0.6149379,0.5357128,0.43007925,0.35839936,0.47157812,1.0148361,1.6033657,1.9127209,2.5238862,3.572676,4.7421894,4.8402777,4.878004,5.0741806,5.462761,5.907931,6.990674,8.224322,8.963757,8.726082,7.17176,6.0512905,5.704209,5.353355,4.5422406,3.1237335,2.4371157,1.5430037,0.76207024,0.32444575,0.36971724,0.33953625,0.22258487,0.090543,0.003772625,0.02263575,0.033953626,0.03772625,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.003772625,0.003772625,0.00754525,0.116951376,0.49044126,0.965792,1.3845534,1.5807298,1.6071383,1.599593,1.5807298,1.5656394,1.5807298,1.5580941,1.5580941,1.6260014,1.7089992,1.6524098,1.3128735,1.2902378,1.5505489,1.841041,1.6750455,1.901403,1.5769572,1.1581959,1.0035182,1.3807807,0.97333723,1.026154,1.5731846,2.1202152,1.6260014,1.6222287,1.2638294,0.95447415,0.80734175,0.663982,0.4640329,1.1355602,1.6939086,1.8976303,2.2183034,1.6222287,1.1695137,1.7240896,2.5880208,1.4826416,2.0108092,1.81086,1.8146327,2.5427492,4.085753,5.4174895,6.1342883,5.6061206,4.425289,4.4215164,3.9725742,4.429062,6.1720147,8.130007,7.756517,9.307066,7.5490227,6.25124,6.387054,6.149379,6.6058664,6.620957,6.300284,6.2323766,7.4735703,8.541223,7.1302614,5.3646727,4.4441524,4.659192,3.229367,2.6446102,2.2107582,1.7354075,1.5128226,1.50905,1.6976813,1.5128226,0.9620194,0.63002837,0.55457586,0.8224323,1.0525624,1.116697,1.1431054,0.9507015,0.84129536,0.70170826,0.46026024,0.090543,0.041498873,0.030181,0.05281675,0.094315626,0.150905,0.08677038,0.056589376,0.03772625,0.03772625,0.056589376,0.23013012,0.392353,0.5357128,0.6149379,0.55080324,0.2678564,0.10940613,0.049044125,0.06413463,0.18485862,0.3169005,0.36971724,0.36971724,0.36594462,0.43007925,0.5357128,0.44516975,0.27540162,0.13204187,0.116951376,0.13958712,0.23390275,0.29049212,0.32067314,0.43385187,0.4640329,0.392353,0.27917424,0.16976812,0.08677038,0.120724,0.29803738,0.4376245,0.43007925,0.23767537,0.28294688,0.36971724,0.5583485,0.7469798,0.6488915,0.32444575,0.23767537,0.15467763,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.041498873,0.071679875,0.08677038,0.094315626,0.13204187,0.15845025,0.07922512,0.0150905,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.026408374,0.056589376,0.06413463,0.026408374,0.011317875,0.00754525,0.00754525,0.0150905,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.060362,0.090543,0.13204187,0.15845025,0.23767537,0.38858038,0.5394854,0.5281675,0.3734899,0.22258487,0.1056335,0.030181,0.011317875,0.003772625,0.0,0.0150905,0.049044125,0.090543,0.08299775,0.06413463,0.0452715,0.026408374,0.0150905,0.011317875,0.0150905,0.0150905,0.011317875,0.0150905,0.026408374,0.033953626,0.03772625,0.030181,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.060362,0.120724,0.21503963,0.331991,0.49421388,0.67152727,0.8639311,1.1242423,1.388326,1.7882242,2.282438,2.7804246,3.1539145,3.4142256,3.731126,4.285702,5.3609,7.333983,11.559323,17.04472,22.39053,26.970495,30.909117,35.326862,40.00869,44.184982,47.68221,50.911575,53.876858,56.41206,56.20834,53.548637,51.3077,50.451313,51.06248,52.13013,52.526257,51.024754,48.930946,47.968925,49.225212,52.281036,55.235004,57.483486,59.060444,60.27523,60.720398,59.25285,59.00763,57.962612,57.766434,59.709335,64.74579,69.61248,73.63787,78.66678,85.084015,91.79551,95.08901,93.71955,89.788475,83.86168,74.9432,69.35594,64.88161,60.92035,57.513668,55.33309,52.74507,49.406296,46.599464,44.879147,44.05294,43.132423,41.49133,39.07685,36.183247,33.41414,31.441057,29.679241,28.5135,28.24187,29.07562,30.562035,31.829638,32.942562,33.761223,33.957397,33.768764,33.440548,33.255688,33.146282,32.67848,31.742867,31.207153,30.920435,31.007204,31.86359,30.909117,30.445084,30.897799,32.025814,32.942562,34.847736,37.548935,40.51422,43.479504,46.441013,48.440506,50.40227,51.7076,52.465897,53.50337,54.446526,54.38239,52.74507,50.119324,48.225464,45.769485,45.810986,47.633163,50.251366,52.450806,52.835613,51.583103,49.100716,46.131657,43.77377,40.865074,39.869102,39.635197,38.982533,36.669914,34.26298,31.176973,28.366367,25.619896,21.537916,20.975796,19.01403,16.935314,15.569623,15.290449,12.381755,11.808316,10.359629,7.8432875,7.115171,7.4396167,7.360391,6.670001,5.6325293,5.0025005,4.7308717,4.938366,5.3948536,5.6513925,5.062863,4.727099,4.5460134,4.644101,4.8855495,4.8553686,4.9760923,5.1081343,5.3684454,5.7796617,6.2436943,6.436098,6.145606,5.5004873,4.821415,4.606375,4.1989317,3.9914372,3.9650288,4.0593443,4.183841,4.2404304,4.1008434,3.8707132,3.5462675,3.029418,2.7540162,2.5616124,3.229367,4.5196047,5.1647234,4.22534,2.8332415,1.4750963,1.1053791,1.5203679,1.3392819,2.4710693,2.505023,2.3088465,2.4899325,3.4066803,5.2137675,4.085753,3.3161373,3.8895764,4.5120597,5.2099953,3.863168,2.4295704,1.6788181,1.1846043,0.5696664,0.331991,0.4678055,0.87147635,1.3430545,0.66020936,0.32444575,0.181086,0.120724,0.08299775,0.060362,0.41498876,0.58475685,0.56212115,0.90920264,0.7394345,0.41121614,1.4977322,3.2935016,2.8106055,1.8787673,2.0787163,1.7882242,0.8299775,0.4979865,2.727608,4.52715,5.0025005,4.349837,3.8254418,2.3314822,1.1129243,0.39989826,0.14335975,0.026408374,0.011317875,0.03772625,0.14335975,0.24899325,0.1659955,0.10940613,0.28294688,0.44139713,0.47535074,0.392353,0.6187105,0.87147635,1.086516,1.2185578,1.2449663,0.9620194,0.58098423,0.38103512,0.32067314,0.041498873,0.150905,0.1056335,0.05281675,0.06413463,0.13958712,0.32067314,0.4979865,0.55457586,0.49044126,0.41498876,0.482896,0.47157812,0.58475685,0.9620194,1.6825907,2.0070364,2.203213,2.5578396,3.1954134,4.0706625,4.285702,3.821669,3.3350005,3.2142766,3.572676,4.5724216,5.462761,6.115425,6.428553,6.3153744,5.27413,4.0895257,3.6858547,3.8707132,3.361409,2.474842,2.1503963,1.9693103,1.5580941,0.59607476,0.3470815,0.29049212,0.24899325,0.16222288,0.0754525,0.030181,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0452715,0.241448,0.5998474,1.1280149,1.8485862,1.9278114,1.6260014,1.327964,1.2298758,1.3468271,1.4637785,1.5203679,1.569412,1.6109109,1.599593,1.3619176,1.3166461,1.388326,1.4750963,1.4750963,1.9127209,1.931584,1.5203679,0.9808825,0.95824677,0.7130261,0.6526641,1.0110635,1.7052265,2.3390274,1.5467763,1.1355602,0.9016574,0.7205714,0.5357128,0.41498876,0.8563859,1.2789198,1.4637785,1.5656394,1.4637785,1.1808317,1.4449154,2.003264,1.599593,2.293756,1.9051756,1.50905,1.6222287,2.1805773,3.482133,4.485651,4.6742826,4.0291634,3.048281,2.8521044,3.9688015,5.6476197,7.413208,9.0543,10.193633,9.948412,8.314865,6.3531003,6.1606965,7.6018395,8.650629,8.518587,7.4396167,6.677546,7.213259,6.0814714,4.878004,4.4177437,4.7233267,3.2482302,2.4333432,2.1843498,2.1202152,1.5882751,1.8863125,1.7919968,1.5656394,1.327964,1.0525624,0.7922512,0.8224323,0.965792,0.98842776,0.6149379,0.60362,0.5583485,0.4678055,0.331991,0.1659955,0.3055826,0.35085413,0.3055826,0.26408374,0.41121614,0.38858038,0.49044126,0.7469798,0.995973,0.86770374,0.95447415,0.9280658,0.7432071,0.452715,0.211267,0.15845025,0.18863125,0.241448,0.35462674,0.66775465,0.694163,0.5394854,0.452715,0.4678055,0.4074435,0.3772625,0.35462674,0.28294688,0.21881226,0.29426476,0.44894236,0.47157812,0.392353,0.30181,0.331991,0.45648763,0.3734899,0.19994913,0.116951376,0.3772625,0.48666862,0.47535074,0.46026024,0.42630664,0.22258487,0.7809334,0.97710985,0.84129536,0.52439487,0.2867195,0.09808825,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0150905,0.05281675,0.071679875,0.08299775,0.124496624,0.15467763,0.090543,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.033953626,0.06790725,0.1056335,0.1056335,0.13958712,0.2867195,0.51684964,0.7092535,0.56212115,0.3961256,0.2263575,0.090543,0.041498873,0.0754525,0.08299775,0.124496624,0.19240387,0.2263575,0.14713238,0.08299775,0.0452715,0.041498873,0.041498873,0.026408374,0.018863125,0.0150905,0.018863125,0.02263575,0.05281675,0.094315626,0.1358145,0.15467763,0.1056335,0.049044125,0.0150905,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.05281675,0.1056335,0.1961765,0.3169005,0.4979865,0.69793564,0.90543,1.1355602,1.3392819,1.599593,1.9164935,2.2748928,2.6521554,3.127506,3.6330378,4.1762958,4.8327327,5.764571,8.050782,11.710228,15.973294,20.036411,23.054512,25.589716,28.807764,32.459667,36.194565,39.555973,43.23051,48.08965,52.760162,56.62333,59.811195,60.644947,61.459835,62.45958,63.18015,62.512398,58.10597,53.201557,49.89674,49.130894,50.666355,53.26192,56.921368,60.04133,61.463608,60.475178,60.46386,59.811195,59.426388,60.475178,64.3723,69.740746,73.01161,75.4525,78.01788,81.37552,83.276924,83.24674,81.86219,79.1044,74.35467,70.02369,65.83985,61.946503,58.63791,56.355473,53.929676,51.100204,48.353733,46.32029,45.731762,44.965916,44.373615,43.170147,40.849983,37.175446,34.040394,31.31656,29.230299,27.932516,27.491117,28.128693,28.977533,29.992369,30.969479,31.5731,32.055996,32.188038,32.097492,31.939043,31.878681,31.27506,31.192064,31.139246,31.12793,31.633461,31.161882,30.51299,30.10932,30.260225,31.154337,32.289898,34.34975,37.19431,40.43122,43.400276,45.19982,47.176674,49.149757,50.956844,52.450806,54.6427,56.81573,57.411808,56.189476,54.2428,50.881393,48.191513,47.19931,47.436985,46.96918,48.538593,50.30418,51.560467,52.39044,53.66182,50.798397,48.34996,46.56551,45.207367,43.543636,41.442287,40.15959,38.40155,35.590942,31.882454,30.067822,26.457418,22.756474,19.908142,18.104828,15.845025,15.294222,13.528633,10.582213,9.4127,9.224068,8.6581745,7.541477,6.1795597,5.342037,5.8211603,6.217286,6.089017,5.564622,5.3571277,5.915476,5.670255,5.696664,6.0324273,5.704209,5.5683947,5.5306683,5.6853456,6.0512905,6.5832305,7.5037513,7.6282477,7.043491,5.9607477,4.7006907,4.402653,4.353609,4.38379,4.4705606,4.749735,4.719554,4.666737,4.52715,4.191386,3.5274043,3.0746894,2.8219235,3.3576362,4.2781568,4.1498876,5.4665337,4.5497856,3.059599,2.4220252,2.6031113,2.1202152,3.127506,3.1954134,2.8445592,2.5314314,2.6408374,3.4783602,2.848332,2.191895,2.071171,2.1768045,3.9159849,3.7047176,3.4066803,3.5047686,3.1124156,1.3770081,1.2261031,2.003264,2.6823363,1.8749946,1.1695137,0.56212115,0.20749438,0.094315626,0.05281675,0.17731337,0.80356914,1.2223305,1.1921495,0.9393836,0.7394345,0.5281675,2.233394,4.738417,3.874486,3.350091,3.6292653,2.9916916,1.5882751,1.4600059,3.2105038,4.9044123,5.028909,3.4444065,1.4034165,0.5470306,0.16222288,0.049044125,0.056589376,0.071679875,0.02263575,0.03772625,0.17731337,0.2867195,0.00754525,0.02263575,0.19240387,0.28294688,0.21503963,0.056589376,0.22258487,0.36971724,0.55457586,0.8186596,1.1846043,1.1732863,0.8563859,0.62248313,0.5017591,0.150905,0.09808825,0.060362,0.0452715,0.06790725,0.13958712,0.27540162,0.3772625,0.3961256,0.38480774,0.47535074,0.58475685,0.6073926,0.84129536,1.3317367,1.8749946,1.901403,2.1164427,2.3880715,2.6295197,2.8256962,2.6936543,2.0372176,1.50905,1.4034165,1.6335466,2.123988,2.546522,3.0218725,3.4972234,3.772625,3.1237335,2.1579416,1.8976303,2.305074,2.263575,1.8334957,2.1315331,2.2899833,1.8184053,0.62625575,0.52439487,0.47157812,0.3772625,0.2263575,0.08677038,0.0754525,0.05281675,0.02263575,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.1358145,0.4640329,1.0487897,1.8938577,1.9994912,1.6373192,1.20724,0.965792,1.0223814,1.2336484,1.3920987,1.4864142,1.5203679,1.5430037,1.4600059,1.3430545,1.1846043,1.0676528,1.1619685,1.5769572,1.7429527,1.478869,0.935611,0.62248313,0.452715,0.35462674,0.47912338,0.9620194,1.9240388,1.0827434,1.1355602,1.1317875,0.7884786,0.47912338,0.4640329,0.58098423,0.73566186,0.87902164,1.0110635,1.2864652,1.2261031,1.2751472,1.5128226,1.6524098,2.04099,1.8825399,1.5958204,1.4222796,1.418507,2.3013012,2.9313297,3.4972234,3.5802212,2.1315331,2.0372176,2.8521044,3.8782585,5.247721,7.914967,8.990166,9.6051035,8.326183,6.013564,5.8437963,6.9680386,8.246958,8.763808,8.096053,6.304056,5.8702044,4.67051,4.036709,4.2706113,4.6516466,3.3953626,2.5804756,2.5201135,2.7502437,2.052308,2.0372176,1.9353566,1.9429018,2.04099,1.961765,1.4034165,1.6675003,1.6410918,1.0789708,0.56589377,0.6375736,0.573439,0.52439487,0.55080324,0.63002837,1.0336993,0.935611,0.7130261,0.6149379,0.7582976,0.77338815,0.84884065,1.0676528,1.2940104,1.1846043,1.2185578,0.965792,0.6073926,0.29049212,0.11317875,0.23390275,0.28294688,0.36971724,0.58098423,0.97333723,0.69793564,0.44516975,0.3772625,0.43385187,0.32821837,0.24899325,0.31312788,0.331991,0.30181,0.3734899,0.5583485,0.56212115,0.4640329,0.35839936,0.35839936,0.55080324,0.44516975,0.21503963,0.1358145,0.56212115,0.8337501,0.72811663,0.52062225,0.35462674,0.25276586,0.754525,0.8601585,0.60362,0.1961765,0.03772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.03772625,0.049044125,0.071679875,0.08299775,0.056589376,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.026408374,0.018863125,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0452715,0.23013012,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.041498873,0.06790725,0.06413463,0.06790725,0.15467763,0.3470815,0.6187105,0.62248313,0.5055317,0.36594462,0.241448,0.12826926,0.181086,0.23390275,0.28294688,0.32444575,0.35839936,0.26408374,0.22258487,0.241448,0.24899325,0.1056335,0.0452715,0.02263575,0.018863125,0.02263575,0.02263575,0.056589376,0.11317875,0.16976812,0.20749438,0.19240387,0.12826926,0.0754525,0.033953626,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.03772625,0.07922512,0.13958712,0.24899325,0.43007925,0.65643674,0.9016574,1.1581959,1.4034165,1.659955,1.9353566,2.2484846,2.6144292,3.2444575,4.014073,4.749735,5.349582,5.772116,6.7831798,8.963757,12.261031,16.109108,19.429018,21.768045,24.261751,27.132719,30.256453,33.191555,36.243607,40.389725,46.214657,53.537323,61.418335,65.56822,67.21309,67.39795,67.133865,67.40926,64.94951,60.973164,55.90653,51.349197,50.096687,50.096687,53.29587,57.562714,61.25234,63.202785,66.20957,66.982956,66.24352,65.496544,67.01314,72.513626,75.59963,76.18816,75.28651,74.96583,74.275444,72.00055,69.1409,66.77169,66.0398,64.50057,62.919838,61.101433,59.011402,56.785553,55.997074,54.77097,53.111015,51.43597,50.56449,48.84795,47.75766,46.486286,44.25289,40.318043,36.858547,34.093212,31.641006,29.437794,27.751429,27.41944,27.615616,28.260735,28.95867,29.011486,29.713194,30.25268,30.29795,30.015005,30.071594,29.988596,30.373404,30.792166,31.143019,31.641006,31.27506,30.637487,29.781101,29.090712,29.283115,29.441565,30.573353,32.62566,35.191048,37.51121,39.3183,41.770504,45.086643,48.666862,51.066254,52.763935,55.29159,57.438217,58.573776,58.63791,56.63842,53.718407,51.183205,48.99131,45.76194,45.120594,45.51672,47.03709,49.45534,52.20936,51.813232,51.330338,50.613537,49.749607,49.03658,47.08236,46.25993,45.26018,43.58891,41.544147,39.25416,35.606033,31.76173,28.328642,25.333178,23.450638,20.734346,17.335213,14.0907545,12.536433,11.732863,10.872705,9.529651,7.9753294,7.1566696,7.0963078,7.1868505,6.696409,5.855114,5.8626595,6.432326,6.405917,6.488915,6.677546,6.2889657,6.066381,6.089017,6.221059,6.40969,6.6850915,7.9300575,8.488406,8.280911,7.2623034,5.4212623,4.9345937,4.7308717,4.7006907,4.8365054,5.2062225,5.342037,5.6287565,5.7004366,5.372218,4.6516466,4.0593443,3.6292653,3.7575345,4.1989317,4.0706625,4.9647746,4.5988297,3.9386206,3.5538127,3.380272,2.7389257,2.2484846,2.2447119,2.2220762,2.2899833,3.138824,2.584248,2.8445592,3.4142256,3.5424948,2.2107582,2.71629,2.938875,3.6594462,4.67051,4.7648253,2.806833,2.8936033,4.1612053,4.90064,2.5314314,2.0636258,1.478869,0.97710985,0.7205714,0.8186596,1.1506506,1.9844007,2.3428001,1.8523588,0.73188925,0.875249,1.2638294,2.6068838,4.112161,3.470815,3.9273026,4.353609,3.731126,2.5201135,2.6483827,2.8521044,2.6898816,1.961765,0.95824677,0.49044126,0.15845025,0.06413463,0.090543,0.14335975,0.16222288,0.05281675,0.1056335,0.21503963,0.241448,0.018863125,0.011317875,0.003772625,0.011317875,0.026408374,0.041498873,0.09808825,0.094315626,0.1659955,0.36971724,0.7092535,0.9016574,0.8299775,0.663982,0.49421388,0.3169005,0.16976812,0.116951376,0.120724,0.15845025,0.23767537,0.3055826,0.23013012,0.2263575,0.38103512,0.6488915,0.7469798,0.73566186,0.88279426,1.1732863,1.297783,1.2525115,1.4411428,1.629774,1.6335466,1.3166461,0.91674787,0.7092535,0.7696155,1.0072908,1.1657411,1.2223305,1.2864652,1.2864652,1.2034674,1.0789708,0.8601585,0.7997965,0.875249,0.98465514,0.9507015,1.3694628,1.841041,1.7354075,1.1506506,0.8903395,1.1431054,0.83752275,0.42630664,0.150905,0.056589376,0.13204187,0.116951376,0.060362,0.003772625,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.211267,0.55457586,1.0412445,1.3392819,1.3996439,1.2261031,0.9393836,0.7696155,0.935611,1.177059,1.3355093,1.388326,1.4373702,1.4260522,1.2223305,0.98465514,0.83752275,0.87147635,1.0186088,1.0601076,1.0525624,0.9922004,0.7922512,0.41876137,0.3055826,0.32444575,0.4074435,0.5319401,0.4376245,1.0487897,1.3091009,0.965792,0.5696664,0.62248313,0.51684964,0.48666862,0.66020936,1.0601076,1.3166461,1.2940104,1.1846043,1.0978339,1.0374719,1.026154,1.327964,1.5430037,1.4826416,1.1695137,1.4675511,2.11267,2.7615614,2.8822856,1.780679,1.841041,1.690136,1.8485862,2.6031113,3.9989824,6.1644692,6.6322746,6.058836,5.1156793,4.4630156,4.4705606,5.172269,6.360646,7.2057137,6.277648,5.2552667,4.1612053,3.6481283,3.7462165,3.832987,3.338773,2.7804246,2.9351022,3.3727267,2.4522061,1.8749946,2.1994405,2.546522,2.6182017,2.6974268,2.2069857,2.727608,2.4371157,1.2562841,0.8337501,0.76584285,0.76584285,0.8224323,0.9280658,1.0789708,1.569412,1.297783,1.0148361,1.0110635,1.1280149,1.146878,1.056335,0.9016574,0.80356914,0.9242931,1.3128735,0.84884065,0.392353,0.2565385,0.241448,0.40367088,0.3470815,0.4074435,0.6488915,0.8601585,0.36594462,0.23013012,0.2565385,0.29049212,0.21881226,0.23013012,0.35462674,0.3772625,0.27917424,0.24899325,0.32821837,0.41876137,0.4979865,0.5583485,0.58475685,0.6451189,0.49044126,0.24899325,0.124496624,0.4074435,0.8262049,0.814887,0.5357128,0.23013012,0.23013012,0.16222288,0.08677038,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.00754525,0.0150905,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.056589376,0.026408374,0.003772625,0.011317875,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09808825,0.49421388,0.09808825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0150905,0.02263575,0.0452715,0.0452715,0.05281675,0.124496624,0.34330887,0.52439487,0.49044126,0.47157812,0.47157812,0.27917424,0.32067314,0.3961256,0.44139713,0.4376245,0.42630664,0.35462674,0.38103512,0.5055317,0.58098423,0.29426476,0.10940613,0.030181,0.018863125,0.026408374,0.018863125,0.03772625,0.0754525,0.120724,0.16976812,0.22258487,0.23767537,0.181086,0.09808825,0.030181,0.018863125,0.00754525,0.00754525,0.011317875,0.018863125,0.00754525,0.03772625,0.018863125,0.018863125,0.056589376,0.08677038,0.16976812,0.31312788,0.5093044,0.76584285,1.0789708,1.4071891,1.7278622,2.052308,2.3918443,2.7615614,3.4179983,4.4215164,5.4438977,6.175787,6.3342376,6.4964604,7.5188417,9.631512,12.694883,16.237377,19.625195,22.575388,25.51049,28.724768,32.387985,35.953117,38.725994,42.034588,47.048405,54.789833,61.64092,65.46636,66.27747,65.526726,66.11148,68.06947,68.774956,66.356705,61.77296,58.788815,54.6012,54.06549,56.82705,62.003094,68.201515,77.037,81.44343,80.84358,76.863464,73.328514,76.66351,79.3383,79.49676,77.19545,74.42258,71.52142,65.69272,59.48675,55.21614,54.94451,55.019962,55.87635,56.59692,56.657284,55.92162,56.82705,57.411808,57.679665,57.59289,57.08736,54.97092,52.38667,49.572292,46.557964,43.192783,40.15582,37.730022,35.334404,32.82561,30.479038,29.124664,28.803991,28.777584,28.434275,27.29117,27.532618,28.090965,28.362595,28.264507,28.219234,28.377686,28.751175,29.456656,30.463947,31.599506,31.150564,30.773302,30.218727,29.501928,28.890762,27.966469,27.970242,28.668177,29.766012,30.92798,32.41062,35.142002,39.197575,43.769997,47.169132,48.168877,49.94578,52.26972,54.846424,57.325035,57.951294,57.951294,57.321266,55.88767,53.30719,49.681698,45.554447,43.011696,42.392986,42.2949,43.785088,46.773006,49.421387,50.926666,51.518967,50.443768,49.187485,48.30469,47.74634,46.86732,45.346954,43.321053,41.110294,38.676952,35.590942,33.768764,28.645542,23.307278,19.40261,17.16167,15.377219,14.071891,12.574159,11.012292,10.306811,8.922258,8.311093,7.8508325,7.356619,7.092535,6.7944975,6.8473144,6.903904,6.8171334,6.643593,6.549277,6.8473144,7.0585814,7.0359454,6.983129,8.047009,8.786444,8.944894,8.360137,6.9567204,6.047518,5.4363527,5.2892203,5.4967146,5.6476197,6.009792,6.628502,6.9680386,6.8058157,6.2021956,5.3873086,4.859141,4.7120085,4.8629136,5.0666356,2.305074,1.7919968,1.9655377,2.3578906,2.6408374,2.6408374,2.444661,2.505023,2.2296214,1.6373192,1.358145,2.1013522,2.9841464,3.399135,3.4330888,3.8593953,3.2482302,2.082489,1.1053791,1.0035182,2.3956168,4.3347464,4.244203,3.1237335,2.1164427,2.516341,3.5538127,4.217795,3.9122121,3.2105038,3.8443048,4.0404816,3.9348478,3.4330888,2.7691069,2.5012503,2.7238352,3.591539,3.9197574,3.712263,4.164978,3.029418,2.2899833,1.7693611,1.3430545,0.91674787,1.8787673,3.4859054,3.6858547,2.1277604,0.1358145,0.0754525,0.08677038,0.1659955,0.24899325,0.19994913,0.1358145,0.23013012,0.2678564,0.17731337,0.030181,0.041498873,0.026408374,0.033953626,0.056589376,0.030181,0.00754525,0.0,0.030181,0.15845025,0.48666862,0.6828451,0.7130261,0.663982,0.56212115,0.36594462,0.20749438,0.13204187,0.14335975,0.2263575,0.33576363,0.47157812,0.3734899,0.33953625,0.43007925,0.5017591,0.49044126,0.35085413,0.29049212,0.32067314,0.26031113,0.38103512,0.45648763,0.47535074,0.422534,0.29049212,0.48666862,0.5885295,0.69793564,0.83752275,0.94692886,0.935611,0.965792,0.965792,0.94692886,1.0072908,1.177059,1.5580941,2.003264,2.3163917,2.2447119,3.3764994,3.361409,2.444661,1.5618668,2.3201644,2.4672968,1.3845534,0.422534,0.07922512,0.030181,0.018863125,0.071679875,0.0754525,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.150905,0.38103512,0.79602385,1.3770081,1.6637276,1.4637785,0.8526133,0.7582976,0.9242931,1.0902886,1.1695137,1.267602,1.4147344,1.2751472,1.0374719,0.8224323,0.70170826,0.7394345,0.77338815,0.84884065,0.91297525,0.83752275,0.44894236,0.20372175,0.1358145,0.21503963,0.33576363,0.29803738,0.47157812,0.97333723,1.4864142,1.267602,0.9507015,0.48666862,0.4979865,0.9507015,1.1431054,1.4977322,1.448688,1.6675003,1.8561316,0.73188925,0.7696155,0.8337501,1.1732863,1.3770081,0.35085413,1.6448646,1.7580433,1.6976813,1.6976813,1.2223305,1.659955,1.4147344,1.2110126,1.4713237,2.2899833,2.4371157,4.06689,5.040227,4.5233774,2.9615107,2.1654868,2.7011995,3.531177,4.115934,4.4101987,4.8138695,4.4177437,3.4557245,2.686109,3.4179983,3.9197574,3.229367,3.4481792,4.146115,2.3654358,2.0372176,2.6031113,2.7691069,2.2598023,1.8297231,2.9916916,2.3578906,1.7655885,1.6524098,1.0525624,0.6752999,0.76207024,0.77338815,0.5772116,0.44139713,0.5017591,0.6488915,0.8601585,1.1280149,1.4335974,1.4826416,1.4034165,1.1355602,0.9016574,1.20724,2.8030603,1.9768555,0.9016574,0.48666862,0.35085413,0.6790725,0.633801,0.62248313,0.6526641,0.33576363,0.24899325,0.32067314,0.35839936,0.27917424,0.120724,0.2678564,0.44139713,0.38103512,0.1358145,0.0754525,0.08677038,0.29426476,0.63002837,0.8903395,0.73188925,0.34330887,0.27917424,0.21503963,0.07922512,0.090543,0.17731337,0.09808825,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.150905,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.060362,0.124496624,0.19994913,0.271629,0.29803738,0.4640329,0.66020936,0.48666862,0.5357128,0.47535074,0.5319401,0.62248313,0.36594462,0.2565385,0.23013012,0.41121614,0.7092535,0.80734175,0.30935526,0.071679875,0.00754525,0.018863125,0.030181,0.030181,0.041498873,0.0754525,0.1358145,0.19994913,0.32067314,0.27917424,0.181086,0.1056335,0.090543,0.041498873,0.030181,0.060362,0.090543,0.030181,0.13958712,0.06790725,0.02263575,0.071679875,0.120724,0.20749438,0.211267,0.271629,0.45648763,0.7469798,1.1280149,1.4675511,1.8146327,2.2258487,2.7615614,3.3463185,4.4818783,5.881522,7.1038527,7.567886,7.250985,7.326438,7.986647,9.276885,11.11038,15.309312,20.29295,25.103046,29.324614,33.09724,37.733795,42.3364,45.5469,47.259674,48.614044,53.27701,60.539314,66.71887,69.895424,69.929375,71.27243,72.8343,75.411,77.61044,75.863716,68.99377,62.83684,59.596157,60.95053,68.05438,82.29981,95.20596,98.92954,92.43308,81.49625,79.26285,80.372,80.74172,78.37628,73.347374,69.03904,63.319736,57.71739,53.32228,50.783306,49.45157,49.345936,50.46263,52.318764,53.95608,54.2843,55.438725,57.72116,60.471405,62.05591,62.252087,59.47166,55.0841,50.74935,48.414097,45.595947,42.07986,39.503155,37.85452,35.462673,32.39553,31.422194,29.969732,27.78161,26.90259,26.936543,26.71773,26.985586,27.743885,28.245644,27.76652,27.559025,27.78161,28.49841,29.63397,30.91289,31.61837,31.954134,32.07863,32.089947,29.916916,28.347504,27.547709,27.340214,27.208172,27.721249,29.294434,31.290152,33.617863,36.74537,40.13696,43.739815,46.225975,47.71616,49.806194,52.2584,54.318256,56.34038,58.128605,58.958584,58.60396,56.18193,52.005634,46.76169,41.487556,38.974987,39.446568,41.238564,43.464413,45.992073,49.394978,51.13416,50.798397,49.029034,47.516212,46.014706,44.833874,44.192528,43.97749,43.74736,41.8535,38.808994,34.84019,30.36963,26.00093,20.934296,16.984358,14.769827,13.905896,13.015556,12.796744,11.917723,11.076427,10.450171,9.703192,9.484379,8.386545,7.643338,7.6093845,7.7678347,7.54525,7.77538,7.914967,7.884786,8.058327,8.98262,9.673011,9.593785,8.89585,8.409182,7.91874,7.194396,6.858632,6.8435416,6.3945994,6.3945994,6.6134114,7.0284004,7.4584794,7.567886,6.56814,6.3908267,6.458734,6.3229194,5.6778007,3.0256453,2.5389767,2.0485353,1.7014539,1.5505489,1.5430037,2.6936543,2.323937,1.9240388,1.9089483,1.5882751,1.690136,2.4710693,2.5729303,1.9429018,1.8334957,1.8863125,3.1614597,3.1463692,1.7769064,1.4298248,1.5354583,1.4034165,1.1242423,0.9393836,1.237421,1.3770081,1.4600059,1.5430037,1.6750455,1.9278114,2.6031113,2.3956168,1.9089483,1.5354583,1.4524606,1.7391801,1.8146327,2.1503963,2.9652832,4.2404304,3.5538127,4.666737,5.1873593,4.13857,1.9655377,1.3166461,1.1129243,1.0638802,0.8563859,0.17354076,0.094315626,0.14335975,0.41498876,0.73188925,0.6752999,0.211267,0.77716076,0.84129536,0.20372175,0.018863125,0.030181,0.23390275,0.32067314,0.19994913,0.030181,0.00754525,0.0,0.00754525,0.049044125,0.18485862,0.27917424,0.331991,0.5055317,0.67152727,0.3772625,0.23767537,0.15467763,0.13204187,0.211267,0.45648763,0.513077,0.35462674,0.3470815,0.5319401,0.62625575,0.51684964,0.44516975,0.3734899,0.29426476,0.23390275,0.36594462,0.33576363,0.2678564,0.26031113,0.39989826,0.41876137,0.3470815,0.3169005,0.43007925,0.77338815,0.5885295,0.5093044,0.48666862,0.49044126,0.543258,0.5394854,0.77338815,0.97333723,1.0827434,1.2411937,2.6898816,2.9615107,2.655928,2.2371666,2.0372176,1.5128226,0.6790725,0.28294688,0.36594462,0.29803738,0.10186087,0.06413463,0.049044125,0.0150905,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.030181,0.003772625,0.011317875,0.0,0.011317875,0.003772625,0.00754525,0.0452715,0.150905,0.271629,0.7997965,1.4034165,1.6976813,1.2449663,0.784706,0.6526641,0.7054809,0.83752275,0.98465514,1.1695137,1.2638294,1.2110126,1.0223814,0.77338815,0.5583485,0.48666862,0.513077,0.56212115,0.5583485,0.422534,0.2263575,0.08677038,0.060362,0.150905,0.19240387,0.1961765,0.29426476,0.7205714,1.8297231,1.5015048,1.0035182,0.8224323,0.9695646,0.9997456,1.5656394,1.3015556,1.0940613,1.0525624,0.47535074,0.58098423,1.0714256,1.6373192,1.7882242,0.83752275,1.9768555,2.1692593,1.6033657,0.8337501,0.7582976,0.9997456,0.875249,1.0714256,1.6675003,2.093807,1.4411428,2.203213,2.9011486,3.0445085,3.1312788,1.9655377,2.4522061,2.969056,2.8143783,2.1881225,3.3048196,3.1237335,2.795515,3.2482302,5.198677,3.5538127,2.3314822,1.7278622,1.5920477,1.448688,1.7844516,2.233394,2.0296721,1.358145,1.3317367,1.4637785,1.1657411,1.7580433,2.5087957,0.6488915,1.1695137,0.8601585,0.67152727,0.8639311,0.9922004,0.7696155,0.935611,1.4864142,1.8938577,1.116697,1.6146835,1.7354075,1.2864652,0.66775465,0.8639311,1.5845025,1.5543215,1.1317875,0.72811663,0.8262049,0.5319401,0.2565385,0.13204187,0.13204187,0.07922512,0.15845025,0.42630664,0.8224323,1.0072908,0.34330887,0.1961765,0.17731337,0.1659955,0.1961765,0.4678055,0.30181,0.35462674,0.4640329,0.46026024,0.14713238,0.06790725,0.056589376,0.041498873,0.0150905,0.018863125,0.033953626,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.011317875,0.011317875,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.06413463,0.1358145,0.19994913,0.23390275,0.27917424,0.32821837,0.29426476,0.24522063,0.20372175,0.19994913,0.21503963,0.18485862,0.181086,0.1659955,0.2263575,0.35085413,0.41876137,0.241448,0.10186087,0.026408374,0.018863125,0.030181,0.041498873,0.05281675,0.0754525,0.09808825,0.10186087,0.25276586,0.36971724,0.41498876,0.39989826,0.3961256,0.47535074,0.47912338,0.36971724,0.20372175,0.150905,0.15467763,0.06413463,0.003772625,0.018863125,0.03772625,0.05281675,0.06790725,0.116951376,0.22258487,0.41876137,0.7092535,1.0487897,1.418507,1.81086,2.2484846,2.8143783,3.6594462,4.859141,6.1003346,6.700182,7.115171,7.492433,7.956466,8.605357,9.495697,11.344283,14.019074,18.12369,23.752447,30.520536,36.945316,42.11381,46.391968,49.84015,52.190495,53.74859,57.019455,61.591877,66.51515,70.32173,72.74753,75.8939,79.27417,82.428085,84.91047,83.088295,77.50481,71.59688,67.97138,68.39769,74.74325,83.98241,89.53194,88.351105,80.94921,76.799324,77.37654,78.72714,78.0443,73.67937,70.47263,66.31898,61.863506,56.993046,50.828575,49.274254,48.697044,48.421642,48.346188,48.93849,49.677925,50.662582,52.696026,55.7594,59.018944,61.606968,62.286037,60.795853,57.479713,53.32228,49.94578,47.15027,45.02628,43.468185,42.136448,39.79742,37.888474,35.88898,33.621635,31.24488,29.29066,28.37014,28.287142,28.717222,29.207663,28.411638,27.928743,27.977787,28.256962,27.947605,28.223007,29.056757,30.19609,31.433512,32.63698,32.146538,31.05625,29.796192,28.558771,27.29117,27.03463,27.498663,28.328642,29.39252,30.799711,33.119873,36.115337,38.771267,40.865074,42.992836,45.26018,47.335125,49.3648,51.424652,53.514687,54.03908,54.348434,54.865284,55.219913,54.2428,50.25514,46.754143,44.388706,43.053196,41.887455,42.521255,44.030308,45.758167,47.09745,47.478485,47.68598,47.048405,46.014706,44.9131,43.96617,41.99686,40.65381,39.39375,37.67343,34.92319,30.950615,26.404602,22.092491,18.780127,17.165443,16.418465,15.011275,13.758763,12.928786,12.242168,11.046246,10.137043,9.899368,10.163452,10.197406,9.390063,9.148616,9.009028,8.854351,8.937348,9.646602,10.884023,11.514051,11.170743,10.26154,9.454198,8.688355,8.160188,7.8432875,7.5301595,7.6848373,7.9526935,8.156415,8.254503,8.326183,8.152642,8.273367,8.526133,8.831716,9.178797,3.651901,5.191132,5.726845,5.4288073,4.5761943,3.5462675,4.7572803,5.9117036,7.326438,7.3377557,2.2975287,3.2557755,3.5651307,2.9501927,1.8146327,1.2525115,1.327964,2.969056,4.6742826,5.1156793,3.138824,2.082489,1.9466745,2.2258487,2.595566,2.8936033,1.539231,1.237421,1.5203679,1.8674494,1.6863633,1.931584,1.931584,2.052308,2.3767538,2.6898816,3.5689032,3.0030096,2.0372176,1.7089992,3.0746894,3.3878171,3.8103511,3.4179983,2.2371666,1.2298758,0.56212115,0.241448,0.21881226,0.3169005,0.24899325,0.6149379,0.41121614,0.33576363,0.6413463,1.1242423,0.44516975,0.6413463,0.6790725,0.3055826,0.05281675,0.049044125,0.1961765,0.3169005,0.2867195,0.02263575,0.011317875,0.03772625,0.03772625,0.018863125,0.05281675,0.0754525,0.094315626,0.19994913,0.32821837,0.25276586,0.23013012,0.18863125,0.15845025,0.16976812,0.2678564,0.35462674,0.33953625,0.33576363,0.36971724,0.362172,0.38858038,0.41121614,0.41876137,0.482896,0.7582976,0.47535074,0.3470815,0.28294688,0.2678564,0.38103512,0.38480774,0.26031113,0.23767537,0.452715,0.9507015,0.5885295,0.41498876,0.331991,0.28294688,0.24522063,0.23013012,0.3734899,0.44516975,0.46026024,0.6790725,1.7957695,2.3465726,2.4899325,2.2786655,1.6561824,0.9695646,0.47157812,0.28294688,0.29426476,0.14713238,0.049044125,0.02263575,0.02263575,0.0150905,0.00754525,0.0,0.003772625,0.003772625,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.0150905,0.003772625,0.003772625,0.0,0.003772625,0.003772625,0.0,0.00754525,0.03772625,0.056589376,0.3169005,0.7884786,1.3091009,1.5882751,1.2600567,0.7922512,0.51684964,0.52062225,0.66020936,0.76584285,0.8337501,0.83752275,0.7809334,0.6828451,0.543258,0.44139713,0.3961256,0.3961256,0.41498876,0.452715,0.38858038,0.23390275,0.071679875,0.071679875,0.071679875,0.056589376,0.16222288,0.4640329,0.98842776,0.91674787,0.9997456,1.0223814,0.9997456,1.1619685,1.9466745,1.7089992,1.2789198,0.9695646,0.59607476,0.7469798,1.0450171,1.20724,1.1619685,1.0638802,1.5882751,1.50905,1.2940104,1.116697,0.8337501,0.73566186,0.59230214,0.6413463,0.95824677,1.448688,0.60362,1.0299267,1.6863633,2.1541688,2.6332922,2.546522,2.2711203,1.871222,1.4222796,0.9922004,1.5543215,1.4939595,1.4562333,1.9730829,3.4481792,2.2899833,1.9278114,1.5807298,1.1619685,1.2864652,3.0445085,2.5540671,1.569412,0.9808825,0.8111144,0.77716076,0.84884065,1.4147344,1.8372684,0.44894236,1.3845534,0.95824677,0.56589377,0.6488915,0.69793564,0.7054809,0.69793564,1.1996948,1.7618159,0.95447415,0.8639311,1.1091517,1.1581959,1.1204696,1.7655885,1.6373192,1.3996439,1.0035182,0.5772116,0.41498876,0.21881226,0.10940613,0.041498873,0.0,0.00754525,0.056589376,0.21503963,0.41121614,0.482896,0.15845025,0.071679875,0.0452715,0.0452715,0.08677038,0.23390275,0.150905,0.15845025,0.17354076,0.14335975,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.003772625,0.0,0.00754525,0.018863125,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.00754525,0.03772625,0.094315626,0.13958712,0.1659955,0.17731337,0.181086,0.18863125,0.18863125,0.16976812,0.14713238,0.14335975,0.18485862,0.18485862,0.16222288,0.181086,0.24899325,0.30181,0.29803738,0.181086,0.071679875,0.026408374,0.030181,0.033953626,0.05281675,0.16222288,0.2867195,0.18485862,0.23390275,0.3772625,0.46026024,0.43007925,0.32821837,0.29049212,0.26408374,0.1961765,0.10940613,0.090543,0.090543,0.041498873,0.00754525,0.00754525,0.00754525,0.0150905,0.026408374,0.060362,0.124496624,0.25276586,0.47157812,0.76584285,1.1091517,1.4750963,1.8372684,2.305074,2.9916916,3.9159849,4.8968673,5.560849,6.0626082,6.752999,7.443389,8.118689,8.937348,10.246449,11.876224,14.25675,17.73511,22.590479,29.24916,37.232037,44.947056,51.258656,55.491543,57.08736,59.464115,61.769188,64.10445,67.526215,71.89491,76.28625,79.73066,81.952736,83.38256,84.79352,84.257805,81.91501,77.91602,72.4344,70.419815,73.78877,77.169044,77.5199,74.12831,71.347885,70.974396,71.347885,71.3177,70.23496,71.261116,69.68038,66.55665,61.36929,51.994316,49.10826,47.338898,46.142975,45.528038,46.026024,46.86732,47.62939,48.93849,50.809715,52.635666,56.008392,59.3283,61.24102,61.056164,58.78127,55.140686,51.786823,48.94981,46.791866,45.392223,44.17744,43.988808,43.094696,40.77076,37.315033,35.209908,33.606544,32.195583,30.969479,30.218727,29.24539,28.709677,28.604042,28.800219,29.064302,28.724768,28.075874,28.064558,28.917171,30.147047,30.675215,31.109066,30.961933,30.120638,28.834173,28.31355,27.555252,27.1629,27.385485,28.121147,29.358568,31.871136,34.444065,36.439785,37.78284,39.559746,41.902546,44.184982,46.06375,47.45962,47.829338,48.463142,49.80242,51.662327,53.224194,53.126106,52.092407,50.11178,47.346443,44.12085,42.200584,41.2612,41.37438,42.11004,42.562756,43.170147,43.985035,44.675426,44.920647,44.40757,42.9287,42.264717,41.717686,40.766987,39.057987,36.2172,32.750156,29.13221,25.816072,23.23937,21.364376,19.57615,17.980331,16.55428,15.147089,13.59654,12.427027,11.759273,11.566868,11.664956,11.159425,11.193378,11.25374,11.234878,11.442371,11.9064045,12.472299,12.830698,12.736382,12.019584,10.95193,10.265312,9.710737,9.186342,8.744945,8.714764,9.012801,9.405154,9.612649,9.303293,10.012547,10.861387,11.491416,11.442371,10.167224,2.4371157,4.568649,5.5570765,5.594803,4.930821,3.85185,4.285702,5.824933,7.911195,8.394091,3.5236318,4.217795,4.2781568,3.8141239,3.1463692,2.8219235,2.6823363,4.142342,6.198423,7.4471617,6.1003346,4.6931453,3.5839937,3.3274553,3.9122121,4.768598,2.8106055,2.7691069,3.8556228,4.8855495,4.2630663,3.8820312,4.4894238,5.1156793,5.138315,4.2781568,4.4516973,3.7537618,2.5012503,1.7052265,3.0746894,3.5953116,2.9200118,1.750498,0.7205714,0.3772625,0.11317875,0.094315626,0.18485862,0.2867195,0.34330887,0.9393836,1.0827434,1.2638294,1.6184561,1.9240388,1.0148361,0.8903395,0.8903395,0.67152727,0.23013012,0.24899325,0.43007925,0.73566186,0.8978847,0.38103512,0.09808825,0.056589376,0.05281675,0.018863125,0.0150905,0.1056335,0.18485862,0.22258487,0.2565385,0.39989826,0.43007925,0.27917424,0.15467763,0.124496624,0.12826926,0.28294688,0.41121614,0.44516975,0.422534,0.48666862,0.5998474,0.52439487,0.5093044,0.66775465,1.0035182,0.5583485,0.38103512,0.30935526,0.27917424,0.32821837,0.271629,0.1961765,0.20372175,0.36594462,0.7130261,0.43007925,0.30181,0.23013012,0.15845025,0.090543,0.090543,0.150905,0.18863125,0.21881226,0.38103512,0.9507015,1.5052774,1.8523588,1.8070874,1.2185578,0.79602385,0.5470306,0.35085413,0.16222288,0.0,0.003772625,0.003772625,0.003772625,0.011317875,0.02263575,0.018863125,0.0150905,0.00754525,0.0,0.0,0.00754525,0.003772625,0.003772625,0.003772625,0.0,0.0,0.011317875,0.033953626,0.06790725,0.090543,0.018863125,0.018863125,0.0754525,0.11317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.30935526,0.8299775,1.6561824,1.81086,1.1959221,0.5772116,0.32067314,0.38480774,0.47912338,0.513077,0.5319401,0.5696664,0.62248313,0.6526641,0.59230214,0.5093044,0.44139713,0.4074435,0.5281675,0.56212115,0.452715,0.26031113,0.18485862,0.241448,0.27917424,0.41121614,0.5319401,0.33576363,0.36594462,0.7922512,0.9997456,0.94692886,1.1431054,1.931584,1.8976303,1.5316857,1.1959221,1.0902886,1.5467763,1.4260522,1.0978339,0.9242931,1.2336484,1.2902378,1.0223814,1.0223814,1.1883769,0.73566186,0.754525,0.63002837,0.44139713,0.38480774,0.7469798,0.3169005,0.4979865,0.9205205,1.4071891,1.9881734,2.6672459,2.4371157,1.8787673,1.4109617,1.2525115,1.0525624,0.84129536,0.88279426,1.3355093,2.252257,1.6109109,1.5052774,1.5467763,1.4637785,1.1091517,3.1765501,2.293756,1.086516,0.633801,0.44516975,0.45648763,0.573439,0.7432071,0.7809334,0.392353,0.98842776,0.6451189,0.3055826,0.27540162,0.24899325,0.5583485,0.63002837,0.9393836,1.3053282,0.91674787,0.362172,0.5093044,0.8601585,1.2034674,1.5882751,1.1581959,0.84129536,0.55457586,0.2678564,0.03772625,0.026408374,0.056589376,0.0452715,0.0,0.0,0.003772625,0.071679875,0.08299775,0.026408374,0.00754525,0.0,0.0,0.003772625,0.0150905,0.033953626,0.030181,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.003772625,0.018863125,0.05281675,0.07922512,0.10186087,0.116951376,0.13204187,0.1659955,0.21503963,0.23013012,0.20372175,0.16976812,0.21503963,0.20749438,0.1961765,0.19994913,0.2263575,0.26408374,0.3470815,0.26031113,0.1358145,0.056589376,0.056589376,0.056589376,0.06413463,0.1659955,0.2867195,0.181086,0.1659955,0.25276586,0.30935526,0.28294688,0.181086,0.090543,0.041498873,0.02263575,0.018863125,0.018863125,0.026408374,0.0150905,0.011317875,0.0150905,0.00754525,0.018863125,0.026408374,0.0452715,0.090543,0.1659955,0.3169005,0.55457586,0.86770374,1.2110126,1.5316857,1.8561316,2.354118,2.9954643,3.7084904,4.4139714,4.927048,5.745708,6.598321,7.424526,8.3525915,9.623966,10.925522,12.423254,14.268067,16.595778,21.835953,29.271797,37.820564,46.674915,55.299137,61.95405,65.60972,66.288795,65.60217,66.745285,71.74401,76.712555,79.88156,80.67381,79.723114,80.636086,82.8808,84.48039,83.54855,78.319695,71.51388,70.34814,71.37052,72.483444,72.93616,71.17057,69.52948,67.66203,65.88889,65.19473,68.4656,69.41253,67.594124,62.708572,54.61252,52.03959,49.244076,46.576828,44.747105,44.837646,45.109276,45.697807,46.158066,46.384426,46.60701,49.130894,52.254627,55.70281,58.634136,59.61502,57.743797,55.84617,53.559956,50.915348,48.346188,47.040863,47.233265,47.052177,45.641216,43.143738,41.268745,39.17871,36.99436,34.91942,33.202873,31.652325,30.690304,30.256453,30.218727,30.39604,29.550972,28.204145,27.317577,27.27608,27.872154,28.60027,29.467974,30.184772,30.520536,30.271544,30.716713,29.724512,28.562544,27.88347,27.725021,28.015512,29.407612,31.05625,32.501163,33.66313,35.67017,38.40155,40.97448,42.807976,43.637955,43.86054,43.958626,44.332115,45.214912,46.663597,49.134666,50.881393,51.141705,49.877876,47.776524,45.354496,43.09847,41.41588,40.276543,39.21644,38.982533,39.684242,40.683987,41.596962,42.302444,42.306217,42.59671,42.460896,41.789368,41.072567,39.284344,37.03586,34.33466,31.339195,28.37014,26.340467,24.623924,22.88097,20.979568,18.99894,17.150352,15.543215,14.2944765,13.494679,13.215506,13.011784,13.091009,13.087236,12.966512,13.038192,13.502225,13.6682205,13.777626,13.875714,13.800262,12.830698,11.955449,11.321648,10.906659,10.521852,10.344538,10.340765,10.525623,10.714255,10.529396,11.619685,13.50977,14.671739,14.056801,11.087745,0.150905,1.0186088,1.4222796,1.720317,1.9240388,1.7052265,1.2864652,1.6675003,2.6936543,3.7688525,3.8443048,3.2746384,3.4783602,4.0216184,4.6290107,5.1760416,4.98741,6.0739264,6.8473144,7.1264887,8.122461,7.2396674,5.1760416,4.063117,4.5912848,6.013564,4.3649273,4.8553686,6.9944468,8.903395,7.2962565,6.4021444,7.3905725,8.171506,7.4509344,4.7610526,3.531177,3.2482302,2.8898308,2.5729303,3.5689032,3.5877664,2.8294687,1.8825399,1.0072908,0.1358145,0.150905,0.241448,0.39989826,0.5357128,0.47912338,0.9318384,1.8825399,2.7917426,3.1614597,2.565385,1.5354583,1.4411428,1.3958713,1.0072908,0.392353,0.482896,0.97333723,1.7240896,2.1654868,1.3355093,0.41498876,0.120724,0.10940613,0.14335975,0.0754525,0.28294688,0.4678055,0.5319401,0.55457586,0.80734175,0.7922512,0.44894236,0.18863125,0.14713238,0.21503963,0.51684964,0.7167987,0.7469798,0.7092535,0.88279426,0.95824677,0.73188925,0.62625575,0.724344,0.7696155,0.60362,0.42630664,0.29426476,0.24522063,0.29426476,0.20749438,0.2263575,0.19994913,0.124496624,0.120724,0.1056335,0.12826926,0.116951376,0.06790725,0.03772625,0.018863125,0.02263575,0.071679875,0.15467763,0.23013012,0.392353,0.724344,1.0336993,1.1317875,0.8224323,0.80356914,0.6526641,0.38480774,0.1056335,0.00754525,0.0150905,0.00754525,0.0,0.00754525,0.026408374,0.03772625,0.033953626,0.018863125,0.00754525,0.00754525,0.0,0.0,0.003772625,0.011317875,0.0,0.003772625,0.02263575,0.071679875,0.1358145,0.19240387,0.056589376,0.06413463,0.19240387,0.28294688,0.0452715,0.011317875,0.003772625,0.003772625,0.003772625,0.0,0.0,0.00754525,0.11317875,0.47157812,1.3015556,2.0070364,1.5958204,0.8563859,0.30935526,0.22258487,0.3470815,0.41498876,0.45648763,0.5093044,0.5998474,0.77716076,0.84129536,0.80356914,0.68661773,0.52062225,0.59607476,0.6375736,0.60362,0.5055317,0.4376245,0.56212115,0.59230214,0.6187105,0.58098423,0.2678564,0.25276586,0.55080324,0.7432071,0.7507524,0.8299775,1.3619176,1.4826416,1.3958713,1.3317367,1.5580941,2.214531,1.81086,1.3694628,1.3128735,1.4449154,1.2864652,1.0487897,0.8639311,0.70170826,0.35085413,0.8186596,0.7507524,0.47157812,0.2565385,0.30935526,0.45648763,0.3734899,0.36971724,0.6526641,1.3128735,1.8184053,2.3088465,2.4484336,2.293756,2.2899833,1.5505489,1.0601076,1.1242423,1.6788181,2.3088465,1.448688,0.8903395,1.1657411,1.7165444,0.875249,2.0070364,1.478869,0.6451189,0.22258487,0.27917424,0.2678564,0.181086,0.08677038,0.094315626,0.362172,0.2867195,0.271629,0.21881226,0.12826926,0.0754525,0.44894236,0.8337501,1.0110635,0.965792,0.90543,0.44139713,0.34330887,0.513077,0.6488915,0.2678564,0.06413463,0.05281675,0.056589376,0.018863125,0.003772625,0.011317875,0.018863125,0.0150905,0.0,0.0,0.011317875,0.07922512,0.094315626,0.049044125,0.030181,0.02263575,0.011317875,0.0150905,0.030181,0.05281675,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.003772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.049044125,0.07922512,0.11317875,0.17731337,0.22258487,0.26408374,0.23767537,0.18863125,0.23767537,0.24899325,0.241448,0.22258487,0.20372175,0.20749438,0.32444575,0.331991,0.26408374,0.18485862,0.16222288,0.120724,0.090543,0.08299775,0.08677038,0.071679875,0.071679875,0.08677038,0.1056335,0.11317875,0.116951376,0.090543,0.0452715,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.02263575,0.030181,0.0452715,0.0754525,0.12826926,0.22258487,0.41498876,0.70170826,1.0450171,1.3656902,1.5807298,1.8599042,2.252257,2.7804246,3.4330888,4.0178456,4.7421894,5.5306683,6.3719635,7.284939,8.43559,9.793735,11.465008,13.268322,14.724555,17.935059,21.624687,27.660887,36.967953,49.519474,62.41808,68.997536,70.82349,69.925606,68.81645,72.20427,76.51261,79.31944,79.674065,78.10465,76.85214,77.78021,80.03624,82.073456,81.6396,75.35064,72.69094,72.33631,73.513374,75.99576,74.6263,72.75884,69.25785,64.82124,61.96914,64.24403,65.86626,64.18367,59.81874,56.691235,56.117798,53.55241,49.911827,46.644737,45.758167,45.135685,45.448814,45.094185,43.985035,43.554955,44.000126,44.48302,46.806957,50.794624,54.29562,55.714127,57.192993,57.223175,55.351955,52.18672,49.94578,48.700817,48.082108,47.693523,47.104996,45.486538,43.585136,41.695053,39.959644,38.367596,36.413376,34.85151,33.82913,33.10856,32.07486,30.811028,29.830147,28.883217,28.05324,27.76652,27.834427,27.740112,28.31355,29.543427,30.558262,32.542664,32.72752,32.097492,31.222244,30.26777,29.747149,29.162392,28.819082,29.04544,30.207409,32.59548,35.33063,38.118603,40.502903,41.898773,42.70989,42.796658,42.38544,41.796913,41.4536,42.483532,44.154804,45.81853,47.10877,47.950066,47.29363,46.29388,44.777287,42.65707,39.948326,38.405323,37.499893,36.89627,36.790638,37.907337,39.34848,40.740578,41.370605,41.385696,41.744095,41.110294,39.81251,37.601753,34.704376,31.837183,30.45263,29.113348,27.453392,25.499172,23.643042,21.737865,20.002459,18.357594,16.890041,15.833707,15.403628,15.030138,14.532151,13.95494,13.577678,14.064346,14.388792,14.596286,14.841507,15.373446,14.822643,13.72481,12.989148,12.845788,12.849561,12.494934,12.064855,11.744182,11.680047,11.993175,12.913695,15.335721,16.7995,15.939341,12.483616,0.090543,0.4074435,0.55080324,0.79602385,0.9620194,0.41121614,0.120724,0.090543,0.21881226,0.36594462,0.36594462,0.392353,0.88279426,1.991946,3.5160866,4.881777,5.2137675,4.8742313,4.349837,4.432834,6.2399216,6.7643166,6.722818,6.7944975,7.194396,7.6584287,5.828706,5.873977,7.809334,9.152389,4.927048,3.5236318,3.3123648,4.08198,4.7120085,3.1727777,2.8332415,3.240685,2.9539654,1.7882242,0.8224323,1.1544232,2.003264,1.9089483,0.8563859,0.32067314,0.5281675,0.5885295,0.69793564,0.8224323,0.68661773,1.0412445,2.071171,2.7691069,2.625747,1.6637276,1.0525624,1.056335,0.94692886,0.5281675,0.1358145,0.28294688,1.3920987,2.8634224,3.7914882,2.9615107,1.177059,0.422534,0.3961256,0.5998474,0.32067314,0.38103512,0.47912338,0.5696664,0.7092535,1.0525624,0.965792,0.72811663,0.48666862,0.38858038,0.5357128,1.20724,1.4449154,1.2261031,0.77338815,0.56589377,0.5998474,0.6375736,0.6451189,0.5998474,0.48666862,0.7432071,0.55080324,0.331991,0.2678564,0.3055826,0.56212115,0.633801,0.4640329,0.16976812,0.060362,0.120724,0.1659955,0.13958712,0.060362,0.0,0.0,0.00754525,0.033953626,0.08677038,0.18485862,0.34330887,0.56589377,0.72811663,0.7582976,0.62625575,0.6375736,0.49421388,0.27917424,0.090543,0.030181,0.030181,0.011317875,0.00754525,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.033953626,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.00754525,0.0452715,0.1056335,0.13958712,0.21503963,0.29049212,0.23013012,0.056589376,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.018863125,0.12826926,0.45648763,1.3505998,1.6071383,1.2298758,0.5394854,0.19994913,0.18485862,0.24899325,0.31312788,0.36971724,0.44139713,0.73566186,1.0186088,1.146878,1.0450171,0.70170826,0.55457586,0.52062225,0.5319401,0.5583485,0.59607476,0.44894236,0.21881226,0.1056335,0.09808825,0.0,0.20749438,0.2678564,0.3055826,0.3772625,0.48666862,0.6111652,0.513077,0.63002837,0.98465514,1.20724,0.9242931,0.7092535,0.8978847,1.3958713,1.6788181,1.1657411,0.9997456,0.7205714,0.30181,0.1659955,0.5470306,0.41121614,0.20372175,0.17354076,0.38103512,0.392353,0.22258487,0.06413463,0.06790725,0.33576363,0.2263575,0.34330887,0.845068,1.6222287,2.305074,1.0450171,0.59607476,0.8337501,1.2449663,0.91674787,0.18485862,0.2565385,1.0072908,1.7542707,1.267602,1.8523588,1.4600059,0.66020936,0.049044125,0.24522063,0.21881226,0.1659955,0.1358145,0.14335975,0.1659955,0.23013012,0.91297525,1.0940613,0.6375736,0.38103512,0.38103512,0.7922512,1.086516,1.0412445,0.7469798,0.6149379,0.46026024,0.23013012,0.0,0.0,0.0,0.026408374,0.0452715,0.041498873,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.011317875,0.041498873,0.090543,0.1056335,0.060362,0.018863125,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.07922512,0.150905,0.18863125,0.18863125,0.18863125,0.2263575,0.33576363,0.38480774,0.27917424,0.20372175,0.1961765,0.120724,0.2678564,0.4074435,0.51684964,0.55080324,0.44139713,0.23390275,0.12826926,0.090543,0.094315626,0.1056335,0.1056335,0.116951376,0.12826926,0.13958712,0.150905,0.116951376,0.060362,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.049044125,0.090543,0.150905,0.23767537,0.4074435,0.66775465,1.0110635,1.388326,1.6448646,1.8372684,2.0673985,2.372981,2.7011995,3.138824,3.6707642,4.304565,5.0515447,5.904158,7.0284004,8.654402,10.133271,11.61214,14.053028,16.825907,19.53088,23.182781,28.754948,37.201855,47.931202,58.98122,67.69221,71.95528,70.21987,70.06142,71.67233,74.13208,76.625786,78.44419,79.37226,77.99525,76.16175,75.10919,75.426094,74.411255,73.13988,70.90649,68.58632,68.63537,70.148186,71.70628,70.25005,66.545334,65.21737,65.851166,63.7385,58.977448,54.06926,53.910812,54.348434,54.559704,53.582592,51.605736,49.9571,49.187485,48.712135,47.519985,45.826077,45.045143,42.9702,41.20461,40.521767,41.57433,44.905556,48.387688,51.700054,54.389935,56.01971,56.16684,54.48425,53.04688,51.349197,49.436478,47.897247,47.323807,47.09745,46.029797,44.445293,44.188755,43.702087,42.35149,40.506676,38.57132,36.971725,35.579628,34.21771,32.867107,31.584417,30.486582,29.13221,28.189054,27.88347,28.249416,29.128437,31.241108,33.738586,36.122883,37.79793,38.05447,36.722733,33.610317,30.343224,27.99665,27.068584,27.826881,29.305752,32.22576,36.062523,39.07685,41.630917,43.47573,44.29439,44.075577,43.136196,40.035095,38.575092,38.09974,38.405323,39.733288,41.72523,44.098213,45.47145,45.18473,43.30596,41.461147,40.076595,38.54491,36.639732,34.515747,34.832645,35.919163,37.303715,38.692043,39.963417,41.038616,41.185745,40.30295,38.2846,35.047688,33.206646,31.939043,30.535627,29.026577,28.181509,27.411894,26.54419,24.601288,21.983086,20.447628,19.078165,18.187824,17.210714,16.105335,15.335721,15.0905,15.230087,15.543215,15.875206,16.143063,15.973294,15.482853,14.924504,14.679284,15.226315,14.154889,13.894578,13.766309,13.58145,13.641812,14.286931,15.230087,16.003475,15.70921,12.985375,0.24899325,0.59607476,0.55080324,0.452715,0.40367088,0.26408374,0.12826926,0.10940613,0.15467763,0.241448,0.3772625,0.41121614,0.4376245,0.95447415,1.9164935,2.746471,1.7089992,1.5769572,2.082489,2.8822856,3.5538127,3.8178966,5.4438977,7.3188925,8.707218,9.258021,7.9828744,8.416726,9.756008,10.831206,10.103089,7.967784,7.6886096,7.997965,7.937603,6.8473144,3.6443558,2.8181508,2.4522061,1.780679,1.177059,2.6408374,5.670255,5.1043615,1.4864142,1.0638802,1.0676528,0.7997965,0.59230214,0.49044126,0.26031113,0.44894236,0.97710985,1.1280149,0.87147635,0.8337501,0.5357128,0.97710985,1.1431054,0.84129536,0.6752999,0.9280658,1.3732355,2.8936033,4.561104,3.6443558,1.5882751,0.6451189,0.35462674,0.32067314,0.23390275,0.2565385,0.2263575,0.18863125,0.32821837,0.9922004,0.94692886,0.8903395,0.95824677,1.0827434,0.97333723,1.2336484,1.5769572,1.4071891,0.8224323,0.6149379,0.7394345,0.8337501,0.90920264,0.935611,0.8526133,0.70170826,0.543258,0.47535074,0.45648763,0.3169005,0.30935526,0.5885295,0.6187105,0.32444575,0.09808825,0.071679875,0.09808825,0.10940613,0.07922512,0.03772625,0.03772625,0.02263575,0.033953626,0.06413463,0.071679875,0.23013012,0.5281675,0.8186596,1.0110635,1.0525624,0.8111144,0.56212115,0.2678564,0.041498873,0.116951376,0.124496624,0.07922512,0.030181,0.00754525,0.026408374,0.018863125,0.02263575,0.030181,0.026408374,0.00754525,0.011317875,0.033953626,0.060362,0.060362,0.011317875,0.0150905,0.02263575,0.018863125,0.018863125,0.0452715,0.06790725,0.056589376,0.06790725,0.116951376,0.14335975,0.090543,0.041498873,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.0452715,0.18863125,0.6790725,1.0072908,0.8978847,0.44894236,0.124496624,0.10186087,0.094315626,0.17354076,0.29803738,0.331991,0.4979865,0.90543,1.1544232,1.086516,0.76207024,0.5281675,0.38103512,0.331991,0.36971724,0.47157812,0.3470815,0.26031113,0.22258487,0.17731337,0.0,0.041498873,0.05281675,0.11317875,0.211267,0.24522063,0.30935526,0.34330887,0.36971724,0.362172,0.241448,0.38858038,0.45648763,0.59607476,0.724344,0.5055317,0.452715,0.5696664,0.5281675,0.3055826,0.19240387,0.20749438,0.18863125,0.11317875,0.06790725,0.23390275,0.41498876,0.33576363,0.26031113,0.2678564,0.26408374,0.17354076,0.3772625,0.62625575,0.9280658,1.5354583,1.1355602,1.026154,1.1016065,1.2525115,1.3430545,1.2826926,1.1883769,1.4562333,1.9051756,1.7655885,1.4750963,1.2261031,0.8563859,0.392353,0.049044125,0.0452715,0.033953626,0.026408374,0.056589376,0.1659955,0.071679875,0.5772116,0.7432071,0.44139713,0.38103512,0.1358145,0.86770374,1.4109617,1.3204187,0.87147635,0.2678564,0.090543,0.0452715,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.003772625,0.0150905,0.041498873,0.056589376,0.033953626,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.049044125,0.030181,0.011317875,0.00754525,0.026408374,0.090543,0.14713238,0.150905,0.13204187,0.124496624,0.17731337,0.24522063,0.1961765,0.16222288,0.17731337,0.16976812,0.3772625,1.5467763,2.252257,2.04099,1.4449154,0.7582976,0.38480774,0.22258487,0.17354076,0.15467763,0.1659955,0.17731337,0.181086,0.17354076,0.17731337,0.15845025,0.10940613,0.05281675,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.011317875,0.030181,0.06413463,0.1056335,0.19994913,0.3470815,0.59607476,0.95447415,1.3996439,1.8146327,2.1541688,2.4710693,2.746471,2.9086938,3.0256453,3.270866,3.6707642,4.22534,4.9044123,5.764571,7.111398,8.6732645,10.370946,12.332711,14.966003,17.674747,20.319359,23.4695,28.400322,34.64779,43.09847,52.333855,60.758125,66.58306,68.642914,69.521935,71.04984,73.38133,75.003555,75.58077,75.40723,74.50557,72.99652,71.129074,70.47641,69.35594,66.61701,62.54635,58.845406,57.449535,57.811707,58.905766,60.644947,63.88563,67.31495,66.40575,61.15048,53.77877,48.757404,47.429443,47.621845,48.44428,49.25539,49.689243,49.15353,49.5572,49.889194,49.52702,48.229237,45.422405,43.05697,41.31402,40.506676,41.087658,41.400787,43.41914,46.331608,49.530792,52.616802,54.4088,54.835106,54.2428,52.937473,51.205837,50.817257,48.83663,47.2144,46.467422,45.652534,44.852737,43.728497,42.619343,41.96668,42.28358,41.057476,40.091686,39.069305,37.74134,35.93048,34.42143,32.399303,31.161882,31.048704,31.459919,31.629688,32.746384,34.61006,36.998135,39.66538,42.211903,42.3364,40.05773,36.33038,33.036877,31.003431,29.996141,29.913143,30.78462,32.802975,35.65885,38.793903,42.117584,45.022507,46.39574,45.50163,44.649017,42.75893,40.05396,38.07333,36.986816,37.341442,38.050697,38.73354,39.703106,40.235046,41.04616,41.098976,39.963417,37.809246,37.190536,36.752914,36.149292,35.40986,34.972233,36.111565,36.579372,36.54919,36.258698,36.00216,34.91942,34.693058,34.55347,33.719723,31.392014,30.486582,28.909626,26.97804,25.329405,24.914415,23.020557,21.1682,20.172226,19.73083,18.421728,18.131235,17.686066,17.440845,17.56157,18.03692,18.470772,17.742655,17.093763,16.818363,16.252468,15.539442,15.584714,15.90916,16.033657,15.460217,15.882751,16.859861,16.886269,15.679029,14.219024,0.116951376,0.2565385,0.21881226,0.14713238,0.1056335,0.090543,0.060362,0.049044125,0.056589376,0.08299775,0.150905,0.181086,0.14713238,0.29049212,0.6149379,0.8865669,0.56589377,0.5281675,0.77716076,1.1808317,1.4562333,1.4977322,2.2220762,3.1954134,4.168751,5.100589,5.50426,6.5756855,8.047009,9.514561,10.484125,9.510788,9.035437,9.175024,9.431562,8.6732645,5.485397,4.112161,3.2520027,2.3277097,1.4864142,2.4559789,4.398881,4.063117,1.6750455,0.9393836,0.965792,0.6526641,0.4979865,0.59230214,0.6375736,0.5281675,0.6752999,0.62248313,0.45648763,0.7922512,1.1921495,1.3770081,1.7467253,2.1994405,2.1277604,1.9391292,2.41448,3.802806,5.1345425,4.244203,1.871222,0.7054809,0.26031113,0.18485862,0.24899325,0.5055317,0.5470306,0.33953625,0.1659955,0.65643674,1.2411937,1.1619685,1.1695137,1.3770081,1.2562841,1.146878,1.2525115,1.2449663,1.0676528,0.965792,0.9280658,0.8941121,0.9808825,1.0412445,0.6451189,0.513077,0.52439487,0.5470306,0.56212115,0.6413463,0.33953625,0.5017591,0.7092535,0.7205714,0.4640329,0.4376245,0.30181,0.181086,0.11317875,0.056589376,0.056589376,0.030181,0.018863125,0.026408374,0.026408374,0.12826926,0.34330887,0.5583485,0.67152727,0.6187105,0.4979865,0.35839936,0.18485862,0.033953626,0.056589376,0.10940613,0.06413463,0.03772625,0.060362,0.08677038,0.06413463,0.03772625,0.018863125,0.011317875,0.0,0.003772625,0.018863125,0.030181,0.030181,0.00754525,0.00754525,0.011317875,0.011317875,0.00754525,0.018863125,0.030181,0.033953626,0.094315626,0.211267,0.3055826,0.22258487,0.124496624,0.049044125,0.018863125,0.026408374,0.011317875,0.003772625,0.0,0.011317875,0.056589376,0.26408374,0.47157812,0.482896,0.30181,0.116951376,0.11317875,0.10186087,0.09808825,0.116951376,0.13958712,0.3055826,0.5394854,0.72811663,0.77716076,0.62248313,0.40367088,0.25276586,0.1961765,0.21881226,0.29426476,0.29049212,0.29426476,0.2678564,0.19240387,0.056589376,0.018863125,0.026408374,0.049044125,0.06790725,0.071679875,0.1358145,0.17354076,0.15467763,0.10186087,0.090543,0.181086,0.18863125,0.2565385,0.36594462,0.32444575,0.48666862,0.7092535,0.60362,0.34330887,0.6375736,0.271629,0.2565385,0.18485862,0.03772625,0.18863125,0.41498876,0.49044126,0.43007925,0.29049212,0.150905,0.17731337,0.26408374,0.38480774,0.6451189,1.297783,1.026154,0.7469798,0.6526641,0.8337501,1.2487389,1.0487897,0.7809334,0.8941121,1.3091009,1.3958713,1.3619176,1.1581959,0.8262049,0.5017591,0.43007925,0.39989826,0.29426476,0.1358145,0.0150905,0.06790725,0.31312788,0.3470815,0.26031113,0.21881226,0.4640329,0.094315626,0.8601585,1.1016065,0.55457586,0.35839936,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.0150905,0.018863125,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.03772625,0.08677038,0.124496624,0.10186087,0.060362,0.033953626,0.056589376,0.0754525,0.08299775,0.08299775,0.09808825,0.1659955,0.24522063,0.23767537,0.21503963,0.2565385,0.45648763,0.633801,1.1280149,1.750498,2.2296214,2.1956677,1.0902886,0.8224323,0.73566186,0.5093044,0.18485862,0.16976812,0.16976812,0.16976812,0.1659955,0.17354076,0.16976812,0.14335975,0.09808825,0.0452715,0.018863125,0.003772625,0.0,0.0,0.0,0.00754525,0.0,0.00754525,0.018863125,0.033953626,0.06413463,0.116951376,0.22258487,0.392353,0.6488915,1.0186088,1.4864142,1.9881734,2.5201135,3.059599,3.5462675,3.5990841,3.6481283,3.7990334,4.104616,4.561104,5.1798143,6.0512905,7.1340337,8.416726,9.9257765,12.113899,14.600059,17.014538,19.447882,22.4358,26.597006,32.16163,39.00517,46.354244,52.794113,57.823025,62.376583,65.58331,67.541306,69.337074,71.449745,73.50583,74.04908,72.78148,70.54809,66.84337,64.61752,62.927383,61.214615,59.316982,55.310455,52.480988,51.892456,53.888176,58.08711,62.135136,62.999065,60.599674,55.84994,50.681446,47.176674,45.086643,44.479248,44.97346,45.758167,45.53181,46.331608,47.6143,48.74986,49.02526,48.13115,45.81476,43.1626,40.982025,39.80874,38.74863,38.77504,39.970963,42.35903,45.897755,49.65529,52.779022,55.04637,56.159294,55.740536,53.903267,50.960617,48.878128,48.078335,47.448303,46.06375,44.592426,43.2041,42.30999,42.547665,42.14022,41.72146,41.359287,40.77076,39.352253,37.99788,36.24738,34.8666,34.112076,33.708405,33.244373,33.07083,33.255688,34.142258,36.34547,40.695305,43.845448,45.51672,45.611034,44.234028,41.91009,37.696068,33.599,30.773302,29.494383,29.93578,31.433512,34.24789,37.8432,40.9028,42.9702,44.686745,45.124367,44.17744,42.547665,40.280315,39.027805,37.386715,35.5419,35.243862,36.386967,37.017,38.29969,39.733288,39.14853,38.888218,37.979015,36.556736,34.945824,33.67445,33.632954,33.436775,33.202873,32.776566,31.727776,31.595734,31.701368,32.53512,33.58768,33.31228,32.46721,31.478783,30.701622,30.343224,30.445084,27.698612,25.42372,23.952396,22.8357,20.8513,20.289177,19.678013,19.134754,18.787672,18.757492,19.893051,20.206179,19.870417,19.017803,17.772837,17.772837,17.689838,17.53516,17.297485,16.976812,17.901106,18.595268,18.874443,19.134754,20.33822,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0150905,0.018863125,0.0150905,0.00754525,0.00754525,0.241448,0.23013012,0.17354076,0.19240387,0.31312788,0.29426476,0.2565385,0.3772625,0.8903395,2.0787163,2.565385,3.2821836,4.353609,5.802297,7.5603404,9.06939,9.322156,9.163706,8.918486,8.405409,6.519096,5.715527,4.768598,3.3538637,2.04099,1.9089483,2.2786655,2.263575,1.6410918,0.86770374,0.724344,0.49044126,0.43007925,0.56589377,0.66775465,0.49421388,0.5583485,0.6111652,0.6413463,0.88279426,1.388326,1.5128226,2.0560806,2.8898308,2.957738,2.372981,2.6068838,3.4972234,4.5196047,4.8063245,3.610402,2.3918443,1.3920987,0.7394345,0.4640329,0.7167987,0.7507524,0.45648763,0.116951376,0.392353,1.2147852,1.2525115,1.2638294,1.50905,1.7693611,2.033445,2.41448,2.493705,2.2183034,1.9278114,1.5505489,1.4260522,1.3845534,1.1996948,0.59607476,0.66775465,0.76207024,0.6488915,0.47157812,0.76207024,0.573439,0.6375736,0.724344,0.7809334,0.94692886,1.086516,0.8111144,0.46026024,0.21503963,0.120724,0.10186087,0.10186087,0.071679875,0.026408374,0.05281675,0.09808825,0.23013012,0.331991,0.33576363,0.211267,0.21881226,0.18485862,0.11317875,0.03772625,0.0,0.12826926,0.071679875,0.030181,0.060362,0.071679875,0.06790725,0.033953626,0.003772625,0.003772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.018863125,0.02263575,0.08299775,0.18485862,0.2678564,0.26408374,0.18485862,0.08677038,0.02263575,0.033953626,0.018863125,0.00754525,0.0,0.0,0.00754525,0.071679875,0.17731337,0.271629,0.3055826,0.23013012,0.15467763,0.1056335,0.05281675,0.003772625,0.018863125,0.12826926,0.19240387,0.27917424,0.38103512,0.4074435,0.23767537,0.13958712,0.094315626,0.10186087,0.150905,0.21881226,0.2678564,0.2678564,0.211267,0.12826926,0.0754525,0.071679875,0.049044125,0.003772625,0.0,0.0452715,0.056589376,0.03772625,0.033953626,0.120724,0.12826926,0.08677038,0.10940613,0.21503963,0.32444575,0.452715,0.6488915,0.573439,0.4678055,1.1883769,0.513077,0.55457586,0.5394854,0.2678564,0.10940613,0.24899325,0.39989826,0.42630664,0.31312788,0.150905,0.181086,0.181086,0.21881226,0.38103512,0.7582976,0.90543,0.60362,0.38858038,0.5017591,0.8865669,0.7054809,0.5281675,0.543258,0.7507524,0.9507015,1.056335,0.8941121,0.573439,0.331991,0.5281675,0.5772116,0.55457586,0.3961256,0.1659955,0.07922512,0.41498876,0.19994913,0.018863125,0.09808825,0.31312788,0.09808825,0.62248313,0.60362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.041498873,0.08677038,0.124496624,0.10940613,0.08299775,0.06790725,0.056589376,0.03772625,0.030181,0.03772625,0.06413463,0.120724,0.17731337,0.20749438,0.23767537,0.31312788,0.513077,0.7130261,0.6375736,0.88279426,1.4562333,1.7693611,0.9808825,0.80734175,0.7394345,0.5357128,0.211267,0.15467763,0.13204187,0.13204187,0.1358145,0.150905,0.15467763,0.150905,0.120724,0.0754525,0.041498873,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.033953626,0.05281675,0.116951376,0.21503963,0.362172,0.5998474,0.97710985,1.4675511,2.0673985,2.746471,3.4783602,3.783943,3.9650288,4.115934,4.3121104,4.606375,5.0439997,5.5570765,6.1908774,6.9869013,8.024373,9.601331,11.5857315,13.754991,15.965749,18.16519,21.187061,24.963459,29.679241,34.92319,39.657833,45.25641,51.183205,56.042343,59.509388,62.3464,65.93794,68.55237,69.68416,69.3484,68.099655,64.210075,62.006863,60.942986,60.67513,61.067482,58.75109,54.778515,51.78305,51.024754,52.394215,53.597683,54.374844,55.008644,54.737015,51.771732,48.76495,45.64876,43.739815,43.253147,43.309734,42.81552,43.1626,44.173668,45.422405,46.256157,47.244583,46.324062,44.762196,43.17392,41.525284,39.631424,38.265736,37.552708,37.831882,39.63897,42.947563,46.84091,50.907803,54.35598,56.03857,55.023735,53.122334,51.541603,50.65881,50.006145,48.240555,46.55042,44.788605,43.23051,42.558983,42.219448,41.683735,41.23479,40.778305,39.85401,38.684498,37.232037,36.115337,35.44004,34.77606,34.368614,33.610317,32.814293,32.516254,33.50091,36.669914,39.9106,43.321053,46.49006,48.497093,49.11958,46.32029,42.15154,37.6093,32.62566,29.550972,28.01174,28.577635,30.894026,33.693314,36.220974,39.284344,41.63469,42.932472,43.743587,42.898518,41.672417,39.16362,35.9418,34.070576,33.670677,33.71595,35.142002,37.318806,38.035606,37.601753,37.952606,37.552708,36.066296,34.372387,33.80649,33.21419,32.49739,31.38824,29.44911,29.63397,29.083166,29.366114,30.663897,31.807001,31.59196,31.671186,32.040905,32.5238,32.776566,30.871391,29.309525,28.072104,26.58946,23.75622,22.790428,21.835953,20.994658,20.345766,19.957186,20.8513,21.60205,21.368149,20.115637,18.648085,18.885761,18.94235,18.731083,18.414183,18.43682,19.496925,19.972277,20.990885,23.654358,29.022804,0.00754525,0.003772625,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.026408374,0.033953626,0.041498873,0.026408374,0.056589376,0.16976812,0.33953625,0.73188925,1.7127718,0.98465514,0.7130261,0.935611,1.8259505,3.682082,6.7756343,8.001738,7.677292,6.7114997,6.598321,5.934339,6.039973,5.4476705,4.006528,2.9086938,1.8863125,1.418507,1.3619176,1.388326,0.9808825,0.56589377,0.41876137,0.3961256,0.40367088,0.392353,0.33576363,0.44516975,0.67152727,0.875249,0.80734175,0.8262049,1.2261031,1.9240388,2.6898816,3.1463692,2.4672968,2.3428001,2.7238352,3.7047176,5.5193505,6.488915,5.6023483,3.8292143,2.071171,1.1581959,1.1846043,0.97710985,0.573439,0.2263575,0.41876137,1.0186088,1.478869,1.6863633,1.7995421,2.2673476,3.0520537,3.9386206,4.146115,3.663219,3.2482302,2.6219745,2.4031622,2.1277604,1.6712729,1.2223305,1.4298248,1.358145,0.86770374,0.331991,0.62248313,0.9242931,1.0978339,0.91674787,0.694163,1.2826926,1.7542707,1.6675003,1.1204696,0.44894236,0.19994913,0.150905,0.1961765,0.16222288,0.06413463,0.094315626,0.124496624,0.24899325,0.29426476,0.23013012,0.15467763,0.1659955,0.14713238,0.094315626,0.033953626,0.0,0.15467763,0.094315626,0.0150905,0.003772625,0.0150905,0.02263575,0.02263575,0.011317875,0.011317875,0.049044125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.06790725,0.02263575,0.003772625,0.0,0.003772625,0.02263575,0.17354076,0.211267,0.13958712,0.030181,0.018863125,0.0150905,0.003772625,0.0,0.0,0.0,0.02263575,0.1056335,0.25276586,0.39989826,0.38858038,0.18863125,0.0754525,0.018863125,0.003772625,0.0,0.0,0.00754525,0.026408374,0.07922512,0.1961765,0.08677038,0.049044125,0.030181,0.030181,0.071679875,0.124496624,0.18863125,0.23390275,0.241448,0.19994913,0.16222288,0.13958712,0.08677038,0.018863125,0.003772625,0.0,0.0,0.011317875,0.030181,0.060362,0.10186087,0.17731337,0.19240387,0.15467763,0.20372175,0.15845025,0.26408374,0.331991,0.5281675,1.3505998,0.6451189,0.7469798,0.94315624,0.8111144,0.21503963,0.2263575,0.2678564,0.32444575,0.3470815,0.2678564,0.26031113,0.27917424,0.2678564,0.21503963,0.181086,0.8224323,0.754525,0.543258,0.47535074,0.56589377,0.8111144,0.87902164,0.73188925,0.543258,0.7092535,0.58475685,0.47535074,0.25276586,0.03772625,0.1961765,0.35085413,0.52062225,0.51684964,0.34330887,0.1961765,0.271629,0.17354076,0.1358145,0.17731337,0.07922512,0.15467763,0.30181,0.23390275,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.056589376,0.030181,0.02263575,0.05281675,0.090543,0.071679875,0.033953626,0.011317875,0.003772625,0.0150905,0.02263575,0.03772625,0.09808825,0.19994913,0.29803738,0.2867195,0.5055317,0.52062225,0.44516975,0.40367088,0.52062225,0.5281675,0.362172,0.23390275,0.21503963,0.2263575,0.15845025,0.10940613,0.090543,0.10186087,0.120724,0.1358145,0.14335975,0.13204187,0.1056335,0.07922512,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.060362,0.11317875,0.1961765,0.3169005,0.5281675,0.845068,1.297783,1.8825399,2.5691576,3.229367,3.7537618,4.146115,4.4441524,4.7044635,5.0553174,5.4401255,5.87775,6.398372,7.020855,7.967784,9.265567,10.8576145,12.679792,14.641558,16.859861,20.006231,23.839218,27.864609,31.339195,35.247635,39.156075,44.117077,49.61002,53.529778,57.683437,59.58484,60.95053,62.425625,63.56496,63.919586,63.474415,61.976685,60.38841,60.90526,62.455807,60.056416,56.261158,52.64698,49.79865,46.44856,45.045143,46.561737,49.361027,49.198803,48.61027,46.5806,45.02628,44.332115,43.351234,42.177948,41.41588,41.083885,41.095203,41.27629,43.023014,43.909584,44.471703,44.660336,43.837902,41.845955,40.231274,38.495865,36.817047,36.07007,37.330124,39.684242,43.279552,47.561485,51.29261,53.571274,54.4503,54.476704,54.0504,53.412827,51.749096,50.183456,48.39146,46.471195,44.943283,43.660587,42.521255,41.51774,40.578354,39.540882,38.04315,36.383194,35.364586,35.047688,34.745876,34.670425,34.03285,33.391502,33.104786,33.30096,33.68954,34.598743,36.398285,39.273026,43.23051,47.5728,49.745834,49.617565,46.889957,41.10275,35.88898,31.569326,29.124664,28.551226,28.856808,29.501928,31.67496,33.798946,35.76071,38.884445,40.89903,41.14802,40.208637,38.609043,36.851,34.172436,33.568817,33.753677,34.161118,34.949596,33.719723,35.81353,37.371624,36.930225,35.40986,35.198593,34.64779,33.565044,32.04845,30.475266,30.607307,29.252934,28.057013,27.826881,28.532362,29.094484,29.833918,30.584671,31.207153,31.58819,32.055996,31.822092,31.354286,30.241362,27.189308,25.736847,24.473019,23.431774,22.662159,22.232079,22.326395,22.503708,22.013268,20.760756,19.319613,19.01403,19.270569,19.410156,19.312067,19.40261,20.085455,20.526854,22.167944,26.566826,35.417404,0.0452715,0.02263575,0.00754525,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.10940613,0.150905,0.124496624,0.0150905,0.0150905,0.02263575,0.041498873,0.0754525,0.1358145,0.211267,0.29426476,0.63002837,1.2638294,2.0447628,1.9957186,2.003264,2.5993385,3.7047176,4.610148,3.9725742,3.3123648,2.7313805,2.674791,3.9197574,2.8596497,1.9353566,1.1883769,0.7092535,0.62625575,0.41876137,0.32067314,0.39989826,0.663982,1.0525624,0.8224323,0.56212115,0.60362,0.8186596,0.6111652,0.56212115,0.9507015,1.7580433,2.8898308,4.195159,3.6330378,4.3083377,5.070408,5.666483,6.730363,8.29223,8.314865,6.458734,3.7914882,2.7917426,2.8785129,2.1956677,1.3204187,0.73566186,0.80734175,1.6146835,2.7879698,3.2029586,2.6597006,1.8749946,1.3996439,1.6222287,2.4371157,3.482133,4.104616,3.7990334,3.1463692,2.7087448,2.6597006,2.806833,2.8181508,2.2107582,1.2826926,0.52439487,0.6111652,1.2940104,1.841041,1.8334957,1.3920987,1.1581959,2.0636258,2.9011486,2.425798,0.90543,0.1358145,0.10186087,0.14713238,0.150905,0.094315626,0.0452715,0.1056335,0.331991,0.36971724,0.21503963,0.23013012,0.19240387,0.1659955,0.1056335,0.02263575,0.0,0.0,0.0,0.0,0.0150905,0.0754525,0.0150905,0.06413463,0.06413463,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.090543,0.018863125,0.0,0.0,0.0,0.0,0.060362,0.26031113,0.29426476,0.13958712,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.124496624,0.26408374,0.35085413,0.19240387,0.07922512,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.033953626,0.0452715,0.071679875,0.120724,0.17731337,0.22258487,0.26031113,0.22258487,0.21503963,0.14713238,0.041498873,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.30181,0.32067314,0.071679875,0.1659955,0.033953626,0.03772625,0.06790725,0.15467763,0.47157812,0.30181,0.23013012,0.8299775,1.6222287,1.0827434,1.1317875,0.79602385,0.4376245,0.2678564,0.36594462,0.6111652,0.7167987,0.7054809,0.694163,0.9016574,0.694163,0.6790725,0.69039035,0.663982,0.62625575,1.2713746,1.2525115,0.8978847,0.5281675,0.44139713,0.44139713,0.34330887,0.1659955,0.0,0.0,0.0,0.0,0.0,0.03772625,0.18485862,0.23013012,0.3734899,0.5055317,0.543258,0.3961256,0.43385187,0.35085413,0.17354076,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.030181,0.00754525,0.0,0.018863125,0.0452715,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.011317875,0.07922512,0.15845025,0.19994913,0.150905,0.12826926,0.1659955,0.16222288,0.1056335,0.1056335,0.19240387,0.17731337,0.1056335,0.06790725,0.21503963,0.21503963,0.13204187,0.071679875,0.071679875,0.1056335,0.14335975,0.16976812,0.18485862,0.17731337,0.150905,0.1056335,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.056589376,0.10940613,0.18485862,0.3169005,0.4979865,0.77716076,1.177059,1.6788181,2.2899833,2.916239,3.5236318,4.0593443,4.485651,4.8629136,5.2326307,5.624984,6.043745,6.470052,6.971811,7.6282477,8.488406,9.623966,11.140562,13.091009,15.513034,18.440592,21.794455,25.344494,28.777584,31.757957,34.859055,38.10351,40.970707,45.037598,48.37637,52.03959,56.58183,62.089863,67.96007,69.84638,67.54885,63.22542,61.433426,60.773216,59.965874,58.143696,55.182186,51.72646,46.89373,43.185238,41.95159,43.132423,45.241318,44.362297,43.73227,43.89072,44.18121,42.74007,41.468693,39.688015,37.892246,36.930225,37.979015,39.835148,40.38218,40.31427,40.408585,41.51774,41.76296,40.853756,39.39375,37.745113,36.009705,36.205883,36.66614,37.937515,40.608536,45.335636,49.900513,53.5675,55.680172,56.53656,57.404263,56.415833,55.076553,53.541096,51.888683,50.15705,47.79916,46.73528,46.339153,45.682716,43.53232,40.38218,38.26951,36.424694,34.96846,34.88169,35.236317,34.745876,34.428974,34.557243,34.666653,34.37616,34.281845,33.995125,33.949852,35.417404,38.578865,41.80446,45.241318,48.22169,49.27048,46.644737,41.55924,36.021023,31.226017,27.525072,27.528845,27.728794,28.230553,29.388748,31.829638,35.100502,36.681232,38.522274,40.57458,40.75567,38.303463,35.719215,33.40282,31.776821,31.312788,30.335678,31.47501,33.463184,35.092957,35.202362,34.73833,33.734814,32.42194,31.109066,30.181,31.278833,30.878935,29.754694,28.788902,28.947351,29.226526,29.252934,29.264252,29.56229,30.501673,32.55398,32.587936,31.90509,31.109066,30.120638,28.132465,27.559025,26.895044,25.79721,25.099274,25.661396,25.344494,24.552244,23.420456,21.835953,20.406128,19.80251,19.308294,18.806536,18.76881,19.353567,19.794964,21.251196,24.944597,32.13522,0.52062225,0.362172,0.24522063,0.3734899,0.513077,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.00754525,0.02263575,0.060362,0.094315626,0.06413463,0.0150905,0.026408374,0.060362,0.094315626,0.124496624,0.150905,0.15467763,0.1961765,0.3055826,0.47157812,0.6149379,0.9205205,1.3053282,1.7316349,2.214531,2.7917426,2.9728284,2.727608,2.3428001,2.444661,1.9391292,1.5203679,1.086516,0.694163,0.5394854,0.3734899,0.38480774,0.5885295,0.84129536,0.87147635,1.9089483,1.0714256,0.29049212,0.23013012,0.3055826,0.9393836,1.0902886,1.418507,1.9051756,1.8636768,4.6818275,5.138315,5.451443,6.168242,6.168242,5.7004366,5.9682927,6.145606,5.772116,4.7836885,5.80607,5.194905,4.244203,3.500996,2.7728794,2.9841464,3.2369123,3.4481792,3.3425457,2.463524,1.9768555,2.003264,2.3616633,2.7653341,2.8219235,3.1614597,3.5349495,3.9197574,4.0291634,3.308592,2.323937,1.539231,0.9922004,0.724344,0.7696155,1.2298758,1.9240388,2.384299,2.293756,1.4637785,1.0299267,1.388326,1.4750963,0.9507015,0.211267,0.18485862,0.23013012,0.31312788,0.3772625,0.38858038,0.271629,0.2867195,0.27917424,0.20372175,0.1056335,0.2263575,0.3169005,0.23013012,0.02263575,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.041498873,0.041498873,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.00754525,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.08677038,0.1358145,0.11317875,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.011317875,0.018863125,0.056589376,0.13204187,0.23013012,0.12826926,0.08299775,0.060362,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.02263575,0.026408374,0.05281675,0.090543,0.14335975,0.211267,0.241448,0.21503963,0.120724,0.030181,0.06413463,0.23767537,0.25276586,0.13958712,0.0,0.0,0.0,0.060362,0.08677038,0.06413463,0.033953626,0.0452715,0.08677038,0.18485862,0.27917424,0.20372175,0.20749438,0.41121614,0.77338815,1.146878,1.2525115,1.7731338,1.2525115,0.63002837,0.33953625,0.32821837,0.38858038,0.5017591,0.5319401,0.52439487,0.694163,0.6526641,0.5470306,0.44516975,0.36594462,0.26031113,0.84884065,0.8639311,0.6111652,0.331991,0.19994913,0.21881226,0.32821837,0.23767537,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.18485862,0.331991,0.39989826,0.3772625,0.3470815,0.27540162,0.18863125,0.08677038,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.094315626,0.3772625,0.0754525,0.0,0.0,0.00754525,0.03772625,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.049044125,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.030181,0.05281675,0.049044125,0.030181,0.056589376,0.1056335,0.116951376,0.08299775,0.094315626,0.20749438,0.19994913,0.13204187,0.08299775,0.150905,0.19994913,0.17354076,0.12826926,0.09808825,0.1056335,0.11317875,0.19240387,0.271629,0.30181,0.23767537,0.16976812,0.14335975,0.116951376,0.071679875,0.02263575,0.003772625,0.00754525,0.011317875,0.011317875,0.0,0.003772625,0.011317875,0.02263575,0.041498873,0.08677038,0.16976812,0.29426476,0.48666862,0.76584285,1.1280149,1.6033657,2.1692593,2.7917426,3.4330888,4.032936,4.5799665,5.093044,5.5759397,6.0286546,6.4436436,6.749226,7.073672,7.4999785,8.09228,8.892077,10.26154,11.917723,13.853079,16.06761,18.595268,20.922977,23.480818,26.514008,29.849009,32.91238,35.73053,38.03938,40.751896,44.528294,49.809967,57.166588,61.278748,62.584076,62.467125,63.25183,63.187695,63.606457,64.80615,65.74554,64.06672,57.55517,50.93044,46.69378,45.18473,44.58488,43.234283,42.317535,41.638462,40.800938,39.223984,37.8847,36.54919,35.55322,35.02128,34.828873,35.319317,35.692806,36.322834,37.40935,38.97876,39.499382,39.75592,39.295662,38.14124,36.77932,36.594463,37.620617,38.337414,38.79013,40.57458,42.951336,46.365562,50.17214,53.959854,57.551395,58.758633,58.901993,58.40778,57.54385,56.415833,53.601456,51.40579,49.87033,48.685726,47.169132,46.06375,44.15103,41.72146,39.36734,37.994106,37.360306,37.39426,37.907337,38.435505,38.2431,37.356533,36.164383,35.183502,34.727013,34.904327,36.092705,37.805473,39.92569,42.238308,44.460384,45.995846,46.20334,44.335888,40.567036,35.998386,31.867363,29.20389,28.151327,28.362595,28.996395,30.705395,31.682505,32.474754,33.62541,35.65508,36.813274,37.088676,36.424694,35.013733,33.289642,31.71646,31.41842,31.105293,30.74312,31.51651,33.433002,34.285618,34.183754,32.87088,29.705648,28.890762,28.558771,28.728539,29.20389,29.569836,29.66415,29.400066,29.007713,28.803991,29.207663,29.716967,30.509218,31.59196,32.606796,32.818066,31.267515,29.268024,28.019285,27.498663,26.480055,26.483828,26.585688,26.642279,26.185791,24.423975,22.654613,21.03993,19.57615,18.52736,18.463226,18.395319,18.391546,19.47429,21.383238,22.57916,1.327964,1.1695137,0.91297525,0.66775465,0.44516975,0.14335975,0.049044125,0.094315626,0.10940613,0.056589376,0.026408374,0.033953626,0.116951376,0.10186087,0.003772625,0.018863125,0.011317875,0.026408374,0.1056335,0.181086,0.056589376,0.041498873,0.08677038,0.24899325,0.44516975,0.422534,0.29049212,0.19994913,0.21503963,0.2867195,0.241448,0.45648763,0.52439487,0.60362,0.98465514,2.0749438,2.1843498,2.5238862,2.6182017,2.3692086,2.0372176,1.7014539,1.3619176,0.98842776,0.6375736,0.44516975,0.32444575,0.29803738,0.35462674,0.4376245,0.44894236,1.2336484,0.9507015,0.4979865,0.29803738,0.27540162,0.814887,1.1280149,1.4637785,1.9768555,2.7200627,5.070408,5.745708,5.956975,6.4474163,7.4735703,8.386545,8.560086,8.088508,6.828451,4.38379,4.6742826,4.0593443,3.2520027,2.655928,2.3503454,2.1315331,2.0862615,3.482133,5.511805,5.281675,5.0062733,4.221567,3.519859,3.1425967,2.9766011,3.5953116,3.308592,3.169005,3.308592,2.9464202,3.3840446,2.3956168,1.3619176,0.8941121,0.8262049,1.267602,2.2107582,2.7879698,2.5578396,1.5241405,1.0035182,1.2638294,1.3317367,0.88279426,0.23767537,0.3169005,0.41121614,0.452715,0.43007925,0.4074435,0.331991,0.3169005,0.30181,0.24522063,0.13204187,0.120724,0.15845025,0.124496624,0.03772625,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.026408374,0.0,0.0,0.0,0.0,0.0150905,0.030181,0.00754525,0.0,0.0,0.0452715,0.08677038,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.060362,0.090543,0.03772625,0.030181,0.011317875,0.02263575,0.0452715,0.00754525,0.00754525,0.00754525,0.02263575,0.0754525,0.181086,0.18863125,0.13204187,0.06790725,0.02263575,0.018863125,0.011317875,0.003772625,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0150905,0.033953626,0.0754525,0.124496624,0.18863125,0.21503963,0.1358145,0.026408374,0.1056335,0.44139713,0.4376245,0.30181,0.21503963,0.33953625,0.362172,0.21881226,0.08299775,0.0452715,0.10186087,0.150905,0.15467763,0.14713238,0.124496624,0.056589376,0.0754525,0.25276586,0.41121614,0.482896,0.52062225,0.9280658,0.7507524,0.44139713,0.2867195,0.41121614,0.32067314,0.24522063,0.2867195,0.44139713,0.5772116,0.4376245,0.26408374,0.20372175,0.2565385,0.24899325,0.43007925,0.35462674,0.31312788,0.31312788,0.056589376,0.06413463,0.12826926,0.10186087,0.0,0.0,0.0,0.0,0.056589376,0.10940613,0.0,0.06790725,0.35085413,0.47157812,0.36971724,0.27917424,0.124496624,0.060362,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05281675,0.1358145,0.17354076,0.033953626,0.0,0.0,0.0,0.0,0.02263575,0.056589376,0.049044125,0.10186087,0.45648763,0.38480774,0.18485862,0.20749438,0.38103512,0.21881226,0.211267,0.14713238,0.0754525,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.011317875,0.003772625,0.00754525,0.02263575,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.011317875,0.02263575,0.018863125,0.0,0.02263575,0.071679875,0.090543,0.06413463,0.0452715,0.094315626,0.14335975,0.150905,0.124496624,0.10186087,0.15467763,0.1961765,0.21503963,0.20749438,0.16976812,0.16222288,0.18863125,0.20372175,0.19994913,0.18485862,0.15845025,0.16222288,0.16976812,0.15845025,0.11317875,0.08677038,0.05281675,0.02263575,0.003772625,0.0,0.0,0.003772625,0.00754525,0.011317875,0.033953626,0.071679875,0.14335975,0.26408374,0.4376245,0.6790725,1.0450171,1.5241405,2.1013522,2.7502437,3.4255435,4.093298,4.7610526,5.409944,6.006019,6.5040054,6.802043,7.3868,8.239413,9.242931,10.170997,10.484125,10.944386,11.5857315,12.468526,13.694629,15.158407,17.003222,19.312067,22.164171,25.634987,28.290915,30.4979,32.418167,34.666653,38.326096,42.762703,47.81425,52.75639,56.721416,58.70582,60.052647,61.203297,63.893177,67.13009,67.20931,62.071,56.47997,51.847187,48.81777,47.29363,45.577084,44.192528,42.45335,40.118095,37.401806,35.65885,34.659107,34.025307,33.380184,32.32008,31.788137,32.044678,33.101013,34.757195,36.632187,37.299942,37.307487,37.32258,37.696068,38.492092,37.096222,37.48103,38.782585,40.20109,40.993343,40.929207,42.4873,44.947056,48.123604,52.36781,55.465134,58.143696,60.237503,61.55415,61.863506,61.161797,59.735744,57.6193,54.853966,51.52274,50.624855,48.889446,46.81073,44.758423,43.00038,42.362804,40.936752,40.64249,41.525284,41.747868,41.412106,40.065277,38.533592,37.36785,36.86232,36.971725,37.15281,38.095966,39.661606,40.842438,42.46467,44.543385,46.00716,46.124115,44.532066,40.389725,36.141747,32.59548,30.192318,29.049213,29.00394,29.29066,29.799965,30.509218,31.47501,32.908607,34.34975,35.16841,35.145775,34.470474,32.814293,31.161882,29.716967,28.954897,29.63397,31.89,33.06706,33.21419,32.403076,30.686531,29.369886,28.732311,28.192827,27.747658,27.966469,28.34373,28.736084,29.467974,30.165909,29.747149,29.158619,29.226526,29.924461,31.093975,32.44835,32.07863,31.199608,30.230043,29.162392,27.56657,27.272306,27.336441,28.000423,28.626678,27.698612,25.182272,23.250689,21.579414,20.168453,19.349794,18.689585,17.818108,17.565342,17.855835,17.697384,1.1280149,1.7354075,2.425798,2.1994405,1.1695137,0.55080324,0.21503963,0.14335975,0.20749438,0.271629,0.17354076,0.06413463,0.11317875,0.116951376,0.049044125,0.071679875,0.026408374,0.10940613,0.2678564,0.36971724,0.19994913,0.21503963,0.24899325,0.3772625,0.51684964,0.392353,0.24899325,0.181086,0.241448,0.33576363,0.23013012,0.4376245,0.49421388,0.6413463,1.0751982,1.9768555,2.3314822,2.8634224,3.2029586,3.097325,2.4182527,2.9426475,1.931584,1.0336993,0.77716076,0.55457586,0.38103512,0.2565385,0.1659955,0.116951376,0.14335975,0.41876137,1.7089992,2.1088974,1.3317367,0.7092535,0.845068,1.1581959,1.5279131,2.0070364,2.8294687,4.496969,5.172269,5.349582,5.764571,7.3868,9.178797,9.805053,9.26934,7.488661,4.285702,3.1350515,2.4408884,1.9391292,1.5467763,1.3430545,1.0072908,0.87147635,2.142851,4.13857,4.2630663,4.217795,3.5575855,2.987919,3.078462,4.2781568,6.326692,6.5455046,5.281675,3.3953626,2.282438,3.1463692,2.4371157,1.7165444,1.4901869,1.1921495,2.1503963,2.595566,2.5201135,1.9881734,1.1317875,0.7922512,1.2110126,1.3128735,0.8601585,0.4376245,0.5357128,0.5470306,0.48666862,0.42630664,0.47535074,0.5394854,0.49421388,0.38480774,0.25276586,0.14335975,0.03772625,0.02263575,0.030181,0.033953626,0.026408374,0.003772625,0.003772625,0.003772625,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.0,0.003772625,0.003772625,0.0150905,0.030181,0.0,0.003772625,0.00754525,0.049044125,0.094315626,0.030181,0.0150905,0.018863125,0.0150905,0.00754525,0.030181,0.026408374,0.011317875,0.02263575,0.060362,0.071679875,0.056589376,0.03772625,0.041498873,0.0452715,0.00754525,0.0,0.0,0.00754525,0.041498873,0.1358145,0.3470815,0.29049212,0.15845025,0.09808825,0.21503963,0.12826926,0.041498873,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.00754525,0.033953626,0.08677038,0.11317875,0.1358145,0.08677038,0.018863125,0.08677038,0.32444575,0.31312788,0.25276586,0.29803738,0.5357128,0.482896,0.331991,0.28294688,0.34330887,0.331991,0.3772625,0.331991,0.241448,0.14335975,0.08677038,0.14713238,0.15467763,0.1358145,0.1056335,0.056589376,0.1659955,0.23013012,0.27540162,0.34330887,0.5017591,0.23390275,0.24899325,0.38103512,0.46026024,0.32067314,0.181086,0.14335975,0.211267,0.3169005,0.31312788,0.15845025,0.049044125,0.116951376,0.24522063,0.060362,0.16222288,0.2263575,0.20749438,0.124496624,0.056589376,0.011317875,0.0754525,0.26031113,0.42630664,0.27917424,0.094315626,0.31312788,0.49421388,0.43385187,0.14713238,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.18485862,0.19994913,0.0754525,0.018863125,0.0,0.0,0.0,0.026408374,0.18485862,0.3055826,0.33953625,0.38103512,0.7054809,0.6488915,0.58098423,0.55457586,0.32821837,0.47535074,0.362172,0.17354076,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.003772625,0.011317875,0.0150905,0.0,0.00754525,0.05281675,0.0754525,0.06413463,0.033953626,0.0150905,0.071679875,0.12826926,0.14335975,0.11317875,0.14335975,0.1961765,0.23390275,0.241448,0.21503963,0.19240387,0.18863125,0.17731337,0.15467763,0.150905,0.150905,0.15467763,0.15845025,0.15845025,0.124496624,0.10940613,0.13204187,0.09808825,0.0150905,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.05281675,0.10940613,0.19994913,0.331991,0.58098423,0.9318384,1.4034165,1.9806281,2.6219745,3.350091,4.13857,4.9685473,5.87775,6.960493,8.412953,10.155907,11.378237,11.744182,11.41219,10.804798,10.423763,10.295494,10.438853,10.880251,11.732863,12.872196,14.317112,16.25624,19.017803,21.330421,23.48459,25.46522,27.562798,30.39604,32.75393,37.07736,42.34017,47.104996,49.50816,50.983253,52.016953,55.050144,59.433933,61.429653,59.192486,56.540333,53.88063,51.424652,49.202576,47.406807,46.275017,45.305454,43.468185,39.19003,36.503918,35.37213,34.617607,33.60277,32.229534,31.324106,31.286379,32.029587,33.421684,35.289135,36.190792,35.836166,35.651306,36.37942,38.08465,36.915134,36.47374,37.401806,39.125893,39.842693,39.46166,40.08414,41.17066,42.82684,45.807213,48.968674,52.488533,56.359245,60.169598,63.13488,65.19473,66.16052,65.27773,62.350174,57.74757,55.627357,54.529522,52.84693,50.349453,48.176422,47.387943,45.150776,43.698315,43.40782,42.78534,43.207874,42.906063,42.374123,41.668644,40.401043,39.07685,37.78284,37.590435,38.33364,38.627907,39.069305,40.91412,43.249374,45.44127,47.146496,46.286335,43.600227,39.933235,36.08516,32.81052,30.475266,29.230299,28.977533,29.328386,29.607561,30.075367,30.901571,31.780594,32.587936,33.372643,33.161373,31.859818,30.433765,29.445337,29.04544,29.279343,29.600016,29.781101,29.856554,30.12441,29.20389,29.120892,28.664404,27.755201,27.442074,27.438301,28.464457,29.830147,30.690304,30.048958,30.184772,29.317068,29.120892,30.101774,31.61837,31.946589,32.5238,32.686024,32.01827,30.343224,29.849009,28.766266,28.649315,29.298206,28.78513,27.408121,25.665169,23.605314,21.553007,20.111864,19.327158,18.229324,17.195625,16.4826,16.218515,0.14335975,1.4939595,3.3161373,3.6368105,2.3201644,1.0638802,0.44516975,0.28294688,0.3734899,0.4678055,0.29426476,0.1056335,0.06790725,0.11317875,0.16976812,0.1358145,0.08677038,0.20372175,0.3772625,0.5055317,0.482896,0.4640329,0.41876137,0.3734899,0.29426476,0.08677038,0.060362,0.124496624,0.211267,0.26031113,0.23390275,0.452715,0.9016574,1.4449154,1.8485862,1.7995421,3.1652324,3.9386206,4.2064767,3.9197574,2.9011486,4.285702,2.535204,1.0940613,0.9922004,0.88279426,0.9620194,1.1204696,1.3468271,1.7693611,2.6483827,1.3355093,3.1237335,4.074435,3.1539145,2.252257,2.505023,2.8521044,2.7011995,2.1843498,2.161714,3.3953626,3.7575345,4.036709,4.644101,5.621211,6.598321,8.197914,9.035437,8.326183,5.885295,3.5236318,2.505023,2.0900342,1.8334957,1.5807298,1.2638294,0.77716076,0.40367088,0.24899325,0.26031113,0.422534,0.7205714,1.116697,2.1013522,4.689373,7.9489207,9.578695,8.096053,4.5837393,2.6898816,2.8898308,2.5427492,2.2786655,2.214531,1.9579924,3.0746894,2.6823363,1.8863125,1.3204187,1.1393328,0.58475685,0.935611,1.1053791,0.8262049,0.6752999,0.65643674,0.5281675,0.41876137,0.4074435,0.5357128,0.7167987,0.62248313,0.39989826,0.18485862,0.08677038,0.018863125,0.0150905,0.033953626,0.03772625,0.003772625,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.003772625,0.003772625,0.011317875,0.018863125,0.0150905,0.018863125,0.06790725,0.033953626,0.0452715,0.033953626,0.011317875,0.060362,0.05281675,0.030181,0.011317875,0.02263575,0.10940613,0.08677038,0.23767537,0.32821837,0.2678564,0.10186087,0.030181,0.003772625,0.0,0.018863125,0.08677038,0.49044126,0.5470306,0.44139713,0.36971724,0.5093044,0.2867195,0.094315626,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.018863125,0.08677038,0.049044125,0.0150905,0.003772625,0.011317875,0.03772625,0.02263575,0.033953626,0.10186087,0.241448,0.4376245,0.26408374,0.25276586,0.46026024,0.70170826,0.56589377,0.63002837,0.63002837,0.543258,0.38103512,0.19240387,0.3470815,0.21881226,0.08299775,0.06790725,0.1358145,0.060362,0.090543,0.26408374,0.4640329,0.4376245,0.15845025,0.47535074,0.69793564,0.513077,0.0,0.0,0.16976812,0.32067314,0.35462674,0.2565385,0.05281675,0.00754525,0.041498873,0.094315626,0.120724,0.32821837,0.52439487,0.513077,0.30181,0.12826926,0.026408374,0.15467763,0.43385187,0.6752999,0.56212115,0.18863125,0.18485862,0.392353,0.5017591,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.09808825,0.049044125,0.1056335,0.09808825,0.06790725,0.03772625,0.00754525,0.018863125,0.28294688,0.5696664,0.66775465,0.3772625,0.875249,1.0412445,0.7997965,0.3734899,0.2867195,0.5885295,0.5055317,0.2867195,0.09808825,0.018863125,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.02263575,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.026408374,0.0150905,0.003772625,0.003772625,0.00754525,0.00754525,0.003772625,0.030181,0.060362,0.06790725,0.05281675,0.011317875,0.030181,0.071679875,0.11317875,0.15467763,0.1961765,0.2263575,0.21503963,0.17731337,0.18485862,0.16976812,0.19994913,0.2263575,0.21503963,0.17731337,0.17731337,0.15845025,0.13204187,0.09808825,0.071679875,0.060362,0.18485862,0.19240387,0.056589376,0.00754525,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.02263575,0.049044125,0.09808825,0.2263575,0.43007925,0.7432071,1.1695137,1.6788181,2.4974778,3.7273536,5.3986263,7.443389,9.669238,11.846043,13.79649,14.283158,13.079691,10.967021,10.163452,9.733373,9.627739,9.774872,10.087999,10.529396,11.121698,11.868678,12.796744,13.947394,15.422491,17.195625,19.591242,22.499935,25.382221,27.657114,30.116865,32.746384,35.39854,37.786613,38.548683,39.310753,41.9365,46.093933,49.24785,49.90428,50.179684,50.30418,49.821285,47.58789,46.444786,46.282562,47.31626,47.489803,42.517483,39.07685,37.435757,36.254925,34.976006,33.825356,33.304733,33.104786,33.255688,33.968716,35.65508,36.726505,36.398285,35.606033,35.217453,36.039886,36.56051,36.02857,35.70035,35.98707,36.469967,37.2094,37.94506,38.710907,39.574837,40.65758,42.37035,44.758423,48.542366,53.571274,58.803905,63.09338,67.17536,69.56721,69.25785,65.70781,61.701283,60.543087,58.44928,54.876602,52.51494,50.900257,49.085625,47.195538,45.16964,42.72498,42.664616,43.37387,44.577335,45.29791,43.886948,41.329105,38.858036,37.45462,37.186764,37.2094,37.145267,38.077103,39.227757,40.710396,43.539864,46.312744,47.187992,46.414604,44.0454,39.92569,35.68526,32.21067,30.060276,29.317068,29.566063,29.34725,28.928488,28.834173,29.384975,30.705395,32.214443,32.520027,32.025814,30.988342,29.486837,27.310032,26.325377,26.1292,26.461191,27.196854,26.868635,27.928743,28.736084,28.664404,28.132465,27.85329,28.981306,29.87919,29.939552,29.554745,31.290152,30.158363,29.63397,30.716713,31.927725,31.71646,32.663387,33.97626,34.81001,34.240345,34.096985,32.188038,30.663897,30.011232,29.041668,29.41893,27.8382,25.329405,22.797974,21.047476,20.470263,19.595015,18.391546,17.240896,16.935314,0.1659955,0.033953626,0.19994913,0.98465514,1.7957695,1.1581959,0.56212115,0.935611,0.8601585,0.18485862,0.0,0.24522063,0.34330887,0.40367088,0.392353,0.120724,0.27917424,0.18485862,0.12826926,0.2867195,0.70170826,0.5055317,0.36594462,0.34330887,0.36594462,0.24522063,0.16976812,0.32821837,0.46026024,0.5885295,0.9922004,1.3958713,2.191895,2.9464202,3.410453,3.5085413,4.376245,4.749735,4.304565,3.2670932,2.425798,2.1579416,1.3317367,0.77338815,0.80734175,1.237421,2.8106055,4.402653,6.0739264,8.507269,13.000465,6.092789,3.229367,3.4368613,5.1081343,6.009792,8.099826,9.461743,7.541477,3.9688015,4.5912848,2.9313297,3.1237335,4.055572,4.851596,4.851596,4.851596,7.020855,9.133525,9.95973,9.276885,6.858632,4.938366,3.6934,3.4972234,4.9119577,4.255521,2.6446102,1.3807807,0.95447415,1.0525624,1.5279131,1.841041,1.5467763,0.8224323,0.44139713,0.41876137,0.9695646,2.4559789,4.568649,6.3644185,8.047009,6.820906,4.1574326,2.0296721,2.8822856,1.6863633,1.7995421,2.0258996,2.252257,3.4481792,1.9353566,1.1883769,0.7809334,0.51684964,0.44139713,0.24899325,0.27917424,0.3169005,0.2565385,0.120724,0.24522063,0.23767537,0.150905,0.05281675,0.0150905,0.003772625,0.0,0.06790725,0.1358145,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.030181,0.030181,0.018863125,0.033953626,0.026408374,0.0,0.0,0.0,0.056589376,0.056589376,0.0,0.0,0.1358145,0.90920264,1.4637785,1.3505998,0.52062225,0.150905,0.02263575,0.0,0.011317875,0.060362,0.42630664,0.83752275,1.0299267,0.91297525,0.59607476,0.26408374,0.08299775,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.011317875,0.03772625,0.060362,0.08677038,0.1659955,0.29426476,0.3734899,0.23013012,0.094315626,0.124496624,0.181086,0.26408374,0.52062225,0.6790725,0.97333723,0.90543,0.46026024,0.1056335,0.25276586,0.25276586,0.1358145,0.026408374,0.1358145,0.18485862,0.19994913,0.27917424,0.3169005,0.0,0.35462674,0.55080324,0.58475685,0.41498876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.03772625,0.0,0.0,0.0,0.36594462,0.49421388,0.27540162,0.090543,0.018863125,0.0,0.10940613,0.21881226,0.0,0.0,0.0,0.23013012,0.5017591,0.19994913,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14713238,0.32067314,0.33953625,0.19240387,0.0452715,0.0452715,0.10186087,0.241448,0.4640329,0.73188925,0.7696155,0.5583485,0.28294688,0.1056335,0.150905,0.18863125,0.362172,0.4678055,0.38480774,0.090543,0.041498873,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.05281675,0.1358145,0.0754525,0.02263575,0.018863125,0.041498873,0.030181,0.018863125,0.00754525,0.0,0.003772625,0.0150905,0.003772625,0.0,0.011317875,0.0452715,0.1056335,0.30181,0.38858038,0.30181,0.124496624,0.0754525,0.1358145,0.18863125,0.20749438,0.19994913,0.21503963,0.21503963,0.1961765,0.17731337,0.15467763,0.1056335,0.056589376,0.10186087,0.150905,0.13958712,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.13204187,0.25276586,0.45648763,0.76207024,1.8863125,4.640329,9.167479,14.396337,18.02183,16.346785,13.551269,11.027383,9.529651,9.125979,9.393836,9.789962,10.242677,10.661438,10.955703,11.053791,11.287694,11.5857315,11.921495,12.298758,13.140053,14.2944765,15.7657995,17.471025,19.240387,20.511763,21.41342,22.499935,24.054256,26.095247,28.290915,30.331905,32.206898,33.90458,35.417404,37.431984,38.858036,39.676697,40.21241,41.151794,42.128902,42.747612,43.724724,44.117077,41.32156,38.963673,36.99436,35.481537,34.447838,33.8744,34.398796,35.02505,35.67017,36.583145,38.32987,38.990078,38.778812,37.620617,36.285107,36.40583,37.873383,38.786358,38.52982,37.348988,36.36056,35.847485,35.481537,36.13043,37.58289,38.56,39.45034,40.89903,43.011696,45.841167,49.394978,54.921875,61.35043,68.22792,73.5926,73.95854,68.52596,63.817726,59.679153,56.604465,55.725445,52.684708,51.04739,50.300407,49.391205,46.690006,42.9702,41.9365,42.52503,43.788857,44.935738,43.728497,40.733032,37.963924,36.232292,35.172184,36.368107,37.22449,38.035606,38.778812,39.10703,40.75567,43.07206,46.15052,48.863037,48.874355,45.309227,39.948326,34.693058,30.822346,28.992622,29.309525,29.37743,29.294434,29.21898,29.388748,29.366114,29.98105,30.863846,31.441057,30.91289,30.241362,28.592726,26.491373,24.510744,23.254461,22.828154,23.8279,25.042685,26.008476,27.008223,29.241617,29.83769,29.988596,29.984823,29.188799,30.143274,29.920689,30.162136,31.5731,33.964943,31.693823,31.282606,32.12013,33.80272,36.1342,37.952606,39.039124,38.190285,35.84371,34.07435,31.995632,29.66415,27.826881,26.321604,24.061802,23.36764,21.711456,19.549744,17.972786,18.693357,1.0940613,0.76584285,0.5696664,0.58098423,0.6828451,0.573439,1.4222796,2.5502944,3.350091,3.180323,1.3656902,0.73188925,0.8601585,0.8903395,0.5885295,0.32821837,0.47912338,0.5696664,0.69039035,0.7884786,0.663982,0.754525,0.90920264,1.6788181,2.927557,3.8707132,2.4597516,1.8749946,2.3088465,3.127506,2.897376,3.0256453,3.9310753,5.1647234,5.8890676,4.8629136,4.402653,4.327201,4.285702,3.9386206,2.938875,1.9278114,1.1204696,0.68661773,0.5998474,0.62625575,1.0487897,1.5052774,1.901403,2.3163917,2.9803739,1.6373192,1.1959221,1.5769572,2.305074,2.546522,2.191895,2.4899325,2.7125173,3.0633714,4.689373,8.937348,6.9265394,4.3007927,3.6594462,4.5460134,4.0782075,5.1043615,7.2358947,9.476834,10.227587,8.084735,6.349328,4.919503,4.063117,4.4139714,4.398881,3.62172,4.908185,7.9526935,9.329701,6.779407,5.13077,4.187614,3.5424948,2.5804756,1.9391292,1.8334957,1.8297231,1.7693611,1.7354075,2.5993385,3.4255435,3.9725742,4.0216184,3.3727267,1.8825399,1.5920477,1.9957186,2.8558772,4.2291126,4.4441524,2.4182527,0.8601585,0.5998474,0.56589377,0.51684964,0.31312788,0.15467763,0.11317875,0.1358145,0.090543,0.13204187,0.14713238,0.10186087,0.0150905,0.02263575,0.011317875,0.018863125,0.03772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.018863125,0.033953626,0.05281675,0.05281675,0.041498873,0.018863125,0.02263575,0.056589376,0.1056335,0.16976812,0.1659955,0.10186087,0.02263575,0.02263575,0.06413463,0.06790725,0.041498873,0.0,0.0,0.14335975,0.39989826,0.69039035,0.8299775,0.56589377,0.14335975,0.0150905,0.0,0.003772625,0.011317875,0.20372175,0.79602385,1.3317367,1.5015048,1.1431054,0.482896,0.14335975,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.10186087,0.14335975,0.18863125,0.2565385,0.16222288,0.11317875,0.08677038,0.06790725,0.071679875,0.060362,0.09808825,0.10940613,0.0754525,0.0452715,0.018863125,0.120724,0.23767537,0.41498876,0.83752275,1.1506506,1.3015556,1.0902886,0.6451189,0.4376245,0.67152727,0.663982,0.45648763,0.26408374,0.49044126,0.27540162,0.19994913,0.20372175,0.20372175,0.120724,0.094315626,0.16976812,0.2867195,0.36971724,0.3055826,0.1961765,0.17731337,0.26031113,0.39989826,0.48666862,0.59607476,0.62248313,0.48666862,0.23767537,0.060362,0.12826926,0.26408374,0.35839936,0.3772625,0.35839936,0.13958712,0.033953626,0.05281675,0.1358145,0.16976812,0.033953626,0.0,0.1961765,0.40367088,0.041498873,0.124496624,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.06413463,0.120724,0.1961765,0.25276586,0.1659955,0.13204187,0.14713238,0.19994913,0.29426476,0.20372175,0.1961765,0.18863125,0.13958712,0.030181,0.06790725,0.1961765,0.26031113,0.22258487,0.150905,0.11317875,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.018863125,0.011317875,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.05281675,0.030181,0.018863125,0.0150905,0.02263575,0.018863125,0.00754525,0.0,0.0,0.0,0.003772625,0.0,0.0150905,0.02263575,0.030181,0.071679875,0.2565385,0.35462674,0.27917424,0.10186087,0.06413463,0.08677038,0.1358145,0.17731337,0.20372175,0.2263575,0.23390275,0.21881226,0.23013012,0.26031113,0.241448,0.24899325,0.20749438,0.16976812,0.14713238,0.06790725,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.090543,0.32821837,1.0902886,2.9464202,6.8246784,10.310584,13.924759,17.13149,18.327412,12.872196,8.488406,6.1644692,5.873977,6.537959,7.3905725,8.431817,9.4127,10.238904,10.993429,11.431054,11.819634,12.166716,12.47607,12.736382,13.102326,13.7700815,14.641558,15.645076,16.750456,17.757746,18.255732,18.757492,19.557287,20.745665,22.160398,23.692085,25.201136,26.729048,28.505955,30.275316,31.659868,32.919926,34.06303,34.817554,35.61735,36.413376,37.2094,37.586662,36.696323,35.13823,34.50443,33.50091,32.003178,31.02984,30.35454,29.867872,29.63397,29.849009,30.822346,32.331398,33.74613,34.693058,35.225,35.847485,37.2509,38.34496,38.84295,38.72222,38.194054,36.9755,35.73053,35.02128,35.002415,35.421177,36.096478,37.530075,39.310753,41.151794,42.8872,46.856003,53.250603,60.87885,68.084564,72.73998,75.0111,75.50909,73.256836,68.63914,63.402737,59.162304,55.385906,52.39044,50.22873,48.681953,46.9805,45.192276,43.686996,42.94379,43.581364,44.071804,43.788857,42.5703,40.446312,37.62439,36.349243,36.941544,38.197826,39.3598,40.11055,40.13696,40.766987,41.913864,43.637955,46.139202,47.595436,46.63342,43.554955,39.125893,34.56856,32.387985,31.795683,31.38824,30.788393,30.645033,29.76224,29.467974,29.667923,29.898052,29.317068,29.366114,29.07562,28.562544,27.63825,25.804754,24.118391,23.156372,22.975286,23.544952,24.76351,26.996904,28.747402,30.384722,31.535372,31.082657,30.35454,30.46772,31.048704,31.939043,33.21042,32.79543,32.493618,33.051968,34.432747,35.82862,37.616844,39.729515,41.845955,43.441776,43.788857,41.94782,38.12992,33.70463,29.584925,26.223516,24.657877,23.495909,22.043447,20.440083,19.655376,1.0638802,0.91674787,1.3317367,1.3505998,0.8262049,0.41876137,1.6788181,2.7238352,4.346064,5.7796617,4.6856003,2.6710186,1.6486372,1.388326,1.4826416,1.3430545,1.0336993,0.965792,1.1695137,1.7429527,2.8256962,3.380272,2.7917426,2.7087448,3.8405323,5.96452,4.727099,3.6745367,3.7688525,4.67051,4.727099,4.085753,4.851596,7.6131573,9.771099,5.5495315,6.009792,8.820397,9.276885,6.360646,2.7389257,1.6071383,1.6561824,1.6637276,1.1883769,0.56589377,0.5017591,0.4678055,0.44139713,0.40367088,0.34330887,0.4074435,1.3430545,2.2220762,2.4220252,1.6222287,3.9197574,4.3007927,3.0256453,1.5015048,2.2975287,4.7346444,3.6368105,2.2258487,1.9504471,2.4861598,2.938875,4.08198,6.1305156,8.699674,10.816116,9.646602,8.216777,6.749226,5.379763,4.1762958,4.244203,3.6669915,4.236658,5.594803,5.2099953,5.8626595,8.805306,8.43559,5.247721,5.8136153,3.9574835,3.240685,2.6219745,1.7429527,0.90920264,1.3204187,1.8297231,2.1994405,2.2409391,1.8372684,1.0789708,0.9016574,1.7769064,3.531177,5.3571277,4.7610526,2.6634734,1.026154,0.5357128,0.6149379,0.724344,0.73188925,0.6790725,0.5394854,0.21881226,0.14335975,0.211267,0.27917424,0.2565385,0.1056335,0.05281675,0.0150905,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.011317875,0.02263575,0.041498873,0.071679875,0.071679875,0.0452715,0.041498873,0.08299775,0.15845025,0.22258487,0.19994913,0.120724,0.056589376,0.120724,0.090543,0.090543,0.1056335,0.124496624,0.14713238,0.13204187,0.13204187,0.1961765,0.2867195,0.2678564,0.06413463,0.003772625,0.0,0.0,0.0,0.060362,0.4678055,1.0978339,1.6410918,1.6109109,0.7696155,0.26408374,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.13958712,0.27540162,0.44139713,0.573439,0.513077,0.44139713,0.30935526,0.19994913,0.14335975,0.120724,0.1358145,0.124496624,0.06790725,0.0,0.0,0.071679875,0.22258487,0.42630664,0.66775465,0.94315624,0.95447415,0.87147635,0.73566186,0.6073926,0.59230214,0.38858038,0.41498876,0.38480774,0.29049212,0.4074435,0.35839936,0.33576363,0.2263575,0.071679875,0.060362,0.011317875,0.030181,0.116951376,0.23013012,0.26408374,0.20749438,0.22258487,0.29426476,0.392353,0.42630664,0.6187105,0.80356914,0.814887,0.6375736,0.3961256,0.28294688,0.26031113,0.32067314,0.4074435,0.41876137,0.30935526,0.29426476,0.32444575,0.36971724,0.41498876,0.08299775,0.1961765,0.3734899,0.392353,0.211267,0.10186087,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026408374,0.07922512,0.120724,0.07922512,0.056589376,0.049044125,0.05281675,0.071679875,0.060362,0.11317875,0.124496624,0.06413463,0.0,0.02263575,0.06413463,0.16222288,0.2263575,0.06790725,0.0754525,0.10186087,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.00754525,0.0,0.0150905,0.026408374,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.00754525,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.049044125,0.011317875,0.00754525,0.00754525,0.00754525,0.00754525,0.0150905,0.003772625,0.0,0.003772625,0.00754525,0.0,0.0150905,0.026408374,0.02263575,0.02263575,0.05281675,0.2263575,0.3055826,0.241448,0.1056335,0.060362,0.0452715,0.07922512,0.14335975,0.21503963,0.27540162,0.271629,0.271629,0.271629,0.271629,0.27540162,0.34330887,0.33576363,0.27540162,0.17731337,0.0754525,0.056589376,0.03772625,0.0150905,0.0,0.00754525,0.00754525,0.00754525,0.011317875,0.018863125,0.026408374,0.23013012,0.8563859,2.372981,5.0854983,9.125979,13.215506,15.939341,15.588487,12.645839,9.797507,6.1531515,3.863168,3.0030096,3.2633207,3.9574835,4.768598,5.753253,6.809588,7.884786,8.9788475,9.906913,10.808571,11.691365,12.468526,12.992921,13.2607765,13.641812,14.188843,14.894323,15.690348,16.467508,16.897587,17.229578,17.63325,18.199142,18.908396,19.844007,20.934296,22.228306,23.903353,25.54067,26.868635,28.045694,29.06053,29.747149,30.860073,31.795683,33.078377,34.73833,36.31529,35.443813,34.127167,32.844475,31.742867,30.64126,29.524563,28.309778,27.29117,26.676231,26.600779,27.487347,28.430502,29.5472,30.939297,32.701115,34.45161,35.95689,36.858547,37.31126,38.009197,38.069557,37.299942,36.469967,35.715443,34.55347,33.93099,34.455383,35.61735,37.10754,38.80522,41.51774,45.705353,50.37209,54.948284,59.305664,66.53779,73.86423,79.01763,80.903946,79.60239,76.10894,70.616,64.52321,59.06799,55.321774,52.763935,50.108006,47.478485,45.21114,43.856766,43.671906,44.42266,44.988552,44.62638,42.962654,40.21241,38.925945,38.541138,38.756176,39.518246,40.08414,40.19732,40.506676,41.43097,43.14751,44.81124,46.49383,47.15027,46.010933,42.574074,39.2768,37.111313,35.02505,33.078377,32.433258,30.939297,30.230043,30.158363,30.471493,30.818573,30.056503,29.17371,28.407866,27.69484,26.698868,26.20088,25.125683,24.091984,23.654358,24.348522,25.363358,27.079903,29.21898,31.022295,31.263742,31.067568,31.207153,31.56178,32.146538,33.11233,33.365097,33.436775,33.847992,34.6742,35.549446,36.971725,38.484547,41.049934,44.732014,48.670635,49.46666,47.70107,44.07935,38.835403,31.724003,29.158619,28.064558,27.083675,25.442583,22.971514,1.3053282,1.1317875,1.8863125,2.252257,1.750498,0.7469798,1.3807807,2.003264,3.7462165,5.7796617,5.3194013,8.409182,5.4288073,2.7389257,2.625747,3.2972744,2.4559789,1.9655377,1.6750455,1.8184053,2.9841464,3.4217708,2.9351022,2.5427492,3.169005,5.6551647,5.8513412,5.149633,6.255012,8.43559,7.541477,4.447925,4.738417,7.726336,10.216269,6.515323,6.428553,8.858124,8.956212,5.723072,2.0372176,1.1506506,1.5920477,1.9278114,1.5580941,0.7054809,0.5394854,0.362172,0.24522063,0.22258487,0.29049212,0.23767537,1.0751982,1.7844516,1.7919968,0.995973,3.6707642,4.06689,2.7879698,1.2751472,1.7957695,1.7731338,1.6033657,1.7316349,2.203213,2.6672459,3.5500402,4.4215164,5.7419353,7.6584287,10.005001,9.910686,9.020347,7.7829256,6.379509,4.708236,4.610148,4.112161,3.6028569,3.0407357,1.9542197,5.4212623,8.827943,9.906913,9.397609,11.068882,7.281166,6.1003346,5.0968165,3.3463185,1.4298248,1.086516,0.90920264,0.83752275,0.845068,0.90920264,0.724344,0.56212115,1.1619685,2.5804756,4.1612053,3.7009451,2.5012503,1.327964,0.6451189,0.63002837,0.69039035,0.7997965,0.875249,0.7884786,0.3734899,0.19240387,0.23013012,0.32821837,0.3470815,0.181086,0.11317875,0.03772625,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.06413463,0.0754525,0.0754525,0.11317875,0.19994913,0.27917424,0.2565385,0.17731337,0.090543,0.049044125,0.10940613,0.06413463,0.090543,0.1358145,0.16222288,0.14713238,0.071679875,0.033953626,0.030181,0.056589376,0.090543,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.1659955,0.65643674,1.3656902,1.9278114,1.1317875,0.44894236,0.08299775,0.0150905,0.00754525,0.011317875,0.030181,0.05281675,0.07922512,0.12826926,0.28294688,0.43007925,0.6526641,0.8903395,0.9393836,0.784706,0.5319401,0.33953625,0.24899325,0.18485862,0.20372175,0.181086,0.10940613,0.049044125,0.10186087,0.32444575,0.44516975,0.6752999,0.9695646,1.0223814,0.77716076,0.6375736,0.6187105,0.6187105,0.422534,0.11317875,0.14713238,0.19240387,0.15845025,0.17354076,0.26408374,0.35085413,0.23390275,0.0,0.0,0.0,0.0,0.033953626,0.08677038,0.10940613,0.10940613,0.13204187,0.1659955,0.18863125,0.18485862,0.32067314,0.5319401,0.6451189,0.5998474,0.42630664,0.2867195,0.211267,0.23013012,0.3055826,0.33953625,0.29803738,0.3734899,0.41498876,0.39989826,0.43385187,0.68661773,0.95447415,0.8563859,0.44516975,0.211267,0.041498873,0.0,0.0,0.011317875,0.056589376,0.0754525,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.071679875,0.060362,0.00754525,0.0,0.00754525,0.003772625,0.0754525,0.15467763,0.0,0.02263575,0.08299775,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.003772625,0.018863125,0.030181,0.02263575,0.02263575,0.033953626,0.030181,0.0150905,0.00754525,0.0,0.026408374,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.041498873,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.003772625,0.00754525,0.0,0.0150905,0.02263575,0.033953626,0.06413463,0.11317875,0.29426476,0.30181,0.23013012,0.13958712,0.06790725,0.030181,0.05281675,0.10940613,0.17731337,0.26408374,0.3055826,0.331991,0.331991,0.31312788,0.2867195,0.3470815,0.35462674,0.30935526,0.23013012,0.16222288,0.12826926,0.08677038,0.049044125,0.02263575,0.00754525,0.03772625,0.0452715,0.08677038,0.26408374,0.7092535,2.5201135,5.485397,8.650629,11.370691,13.309821,13.728582,13.196642,10.246449,5.674028,2.5314314,1.4939595,1.1431054,1.2411937,1.5769572,1.9806281,2.5125682,3.1916409,4.032936,5.0138187,6.0739264,7.1679873,8.36391,9.635284,10.861387,11.861133,12.510024,13.094781,13.705947,14.362384,15.00373,15.690348,16.25624,16.65614,16.927769,17.176762,17.448391,17.855835,18.534906,19.549744,20.8513,21.990631,23.378958,24.491882,25.287905,26.212198,27.196854,28.02683,29.17371,30.92798,33.421684,33.410366,32.527573,31.878681,31.599506,30.852528,29.852781,28.611588,27.381712,26.374422,25.778347,26.057522,26.29897,26.664913,27.340214,28.502182,29.709421,31.309015,32.50871,33.25946,34.270527,36.07384,37.00568,37.450848,37.420666,36.537872,34.557243,33.923443,33.98758,34.625153,36.21343,38.31478,40.465176,41.646008,42.2949,44.301937,51.194523,60.524223,70.129326,78.7875,86.24598,89.65643,88.18888,83.04302,75.965576,69.250305,64.10067,59.535793,55.510403,51.915092,48.568775,46.569283,46.474968,47.26722,48.08965,48.255646,46.241066,44.000126,42.057224,40.78585,40.408585,40.502903,40.495358,40.55949,40.733032,40.95939,41.41965,43.37387,45.678944,47.335125,47.45962,46.82582,44.18121,40.668896,37.360306,35.27027,34.15735,32.62566,31.757957,31.901318,32.66716,32.071087,30.558262,28.894535,27.540163,26.619642,26.736593,26.393284,25.842482,25.4954,25.933023,26.034885,26.563053,27.626932,28.966215,29.98105,31.063795,31.908863,32.587936,33.25946,34.142258,35.08541,35.00996,35.119366,35.5834,35.538128,36.941544,37.880928,39.582382,42.691025,47.274765,51.254883,53.111015,52.08109,47.712387,39.88419,36.08516,33.523544,31.64478,29.830147,27.423212,1.9353566,1.5015048,1.9542197,2.516341,2.546522,1.5354583,1.2411937,1.3166461,2.3390274,3.8103511,4.1762958,14.388792,10.106862,4.6818275,3.6783094,4.8855495,3.6669915,3.308592,3.0143273,2.5691576,2.3314822,1.7391801,1.81086,1.9051756,2.4333432,4.859141,6.3455553,6.0512905,8.405409,12.121444,10.174769,4.5761943,4.247976,5.9192486,7.364164,7.4018903,5.3156285,4.304565,3.4934506,2.516341,1.5052774,1.146878,1.3694628,1.6939086,1.6939086,1.0035182,0.80734175,0.5319401,0.32821837,0.26031113,0.27917424,0.07922512,0.02263575,0.0150905,0.033953626,0.1056335,0.08677038,0.13958712,0.754525,1.871222,2.8785129,2.9237845,2.9992368,3.3010468,3.8820312,4.644101,4.7836885,4.727099,5.028909,5.938112,7.4018903,8.14887,8.243186,7.7904706,6.9454026,5.907931,5.5457587,5.13077,4.38379,3.5802212,3.5689032,6.620957,5.938112,8.039464,12.985375,14.369928,10.038955,8.461998,7.2057137,5.3910813,3.6934,1.8372684,0.7394345,0.56589377,0.9808825,1.1280149,0.9620194,0.5998474,0.39989826,0.5885295,1.267602,2.1654868,2.3956168,1.9466745,1.1921495,0.90543,0.62248313,0.5885295,0.7507524,0.8941121,0.6187105,0.21503963,0.14713238,0.23767537,0.32067314,0.23013012,0.20749438,0.10186087,0.02263575,0.011317875,0.00754525,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.018863125,0.03772625,0.0452715,0.071679875,0.1659955,0.29803738,0.362172,0.24899325,0.12826926,0.0452715,0.011317875,0.0,0.0150905,0.06413463,0.09808825,0.08677038,0.011317875,0.026408374,0.056589376,0.08299775,0.10186087,0.10940613,0.05281675,0.026408374,0.011317875,0.0,0.0,0.0,0.02263575,0.2565385,0.8563859,1.9240388,1.539231,0.79602385,0.25276586,0.090543,0.08677038,0.1056335,0.124496624,0.14335975,0.18863125,0.3055826,0.58475685,0.7205714,0.8337501,0.9997456,1.2713746,1.0148361,0.7054809,0.482896,0.36971724,0.27540162,0.27917424,0.24522063,0.17354076,0.12826926,0.241448,0.55457586,0.62248313,0.80356914,1.086516,1.0601076,0.8601585,0.8299775,0.8299775,0.6790725,0.14713238,0.14335975,0.1659955,0.14713238,0.07922512,0.0,0.049044125,0.18485862,0.16222288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0,0.0,0.071679875,0.14335975,0.16222288,0.120724,0.18485862,0.14713238,0.1056335,0.11317875,0.18485862,0.11317875,0.19240387,0.23390275,0.21881226,0.27917424,1.3317367,1.6071383,1.2261031,0.5319401,0.08677038,0.06413463,0.02263575,0.0,0.02263575,0.10940613,0.14713238,0.06413463,0.018863125,0.049044125,0.056589376,0.026408374,0.011317875,0.018863125,0.033953626,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.011317875,0.003772625,0.0,0.011317875,0.02263575,0.02263575,0.056589376,0.049044125,0.026408374,0.00754525,0.0,0.003772625,0.05281675,0.06413463,0.018863125,0.0,0.003772625,0.003772625,0.0,0.003772625,0.011317875,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.00754525,0.0452715,0.11317875,0.20749438,0.3961256,0.32444575,0.22258487,0.16976812,0.08677038,0.041498873,0.056589376,0.08299775,0.10940613,0.17731337,0.29426476,0.362172,0.39989826,0.4074435,0.392353,0.4074435,0.34330887,0.27917424,0.24899325,0.24899325,0.17731337,0.120724,0.08299775,0.060362,0.026408374,0.13958712,0.33953625,0.845068,1.8561316,3.531177,7.250985,11.800771,14.584969,14.43029,11.604594,7.6810646,3.9801195,1.4449154,0.33953625,0.25276586,0.4979865,0.5885295,0.6375736,0.7167987,0.83752275,1.0940613,1.478869,1.9881734,2.5993385,3.2972744,4.1536603,5.2062225,6.4247804,7.748972,9.0957985,10.314357,11.431054,12.408164,13.230596,13.8719425,14.626467,15.414946,16.01102,16.36942,16.618414,16.833452,16.984358,17.372938,18.048239,18.829172,19.18757,20.4514,21.579414,22.413166,23.695858,24.257978,24.793692,25.144547,25.646305,27.128946,27.875927,28.67195,29.422703,29.93578,29.920689,29.528336,28.97376,28.234325,27.479801,27.061039,27.185535,27.083675,26.70264,26.11411,25.484081,25.310541,26.1707,27.19308,27.860836,28.01174,30.456402,32.99915,35.2665,37.130177,38.710907,36.983044,35.98707,35.08164,34.481792,35.277817,37.239582,38.348732,37.560253,35.51549,34.5082,37.15658,42.932472,51.11907,61.91632,76.47111,89.497986,96.23966,96.99419,93.04425,86.65343,79.738205,72.95125,67.069725,62.104954,57.325035,53.26192,51.0323,50.353226,50.839893,52.009407,52.050907,50.594673,48.44428,46.146748,43.9624,42.136448,41.64978,41.40456,40.917892,40.336906,40.231274,40.67644,41.67619,43.483276,46.61833,50.549404,50.18723,47.606754,44.14726,40.42745,39.201347,36.371876,34.4667,34.081894,33.90458,33.983807,32.603024,30.754438,28.966215,27.287397,26.676231,26.853544,27.396803,27.970242,28.336185,28.08342,27.476028,27.155355,27.460938,28.449366,30.51299,32.240852,33.7914,35.108047,35.92671,37.620617,37.239582,37.08113,37.416893,36.5341,37.680977,38.41664,39.054214,40.20109,42.736298,47.821796,51.96791,53.46564,51.700054,47.131405,42.98529,39.012714,35.73053,33.448093,32.23708,1.9240388,1.5580941,1.5656394,1.6524098,1.8787673,2.6710186,2.6219745,1.9579924,1.8146327,3.3312278,7.6886096,11.144334,8.778898,5.847569,4.4215164,3.3727267,2.0070364,3.8895764,6.696409,8.43559,7.4471617,5.0175915,3.4670424,3.180323,4.61392,8.299775,8.360137,6.436098,6.1078796,7.8923316,9.246704,5.523123,4.9044123,5.594803,6.3644185,6.560595,4.768598,4.244203,3.5689032,2.5540671,2.2748928,2.8332415,3.2142766,3.1463692,2.5917933,1.7240896,1.237421,0.59230214,0.16976812,0.056589376,0.0452715,0.033953626,0.02263575,0.02263575,0.041498873,0.090543,0.056589376,0.03772625,0.10940613,0.29049212,0.5357128,2.474842,3.8292143,4.025391,3.4594972,3.5085413,2.252257,1.7278622,1.9655377,2.674791,3.2520027,4.557331,6.3945994,7.6923823,7.9225125,7.0812173,6.3342376,5.7381625,5.100589,4.606375,4.776143,5.1534057,5.6325293,6.1041074,6.507778,6.8359966,7.7037,5.5193505,4.587512,6.6586833,10.955703,6.560595,2.6144292,0.72811663,0.7884786,0.94692886,0.6413463,0.25276586,0.181086,0.422534,0.59607476,1.1317875,2.6936543,3.1765501,2.372981,1.9693103,1.1393328,0.995973,1.3505998,1.6561824,1.0223814,0.3734899,0.150905,0.1358145,0.21503963,0.35085413,0.35085413,0.23013012,0.116951376,0.056589376,0.030181,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.018863125,0.0,0.0,0.0,0.00754525,0.033953626,0.071679875,0.1056335,0.08299775,0.041498873,0.0150905,0.011317875,0.0,0.02263575,0.041498873,0.0452715,0.049044125,0.060362,0.1358145,0.181086,0.120724,0.0,0.0,0.0,0.056589376,0.056589376,0.0,0.0,0.0,0.0,0.07922512,0.422534,1.3128735,1.9353566,1.4864142,0.80734175,0.392353,0.36594462,0.41498876,0.30935526,0.19240387,0.15845025,0.24522063,1.20724,1.5580941,1.358145,0.91674787,0.80734175,0.8337501,0.7205714,0.58475685,0.49421388,0.45648763,0.482896,0.35085413,0.211267,0.14335975,0.1659955,0.27917424,0.38858038,0.4979865,0.63002837,0.83752275,0.97333723,0.9507015,0.7809334,0.5357128,0.36594462,0.34330887,0.45648763,0.52062225,0.40367088,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.2678564,0.29049212,0.15467763,0.0,0.0,0.0,0.0,0.116951376,0.3055826,0.36594462,0.44139713,0.44894236,0.52062225,0.5998474,0.44139713,0.32067314,0.116951376,0.0,0.0,0.0,0.0,0.0,0.090543,0.23767537,0.27540162,0.13958712,0.060362,0.08677038,0.17354076,0.19994913,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.0754525,0.06413463,0.03772625,0.0,0.011317875,0.0150905,0.00754525,0.0,0.0,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.0,0.00754525,0.02263575,0.060362,0.18485862,0.34330887,0.26408374,0.150905,0.11317875,0.1358145,0.041498873,0.05281675,0.08677038,0.1056335,0.090543,0.18863125,0.3055826,0.38480774,0.47535074,0.73188925,0.8186596,0.5998474,0.32821837,0.1358145,0.0754525,0.0754525,0.094315626,0.1056335,0.11317875,0.1358145,0.4074435,1.3241913,3.4745877,6.8397694,10.816116,13.309821,12.400619,8.7600355,4.293247,2.1692593,1.0072908,0.41498876,0.1659955,0.13204187,0.29049212,1.0827434,1.2638294,1.026154,0.63002837,0.3961256,0.47157812,0.62625575,0.8639311,1.1732863,1.5430037,2.052308,2.686109,3.4557245,4.3686996,5.43258,6.700182,8.062099,9.442881,10.710483,11.6875925,12.615658,13.615403,14.50197,15.192361,15.716756,16.252468,16.690092,17.033401,17.30503,17.546478,17.474798,17.738882,18.516043,19.693102,20.889025,21.986858,22.337713,22.450891,22.526344,22.416937,22.990377,23.820354,24.718239,25.5369,26.185791,26.966724,27.543936,27.78161,27.755201,27.755201,27.559025,26.796955,26.4876,26.706413,26.597006,25.631214,24.401339,23.748674,23.58268,22.873425,23.179008,24.793692,27.559025,31.169428,35.172184,37.61307,38.526047,38.163876,37.315033,37.292397,38.90331,39.269253,38.910854,37.288624,32.82184,32.701115,34.315796,37.880928,44.192528,54.6427,68.91454,79.57598,88.10966,94.50426,97.27336,93.3687,86.43084,79.10818,72.57021,66.52647,60.716625,56.464878,54.114532,53.548637,54.18244,54.574795,54.737015,54.133396,52.424397,49.470432,46.576828,44.505657,43.10224,42.230762,41.77805,42.41185,41.38947,40.004917,39.36734,40.40481,44.630154,50.64749,53.971172,53.182693,49.911827,44.369843,40.555717,38.86181,38.065784,35.36836,33.17269,32.39553,32.557755,32.71998,31.463692,30.256453,29.667923,29.64906,29.728285,29.007713,27.98156,28.649315,29.747149,30.143274,28.837946,30.961933,31.769276,33.58768,36.27756,37.232037,38.624134,39.28057,39.5522,39.66915,39.778557,38.593952,38.484547,38.914627,40.061504,42.78534,43.505913,44.758423,46.63719,48.108513,46.99559,45.75062,44.709377,42.392986,39.14853,37.10754,0.55457586,0.784706,1.3091009,1.5203679,1.3166461,1.0827434,1.3845534,1.0299267,1.2411937,2.3201644,3.663219,5.028909,5.43258,6.2814207,7.8923316,9.49947,5.409944,4.164978,5.27413,6.9982195,6.3719635,3.4934506,2.4107075,2.957738,4.727099,7.0548086,5.20245,4.191386,6.043745,10.397354,14.494425,9.337247,5.4967146,3.8895764,4.346064,5.583485,10.401127,11.962994,11.638548,10.33322,8.511042,6.2323766,6.771862,6.296511,4.236658,3.2633207,2.5314314,2.0900342,1.8523588,1.8033148,1.9881734,1.750498,1.6750455,1.5920477,1.3128735,0.6413463,0.38858038,0.18485862,0.116951376,0.20749438,0.41121614,0.84884065,0.97710985,0.94315624,0.91297525,1.0789708,1.0940613,1.0374719,1.3392819,2.0975795,3.0897799,3.9499383,5.081726,6.1418333,7.0548086,8.009283,6.9793563,5.3080835,4.0706625,3.6594462,3.7499893,4.4215164,5.772116,7.4207535,8.990166,10.133271,10.159679,8.111144,5.59103,3.8292143,3.6934,2.9124665,2.6672459,3.0860074,3.4368613,2.142851,1.1355602,1.0450171,1.7165444,2.8256962,3.904667,4.5950575,5.251494,4.5497856,2.7917426,1.9202662,0.875249,0.7054809,1.1393328,1.6637276,1.5354583,0.694163,0.32444575,0.19994913,0.21881226,0.41121614,0.38103512,0.26408374,0.211267,0.23767537,0.21503963,0.10186087,0.05281675,0.02263575,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.018863125,0.0150905,0.02263575,0.0452715,0.03772625,0.00754525,0.00754525,0.02263575,0.03772625,0.033953626,0.03772625,0.36971724,0.35839936,0.011317875,0.0,0.0150905,0.23390275,0.2678564,0.10940613,0.120724,0.07922512,0.049044125,0.03772625,0.060362,0.14713238,0.17731337,0.14335975,0.06790725,0.0,0.0,0.0,0.0,0.0150905,0.21881226,0.935611,1.9278114,2.1881225,1.9391292,1.448688,1.0148361,0.58475685,0.27540162,0.1056335,0.05281675,0.060362,0.5281675,0.7922512,0.8563859,0.72811663,0.392353,0.47535074,0.46026024,0.3734899,0.3055826,0.38480774,0.44894236,0.4074435,0.30935526,0.211267,0.1659955,0.16222288,0.18863125,0.24522063,0.35085413,0.5583485,0.7997965,1.0110635,1.0902886,1.0148361,0.8526133,0.5281675,0.241448,0.20749438,0.31312788,0.14713238,0.1961765,0.2678564,0.271629,0.211267,0.16976812,0.19994913,0.08299775,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0,0.03772625,0.056589376,0.03772625,0.060362,0.3055826,0.11317875,0.056589376,0.030181,0.0,0.0,0.08677038,0.0452715,0.02263575,0.060362,0.071679875,0.1961765,0.3772625,0.513077,0.47157812,0.08677038,0.21881226,0.27540162,0.25276586,0.19994913,0.21881226,0.30935526,0.35839936,0.34330887,0.241448,0.056589376,0.026408374,0.35462674,0.63002837,0.63002837,0.331991,0.25276586,0.094315626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.003772625,0.011317875,0.011317875,0.011317875,0.00754525,0.003772625,0.011317875,0.011317875,0.02263575,0.026408374,0.02263575,0.011317875,0.011317875,0.018863125,0.0452715,0.060362,0.011317875,0.033953626,0.06790725,0.08299775,0.060362,0.011317875,0.033953626,0.026408374,0.00754525,0.0,0.0,0.003772625,0.018863125,0.026408374,0.018863125,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.011317875,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.00754525,0.02263575,0.049044125,0.13958712,0.116951376,0.0754525,0.060362,0.06413463,0.06413463,0.06413463,0.05281675,0.03772625,0.056589376,0.19994913,0.32821837,0.38103512,0.41121614,0.6111652,0.9318384,0.90543,0.6187105,0.2565385,0.08677038,0.049044125,0.10186087,0.17354076,0.4678055,1.4675511,4.0404816,7.4169807,9.797507,10.242677,8.707218,5.904158,4.217795,2.6672459,1.1846043,0.59230214,0.33953625,0.27540162,0.42630664,0.72811663,1.0336993,1.0751982,0.8262049,0.48666862,0.2263575,0.18863125,0.21503963,0.31312788,0.46026024,0.6413463,0.88279426,1.0450171,1.3656902,1.7995421,2.323937,2.9652832,3.7952607,4.727099,5.7494807,6.820906,7.865923,8.959985,10.163452,11.3820095,12.5326605,13.555041,14.524607,15.16218,15.592259,15.984612,16.569368,16.957949,17.21826,17.53516,17.99542,18.606586,19.413929,20.19109,20.900343,21.417192,21.560553,21.647322,21.805773,22.01704,22.299986,22.692339,23.473272,24.333431,25.038912,25.559534,26.046204,26.32915,26.046204,26.087702,27.011995,29.06053,27.747658,25.148317,23.322369,22.684793,22.005722,21.402102,21.481327,22.49239,24.427748,27.015768,30.248907,33.863083,36.439785,37.548935,37.76775,38.84295,39.303207,38.469456,36.42092,33.995125,33.74613,33.036877,34.029076,37.669662,43.70586,53.786316,60.64872,66.41706,72.69471,80.553085,85.45373,86.34407,84.73693,81.601875,77.353905,71.11398,64.90801,59.80365,56.532787,55.47645,56.551647,57.94752,58.76995,58.14747,55.23123,51.183205,47.120087,43.743587,41.67619,41.44983,42.200584,42.219448,41.11784,39.37866,38.367596,38.48832,40.45763,43.426685,47.09745,51.718918,54.4088,52.337627,47.9727,43.151283,39.118347,36.960407,35.523037,34.79115,34.496883,34.138485,33.278324,32.57662,31.67496,30.535627,29.434021,29.513245,30.003687,30.301723,30.573353,31.757957,33.04065,34.315796,35.794666,37.23581,37.963924,37.579117,38.409096,39.903053,41.027298,40.269,40.04264,39.340935,39.246616,39.85024,40.257683,41.370605,43.09847,44.22271,44.184982,43.10224,42.600483,41.3027,39.661606,39.00517,41.529057,0.7092535,0.9242931,1.1544232,1.3958713,1.7693611,2.516341,1.961765,1.267602,1.1883769,1.690136,1.9693103,2.003264,2.9464202,4.29702,5.9418845,8.130007,6.858632,6.387054,5.692891,4.4705606,3.127506,2.6068838,2.7879698,5.251494,8.914713,10.050273,8.492179,5.27413,4.2894745,6.5266414,10.057818,8.722309,6.439871,4.568649,3.772625,4.0216184,7.277394,9.001483,9.348565,8.386545,6.096562,5.070408,4.9760923,4.346064,3.2859564,3.4745877,5.160951,5.704209,5.081726,3.8141239,2.9841464,2.5804756,2.655928,2.4597516,1.7542707,0.80734175,0.58098423,0.3961256,0.3961256,0.5885295,0.8224323,0.633801,0.3734899,0.33953625,0.5583485,0.77338815,1.0186088,1.3392819,1.6146835,1.8297231,2.071171,2.9351022,3.4368613,4.1989317,5.451443,7.032173,7.352846,6.63982,5.4740787,4.2404304,3.1199608,4.436607,4.9987283,5.772116,6.85486,7.484888,6.349328,5.934339,5.1081343,4.0103,4.0480266,4.930821,5.885295,6.270103,5.560849,3.3312278,2.2711203,2.6823363,3.5990841,4.13857,3.5387223,3.482133,3.4179983,3.572676,3.8556228,3.8480775,2.9124665,2.2220762,1.8787673,1.7542707,1.4977322,0.8639311,0.38858038,0.14713238,0.120724,0.21503963,0.181086,0.116951376,0.094315626,0.116951376,0.11317875,0.060362,0.033953626,0.0150905,0.0,0.0,0.0452715,0.07922512,0.06413463,0.011317875,0.026408374,0.0452715,0.03772625,0.030181,0.030181,0.018863125,0.056589376,0.07922512,0.090543,0.090543,0.07922512,0.1056335,0.30181,0.26031113,0.003772625,0.0,0.011317875,0.116951376,0.13958712,0.0754525,0.071679875,0.030181,0.0452715,0.06790725,0.071679875,0.071679875,0.08677038,0.06413463,0.030181,0.0,0.0,0.0,0.0,0.003772625,0.09808825,0.44516975,1.2902378,1.9579924,2.1805773,1.9089483,1.3128735,0.7696155,0.34330887,0.09808825,0.02263575,0.02263575,0.1961765,0.29803738,0.38480774,0.47157812,0.5281675,0.543258,0.44894236,0.2867195,0.16222288,0.21881226,0.29426476,0.30935526,0.25276586,0.150905,0.06790725,0.05281675,0.056589376,0.094315626,0.17731337,0.3055826,0.3772625,0.513077,0.7054809,0.91674787,1.0940613,0.68661773,0.36594462,0.18485862,0.13204187,0.15467763,0.11317875,0.13204187,0.1358145,0.116951376,0.13958712,0.10940613,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.026408374,0.049044125,0.11317875,0.27917424,0.11317875,0.13958712,0.15845025,0.124496624,0.14713238,0.26408374,0.116951376,0.0,0.0,0.0,0.14713238,0.29426476,0.38858038,0.38103512,0.23013012,0.29049212,0.3169005,0.27540162,0.19994913,0.17354076,0.24899325,0.2678564,0.211267,0.09808825,0.0,0.0,0.17354076,0.3055826,0.29803738,0.14713238,0.120724,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.003772625,0.0,0.0,0.003772625,0.0150905,0.0150905,0.02263575,0.02263575,0.018863125,0.0150905,0.02263575,0.02263575,0.03772625,0.049044125,0.0150905,0.0150905,0.0452715,0.08299775,0.10186087,0.060362,0.05281675,0.06790725,0.071679875,0.049044125,0.0150905,0.018863125,0.011317875,0.00754525,0.00754525,0.0,0.0150905,0.05281675,0.05281675,0.018863125,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.094315626,0.08677038,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.033953626,0.38480774,1.6637276,1.5656394,0.18863125,0.03772625,0.09808825,0.10940613,0.07922512,0.033953626,0.03772625,0.150905,0.28294688,0.33953625,0.34330887,0.41498876,0.8299775,1.1016065,1.0336993,0.66775465,0.28294688,0.13204187,0.41121614,1.5128226,3.3312278,5.251494,6.9152217,8.412953,8.737399,7.484888,4.881777,2.1994405,1.0789708,0.5885295,0.29049212,0.25276586,0.26408374,0.32067314,0.41498876,0.55080324,0.7167987,0.5772116,0.43007925,0.30181,0.23013012,0.26408374,0.26408374,0.29426476,0.35085413,0.41121614,0.452715,0.47535074,0.5998474,0.7997965,1.0676528,1.4147344,1.8787673,2.4484336,3.127506,3.8971217,4.7233267,5.6853456,6.752999,7.91874,9.171251,10.469034,11.736636,12.672247,13.3626375,13.95494,14.641558,15.399856,15.961976,16.365646,16.690092,17.067356,17.652113,18.402864,19.229069,19.979822,20.4514,20.560806,20.564579,20.455173,20.300495,20.274086,20.760756,21.477554,22.288668,23.069601,23.714722,23.95617,24.239115,25.03514,26.502691,28.49841,28.332415,26.389511,24.125937,22.450891,21.734093,20.723028,19.994913,19.998686,20.813572,22.130219,24.544699,27.845745,31.508965,34.8666,37.111313,38.194054,37.91111,36.737823,35.25518,34.15735,34.1913,33.93476,34.39125,36.11911,39.22021,43.626637,47.380398,51.288837,56.117798,62.610485,68.948494,73.347374,76.17684,77.863205,78.90068,77.73871,74.40371,69.71056,64.82501,61.274975,60.57327,61.15048,62.440716,63.659275,63.84036,60.992027,55.97821,50.262684,45.233772,42.189266,41.264973,40.917892,40.608536,39.96719,38.808994,37.318806,36.828365,37.6093,40.061504,44.690517,50.02501,53.107243,54.235256,53.21665,49.38366,44.656563,40.567036,38.122375,37.330124,37.19431,35.68526,34.79115,34.440292,34.17998,33.176464,31.90509,32.037132,32.188038,32.199356,33.134964,34.523293,35.911617,37.37917,38.552456,38.593952,37.126404,37.67343,39.12212,40.378407,40.351997,39.831375,39.19003,38.812767,38.79013,38.914627,40.216183,42.249626,43.781315,44.230255,43.67568,42.09118,40.736805,39.10326,37.952606,39.337162,0.9205205,1.0751982,1.1732863,1.4109617,1.961765,2.9992368,3.5387223,4.06689,3.7763977,2.6823363,1.6033657,1.1996948,1.5505489,2.3616633,3.6141748,5.5683947,6.1833324,7.9451485,8.269594,6.1606965,2.1805773,2.2862108,3.7009451,7.0170827,11.027383,12.709973,10.457717,5.8513412,3.0860074,3.5349495,5.7419353,6.255012,6.009792,5.6061206,5.87775,7.8961043,6.749226,5.6363015,4.7836885,4.036709,2.8822856,3.240685,3.0143273,2.493705,2.1164427,2.4597516,4.5950575,5.3609,5.0213637,4.195159,3.8556228,3.904667,3.9801195,3.6443558,2.686109,1.1091517,0.8262049,0.66020936,0.65643674,0.8299775,1.1393328,0.663982,0.36594462,0.362172,0.5885295,0.8111144,1.0374719,1.3053282,1.4260522,1.418507,1.50905,2.11267,2.1881225,2.6446102,3.7348988,5.028909,6.3342376,7.2396674,6.8774953,5.194905,2.9652832,4.146115,4.085753,4.4441524,5.455216,5.915476,5.0175915,5.794752,6.221059,6.009792,6.651138,7.7602897,8.420499,9.122208,9.2995205,7.333983,6.175787,6.1229706,5.696664,4.2819295,2.1164427,1.8636768,1.9579924,2.8030603,3.893349,3.8254418,3.1199608,2.293756,1.6524098,1.2600567,0.9242931,0.77338815,0.5470306,0.39989826,0.33576363,0.22258487,0.11317875,0.0452715,0.02263575,0.030181,0.026408374,0.026408374,0.026408374,0.026408374,0.026408374,0.030181,0.16222288,0.2678564,0.26408374,0.18863125,0.19240387,0.21503963,0.14335975,0.07922512,0.06413463,0.09808825,0.19240387,0.19240387,0.18485862,0.21503963,0.26408374,0.26031113,0.2263575,0.124496624,0.0,0.0,0.056589376,0.03772625,0.02263575,0.026408374,0.02263575,0.003772625,0.03772625,0.060362,0.0452715,0.0,0.0,0.0,0.120724,0.331991,0.4376245,0.31312788,0.120724,0.011317875,0.030181,0.120724,0.59607476,1.2940104,1.8070874,1.8863125,1.4524606,1.0374719,0.5583485,0.19240387,0.0150905,0.018863125,0.1659955,0.1961765,0.18863125,0.23013012,0.41876137,0.49044126,0.44894236,0.2678564,0.060362,0.071679875,0.116951376,0.13958712,0.116951376,0.060362,0.0,0.0,0.0,0.02263575,0.06413463,0.10940613,0.1056335,0.15467763,0.41876137,0.8186596,1.0412445,0.88279426,0.51684964,0.29049212,0.2678564,0.22258487,0.16222288,0.060362,0.0,0.011317875,0.056589376,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.0754525,0.07922512,0.041498873,0.011317875,0.030181,0.08299775,0.12826926,0.08299775,0.13958712,0.15845025,0.16222288,0.32821837,0.32067314,0.14335975,0.02263575,0.018863125,0.0,0.094315626,0.150905,0.20372175,0.24522063,0.23013012,0.21503963,0.18863125,0.14713238,0.10186087,0.06413463,0.094315626,0.090543,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.018863125,0.02263575,0.018863125,0.0150905,0.02263575,0.02263575,0.056589376,0.12826926,0.19240387,0.120724,0.07922512,0.0754525,0.08677038,0.08677038,0.071679875,0.06413463,0.049044125,0.02263575,0.00754525,0.00754525,0.003772625,0.00754525,0.0150905,0.00754525,0.02263575,0.05281675,0.0452715,0.011317875,0.011317875,0.018863125,0.018863125,0.018863125,0.02263575,0.041498873,0.18863125,0.1659955,0.07922512,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.056589376,0.39989826,2.1088974,2.2598023,0.7205714,0.13958712,0.116951376,0.11317875,0.08677038,0.0452715,0.03772625,0.11317875,0.23013012,0.29426476,0.29426476,0.29803738,0.6451189,1.2449663,1.6410918,1.5618668,0.935611,0.55080324,1.8184053,3.7650797,5.4665337,6.039973,6.417235,5.8437963,4.666737,3.2067313,1.7278622,0.67152727,0.29803738,0.23767537,0.26408374,0.32821837,0.3470815,0.38480774,0.3961256,0.3961256,0.46026024,0.4678055,0.7507524,1.1695137,1.5505489,1.6825907,1.5279131,1.4977322,1.4449154,1.3430545,1.2638294,0.97710985,0.7809334,0.633801,0.5583485,0.6413463,0.8563859,1.1544232,1.5241405,1.961765,2.4672968,3.127506,3.8858037,4.772371,5.8098426,7.0284004,8.337502,9.484379,10.461489,11.302785,12.091263,12.974057,13.747445,14.396337,14.93205,15.403628,15.875206,16.535416,17.391802,18.357594,19.25925,19.534653,19.610106,19.500698,19.266796,19.002712,19.051756,19.304522,19.810055,20.52308,21.300241,21.51528,22.077402,23.34123,25.118137,26.680004,27.517527,27.053493,25.363358,23.201643,21.971767,20.870161,19.779873,19.18757,19.229069,19.670467,20.877707,22.956423,26.136745,30.101774,34.01399,35.998386,35.953117,34.97978,33.96117,33.553726,34.161118,35.16841,36.334152,37.503666,38.61659,38.280827,39.00894,41.10652,44.671654,49.572292,54.95583,59.777245,64.10067,68.06193,71.86851,75.04883,76.77669,76.67106,74.50557,70.22742,66.62456,65.341866,65.52295,66.58683,68.220375,69.167305,66.46233,61.373062,55.21614,49.35348,44.93951,41.744095,40.046413,39.40884,38.692043,37.79416,36.90759,36.08516,35.938026,37.616844,41.604507,46.584373,51.635918,55.170868,54.933193,52.254627,48.97622,45.66008,42.679707,40.189774,39.19003,37.48103,36.66237,36.783092,36.349243,34.998642,34.95714,34.72324,34.134712,34.387478,35.590942,36.48883,37.801704,39.261707,39.63897,38.17142,38.12615,38.94481,39.98228,40.495358,39.793648,39.039124,38.54491,38.41664,38.56,40.189774,41.876137,43.33237,44.31325,44.603745,42.796658,42.347717,41.27629,39.356026,38.12992,0.694163,0.94315624,1.4524606,1.9844007,2.2711203,2.0108092,4.274384,6.5002327,6.368191,3.9499383,1.7014539,1.5731846,1.4335974,1.8334957,2.8634224,4.1612053,4.214022,7.1679873,10.461489,10.925522,4.8025517,3.1463692,4.9044123,7.250985,9.159933,11.3971,8.099826,5.1081343,4.172523,5.353355,7.0170827,5.198677,5.1458607,6.304056,8.7751255,13.324911,9.303293,5.2665844,2.8898308,2.3654358,2.425798,3.2821836,3.772625,3.4029078,2.323937,1.3355093,1.3392819,1.3732355,1.7769064,2.7087448,4.172523,4.991183,4.930821,4.557331,3.7047176,1.4449154,1.0223814,0.8262049,0.7809334,0.94692886,1.5165952,0.94692886,0.8639311,0.8224323,0.7130261,0.7432071,0.8186596,0.694163,0.6413463,0.9016574,1.6825907,1.7165444,1.5580941,1.720317,2.2862108,2.9011486,4.06689,5.8588867,6.541732,5.541986,3.4368613,3.4632697,3.4255435,4.304565,5.87775,6.7341356,7.3453007,7.5565677,7.352846,7.375482,8.918486,10.740664,10.499215,11.638548,13.536179,11.536687,9.714509,8.514814,6.3417826,3.2821836,1.0789708,1.2789198,1.9957186,2.6031113,2.6031113,1.6222287,1.1921495,0.7809334,0.5772116,0.5394854,0.36971724,0.6149379,0.814887,0.88279426,0.7582976,0.38480774,0.19240387,0.10186087,0.13204187,0.19994913,0.13204187,0.090543,0.11317875,0.12826926,0.120724,0.124496624,0.30935526,0.5055317,0.5583485,0.47157812,0.422534,0.4376245,0.29426476,0.20749438,0.26031113,0.392353,0.44516975,0.38858038,0.3961256,0.5093044,0.6451189,0.513077,0.2867195,0.10186087,0.02263575,0.041498873,0.120724,0.07922512,0.02263575,0.003772625,0.011317875,0.003772625,0.0,0.0,0.00754525,0.041498873,0.30935526,0.6488915,1.4260522,2.3616633,2.5427492,1.3619176,0.44516975,0.0150905,0.003772625,0.02263575,0.150905,0.5998474,1.1581959,1.5656394,1.5241405,1.3015556,0.8601585,0.3961256,0.0754525,0.02263575,0.23390275,0.27540162,0.18863125,0.060362,0.0150905,0.21881226,0.35085413,0.241448,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.09808825,0.150905,0.124496624,0.1659955,0.16976812,0.40367088,0.7696155,0.77716076,0.9280658,0.55457586,0.46026024,0.66775465,0.4074435,0.38858038,0.23767537,0.11317875,0.060362,0.0,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.060362,0.14713238,0.15845025,0.07922512,0.02263575,0.0,0.0,0.0,0.0,0.0,0.003772625,0.08299775,0.36594462,0.19994913,0.094315626,0.049044125,0.03772625,0.0,0.0,0.0,0.03772625,0.07922512,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.003772625,0.011317875,0.011317875,0.02263575,0.0754525,0.19240387,0.3734899,0.22258487,0.090543,0.041498873,0.07922512,0.13958712,0.14713238,0.11317875,0.056589376,0.011317875,0.02263575,0.030181,0.018863125,0.011317875,0.0150905,0.011317875,0.0150905,0.0150905,0.00754525,0.003772625,0.02263575,0.03772625,0.030181,0.02263575,0.03772625,0.090543,0.21503963,0.17354076,0.0754525,0.003772625,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.10186087,0.95447415,1.4411428,1.1544232,0.482896,0.241448,0.124496624,0.071679875,0.0452715,0.049044125,0.1056335,0.21881226,0.29049212,0.3055826,0.29803738,0.5055317,1.2864652,2.203213,2.7917426,2.5540671,1.9391292,3.6443558,5.1345425,5.0779533,3.3350005,3.127506,2.0900342,1.0186088,0.36594462,0.27540162,0.2263575,0.21881226,0.25276586,0.3169005,0.36971724,0.392353,0.4376245,0.5055317,0.6073926,0.7922512,1.2336484,2.1579416,3.3764994,4.508287,4.98741,4.504514,4.255521,3.9386206,3.5575855,3.3878171,2.7540162,1.9806281,1.2713746,0.7469798,0.45648763,0.55457586,0.6149379,0.7130261,0.875249,1.0940613,1.4373702,1.8599042,2.3805263,3.029418,3.8480775,4.919503,6.058836,7.1793056,8.224322,9.167479,9.982366,10.763299,11.570641,12.385528,13.113645,13.573905,14.249205,15.218769,16.4411,17.765291,18.187824,18.51227,18.685812,18.648085,18.316093,17.927513,17.655886,17.674747,18.074646,18.859352,19.217752,19.772327,21.09652,23.065828,24.865372,26.34424,27.29494,26.740366,24.797464,22.677248,21.349285,20.130728,19.25925,18.848034,18.878216,19.251705,20.315586,22.137764,24.90687,28.90208,31.859818,33.093468,33.02933,32.403076,32.23708,33.30096,35.160866,37.371624,39.125893,39.25416,36.685005,34.93451,35.108047,37.662117,42.430714,47.003136,50.83612,54.495567,58.056927,61.116524,65.26641,70.793304,76.04858,78.979904,77.13886,73.21533,70.41227,68.12606,66.63965,67.10745,71.77796,73.343605,72.208046,68.78627,63.478188,56.385654,49.3233,43.694542,40.02755,37.982788,37.79416,37.71116,36.956635,35.722984,35.191048,36.205883,38.495865,42.260944,46.89373,50.9908,54.43898,55.46136,53.484505,49.130894,44.215164,43.909584,41.083885,38.888218,38.26951,37.96015,37.81679,37.865837,37.371624,36.552963,36.579372,36.726505,36.613327,37.39426,39.080624,40.52554,39.9936,39.804966,40.09923,40.57458,40.47272,40.114323,39.065533,38.480774,38.642998,38.94481,40.631172,41.668644,42.634434,43.739815,44.80747,43.626637,44.166122,44.20762,42.872112,40.638718,0.48666862,0.84129536,2.0749438,3.8103511,4.708236,2.4861598,1.3015556,1.3204187,1.5430037,1.569412,1.5580941,1.9353566,2.7351532,2.9464202,2.5125682,2.305074,2.7691069,3.3425457,6.862405,11.1631975,9.061845,6.5002327,6.820906,6.9793563,5.6815734,3.3878171,3.218049,5.2326307,8.7600355,12.596795,15.015047,9.522105,7.4509344,7.281166,7.4773426,6.5002327,4.561104,4.4139714,5.481624,6.198423,4.014073,6.379509,7.8508325,7.1981683,4.719554,2.2258487,0.9695646,0.4640329,0.3734899,0.7922512,2.2447119,3.0256453,3.0558262,3.006782,2.6898816,1.0676528,0.7507524,0.5998474,0.83752275,1.5882751,2.8822856,2.6634734,3.3123648,3.1916409,2.1353056,1.4637785,0.67152727,0.32821837,0.35839936,0.80356914,1.8146327,1.5958204,1.2562841,1.1242423,1.2789198,1.5731846,1.9730829,2.516341,3.4444065,4.4630156,4.7308717,3.2520027,3.029418,3.7801702,4.9157305,5.5382137,6.9793563,4.115934,2.2673476,4.376245,11.016065,17.399347,16.433554,14.988639,13.879487,7.8734684,4.4818783,3.2029586,2.3088465,1.2600567,0.68661773,0.724344,0.98842776,1.1431054,1.0374719,0.73188925,0.62248313,0.6488915,0.814887,0.9922004,0.9318384,0.8941121,1.0223814,1.0299267,0.7507524,0.150905,0.06790725,0.1358145,0.43007925,0.7167987,0.47157812,0.27917424,0.38480774,0.43385187,0.34330887,0.32067314,0.36971724,0.6187105,0.724344,0.60362,0.45648763,0.38480774,0.32821837,0.44516975,0.7205714,0.97710985,0.80734175,0.7922512,0.94315624,1.1846043,1.3430545,0.91674787,0.38858038,0.10186087,0.11317875,0.19994913,0.11317875,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.041498873,0.21503963,1.5430037,3.2482302,5.915476,8.499724,8.314865,3.6896272,1.0223814,0.00754525,0.0,0.0,0.0,0.18485862,0.63002837,1.1959221,1.5241405,1.3317367,1.0714256,0.7092535,0.32821837,0.1056335,0.0452715,0.011317875,0.0,0.003772625,0.0150905,0.11317875,0.1659955,0.10940613,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1659955,0.482896,0.7582976,0.62625575,0.47912338,0.3055826,0.21881226,0.29049212,0.5357128,0.362172,0.48666862,0.69793564,0.8111144,0.6413463,0.49421388,0.60362,0.573439,0.3055826,0.0,0.09808825,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.02263575,0.00754525,0.0,0.0,0.0,0.018863125,0.018863125,0.0,0.0,0.0,0.00754525,0.033953626,0.056589376,0.030181,0.00754525,0.00754525,0.08677038,0.23767537,0.3961256,0.422534,0.32821837,0.1659955,0.049044125,0.120724,0.10940613,0.071679875,0.033953626,0.011317875,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.011317875,0.00754525,0.02263575,0.056589376,0.030181,0.056589376,0.033953626,0.00754525,0.0150905,0.0754525,0.06413463,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.31312788,1.1883769,0.7130261,0.32067314,0.10186087,0.049044125,0.060362,0.10940613,0.27917424,0.39989826,0.4074435,0.33576363,0.543258,1.0902886,2.2069857,3.8858037,5.873977,5.3382645,3.7386713,2.4031622,1.81086,1.6033657,0.79602385,0.40367088,0.26408374,0.23767537,0.21503963,0.21503963,0.1961765,0.19994913,0.24899325,0.32067314,0.43007925,0.59607476,0.77716076,1.0601076,1.6486372,2.9766011,4.738417,6.820906,8.854351,10.223814,9.26934,8.318638,7.3377557,6.4511886,5.9494295,5.560849,3.9348478,2.4823873,1.5920477,0.6413463,0.7394345,0.47157812,0.29426476,0.33953625,0.41121614,0.5583485,0.7507524,0.98465514,1.2600567,1.6033657,2.214531,3.0331905,4.002755,5.040227,6.043745,6.8359966,7.594294,8.386545,9.220296,10.023865,10.574668,11.306557,12.411936,13.845533,15.335721,15.946886,16.920223,17.591751,17.621931,16.999449,16.316603,15.905387,15.735619,15.773345,15.992157,16.418465,17.056038,18.467,20.802254,23.805264,26.75923,28.532362,28.468227,26.64605,23.850534,21.409647,20.175999,19.50447,19.108345,19.074392,19.281887,19.636513,20.387266,21.749184,23.910898,25.948114,27.823109,29.294434,30.128183,30.090458,30.811028,32.584164,35.16464,37.643253,38.435505,36.86232,34.745876,33.35755,33.798946,37.032085,41.012207,44.618835,48.670635,52.839386,55.6349,58.38137,62.169086,65.730446,68.959816,72.95125,77.35767,75.173325,70.095375,65.61726,65.03251,67.778984,70.73672,74.30185,77.95752,80.27392,76.59938,68.63914,58.50964,48.210377,39.642742,36.40583,36.11911,36.854774,37.548935,38.02429,37.57157,36.583145,36.307743,37.273537,39.261707,44.573563,47.995335,50.639946,52.382896,51.89623,48.36505,45.29791,43.494595,42.366577,39.903053,38.54491,38.74863,39.774784,40.70285,40.434994,38.737312,37.45462,37.37917,38.424187,39.597473,40.25391,41.72146,42.29867,41.37438,39.397522,39.325844,38.601498,37.78284,37.763977,39.763466,40.080368,41.33288,43.170147,45.05269,46.24861,43.845448,42.921154,43.37387,44.445293,44.73956,0.452715,1.2261031,2.0636258,3.519859,5.6551647,8.039464,5.5306683,3.108643,1.7278622,1.2713746,0.56589377,0.76207024,1.6825907,3.2369123,4.738417,4.8930945,4.2706113,4.0970707,4.2064767,4.5120597,4.9987283,5.59103,6.700182,6.115425,3.9650288,2.71629,4.115934,6.277648,7.364164,7.7414265,9.97482,10.748209,10.61994,10.084227,8.793989,5.560849,3.6896272,3.682082,3.3236825,2.8143783,4.768598,5.613666,5.3269467,6.3531003,8.031919,6.598321,3.1237335,2.1881225,2.323937,2.8219235,3.7084904,2.595566,1.9768555,1.9202662,2.0070364,1.3128735,0.8865669,0.5998474,1.1053791,3.5764484,9.695646,11.778135,9.424017,8.265821,8.213005,3.429316,4.991183,9.574923,14.124708,15.113135,8.578949,5.0779533,4.183841,4.659192,5.723072,7.039718,5.624984,4.7233267,5.0138187,6.560595,8.831716,6.466279,4.6214657,4.3347464,5.330719,6.039973,5.613666,5.194905,5.987156,7.986647,9.978593,11.7555,11.921495,13.177779,14.479335,11.012292,6.485142,3.8593953,2.1164427,0.9016574,0.55080324,0.6187105,0.7432071,0.7809334,0.67152727,0.4640329,0.35462674,0.46026024,0.6451189,0.7884786,0.79602385,1.0525624,1.7957695,2.4333432,2.4974778,1.6675003,0.965792,1.3958713,2.2598023,2.886058,2.6332922,1.2185578,0.8526133,1.6260014,2.4974778,1.2600567,1.3468271,1.9957186,2.1051247,1.7882242,2.372981,2.1654868,1.539231,1.056335,0.97333723,1.2562841,1.1355602,0.8978847,0.76207024,0.724344,0.55080324,0.35462674,0.331991,0.35839936,0.35839936,0.29426476,0.19994913,0.150905,0.2263575,0.38103512,0.4376245,0.84884065,1.2147852,1.5430037,2.637065,6.096562,5.1534057,3.9084394,3.1312788,2.704972,1.6637276,0.95447415,0.5093044,0.3734899,0.35085413,0.0,0.0,0.03772625,0.124496624,0.452715,1.3656902,1.3091009,1.3468271,1.1657411,0.8111144,0.6790725,0.21881226,0.049044125,0.124496624,0.30935526,0.38103512,0.24522063,0.19994913,0.19994913,0.1961765,0.14713238,0.030181,0.0,0.0,0.0150905,0.071679875,0.08299775,0.18485862,0.27540162,0.33576363,0.41876137,0.70170826,0.49421388,0.3169005,0.3470815,0.4376245,0.38103512,0.482896,0.5885295,0.573439,0.33576363,0.44139713,0.271629,0.11317875,0.060362,0.0,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.00754525,0.0,0.00754525,0.030181,0.06413463,0.1056335,0.10940613,0.090543,0.049044125,0.018863125,0.060362,0.12826926,0.120724,0.07922512,0.033953626,0.011317875,0.02263575,0.033953626,0.026408374,0.011317875,0.0,0.011317875,0.041498873,0.060362,0.06413463,0.07922512,0.033953626,0.018863125,0.033953626,0.060362,0.06413463,0.033953626,0.011317875,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.120724,0.482896,0.513077,0.31312788,0.14335975,0.094315626,0.09808825,0.14713238,0.26408374,0.422534,0.5319401,0.422534,1.0487897,2.474842,4.085753,5.3986263,6.0701537,5.485397,3.9612563,2.4672968,1.5128226,1.1506506,0.9016574,0.49421388,0.22258487,0.14713238,0.1056335,0.094315626,0.094315626,0.124496624,0.18485862,0.26031113,0.42630664,0.6526641,1.2600567,2.2673476,3.380272,6.168242,8.379,9.484379,9.476834,8.892077,7.2358947,6.3153744,5.4212623,4.504514,4.1800685,4.357382,3.8895764,2.9954643,1.9881734,1.3015556,0.8601585,0.55457586,0.3169005,0.15467763,0.13204187,0.18863125,0.2867195,0.43007925,0.6111652,0.79602385,1.2110126,1.6825907,2.1805773,2.7238352,3.380272,4.134797,4.8666863,5.5985756,6.356873,7.194396,7.967784,8.820397,9.805053,10.880251,11.92904,13.166461,14.407655,14.977322,14.762281,14.226569,13.8870325,13.849306,13.9888935,14.1926155,14.34352,14.535924,15.049001,16.22606,18.41041,21.96045,24.337204,24.971004,24.35984,23.1526,22.152855,21.420965,20.474035,19.595015,19.032892,19.036665,19.76101,20.677757,21.319103,21.794455,22.764019,23.75622,25.091728,26.710184,28.35505,29.57738,31.060022,33.06706,34.843964,35.722984,35.142002,34.278072,34.040394,33.67445,33.123646,33.018013,35.87389,39.02026,42.132675,45.305454,49.07808,53.36001,57.50235,61.173115,64.3723,67.44699,71.27621,71.39316,70.129326,68.83154,67.86575,67.33004,67.137634,68.51842,71.91,76.94269,82.56767,85.66877,84.48039,78.17256,66.850914,54.963375,46.690006,41.43097,38.424187,36.730278,36.52278,36.74914,37.069813,37.26222,37.22072,37.658344,38.563774,40.178455,42.4873,45.180958,47.346443,48.036835,47.161587,45.094185,42.649525,40.318043,39.212666,39.5522,41.03107,42.804203,43.713406,43.800175,43.155056,41.98177,40.5859,40.393497,40.97448,41.510193,41.50642,40.778305,40.246365,38.952354,38.212917,38.541138,39.65406,40.929207,43.094696,45.28659,46.999363,48.067017,45.63367,43.694542,43.139965,44.44152,47.6558,0.2867195,0.7205714,1.0374719,1.6750455,2.9501927,5.0553174,6.0022464,5.2137675,3.429316,1.5656394,0.73188925,0.9242931,1.3958713,2.4899325,3.8367596,4.357382,3.399135,3.187868,3.7348988,4.927048,6.5455046,5.1798143,5.4212623,4.8440504,3.3463185,3.1237335,4.957229,7.01331,7.0548086,5.3382645,4.6290107,5.6098933,6.387054,6.8359966,6.688864,5.5004873,6.205968,5.983383,4.6516466,3.3236825,4.4101987,4.3913355,3.772625,5.0025005,7.6886096,8.631766,7.175533,5.8513412,5.3458095,5.0477724,3.029418,1.5165952,0.98465514,0.8639311,0.784706,0.5772116,0.40367088,0.27540162,0.59230214,2.3088465,6.930312,8.873214,7.779153,6.8925858,6.273875,2.8219235,3.1539145,5.198677,7.61693,8.507269,5.379763,3.1916409,2.5502944,2.9237845,3.6330378,3.8669407,3.7952607,4.4516973,5.160951,6.0701537,8.152642,7.6018395,7.1679873,6.651138,6.0362,5.515578,4.5196047,4.5309224,6.326692,9.590013,12.887287,13.392818,12.566614,12.396846,12.725064,11.219787,8.099826,5.3269467,2.938875,1.1846043,0.5093044,0.47157812,0.4979865,0.47912338,0.38858038,0.2867195,0.27917424,0.33953625,0.43385187,0.513077,0.51684964,0.6111652,1.3543724,2.1353056,2.4786146,2.0636258,1.7429527,2.4220252,3.5839937,4.5196047,4.3347464,2.987919,2.263575,2.5917933,2.9501927,0.8639311,0.8526133,1.2525115,1.4939595,1.4373702,1.3807807,1.1808317,0.935611,0.8526133,1.026154,1.4298248,2.071171,1.8523588,1.2449663,0.6752999,0.51684964,0.7167987,1.1431054,1.5505489,1.7957695,1.8297231,1.7316349,1.6146835,2.2560298,3.4670424,4.08198,2.4559789,2.052308,2.4597516,3.3350005,4.3913355,2.6936543,1.629774,0.97333723,0.5093044,0.03772625,0.24522063,0.35085413,0.35839936,0.2565385,0.0,0.0,0.0,0.00754525,0.150905,0.6790725,0.9620194,1.3656902,1.6712729,1.7542707,1.5920477,0.8978847,0.6073926,0.5055317,0.4678055,0.42630664,0.24522063,0.12826926,0.090543,0.09808825,0.071679875,0.03772625,0.0754525,0.116951376,0.12826926,0.1358145,0.19240387,0.271629,0.26031113,0.18863125,0.2565385,0.6111652,0.5470306,0.42630664,0.35085413,0.1659955,0.15467763,0.26408374,0.33576363,0.3055826,0.1961765,0.18863125,0.0754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.018863125,0.018863125,0.011317875,0.0,0.0,0.003772625,0.011317875,0.0150905,0.02263575,0.0150905,0.011317875,0.00754525,0.003772625,0.026408374,0.060362,0.06413463,0.049044125,0.041498873,0.060362,0.05281675,0.06790725,0.0754525,0.05281675,0.018863125,0.02263575,0.026408374,0.026408374,0.030181,0.0452715,0.0150905,0.00754525,0.0150905,0.030181,0.02263575,0.011317875,0.003772625,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.030181,0.13204187,0.1961765,0.13204187,0.071679875,0.056589376,0.071679875,0.120724,0.20749438,0.3169005,0.52062225,0.95447415,2.5012503,3.4896781,3.9084394,3.9499383,4.0216184,5.05909,4.9119577,4.1197066,2.9426475,1.3656902,0.79602385,0.41121614,0.19994913,0.116951376,0.0754525,0.06413463,0.124496624,0.16222288,0.21503963,0.47157812,1.5920477,2.5616124,3.6443558,4.817642,5.7570257,7.0246277,7.937603,7.7829256,6.719045,5.775889,4.9345937,4.61392,4.3875628,4.1272516,3.983892,4.3611546,4.22534,3.5538127,2.5389767,1.6033657,0.814887,0.5017591,0.35085413,0.21881226,0.124496624,0.10940613,0.1056335,0.14713238,0.24899325,0.40367088,0.6526641,0.9620194,1.20724,1.3656902,1.5430037,2.0258996,2.6031113,3.2444575,3.942393,4.719554,5.481624,6.258785,6.9793563,7.6093845,8.137552,9.186342,10.408672,11.291467,11.668729,11.747954,11.838497,12.049765,12.359119,12.67602,12.868423,12.958967,13.287186,14.162435,15.769572,18.168962,19.68933,19.828917,19.557287,19.470518,19.768555,19.821371,19.478064,19.319613,19.425245,19.383747,19.998686,20.987112,21.83218,22.322622,22.575388,23.073374,24.148573,25.563307,27.1629,28.90208,31.218472,33.05574,33.821583,33.289642,31.580645,30.36963,30.682758,31.433512,32.07486,32.606796,33.85931,35.017506,36.568054,38.895763,42.26849,46.901276,51.37938,55.9518,60.53177,64.67788,67.75635,69.12203,69.6087,69.42384,68.133606,67.167816,66.77169,66.99805,67.929886,69.71056,74.70929,80.22487,85.07647,87.83803,86.81942,80.91904,72.99275,64.14217,55.412315,47.78784,42.264717,39.039124,37.02077,35.572083,34.53461,34.527065,35.089184,35.575855,36.122883,37.605526,41.06502,44.31325,46.316517,46.788094,46.199566,43.339916,41.038616,40.280315,41.04239,42.306217,45.460133,48.100967,49.342163,48.813995,46.663597,44.071804,42.962654,42.362804,41.717686,40.883938,40.480267,39.80874,39.340935,39.23907,39.3598,40.551945,42.389214,44.015217,45.120594,45.924164,44.49811,43.336143,43.083378,43.841675,45.162094,0.17731337,0.3734899,0.4376245,0.4979865,0.7696155,1.5807298,3.8443048,4.496969,3.4481792,1.9429018,2.5691576,4.183841,3.361409,3.2067313,4.2894745,4.6327834,3.500996,3.5764484,4.689373,6.1342883,6.700182,4.9345937,5.0968165,4.98741,4.285702,4.52715,5.915476,7.5716586,7.877241,6.458734,4.214022,3.3010468,3.9197574,5.66271,6.8133607,4.346064,5.802297,5.6815734,4.644101,3.5953116,3.7273536,4.093298,3.3538637,3.6443558,5.3344917,7.009537,7.2094865,5.9796104,4.949684,4.1310244,1.9391292,1.3091009,1.237421,1.1016065,0.7922512,0.724344,0.8978847,0.83752275,0.8865669,1.4977322,3.2520027,3.5538127,3.572676,3.2331395,2.5125682,1.448688,1.7957695,1.6976813,1.81086,2.5276587,3.9461658,4.044254,3.7273536,3.904667,4.4403796,4.115934,4.8930945,5.409944,4.98741,4.29702,5.3609,6.7114997,7.1340337,7.594294,8.047009,7.443389,5.4174895,4.4630156,5.96452,9.593785,13.309821,13.151371,12.038446,11.536687,12.004493,12.596795,10.842525,7.8734684,4.930821,2.704972,1.3505998,1.3241913,1.5807298,1.3958713,0.73566186,0.26408374,0.28294688,0.35462674,0.6187105,0.845068,0.44894236,0.2867195,0.9507015,1.5580941,1.7089992,1.4901869,1.5241405,2.2069857,3.3764994,4.5196047,4.776143,3.9688015,3.059599,2.6144292,2.2107582,0.422534,0.55457586,1.1129243,1.6825907,1.9881734,1.8787673,1.327964,1.0299267,1.026154,1.2336484,1.4222796,2.9049213,2.746471,1.841041,1.0525624,1.2185578,1.8749946,2.1994405,2.2748928,2.2598023,2.3805263,2.4107075,2.463524,3.1765501,4.255521,4.4743333,3.048281,2.2673476,2.3993895,2.757789,1.7240896,0.55080324,0.15467763,0.06790725,0.06413463,0.13958712,0.23013012,0.26408374,0.20372175,0.07922512,0.0,0.0,0.0,0.018863125,0.124496624,0.42630664,1.0827434,1.6184561,2.474842,3.4066803,3.5085413,2.3277097,1.4562333,0.8262049,0.41876137,0.26408374,0.52062225,0.69793564,0.6187105,0.32067314,0.06790725,0.06413463,0.16222288,0.27540162,0.3470815,0.34330887,0.29803738,0.24522063,0.16976812,0.094315626,0.10940613,0.30935526,0.32821837,0.29049212,0.211267,0.03772625,0.056589376,0.14713238,0.17354076,0.13958712,0.17731337,0.094315626,0.060362,0.056589376,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.00754525,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.02263575,0.018863125,0.018863125,0.0150905,0.00754525,0.0,0.0,0.003772625,0.0150905,0.026408374,0.0150905,0.003772625,0.00754525,0.00754525,0.0,0.00754525,0.018863125,0.030181,0.0452715,0.06790725,0.09808825,0.071679875,0.10186087,0.120724,0.09808825,0.030181,0.02263575,0.00754525,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.00754525,0.00754525,0.00754525,0.011317875,0.018863125,0.033953626,0.08299775,0.18863125,0.44516975,1.0638802,2.384299,3.7877154,3.6443558,2.8634224,2.203213,2.282438,4.085753,5.3344917,5.6400743,4.768598,2.674791,1.3392819,0.60362,0.241448,0.094315626,0.06413463,0.08299775,0.17354076,0.5093044,1.1506506,2.0598533,3.361409,4.2706113,5.028909,5.66271,5.983383,5.847569,5.794752,5.3458095,4.6252384,4.3686996,4.3121104,4.353609,4.4894238,4.538468,4.168751,4.2630663,4.032936,3.4217708,2.5314314,1.6260014,1.2223305,1.2223305,1.0638802,0.66775465,0.43007925,0.35839936,0.23390275,0.14335975,0.120724,0.18485862,0.33953625,0.59607476,0.7092535,0.633801,0.5017591,0.7130261,1.0676528,1.5430037,2.1088974,2.704972,3.308592,3.9348478,4.478106,4.881777,5.160951,5.8966126,6.94163,7.9941926,8.858124,9.435335,9.842778,10.242677,10.661438,11.057564,11.314102,11.446144,11.717773,12.381755,13.460726,14.750964,15.448899,15.520579,15.724301,16.32792,17.13149,17.293713,17.554024,18.41041,19.628967,20.270313,20.568352,21.326649,22.213217,22.869654,22.926243,23.250689,24.114618,25.306768,26.763002,28.57009,30.799711,31.984314,31.927725,30.701622,28.65686,27.426983,27.498663,28.468227,29.924461,31.448603,31.874908,31.697596,32.089947,33.632954,36.34547,40.193546,44.286846,49.11958,54.672882,60.38841,64.296844,66.98673,68.45805,68.80136,68.201515,67.458305,66.93768,66.46611,65.968124,65.45882,67.20931,70.15573,74.79229,80.64363,86.24221,88.652916,87.68335,84.29931,78.606415,69.86147,59.87533,51.371834,44.32457,38.8769,35.349495,34.213936,33.991352,33.851765,33.644268,33.915897,36.183247,38.967445,41.54792,43.596455,45.180958,44.56225,43.31728,42.18172,41.81955,42.830612,45.705353,49.417614,52.752617,54.665337,54.291847,51.213383,48.810223,46.501377,44.15103,42.060997,40.774532,40.129414,39.642742,39.23907,39.295662,40.076595,40.93298,41.800686,42.51371,42.804203,41.446056,41.427197,41.446056,41.114067,40.96316,0.1358145,0.3772625,0.47535074,0.452715,0.4376245,0.66775465,1.026154,1.5203679,1.5807298,1.8221779,4.0480266,7.073672,5.2892203,4.402653,5.553304,5.3382645,4.0480266,4.3649273,5.040227,5.0741806,3.731126,3.904667,4.7836885,5.2062225,5.0439997,5.198677,5.6589375,6.670001,7.9036493,8.582722,7.5112963,5.3609,5.5985756,7.9451485,9.020347,2.3390274,2.5125682,2.9803739,2.9351022,2.6710186,3.5689032,4.395108,3.500996,2.6483827,2.6332922,3.3161373,3.2482302,2.5125682,1.6109109,1.0601076,1.3845534,1.8825399,2.1843498,2.1088974,1.7957695,1.7052265,2.2296214,2.5238862,2.686109,2.6068838,1.9844007,0.7809334,0.7394345,0.65643674,0.29426476,0.392353,2.1692593,2.535204,2.463524,3.0369632,5.451443,6.620957,6.4964604,6.692637,7.488661,7.805561,8.16396,6.9680386,4.8138695,2.8747404,2.897376,4.538468,4.285702,5.7117543,8.66572,9.273112,6.6020937,4.9119577,5.7796617,8.590267,10.533169,10.650121,10.446399,11.02361,12.630749,14.671739,13.687083,10.978339,8.107371,5.6891184,3.4029078,3.0860074,3.531177,3.2105038,1.9693103,1.0186088,0.9280658,0.95824677,1.4826416,2.071171,1.4864142,1.1091517,1.3619176,1.4071891,1.0336993,0.6451189,0.7167987,1.0902886,1.8674494,2.8521044,3.5764484,3.3651814,2.7728794,2.161714,1.659955,1.1619685,1.6373192,2.2409391,2.886058,3.6858547,4.9421387,3.6330378,2.1654868,1.4335974,1.4411428,1.3166461,2.848332,2.8709676,2.335255,1.9542197,2.203213,2.8332415,2.7502437,2.2748928,1.8221779,1.8749946,1.8825399,2.0862615,2.3314822,2.3692086,1.8599042,2.6295197,2.04099,1.6976813,1.7655885,0.95824677,0.87902164,0.73188925,0.5281675,0.3772625,0.482896,0.38858038,0.28294688,0.24899325,0.3055826,0.4376245,0.32821837,0.19240387,0.1358145,0.26408374,0.6752999,1.5015048,1.9994912,3.1652324,4.7535076,5.311856,4.0593443,2.7389257,1.7089992,1.0336993,0.5093044,0.97710985,1.4109617,1.3053282,0.7092535,0.2565385,0.116951376,0.18863125,0.3470815,0.47912338,0.5017591,0.29426476,0.09808825,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.071679875,0.11317875,0.150905,0.12826926,0.08677038,0.19240387,0.15467763,0.124496624,0.10940613,0.08677038,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.003772625,0.0,0.0,0.003772625,0.0150905,0.033953626,0.018863125,0.00754525,0.011317875,0.011317875,0.02263575,0.02263575,0.018863125,0.0150905,0.02263575,0.011317875,0.011317875,0.011317875,0.003772625,0.003772625,0.0,0.0150905,0.041498873,0.06413463,0.041498873,0.011317875,0.003772625,0.0,0.0,0.003772625,0.003772625,0.011317875,0.026408374,0.033953626,0.0150905,0.003772625,0.0150905,0.0150905,0.0,0.0,0.02263575,0.060362,0.1056335,0.13204187,0.08677038,0.08299775,0.12826926,0.16222288,0.1358145,0.041498873,0.011317875,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.00754525,0.0150905,0.0150905,0.090543,0.4376245,1.3355093,2.7502437,4.349837,4.221567,2.9652832,1.8448136,1.4901869,1.9089483,3.108643,5.0779533,6.3719635,6.270103,4.7874613,2.9086938,1.5052774,0.59230214,0.13958712,0.06790725,0.16222288,0.32821837,1.1242423,2.5880208,4.255521,5.010046,5.1043615,5.040227,4.90064,4.327201,3.7952607,3.7575345,4.0404816,4.5497856,5.2892203,5.379763,5.3458095,5.27413,5.0025005,4.0970707,3.7084904,3.399135,2.969056,2.4333432,2.003264,2.4182527,2.7653341,2.625747,1.9391292,1.0148361,0.9016574,0.7167987,0.55080324,0.44516975,0.38858038,0.362172,0.5281675,0.58475685,0.4376245,0.21881226,0.20372175,0.29803738,0.5394854,0.8903395,1.2449663,1.6486372,2.1390784,2.6219745,3.0445085,3.380272,3.9461658,4.727099,5.621211,6.515323,7.284939,7.8395147,8.397863,8.948667,9.420244,9.654147,9.839006,10.163452,10.733118,11.52537,12.3893,12.679792,13.034419,13.59654,14.2944765,14.822643,14.894323,15.539442,17.154125,19.425245,21.31533,21.492645,21.93027,22.496162,22.982832,23.129965,23.511,24.242887,25.344494,26.755457,28.321096,29.566063,29.882963,29.388748,28.290915,26.895044,26.340467,25.963205,26.223516,27.189308,28.505955,28.736084,28.483318,28.58518,29.622652,31.92018,34.685513,37.677204,41.51774,46.573055,52.929928,58.72468,63.01793,65.74176,67.220634,68.19774,67.7073,66.899956,66.21712,65.86626,65.8059,65.27396,64.64393,64.97592,66.783005,70.05765,75.8939,82.36395,88.656685,92.50099,90.158195,81.99423,72.109955,61.622055,51.760414,43.856766,38.725994,35.651306,34.345978,34.24789,34.49311,35.115593,35.65885,36.43224,37.745113,39.91437,42.562756,44.083122,43.985035,43.34369,44.81124,45.494083,48.11983,52.18672,56.574284,59.516933,59.034035,57.253357,54.163578,50.134415,45.912846,42.374123,40.31427,39.069305,38.567547,39.30698,39.959644,39.91437,40.182228,40.721714,40.44254,38.31101,38.820312,39.197575,38.86181,39.439022,0.0150905,0.041498873,0.10186087,0.25276586,0.41121614,0.35085413,0.38858038,0.55080324,0.6073926,0.5470306,0.59607476,0.8639311,1.1317875,1.6033657,2.04099,1.7844516,0.663982,0.7922512,1.478869,1.9089483,1.1921495,0.5055317,0.482896,1.0072908,1.6712729,1.7542707,1.327964,1.6071383,3.218049,5.5683947,6.851087,5.6778007,6.9793563,8.311093,7.356619,1.9240388,2.7389257,3.8971217,3.6028569,2.7389257,4.851596,3.2520027,2.9351022,2.2296214,1.2789198,2.0598533,1.2789198,0.8262049,0.80734175,1.1431054,1.5580941,1.5580941,1.5656394,1.5543215,1.5354583,1.5731846,2.535204,4.617693,5.80607,4.82896,1.1280149,0.8865669,1.9693103,1.7165444,0.15845025,0.0,0.14713238,0.120724,0.10186087,0.21503963,0.52062225,0.7507524,1.0638802,1.4750963,2.0447628,2.9011486,3.6556737,4.1310244,4.1762958,3.7763977,3.006782,2.5314314,1.6863633,1.2223305,1.4826416,2.4107075,2.9351022,3.3689542,4.847823,7.322665,9.582467,14.305794,14.332202,12.826925,11.853588,12.3893,13.072145,13.309821,12.355347,9.993684,6.515323,4.5497856,4.104616,4.134797,4.0593443,3.7537618,3.4368613,2.9728284,3.1539145,4.063117,5.0515447,4.4403796,2.9049213,1.6712729,1.1242423,0.7922512,0.98842776,0.7809334,0.55457586,0.5357128,0.7922512,1.1959221,2.0108092,2.867195,3.591539,4.22534,4.7874613,3.2520027,2.7540162,4.5988297,8.284684,6.2361493,2.516341,0.5885295,0.98842776,1.3430545,1.026154,1.7165444,2.8747404,3.5953116,2.595566,1.7391801,1.8938577,2.4371157,2.8294687,2.6106565,1.7655885,1.1996948,1.297783,2.082489,3.2029586,2.9954643,1.9655377,1.4034165,1.4713237,1.1883769,1.629774,2.123988,1.9579924,1.3355093,1.3732355,1.0450171,0.7507524,0.90920264,1.5241405,2.1805773,1.6448646,0.9620194,0.5583485,0.51684964,0.56589377,1.0789708,1.7995421,2.6597006,3.5047686,4.0895257,4.9685473,4.98741,4.7308717,4.0970707,2.305074,1.0336993,0.5055317,0.32821837,0.34330887,0.6111652,0.15845025,0.10940613,0.15845025,0.150905,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.1056335,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.041498873,0.030181,0.018863125,0.00754525,0.00754525,0.0150905,0.0150905,0.0150905,0.0150905,0.033953626,0.060362,0.060362,0.071679875,0.056589376,0.033953626,0.02263575,0.0452715,0.0452715,0.06413463,0.05281675,0.0150905,0.0150905,0.003772625,0.03772625,0.12826926,0.19994913,0.0754525,0.041498873,0.011317875,0.0,0.003772625,0.0150905,0.0150905,0.02263575,0.018863125,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.02263575,0.1056335,0.20749438,0.23390275,0.0150905,0.0754525,0.15467763,0.19994913,0.17354076,0.0754525,0.026408374,0.00754525,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.00754525,0.0150905,0.0150905,0.19994913,1.3317367,3.6971724,6.058836,5.692891,3.5424948,1.9806281,1.448688,1.8334957,2.4559789,3.187868,5.093044,6.722818,7.303802,6.730363,5.3873086,3.5387223,1.7089992,0.4074435,0.150905,0.38480774,0.8639311,1.7052265,2.9237845,4.425289,5.670255,5.753253,5.832478,5.7683434,4.1197066,2.8747404,3.0746894,3.9989824,5.1534057,6.300284,6.217286,6.058836,5.613666,4.8063245,3.7084904,3.3312278,3.410453,3.682082,3.9197574,3.9197574,4.4705606,4.323428,4.678055,4.749735,1.7693611,1.659955,1.6033657,1.629774,1.7052265,1.7542707,1.0827434,0.9507015,0.98842776,0.9393836,0.67152727,0.3055826,0.11317875,0.094315626,0.21881226,0.42630664,0.73188925,1.1091517,1.5316857,1.9655377,2.3805263,2.757789,3.2029586,3.7688525,4.5007415,5.4174895,6.0512905,6.722818,7.4811153,8.107371,8.118689,8.058327,8.333729,8.835487,9.461743,10.133271,10.902886,11.9064045,12.989148,13.747445,13.5663595,14.079436,14.728328,16.388283,19.010258,21.620914,22.209444,22.499935,22.439573,22.213217,22.26226,22.945105,23.922215,25.046457,26.159382,27.098766,27.513754,27.362848,26.868635,26.393284,26.44233,26.600779,26.212198,25.767029,25.63876,26.076384,25.174726,25.114365,25.74062,27.027086,29.052984,32.07863,33.97249,35.779575,38.537365,43.27578,49.19503,54.65779,59.67538,63.78,66.02471,66.745285,67.895935,68.103424,67.37908,67.12254,65.09664,64.194984,63.82527,63.22165,61.463608,63.734726,67.60544,71.43843,75.98821,84.39739,88.7925,90.05256,86.03094,76.7201,64.26667,53.06197,44.400024,38.737312,35.95689,35.38345,36.00593,36.89627,37.55648,37.533848,36.424694,37.545162,40.34445,42.932472,44.48302,45.226227,45.177185,45.89021,48.45937,52.865795,57.966385,62.03327,64.651474,64.19876,60.196003,53.299644,47.03709,42.185493,39.065533,37.877155,38.695816,40.01623,39.99737,39.789875,39.72197,39.30698,37.779068,37.635708,40.031322,43.830357,45.637444,0.026408374,0.05281675,0.09808825,0.12826926,0.13204187,0.120724,0.17354076,0.20749438,0.23013012,0.35462674,0.754525,0.9620194,1.0940613,1.6675003,2.293756,1.6863633,0.8299775,0.935611,1.5430037,2.4408884,3.6934,4.8440504,4.2328854,3.0633714,2.2862108,2.595566,3.1765501,2.8709676,2.425798,2.2069857,2.1881225,3.0558262,5.330719,6.688864,6.790725,7.2585306,9.461743,8.114917,5.2062225,2.9803739,3.9499383,5.4740787,6.3417826,6.579458,6.277648,5.564622,5.7796617,6.439871,6.930312,6.515323,4.3649273,3.0860074,2.8256962,2.9237845,3.1463692,3.6707642,3.9122121,5.828706,6.670001,5.5268955,3.3010468,5.7419353,6.488915,4.274384,0.77716076,0.5998474,1.1431054,1.6561824,3.4066803,6.119198,7.9753294,4.274384,3.470815,4.1498876,4.5761943,2.71629,2.584248,3.4594972,4.5837393,5.847569,7.752744,8.303548,7.3792543,6.0626082,5.270357,5.7796617,5.523123,5.50426,5.492942,5.828706,7.4207535,9.774872,10.687846,11.45369,12.057309,11.170743,14.879233,13.060828,9.876732,7.462252,5.904158,5.5004873,4.8968673,4.025391,3.0860074,2.546522,2.6974268,4.025391,6.085244,7.9753294,8.360137,8.66572,6.3116016,5.511805,6.1606965,3.8556228,2.04099,3.1312788,5.409944,7.2660756,7.1906233,5.1798143,4.06689,3.3312278,2.7238352,2.2748928,2.2409391,1.5279131,1.0714256,1.2600567,1.9391292,1.539231,0.84129536,0.6790725,1.026154,0.98842776,0.6111652,1.6109109,2.7841973,3.591539,4.142342,3.7084904,3.482133,2.8898308,2.0900342,1.9994912,2.0145817,2.2484846,2.565385,2.5540671,1.50905,0.87902164,0.52062225,0.392353,0.41498876,0.44516975,0.56212115,1.6788181,2.6898816,3.4066803,4.5460134,3.651901,2.0296721,4.014073,8.141325,7.149124,3.429316,1.4675511,0.69793564,0.66775465,1.0299267,1.7052265,2.252257,2.8143783,3.5802212,4.7610526,6.643593,7.8244243,7.5565677,5.794752,3.169005,1.1016065,0.31312788,0.11317875,0.08677038,0.120724,0.030181,0.02263575,0.030181,0.030181,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.018863125,0.00754525,0.00754525,0.0150905,0.02263575,0.05281675,0.060362,0.049044125,0.049044125,0.060362,0.049044125,0.041498873,0.03772625,0.02263575,0.003772625,0.00754525,0.03772625,0.041498873,0.041498873,0.041498873,0.041498873,0.0452715,0.049044125,0.05281675,0.05281675,0.026408374,0.030181,0.026408374,0.0452715,0.06790725,0.041498873,0.030181,0.03772625,0.0452715,0.041498873,0.0150905,0.003772625,0.00754525,0.00754525,0.003772625,0.011317875,0.026408374,0.05281675,0.08299775,0.10940613,0.11317875,0.1659955,0.1659955,0.14335975,0.09808825,0.041498873,0.06790725,0.06790725,0.03772625,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.011317875,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.00754525,0.026408374,0.56212115,1.871222,3.2821836,4.0404816,3.3236825,2.2598023,1.4864142,1.2110126,1.5203679,2.4069347,3.1312788,4.323428,6.013564,7.756517,8.60913,8.035691,6.851087,5.0062733,2.848332,1.1280149,0.9318384,1.8146327,2.7313805,3.0709167,2.6672459,2.886058,3.3727267,4.3611546,5.617439,6.439871,4.5799665,4.217795,4.357382,4.61392,5.20245,6.307829,6.858632,6.730363,6.058836,5.2326307,3.99521,3.6783094,3.9989824,4.5535583,4.7874613,4.82896,4.564876,4.696918,4.930821,3.942393,4.3913355,4.715781,4.9459114,5.032682,4.8553686,3.482133,3.078462,2.4182527,1.3920987,1.026154,0.66020936,0.39989826,0.2565385,0.21881226,0.27917424,0.41121614,0.6111652,0.87902164,1.1695137,1.4298248,1.7089992,2.0447628,2.505023,3.1350515,3.9650288,4.727099,6.0286546,7.224577,7.77538,7.250985,6.8963585,7.0510364,7.492433,8.043237,8.5563135,9.190115,9.955957,11.038701,12.313848,13.381501,13.924759,14.324657,15.154634,16.735365,19.1423,20.82489,21.21347,20.836208,20.258997,20.115637,21.100292,22.066084,22.847017,23.533634,24.476791,25.242634,25.442583,25.634987,26.182018,27.238352,27.279852,27.10631,26.729048,26.1707,25.46522,23.850534,23.371412,23.303505,23.624178,24.989868,27.819336,30.78462,33.88572,36.869865,39.2353,41.510193,44.996098,49.538338,54.42766,58.370052,60.9958,63.84413,65.96058,66.97919,67.12254,64.851425,63.10847,61.373062,59.91306,59.777245,61.354202,62.470898,62.527485,62.614258,65.489,69.367256,73.158745,75.576996,76.05989,74.780975,71.755325,66.27747,59.022717,51.22093,44.660336,41.10652,39.56352,39.227757,39.288116,38.94858,37.514984,38.390232,39.80874,41.77805,46.10525,49.02526,50.553177,50.84744,50.522995,50.655037,52.828068,56.363018,59.3698,60.50536,58.988766,55.17464,50.077824,45.045143,41.01598,38.51473,38.122375,37.126404,36.775547,36.722733,35.047688,33.11233,31.508965,32.06354,34.715694,37.560253,1.1016065,0.62625575,0.29426476,0.16976812,0.25276586,0.47157812,0.4678055,0.331991,0.24899325,0.36971724,0.8299775,0.8941121,0.9205205,1.3543724,1.9202662,1.6373192,1.4222796,1.690136,2.2296214,3.029418,4.3007927,5.794752,7.6584287,8.6581745,8.311093,6.888813,6.5266414,6.047518,5.1043615,4.085753,4.0895257,4.3611546,5.100589,5.2967653,5.2175403,6.4134626,5.873977,4.5724216,2.8294687,1.4411428,1.7089992,2.8898308,3.4670424,3.610402,3.3878171,2.7691069,2.9086938,3.270866,3.5274043,3.3123648,2.1994405,1.5316857,1.4260522,1.5618668,1.841041,2.4031622,2.969056,5.451443,6.7756343,6.2663302,5.6476197,7.7150183,7.5188417,5.2364035,2.4031622,1.9202662,2.003264,1.8938577,2.5389767,4.032936,5.613666,3.7801702,3.3425457,4.1008434,5.062863,4.45547,4.1083884,4.8327327,4.7421894,3.9122121,4.353609,4.7006907,4.5535583,4.2064767,3.9273026,3.9499383,3.4896781,3.380272,3.380272,3.6066296,4.538468,5.9682927,7.6508837,9.695646,11.442371,11.487643,12.887287,10.0276375,6.9454026,5.2665844,4.1762958,3.7198083,3.270866,2.505023,1.5505489,0.98842776,1.116697,2.3805263,4.5535583,6.8963585,8.13378,8.963757,7.6093845,6.6020937,6.8963585,7.865923,5.772116,5.036454,5.4891696,6.5341864,7.149124,4.9421387,4.851596,4.5309224,3.289729,2.123988,1.8372684,1.4562333,1.0638802,0.7205714,0.47912338,0.4979865,0.73566186,1.3505998,2.3805263,3.712263,2.6106565,2.2371666,2.5012503,2.8596497,2.3428001,2.0598533,2.1051247,1.8787673,1.3430545,1.0412445,1.3091009,1.9429018,2.4672968,2.4710693,1.6222287,1.6146835,2.1277604,2.3126192,2.033445,1.8334957,1.6146835,1.9051756,2.625747,3.4934506,4.032936,3.8858037,2.746471,4.134797,7.2472124,6.9189944,3.7499893,1.9994912,1.2298758,1.0638802,1.2185578,1.9466745,2.4861598,2.8445592,3.338773,4.5912848,6.1833324,7.0812173,6.6247296,4.8100967,2.3163917,0.7432071,0.17354076,0.05281675,0.041498873,0.018863125,0.003772625,0.033953626,0.06413463,0.0754525,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.003772625,0.00754525,0.011317875,0.033953626,0.03772625,0.033953626,0.030181,0.033953626,0.026408374,0.02263575,0.033953626,0.030181,0.0150905,0.00754525,0.030181,0.0452715,0.05281675,0.049044125,0.026408374,0.033953626,0.030181,0.02263575,0.018863125,0.02263575,0.030181,0.026408374,0.03772625,0.06413463,0.071679875,0.060362,0.0452715,0.030181,0.02263575,0.0150905,0.003772625,0.00754525,0.00754525,0.0,0.00754525,0.011317875,0.02263575,0.03772625,0.060362,0.10186087,0.1358145,0.13958712,0.16222288,0.18863125,0.13204187,0.07922512,0.0452715,0.02263575,0.0150905,0.033953626,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.011317875,0.056589376,0.694163,1.6486372,2.2862108,2.3578906,1.9994912,1.5656394,1.0487897,0.7205714,0.7997965,1.4524606,2.2258487,3.1199608,4.4705606,6.3644185,8.612903,10.431308,10.544487,9.955957,9.574923,10.18986,9.963503,8.710991,6.4134626,3.6783094,1.750498,1.4864142,1.8033148,2.516341,3.3312278,3.8443048,3.410453,3.663219,3.863168,3.8707132,4.168751,5.142088,5.4288073,5.119452,4.38379,3.482133,3.0030096,3.3274553,4.142342,5.2288585,6.488915,6.85486,6.820906,6.488915,6.009792,5.6023483,6.1305156,6.470052,6.3945994,5.9607477,5.492942,4.0291634,2.8181508,1.9089483,1.2751472,0.8111144,0.5055317,0.30935526,0.22258487,0.19994913,0.18863125,0.18863125,0.27540162,0.422534,0.59607476,0.7432071,0.9016574,1.1506506,1.5316857,2.0560806,2.7313805,3.5047686,4.7120085,5.8098426,6.3908267,6.2021956,6.0739264,6.326692,6.6586833,6.9491754,7.2472124,7.6848373,8.280911,9.333474,10.944386,13.041965,14.083209,14.120935,13.973803,14.347293,15.833707,17.448391,18.010511,17.840744,17.542706,17.991648,19.979822,21.1682,21.466236,21.353058,21.90386,22.899834,23.616632,24.299479,25.19359,26.529099,27.442074,28.200373,28.434275,27.898561,26.438557,23.488363,22.152855,21.752956,22.013268,23.046967,24.650331,27.581661,31.678732,35.95689,38.627907,38.63168,40.216183,43.438004,47.546394,51.002117,54.276756,57.713615,60.441227,62.184177,63.240513,62.82175,61.6296,59.48298,56.940228,55.272728,55.672626,55.480225,54.714382,54.14094,55.25009,56.989273,59.188713,61.701283,64.17235,66.0398,68.216606,69.10694,68.36374,65.96058,62.18795,56.619556,50.738033,46.120342,43.294643,41.77805,39.00894,38.454365,38.725994,39.937008,43.736042,48.538593,52.54512,54.133396,53.058197,50.428677,48.99885,49.911827,51.647236,53.197784,54.06549,53.797634,51.130386,47.78407,44.43775,40.710396,38.692043,37.17922,35.783348,34.236572,32.414394,30.056503,28.35505,27.977787,28.822855,30.026323,1.2185578,0.72811663,0.32444575,0.17731337,0.36971724,0.875249,0.97333723,0.91297525,0.70170826,0.52062225,0.69039035,0.7054809,0.7092535,0.9242931,1.3015556,1.5128226,1.9278114,2.5125682,3.4934506,4.6252384,5.198677,4.708236,6.6322746,8.186596,8.043237,6.319147,5.451443,5.160951,4.617693,3.8669407,3.8443048,3.4783602,3.199186,2.867195,2.6446102,3.0256453,1.4600059,0.98465514,0.69793564,0.331991,0.23013012,0.48666862,1.0299267,1.237421,1.0186088,0.814887,0.6111652,0.56589377,0.633801,0.7507524,0.87147635,1.0072908,1.1242423,1.2562841,1.5467763,2.2748928,3.3236825,5.621211,6.930312,6.647365,5.794752,6.1229706,5.6815734,4.727099,3.6745367,3.1048703,2.987919,2.1579416,1.388326,1.1883769,1.8221779,1.8372684,1.9504471,2.8181508,4.183841,4.90064,4.255521,4.425289,3.610402,1.8674494,1.0940613,1.2298758,1.4562333,1.6750455,1.7957695,1.7467253,1.6675003,1.8334957,2.565385,3.5274043,3.712263,3.9801195,5.3684454,7.326438,9.092027,9.691874,9.103344,6.971811,5.221313,4.564876,4.508287,3.5123138,2.8785129,2.867195,3.1312788,2.704972,2.2862108,2.335255,3.218049,4.821415,6.5341864,8.001738,8.684583,8.778898,8.98262,10.484125,8.428044,6.466279,5.7494807,6.1116524,6.039973,5.010046,5.613666,5.5382137,4.3347464,3.4066803,3.6707642,3.0822346,2.1390784,1.3053282,0.98465514,0.8978847,1.2789198,2.4371157,4.266839,6.25124,4.587512,2.7992878,2.0145817,2.1013522,1.6825907,0.8337501,0.8224323,1.0110635,1.0601076,0.935611,1.5618668,2.1579416,2.4107075,2.3088465,2.1466236,2.7011995,3.1765501,3.048281,2.4597516,2.2371666,2.052308,2.2220762,2.71629,3.2218218,3.1652324,3.5538127,3.1312788,3.2935016,4.285702,5.2099953,4.0782075,2.957738,2.0900342,1.6222287,1.6071383,2.5201135,3.2067313,3.361409,3.2369123,3.6669915,4.4516973,4.768598,4.1272516,2.6710186,1.1619685,0.46026024,0.1961765,0.18485862,0.24522063,0.19994913,0.116951376,0.071679875,0.06413463,0.0754525,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.03772625,0.026408374,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.018863125,0.02263575,0.0150905,0.00754525,0.0150905,0.03772625,0.049044125,0.041498873,0.00754525,0.00754525,0.011317875,0.0150905,0.018863125,0.02263575,0.018863125,0.0150905,0.018863125,0.033953626,0.056589376,0.056589376,0.049044125,0.026408374,0.00754525,0.00754525,0.0,0.00754525,0.0150905,0.0150905,0.018863125,0.0150905,0.011317875,0.0150905,0.033953626,0.056589376,0.090543,0.09808825,0.1358145,0.181086,0.15467763,0.071679875,0.02263575,0.00754525,0.0150905,0.041498873,0.056589376,0.049044125,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.033953626,0.13958712,0.41121614,1.0035182,1.50905,1.7052265,1.6335466,1.6260014,1.3543724,0.73188925,0.29426476,0.26408374,0.573439,1.1695137,1.8976303,2.9086938,4.5120597,7.183078,10.785934,13.656902,16.822134,20.055275,21.907633,18.161417,12.875969,7.515069,3.3727267,1.5731846,1.358145,1.3430545,1.4411428,1.5241405,1.3996439,1.8900851,2.776652,3.1312788,2.8596497,2.704972,3.0030096,2.8936033,2.5427492,2.1202152,1.8221779,2.8709676,4.1762958,5.66271,7.2396674,8.7751255,8.684583,8.043237,6.964266,5.824933,5.2628117,5.194905,5.119452,4.666737,3.9122121,3.3953626,2.5578396,1.4939595,0.87147635,0.7092535,0.392353,0.211267,0.124496624,0.10940613,0.124496624,0.09808825,0.056589376,0.094315626,0.1659955,0.24522063,0.30935526,0.3772625,0.5394854,0.814887,1.2034674,1.6825907,2.3201644,3.187868,4.055572,4.745962,5.1345425,5.323174,5.6363015,5.9230213,6.1305156,6.319147,6.677546,7.224577,8.22055,9.831461,12.113899,13.483362,13.309821,12.657157,12.344029,12.96274,14.000212,14.68683,14.966003,15.230087,16.33924,19.232841,21.051247,21.27006,20.421219,20.074137,20.994658,22.100037,23.00924,23.869398,25.344494,26.921452,28.287142,28.954897,28.479546,26.457418,23.182781,21.73032,21.228561,21.202152,21.55678,22.171717,24.401339,28.389004,33.187782,36.76046,36.654823,37.205627,39.60879,43.524776,47.074814,49.485523,52.26972,54.631382,56.33661,57.713615,58.547367,57.740025,55.815987,53.197784,50.206093,48.878128,47.840656,47.22572,47.278538,48.346188,48.681953,49.68547,51.00589,52.424397,53.85045,57.623074,61.59565,65.511635,68.824,70.71031,68.488235,63.614002,58.026745,52.895977,48.632908,44.362297,41.8535,40.597218,40.61608,42.475986,46.65605,51.526512,54.978466,55.785805,53.62032,50.496586,48.930946,48.214146,47.984016,48.244328,49.579838,48.878128,47.557713,45.901527,43.07206,40.634945,38.80522,36.76046,34.330887,32.014496,29.969732,29.079393,28.619133,28.215462,27.841972,0.26408374,0.26408374,0.17354076,0.1358145,0.3169005,0.8903395,1.1317875,1.2713746,1.026154,0.5394854,0.35462674,0.41876137,0.47535074,0.56589377,0.7922512,1.3430545,2.071171,2.8332415,4.183841,5.6023483,5.50426,2.6898816,2.1805773,2.0862615,1.6561824,1.3015556,0.8639311,0.87147635,0.9016574,0.7432071,0.41121614,0.33576363,0.26031113,0.21503963,0.20372175,0.18485862,0.19240387,0.24899325,0.29426476,0.26031113,0.060362,0.06413463,0.9318384,1.4600059,1.3732355,1.3317367,1.0148361,1.0110635,1.1808317,1.4260522,1.7052265,2.0862615,2.4823873,2.927557,3.4142256,3.904667,4.647874,6.066381,7.220804,7.5527954,6.858632,7.032173,6.587003,5.855114,5.168496,4.8402777,4.6327834,3.2557755,1.9994912,1.2902378,0.694163,0.46026024,0.5885295,1.3505998,2.4672968,3.1010978,2.2598023,2.003264,1.7882242,1.4600059,1.2600567,1.7618159,2.2371666,2.142851,1.7354075,2.0673985,2.1768045,2.7992878,4.266839,5.6287565,4.689373,3.4444065,3.6707642,4.7610526,5.9682927,6.432326,6.0739264,5.6513925,5.330719,5.5306683,6.9567204,6.537959,6.2021956,6.628502,7.213259,6.058836,5.828706,5.692891,5.6400743,5.9305663,7.111398,8.616675,10.193633,11.348056,11.491416,9.940866,7.8810134,6.560595,6.741681,7.3792543,5.617439,6.017337,6.417235,6.2399216,5.6853456,5.704209,6.7680893,5.96452,4.3121104,2.7992878,2.3918443,1.9353566,2.1390784,3.531177,5.6061206,6.820906,4.908185,2.6597006,1.3543724,1.3996439,2.3277097,0.9695646,0.65643674,0.94692886,1.4034165,1.6033657,2.4295704,2.6823363,2.5540671,2.3013012,2.2598023,2.6446102,2.3692086,1.7240896,1.1695137,1.327964,1.5165952,2.3993895,3.0935526,3.2784111,3.1916409,3.3727267,3.187868,2.5201135,2.1805773,3.92353,4.738417,4.2027044,3.270866,2.625747,2.7011995,3.5123138,4.002755,3.8103511,3.0671442,2.3880715,2.3314822,2.293756,1.7618159,0.9393836,0.7582976,0.55080324,0.38103512,0.3772625,0.47535074,0.38103512,0.241448,0.094315626,0.011317875,0.003772625,0.02263575,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.08677038,0.094315626,0.06413463,0.033953626,0.026408374,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.041498873,0.056589376,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.02263575,0.018863125,0.0,0.003772625,0.00754525,0.011317875,0.011317875,0.011317875,0.003772625,0.00754525,0.00754525,0.0,0.003772625,0.02263575,0.041498873,0.03772625,0.0150905,0.0,0.0,0.00754525,0.018863125,0.030181,0.041498873,0.030181,0.011317875,0.003772625,0.011317875,0.03772625,0.071679875,0.060362,0.049044125,0.056589376,0.07922512,0.06413463,0.03772625,0.018863125,0.011317875,0.02263575,0.0754525,0.08677038,0.06413463,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.02263575,0.116951376,0.2565385,0.4979865,0.97710985,1.6448646,2.003264,2.033445,1.8334957,1.6410918,1.2034674,0.5017591,0.116951376,0.1358145,0.181086,0.4074435,0.90920264,1.6410918,2.837014,5.0062733,9.578695,16.878725,25.242634,31.369377,30.35454,20.700394,12.294985,6.466279,3.5123138,2.674791,2.4333432,2.11267,1.7769064,1.4713237,1.2110126,1.3732355,2.2183034,2.4786146,1.9127209,1.3241913,1.0374719,0.8224323,0.76584285,1.1204696,2.2748928,4.429062,6.089017,7.598067,8.858124,9.35611,8.07719,6.40969,4.8365054,3.6443558,2.9313297,2.203213,1.720317,1.1959221,0.62625575,0.31312788,0.32821837,0.24899325,0.15845025,0.090543,0.06790725,0.018863125,0.011317875,0.018863125,0.02263575,0.0150905,0.003772625,0.033953626,0.06413463,0.08677038,0.09808825,0.11317875,0.19240387,0.35085413,0.5772116,0.86770374,1.2864652,1.8372684,2.5125682,3.270866,4.0216184,4.4403796,4.7874613,5.160951,5.5382137,5.772116,6.175787,6.7567716,7.6622014,8.952439,10.597303,11.815862,11.668729,11.148107,10.872705,11.117926,11.548005,12.253486,12.970284,13.79649,15.181043,18.327412,20.92675,21.734093,20.73812,19.15739,19.678013,20.877707,21.964222,22.854563,24.197617,25.71044,26.845999,27.189308,26.438557,24.412657,22.137764,21.462463,21.277605,20.979568,20.485353,20.387266,21.481327,24.156118,28.019285,31.89,33.206646,33.780083,35.998386,40.333134,45.324318,47.308716,48.666862,49.892967,51.20961,52.552666,53.19024,52.15654,50.685215,48.972446,46.16561,43.283325,41.438515,40.6274,40.84621,42.04968,42.506165,43.69077,44.743332,45.33941,45.69026,48.829086,51.98677,55.551903,59.788563,64.84765,68.83532,70.12556,68.608955,64.67788,59.21135,53.910812,49.45534,46.3052,44.690517,44.607517,46.086388,49.017715,52.737526,55.86126,56.26493,54.506886,53.148743,51.46238,49.304436,47.104996,47.39926,46.886185,46.139202,45.30168,44.090668,42.781567,41.35174,39.72197,37.552708,34.2328,32.62566,32.33517,32.33517,32.037132,31.309015,0.030181,0.090543,0.150905,0.18863125,0.1961765,0.18485862,0.120724,0.08677038,0.0452715,0.0,0.0,0.02263575,0.1659955,0.392353,0.73188925,1.2826926,1.7957695,2.04099,2.0296721,1.7693611,1.2826926,0.58475685,0.5055317,0.8526133,1.2298758,1.0223814,0.5357128,0.44894236,0.47157812,0.46026024,0.41121614,0.91297525,0.6451189,0.25276586,0.1358145,0.42630664,0.52439487,0.45648763,0.34330887,0.24522063,0.18485862,0.1961765,0.25276586,0.35085413,0.44139713,0.42630664,0.452715,0.694163,0.9997456,1.2902378,1.5731846,1.8146327,2.867195,4.6214657,5.8211603,4.014073,2.6597006,4.112161,7.01331,11.144334,17.455936,23.254461,20.821117,14.698147,9.393836,9.367428,7.745199,5.481624,4.5950575,4.5007415,1.9994912,1.1317875,0.5583485,0.29049212,0.2678564,0.36594462,0.56212115,0.9205205,1.5015048,2.2748928,3.127506,4.508287,6.930312,6.9491754,5.093044,5.873977,4.4215164,5.2854476,6.8246784,7.1566696,4.164978,2.516341,2.0975795,3.048281,4.919503,6.651138,6.858632,6.828451,6.8963585,7.356619,8.469543,11.812089,14.554788,13.50977,8.865668,4.164978,7.413208,11.759273,14.290704,14.607604,14.815099,13.788944,11.548005,9.0957985,6.9265394,5.0213637,3.6028569,3.6254926,4.5912848,5.3382645,4.044254,4.678055,6.145606,7.3415284,7.9753294,8.560086,9.0957985,9.193887,8.182823,6.458734,5.492942,4.236658,3.5651307,4.0103,5.0515447,5.111907,2.7313805,1.3317367,0.58475685,0.241448,0.1056335,0.29049212,0.59230214,1.4109617,2.2409391,1.6788181,1.3015556,1.2336484,1.8146327,2.4672968,1.7089992,0.9507015,0.69793564,0.72811663,0.98465514,1.5731846,2.022127,2.546522,3.0746894,3.410453,3.2670932,2.9954643,2.7011995,1.8636768,1.3015556,3.1425967,4.927048,5.0779533,4.8025517,4.749735,5.0213637,4.3347464,3.3312278,2.5012503,1.9579924,1.4335974,0.7130261,0.4979865,0.7167987,1.2223305,1.7693611,1.086516,0.60362,0.35462674,0.24899325,0.0754525,0.05281675,0.08299775,0.06413463,0.02263575,0.120724,0.10940613,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.090543,0.090543,0.071679875,0.060362,0.06413463,0.0754525,0.041498873,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.08299775,0.20372175,0.29049212,0.15467763,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.02263575,0.02263575,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.03772625,0.060362,0.03772625,0.011317875,0.0,0.00754525,0.030181,0.056589376,0.060362,0.049044125,0.02263575,0.0,0.011317875,0.0150905,0.02263575,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.049044125,0.0,0.060362,0.52439487,0.95824677,1.1732863,1.2223305,2.516341,3.361409,3.2557755,2.263575,1.0072908,0.3734899,0.1961765,0.23767537,0.27917424,0.1056335,0.120724,0.22258487,0.49044126,1.2336484,2.9916916,9.544742,22.537663,34.244118,38.178967,29.098257,17.255987,11.642321,9.390063,8.182823,6.2399216,4.689373,4.055572,3.6481283,3.1048703,2.3956168,2.0296721,1.9730829,1.9240388,1.7655885,1.5580941,1.2525115,1.2110126,1.5731846,2.7653341,5.523123,6.8171334,7.001992,6.428553,5.342037,3.874486,2.4107075,1.3392819,0.5998474,0.18485862,0.1358145,0.10186087,0.1358145,0.16222288,0.13204187,0.0452715,0.056589376,0.071679875,0.08677038,0.1056335,0.090543,0.056589376,0.018863125,0.0,0.003772625,0.0150905,0.003772625,0.018863125,0.03772625,0.049044125,0.060362,0.049044125,0.056589376,0.120724,0.2565385,0.42630664,0.67152727,1.0148361,1.4750963,2.033445,2.655928,3.2784111,3.9197574,4.5422406,5.089271,5.492942,5.8966126,6.48137,7.2283497,8.069645,8.91094,9.533423,9.57115,9.540969,9.725827,10.178542,10.336992,10.944386,11.891314,13.023102,14.143571,16.539188,19.425245,21.439827,21.50019,18.814081,18.742401,19.711966,21.420965,23.013012,23.088465,23.952396,24.005213,22.865881,21.179516,20.628714,19.651604,19.794964,20.836208,21.90386,21.439827,19.73083,19.28566,20.017548,21.952906,25.22377,27.41944,28.709677,30.290405,33.54618,40.038868,46.252384,46.433468,45.86003,47.01068,49.560974,49.534565,48.319782,47.07104,45.935482,44.06803,41.32156,38.85049,36.858547,35.775803,36.239838,37.58289,37.75266,38.820312,40.61231,40.710396,44.384933,48.051926,49.90428,50.17591,51.103977,55.96312,60.939213,65.37582,68.45428,69.19749,65.986984,61.678646,56.717644,52.28481,50.307953,49.30821,48.380142,49.485523,52.27349,54.091896,55.46136,58.38137,59.011402,56.321518,52.1075,50.3155,48.731,46.82582,44.675426,42.95511,43.879402,44.8716,44.762196,42.921154,39.261707,36.209656,34.50443,34.960915,36.52278,36.254925,0.17731337,0.23013012,0.17731337,0.1056335,0.060362,0.049044125,0.026408374,0.018863125,0.00754525,0.0,0.0,0.0150905,0.0452715,0.094315626,0.18863125,0.3772625,0.6752999,1.0751982,1.6825907,2.123988,1.539231,1.2525115,0.87147635,0.573439,0.422534,0.362172,0.3055826,0.41498876,0.5772116,0.66775465,0.5583485,0.6790725,0.482896,0.40367088,0.44139713,0.15845025,0.2867195,0.4678055,0.52062225,0.4640329,0.5017591,0.55080324,0.5772116,0.56212115,0.49421388,0.36594462,0.34330887,0.49421388,0.8601585,1.5165952,2.546522,3.2218218,3.6481283,5.0779533,9.042982,17.354074,13.226823,7.677292,3.9348478,3.0709167,3.9914372,5.1232247,4.8930945,4.146115,3.640583,4.0480266,3.6330378,3.6556737,6.066381,10.834979,15.950659,8.578949,6.9227667,5.0175915,2.3277097,3.7348988,4.183841,4.2706113,4.859141,5.6287565,5.0553174,3.2331395,2.6295197,2.425798,2.5389767,3.6028569,4.9647746,5.0515447,4.112161,2.9916916,3.1161883,4.768598,3.9273026,3.742444,4.9987283,6.126743,7.0963078,7.4094353,7.066127,6.477597,6.466279,8.122461,9.574923,9.616421,8.182823,6.375736,7.6282477,7.3453007,7.4094353,8.805306,11.631002,12.264804,13.053283,14.245432,15.128226,14.015302,12.287439,11.570641,11.370691,11.02361,9.718282,8.929804,9.314611,9.533423,9.133525,8.548768,8.412953,9.152389,9.507015,8.948667,7.7037,6.2021956,5.1835866,4.6290107,4.195159,3.2331395,2.746471,2.6332922,2.3013012,1.9466745,2.535204,2.9351022,1.9844007,1.7165444,2.203213,1.5920477,0.8941121,0.55457586,0.5319401,0.67152727,0.694163,0.62248313,0.8262049,0.97710985,0.9318384,0.7167987,1.2864652,2.4107075,3.3123648,3.6028569,3.289729,2.6597006,2.7200627,2.7351532,2.5238862,2.4823873,3.259548,3.7914882,5.2099953,7.2623034,8.29223,8.016829,7.4396167,7.254758,7.175533,5.938112,1.7995421,0.65643674,0.95447415,1.5731846,1.8184053,1.4298248,1.3770081,1.6637276,1.9240388,1.4298248,1.2902378,1.0412445,0.6828451,0.32444575,0.20749438,0.24522063,0.38103512,0.52062225,0.6111652,0.62248313,0.7205714,0.77338815,0.754525,0.6790725,0.6149379,0.34330887,0.18863125,0.11317875,0.0754525,0.041498873,0.10940613,0.10940613,0.060362,0.0,0.0,0.0,0.0,0.02263575,0.056589376,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18485862,0.1961765,0.24899325,0.3470815,0.27917424,0.08299775,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.018863125,0.030181,0.026408374,0.0150905,0.026408374,0.026408374,0.018863125,0.0150905,0.0150905,0.0,0.0,0.00754525,0.018863125,0.026408374,0.026408374,0.0452715,0.05281675,0.041498873,0.033953626,0.049044125,0.033953626,0.018863125,0.00754525,0.0,0.00754525,0.011317875,0.011317875,0.011317875,0.003772625,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.03772625,0.116951376,0.30181,0.56589377,1.1053791,2.3088465,4.38379,6.881268,7.073672,4.745962,2.1805773,1.4864142,0.84129536,0.41498876,0.23013012,0.15467763,0.392353,1.4600059,3.2520027,5.692891,8.741172,14.554788,21.477554,24.642786,22.447119,16.550507,12.804289,10.970794,11.32542,12.770335,12.830698,10.042727,7.8017883,6.560595,6.1342883,5.6778007,4.617693,3.9310753,3.651901,3.5538127,3.1312788,3.4330888,4.459243,5.462761,6.319147,7.5263867,6.2323766,4.8553686,3.6858547,2.7879698,1.9957186,1.2034674,0.7130261,0.51684964,0.5017591,0.44139713,0.30935526,0.34330887,0.32444575,0.19240387,0.056589376,0.12826926,0.16976812,0.15845025,0.11317875,0.090543,0.056589376,0.041498873,0.026408374,0.011317875,0.0150905,0.011317875,0.02263575,0.03772625,0.0452715,0.049044125,0.06413463,0.124496624,0.17731337,0.211267,0.2565385,0.43385187,0.6149379,0.83752275,1.146878,1.6071383,2.3163917,3.169005,3.99521,4.67051,5.1043615,5.330719,5.6363015,6.1003346,6.722818,7.4584794,8.09228,8.333729,8.337502,8.333729,8.627994,8.884532,10.065364,11.717773,13.230596,13.826671,14.403882,16.51278,18.94235,20.515535,20.096773,19.670467,18.591496,18.474545,19.583696,20.828663,22.04722,22.684793,21.839725,19.647831,17.274849,17.037174,17.48989,18.45568,19.610106,20.474035,19.08571,17.410664,16.690092,17.670975,20.621168,23.41291,23.907125,24.091984,26.223516,32.82561,45.26018,47.761433,45.335636,42.65707,44.10576,46.5391,46.467422,45.426178,44.528294,44.45661,43.430458,41.306473,38.808994,36.439785,34.481792,34.17621,34.576107,35.304226,36.326607,37.98656,40.19732,42.98529,45.614807,47.22572,46.803185,47.19931,49.032806,51.933956,55.53304,59.48298,62.685936,64.60243,65.21359,64.52698,62.58785,61.41079,57.494804,54.28053,53.039333,52.88466,54.963375,56.40452,57.189224,57.498577,57.709846,56.921368,54.778515,52.17163,49.576065,47.05595,44.271755,43.649273,43.947308,44.39248,44.656563,42.981518,39.223984,36.220974,34.783604,33.70463,0.35839936,0.26408374,0.181086,0.1056335,0.049044125,0.0150905,0.011317875,0.0150905,0.026408374,0.033953626,0.026408374,0.011317875,0.00754525,0.08299775,0.271629,0.573439,0.73566186,0.784706,1.026154,1.418507,1.5845025,1.327964,1.0148361,0.8639311,0.80734175,0.52062225,0.56212115,0.513077,0.52062225,0.60362,0.694163,0.573439,0.41498876,0.38858038,0.422534,0.19994913,0.31312788,0.41498876,0.46026024,0.4640329,0.4979865,0.55080324,0.482896,0.392353,0.33576363,0.31312788,0.34330887,0.45648763,0.663982,1.026154,1.6373192,2.2899833,3.1124156,4.719554,7.4094353,11.159425,7.3000293,3.942393,1.780679,0.8299775,0.43385187,0.58098423,1.2110126,1.4750963,1.2600567,1.177059,1.0902886,1.3241913,2.6483827,5.138315,8.152642,5.7117543,7.54525,8.080963,7.6207023,12.340257,9.695646,8.748717,8.533678,8.314865,7.598067,5.832478,3.7952607,2.282438,1.7052265,2.093807,3.5500402,3.904667,3.0331905,1.7391801,1.7655885,2.5276587,2.5880208,2.9200118,3.9197574,5.409944,7.9036493,9.774872,9.797507,8.333729,7.3377557,7.816879,9.001483,9.952185,10.431308,10.917976,12.019584,9.480607,7.3188925,7.1793056,8.314865,9.0807085,10.729345,12.306303,12.909923,11.680047,11.057564,11.604594,11.861133,11.234878,9.986138,9.088254,8.643084,8.088508,7.213259,6.175787,5.3910813,5.2099953,5.3986263,5.73439,6.013564,5.9494295,5.3684454,4.7950063,4.5007415,4.5120597,5.281675,5.3684454,5.028909,4.772371,5.3571277,5.349582,3.8858037,2.425798,1.5882751,1.1506506,0.69793564,0.573439,0.8299775,1.297783,1.5769572,1.4864142,1.3166461,1.0148361,0.63002837,0.31312788,0.90920264,2.282438,3.5689032,4.134797,3.5990841,3.9159849,4.881777,5.3080835,5.0439997,4.957229,5.87775,6.436098,6.8963585,7.1340337,6.6549106,5.4891696,4.659192,4.4705606,4.568649,3.904667,1.4260522,0.6488915,0.7469798,1.1053791,1.3355093,1.478869,2.191895,3.0030096,3.5424948,3.5462675,3.199186,3.1350515,2.9803739,2.8294687,3.2331395,3.308592,2.806833,2.2711203,2.0598533,2.335255,2.6823363,2.8256962,2.776652,2.5616124,2.1843498,1.5882751,1.116697,0.8111144,0.6111652,0.3772625,0.29426476,0.19994913,0.13204187,0.10186087,0.06413463,0.094315626,0.12826926,0.16222288,0.18863125,0.19994913,0.120724,0.090543,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.056589376,0.10186087,0.24522063,0.31312788,0.32444575,0.27540162,0.1358145,0.033953626,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.018863125,0.018863125,0.030181,0.030181,0.02263575,0.011317875,0.003772625,0.0,0.0,0.003772625,0.00754525,0.011317875,0.011317875,0.030181,0.033953626,0.033953626,0.030181,0.03772625,0.030181,0.033953626,0.026408374,0.0150905,0.0,0.0,0.0,0.00754525,0.018863125,0.026408374,0.026408374,0.0150905,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.018863125,0.060362,0.10186087,0.19240387,0.452715,1.0789708,2.2484846,3.9461658,4.5309224,3.6594462,2.2899833,1.8900851,1.2298758,0.9997456,1.4562333,2.4182527,3.1010978,4.8100967,6.590776,7.8923316,8.5563135,10.963248,13.570132,14.305794,12.951422,11.159425,11.042474,10.804798,11.02361,11.747954,12.494934,12.351574,11.7555,10.853842,9.789962,8.695901,7.164215,5.692891,4.636556,4.187614,4.3385186,5.2665844,6.360646,6.8246784,6.5945487,6.3417826,4.6290107,2.987919,1.841041,1.2826926,1.086516,0.8903395,0.9280658,1.0450171,1.0638802,0.784706,0.8978847,1.1959221,1.1883769,0.7582976,0.16976812,0.18485862,0.29049212,0.35839936,0.29803738,0.056589376,0.033953626,0.02263575,0.0150905,0.00754525,0.0150905,0.060362,0.07922512,0.0754525,0.071679875,0.10940613,0.120724,0.124496624,0.14713238,0.17354076,0.18485862,0.24899325,0.32821837,0.43007925,0.60362,0.9318384,1.5958204,2.4559789,3.308592,3.99521,4.3913355,4.538468,4.7006907,4.979865,5.4212623,6.0324273,6.5228686,6.832224,6.9454026,6.94163,6.9869013,7.624475,9.110889,10.921749,12.434572,12.943876,12.932558,13.932304,15.596032,17.365393,18.45568,18.055782,17.048492,16.795727,17.667202,19.081938,19.383747,20.043957,19.579924,17.825653,15.939341,15.056546,15.165953,15.924251,17.184307,18.987621,18.568861,17.086218,15.667711,15.369675,17.199398,20.14959,21.654867,22.303759,23.590223,27.917425,37.08113,40.634945,41.008434,40.650036,42.027042,44.26421,43.769997,42.85325,42.906063,44.38116,43.909584,42.355263,40.174683,37.809246,35.662624,34.95714,34.459156,34.070576,34.172436,35.61358,36.960407,38.75995,40.83112,42.72498,43.724724,44.022762,44.98478,46.339153,48.134922,50.73426,55.027508,58.890675,62.9387,66.95655,69.895424,72.34386,69.386116,64.45152,59.928146,57.151497,56.63842,56.144207,55.9933,56.27625,56.834595,56.634647,55.502857,54.171124,52.877113,51.356743,47.221947,44.218937,43.192783,44.0039,45.520493,45.05269,42.66839,39.929462,37.458393,34.960915,0.3734899,0.21503963,0.14335975,0.09808825,0.049044125,0.0150905,0.018863125,0.02263575,0.030181,0.041498873,0.026408374,0.003772625,0.003772625,0.10940613,0.3772625,0.83752275,0.9016574,0.84129536,0.94315624,1.2562841,1.6033657,1.3166461,1.237421,1.2298758,1.1808317,0.995973,0.9695646,0.9393836,0.814887,0.663982,0.7394345,0.56212115,0.392353,0.36971724,0.44516975,0.35839936,0.36971724,0.35462674,0.362172,0.41498876,0.49044126,0.543258,0.4376245,0.33576363,0.31312788,0.331991,0.44894236,0.65643674,0.9507015,1.2449663,1.3770081,1.5467763,2.2371666,3.2633207,3.9801195,3.2670932,1.1883769,0.7092535,0.79602385,0.8903395,0.9205205,0.83752275,1.3317367,1.3694628,0.84129536,0.5357128,0.58475685,0.46026024,0.331991,0.31312788,0.47157812,1.6071383,4.214022,5.7192993,6.700182,10.914205,8.322411,7.914967,8.827943,10.11818,10.767072,8.873214,6.3531003,4.006528,2.3314822,1.5430037,1.9693103,2.2748928,1.9806281,1.2261031,0.80734175,0.45648763,0.95447415,1.7957695,2.806833,4.142342,6.405917,9.005256,9.971047,9.34102,9.163706,9.325929,10.20495,11.400873,12.823153,14.683057,15.184815,12.034674,9.039209,7.8696957,8.039464,8.7751255,9.876732,10.450171,10.152134,9.175024,10.514306,10.789707,10.303039,9.318384,8.073418,7.092535,6.1342883,5.2326307,4.3724723,3.5123138,2.6483827,1.9127209,1.7731338,2.3163917,3.2520027,3.640583,3.5387223,3.4745877,3.6934,4.1574326,5.2552667,5.572167,5.4703064,5.270357,5.2552667,4.851596,3.7613072,2.3880715,1.2751472,1.1091517,1.1393328,1.4411428,1.7429527,1.8184053,1.5165952,1.4373702,1.3091009,1.1581959,1.146878,1.5731846,1.9542197,2.5238862,3.1614597,3.561358,3.2633207,3.7877154,4.7912335,5.2854476,5.270357,5.7419353,6.7454534,7.073672,6.579458,5.4401255,4.164978,2.71629,1.7542707,1.358145,1.327964,1.20724,0.7054809,0.45648763,0.4074435,0.49421388,0.663982,1.0374719,2.0485353,3.180323,4.22534,5.2779026,5.726845,6.432326,6.72659,6.6662283,7.0284004,7.3905725,6.6850915,5.5382137,4.647874,4.776143,5.2665844,5.4665337,5.353355,4.98741,4.534695,3.8820312,3.2331395,2.6672459,2.173032,1.6675003,1.1846043,0.784706,0.52439487,0.39989826,0.32067314,0.32444575,0.32067314,0.31312788,0.31312788,0.34330887,0.24522063,0.17354076,0.116951376,0.06790725,0.041498873,0.03772625,0.02263575,0.05281675,0.09808825,0.018863125,0.018863125,0.00754525,0.0,0.003772625,0.011317875,0.018863125,0.030181,0.03772625,0.030181,0.00754525,0.0,0.003772625,0.026408374,0.06790725,0.11317875,0.15845025,0.21503963,0.20749438,0.124496624,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.026408374,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.018863125,0.02263575,0.02263575,0.02263575,0.02263575,0.030181,0.060362,0.0754525,0.060362,0.060362,0.071679875,0.041498873,0.033953626,0.056589376,0.071679875,0.0452715,0.02263575,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.0150905,0.0,0.011317875,0.011317875,0.02263575,0.056589376,0.10186087,0.40367088,0.9507015,1.5882751,2.0787163,2.0862615,2.595566,3.1576872,4.0178456,5.028909,5.6551647,5.1798143,6.096562,6.8473144,6.6360474,5.4250345,5.3910813,5.8136153,6.296511,6.934085,8.322411,10.31813,11.393328,11.7555,11.91395,12.657157,13.65313,13.947394,13.411682,12.170488,10.582213,9.793735,8.371455,7.001992,6.2361493,6.511551,7.1566696,7.515069,6.9793563,5.6476197,4.304565,2.927557,1.6712729,0.8941121,0.69039035,0.90920264,1.086516,1.659955,2.425798,3.0218725,2.9086938,2.6106565,2.5389767,2.173032,1.4109617,0.58475685,0.49421388,0.51684964,0.48666862,0.33953625,0.07922512,0.05281675,0.018863125,0.003772625,0.00754525,0.0150905,0.10940613,0.15467763,0.1659955,0.15845025,0.14713238,0.13204187,0.094315626,0.08677038,0.11317875,0.124496624,0.13958712,0.181086,0.24522063,0.35839936,0.5772116,1.1280149,1.9089483,2.7125173,3.350091,3.6707642,3.7801702,3.8820312,4.036709,4.3385186,4.9232755,5.240176,5.4476705,5.583485,5.666483,5.6778007,6.439871,7.805561,9.480607,11.068882,12.095036,12.31762,12.728837,13.521088,14.758509,16.388283,16.433554,15.992157,15.920478,16.373192,16.776863,16.720274,17.629477,17.769064,16.791954,15.724301,14.392565,14.200161,14.600059,15.494171,17.225805,18.16519,17.512526,16.305285,15.448899,15.705438,18.61036,21.918951,23.75622,23.94485,24.012758,27.774065,31.59196,35.15332,38.33364,41.197063,42.5703,41.657326,40.182228,39.548428,40.853756,41.355515,40.631172,39.397522,38.261963,37.688522,37.17922,36.077614,34.817554,34.021534,34.527065,35.15332,36.209656,37.514984,39.00894,40.748123,42.238308,43.604,44.61129,45.290363,45.969437,48.802677,51.6246,55.74808,61.320248,67.30363,72.600395,73.73973,71.66856,67.80539,64.01768,60.618538,58.053154,56.28379,55.035053,53.782543,53.371326,53.024246,52.77525,52.62812,52.541348,49.85524,46.32029,43.996353,43.41914,43.566273,43.649273,42.721207,41.24611,39.371113,36.94909,0.21503963,0.124496624,0.08299775,0.05281675,0.02263575,0.011317875,0.02263575,0.018863125,0.0150905,0.011317875,0.0,0.011317875,0.041498873,0.13958712,0.36594462,0.7922512,0.7205714,0.8601585,1.1996948,1.5354583,1.4637785,1.2826926,1.418507,1.4260522,1.3015556,1.4675511,1.2562841,1.3694628,1.2261031,0.80734175,0.66775465,0.6187105,0.513077,0.5281675,0.6187105,0.5281675,0.38480774,0.362172,0.38103512,0.41876137,0.5357128,0.62248313,0.59230214,0.5583485,0.56589377,0.5772116,0.8563859,1.1581959,1.6071383,2.0145817,1.8863125,1.5165952,1.448688,1.3996439,1.2487389,1.0450171,0.76207024,0.70170826,0.8563859,1.177059,1.5731846,1.0412445,1.0110635,1.0751982,1.0601076,1.0638802,1.2487389,0.965792,0.63002837,0.44894236,0.41498876,0.35085413,0.4678055,0.5998474,0.73566186,1.0299267,1.478869,2.493705,5.2175403,8.926031,11.027383,8.571404,6.5228686,4.640329,2.8785129,1.3656902,0.9393836,0.88279426,0.87147635,0.73188925,0.47157812,0.17731337,0.2678564,0.8978847,1.8033148,2.3126192,2.927557,4.8968673,6.590776,7.6923823,9.1825695,9.759781,10.27663,11.16697,12.596795,14.468017,13.7851715,11.212241,8.918486,8.103599,8.993938,9.910686,10.26154,10.050273,9.510788,9.0957985,11.404645,9.940866,7.884786,6.5455046,5.3910813,4.3007927,3.3463185,2.5993385,2.0636258,1.6825907,1.2110126,0.77716076,0.66020936,0.87902164,1.1959221,0.94315624,1.086516,1.4826416,1.8448136,1.7316349,2.595566,3.531177,4.036709,3.874486,3.0709167,2.3277097,1.931584,1.6486372,1.4562333,1.5015048,1.7995421,2.1843498,2.022127,1.2223305,0.23390275,0.34330887,0.6790725,1.2487389,2.1088974,3.3764994,3.350091,2.848332,2.3993895,2.2447119,2.3314822,2.1503963,2.5087957,3.3312278,4.285702,4.7610526,4.5912848,4.425289,3.8858037,3.029418,2.3465726,1.629774,0.98465514,0.5357128,0.31312788,0.26408374,0.27917424,0.20372175,0.13204187,0.1056335,0.120724,0.36971724,1.0638802,2.1994405,3.8141239,5.987156,8.009283,9.948412,11.057564,11.408418,11.898859,12.838243,12.064855,10.042727,7.914967,7.533932,8.246958,8.390318,7.9828744,7.3113475,6.9227667,6.488915,5.855114,5.111907,4.3385186,3.6066296,2.7125173,1.8976303,1.2864652,0.91674787,0.7582976,0.67152727,0.56212115,0.47157812,0.4074435,0.3772625,0.3169005,0.241448,0.22258487,0.24899325,0.21503963,0.20749438,0.1659955,0.20749438,0.271629,0.10186087,0.090543,0.05281675,0.03772625,0.06413463,0.1358145,0.22258487,0.20749438,0.2678564,0.32821837,0.060362,0.026408374,0.03772625,0.056589376,0.06413463,0.06790725,0.03772625,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.033953626,0.026408374,0.0150905,0.00754525,0.00754525,0.00754525,0.011317875,0.0150905,0.0150905,0.033953626,0.030181,0.02263575,0.0150905,0.0150905,0.026408374,0.07922512,0.10940613,0.11317875,0.150905,0.1659955,0.09808825,0.06413463,0.08299775,0.08677038,0.03772625,0.011317875,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.00754525,0.0,0.00754525,0.02263575,0.056589376,0.08299775,0.13204187,0.20372175,0.2565385,0.32821837,0.32821837,0.69793564,1.4864142,2.3465726,3.9763467,6.221059,8.118689,8.941121,8.186596,6.039973,5.1232247,4.29702,3.1425967,1.961765,1.8825399,2.1202152,2.6898816,3.9310753,6.488915,9.691874,12.00072,13.45318,14.25675,14.796235,14.78869,14.600059,14.124708,13.215506,11.691365,12.3289385,11.846043,10.989656,10.257768,9.903141,8.986393,7.8319697,6.2436943,4.357382,2.637065,1.6335466,0.9393836,0.633801,0.754525,1.2864652,1.8900851,2.987919,4.4516973,5.723072,5.8173876,4.6856003,3.8895764,3.059599,2.1768045,1.599593,1.5052774,1.0714256,0.56212115,0.20749438,0.181086,0.10940613,0.03772625,0.00754525,0.0150905,0.0150905,0.14335975,0.23013012,0.26031113,0.23390275,0.13958712,0.09808825,0.056589376,0.041498873,0.0452715,0.05281675,0.08299775,0.13204187,0.19994913,0.30181,0.4376245,0.8526133,1.5165952,2.214531,2.7615614,3.0143273,3.1124156,3.2105038,3.308592,3.5387223,4.1272516,4.357382,4.425289,4.485651,4.61392,4.8138695,5.3344917,6.2399216,7.567886,9.21275,10.917976,11.706455,12.234623,12.653384,13.264549,14.48688,15.105591,15.041456,14.966003,14.898096,14.2077055,14.656648,15.848798,16.350557,15.82239,15.007503,14.143571,14.1058445,14.215251,14.460471,15.471535,17.557796,17.984104,17.512526,16.686321,15.860115,18.293459,23.00924,25.850027,25.054003,21.266287,21.824636,25.182272,29.769783,34.55347,39.012714,40.00869,39.34848,37.31126,35.2665,35.677715,37.175446,37.03586,36.647278,36.881184,38.08465,38.009197,37.303715,36.137974,35.02505,34.81001,34.81001,35.45136,36.281334,37.099995,37.941288,39.774784,41.596962,43.219193,44.426434,44.947056,46.16561,46.984272,48.844177,52.364037,57.362762,62.62935,67.75635,70.7254,70.98949,69.44271,65.82476,62.233223,58.894447,55.695263,52.18672,50.636173,49.76847,49.35348,49.368572,50.006145,49.960873,48.11983,45.735535,43.3701,40.906574,40.44254,39.703106,38.974987,38.239326,37.13395,0.1056335,0.033953626,0.033953626,0.033953626,0.011317875,0.0,0.011317875,0.0150905,0.00754525,0.0,0.0,0.060362,0.1659955,0.33953625,0.55080324,0.73188925,0.36594462,0.40367088,0.44516975,0.452715,0.73188925,0.84129536,1.0450171,1.4600059,1.8825399,1.7844516,1.2110126,0.9507015,0.76584285,0.59607476,0.5357128,0.7167987,1.0450171,1.0714256,0.79602385,0.68661773,0.4678055,0.55080324,0.60362,0.52062225,0.41121614,0.6073926,0.7922512,0.8978847,0.9922004,1.297783,1.9542197,2.0108092,1.8636768,1.5807298,0.8865669,0.70170826,0.63002837,0.7922512,1.1280149,1.3732355,1.4335974,1.569412,1.4826416,1.0827434,0.47157812,0.25276586,0.21503963,0.3772625,0.6488915,0.8563859,0.8563859,0.6451189,0.6073926,0.8299775,1.0978339,1.026154,1.5920477,1.8297231,1.5052774,1.1129243,0.784706,0.4074435,0.3470815,0.69793564,1.297783,0.79602385,0.80734175,0.77716076,0.513077,0.18485862,0.08677038,0.72811663,1.1506506,0.995973,0.52062225,0.27540162,0.120724,0.041498873,0.06790725,0.27540162,0.995973,1.9429018,2.7804246,3.3727267,3.7990334,4.9232755,6.047518,6.760544,6.9869013,6.9755836,6.5341864,5.553304,4.6554193,4.221567,4.3800178,5.062863,6.1229706,6.6850915,6.398372,5.4476705,4.6290107,3.6028569,2.7351532,2.1051247,1.4939595,1.4713237,1.3920987,1.2449663,1.0450171,0.83752275,0.5470306,0.27917424,0.17731337,0.27917424,0.55080324,1.0487897,1.3958713,1.4977322,1.3770081,1.1431054,2.2560298,3.7763977,4.8402777,4.9119577,3.8141239,2.252257,1.569412,1.4901869,1.659955,1.6486372,1.4298248,0.68661773,0.14335975,0.0150905,0.0150905,0.0150905,0.02263575,0.6488915,1.7014539,2.2296214,1.9089483,2.3163917,2.5917933,2.3805263,1.8297231,1.7580433,2.546522,5.1043615,7.835742,6.651138,2.867195,1.8599042,1.3355093,0.5281675,0.19994913,0.124496624,0.08677038,0.06413463,0.0452715,0.0452715,0.31312788,0.16976812,0.030181,0.02263575,0.0,0.21881226,0.4678055,1.237421,2.8634224,5.523123,8.356364,11.619685,14.475562,17.086218,20.613623,22.284895,19.681786,14.905642,10.63503,10.148361,11.808316,11.634775,10.378491,8.888305,8.13378,7.8508325,7.213259,6.48137,5.7683434,5.036454,4.1197066,3.1124156,2.2258487,1.5882751,1.237421,1.0412445,0.8903395,0.7130261,0.5017591,0.3055826,0.29426476,0.34330887,0.44894236,0.56589377,0.6413463,0.663982,0.6073926,0.5017591,0.3961256,0.33576363,0.27540162,0.1961765,0.18485862,0.29426476,0.55080324,0.9393836,0.754525,0.9808825,1.3317367,0.24522063,0.120724,0.14713238,0.18863125,0.19994913,0.21503963,0.116951376,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.030181,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.0452715,0.041498873,0.030181,0.030181,0.030181,0.030181,0.02263575,0.0150905,0.0150905,0.05281675,0.033953626,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.056589376,0.1056335,0.150905,0.12826926,0.094315626,0.056589376,0.026408374,0.0150905,0.003772625,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.049044125,0.018863125,0.00754525,0.033953626,0.1056335,0.23013012,0.35085413,0.47912338,0.6111652,0.73188925,0.694163,0.56589377,0.7884786,1.7618159,3.8593953,5.764571,7.8432875,8.616675,8.122461,7.9036493,7.575431,5.6778007,3.1576872,1.0336993,0.41121614,1.9240388,3.31991,4.564876,5.7683434,7.17176,8.929804,10.906659,12.702429,13.966258,14.403882,15.39231,16.143063,15.886524,14.7170105,13.59654,14.290704,14.7321005,14.962231,14.7736,13.687083,10.121953,6.5568223,3.9159849,2.3918443,1.4637785,0.84129536,0.59607476,0.663982,1.1053791,2.1051247,3.85185,5.3948536,6.462507,6.719045,5.7683434,4.851596,4.4403796,3.9876647,3.5160866,3.5990841,3.821669,2.3277097,0.83752275,0.181086,0.29049212,0.13204187,0.03772625,0.00754525,0.0150905,0.0150905,0.17354076,0.29426476,0.26031113,0.12826926,0.150905,0.07922512,0.033953626,0.02263575,0.026408374,0.0150905,0.026408374,0.08677038,0.1659955,0.2565385,0.36594462,0.67152727,1.1053791,1.5882751,2.0145817,2.2598023,2.4031622,2.5427492,2.7087448,2.9539654,3.3576362,3.6858547,3.8593953,3.8858037,3.9008942,4.1800685,4.425289,4.851596,5.541986,6.5832305,8.073418,9.193887,10.054046,10.767072,11.299012,11.461235,12.106354,12.5326605,12.593022,12.54775,13.060828,13.634267,13.981348,13.521088,12.393073,11.427281,11.808316,12.525115,12.883514,13.057055,14.068119,16.094019,17.89356,17.746428,16.263786,16.373192,17.20317,21.583187,24.556017,24.133482,21.300241,22.156626,23.933533,26.566826,29.63397,32.39553,33.821583,33.8329,33.21419,33.1991,35.447586,35.55699,34.730785,33.821583,33.44432,33.980034,34.542156,35.19482,35.549446,35.590942,35.673943,35.492855,35.8588,36.37565,36.711414,36.5756,36.711414,37.541393,39.095715,41.344196,44.188755,45.592175,46.24484,46.77678,47.840656,50.11178,52.85825,56.15552,59.539566,63.255604,68.220375,69.95579,68.42033,64.61752,59.709335,55.008644,51.503876,48.47823,46.712643,46.15052,45.867577,45.992073,46.241066,45.667625,43.67568,40.038868,37.57157,36.36056,35.56831,34.68174,33.508453,0.02263575,0.00754525,0.0150905,0.02263575,0.026408374,0.02263575,0.00754525,0.011317875,0.00754525,0.0,0.0,0.011317875,0.033953626,0.28294688,0.724344,1.0751982,0.9016574,0.7922512,0.8111144,0.965792,1.1959221,1.0223814,0.935611,1.0412445,1.237421,1.1996948,1.1129243,1.1280149,1.1431054,1.0676528,0.80356914,0.55457586,0.44139713,0.33953625,0.241448,0.26031113,0.43007925,0.51684964,0.51684964,0.52439487,0.7167987,0.8526133,0.95824677,1.0676528,1.2261031,1.4939595,2.082489,2.4710693,2.493705,2.1390784,1.5807298,1.7391801,1.7882242,1.7618159,1.841041,2.3503454,2.0787163,1.9693103,1.7316349,1.2940104,0.80356914,0.5055317,0.3961256,0.48666862,0.66775465,0.7092535,0.42630664,0.24522063,0.20749438,0.30935526,0.5017591,0.41876137,0.8563859,1.3807807,1.6033657,1.2110126,0.814887,0.49421388,0.33576363,0.32821837,0.36971724,0.19240387,0.241448,0.362172,0.4376245,0.40367088,0.7054809,0.965792,0.9242931,0.6413463,0.5055317,0.28294688,0.120724,0.030181,0.0150905,0.06790725,0.22258487,0.5093044,0.91674787,1.4373702,2.0900342,3.2142766,4.666737,5.4438977,5.353355,5.0213637,4.4743333,3.7688525,3.0256453,2.3805263,1.961765,1.9051756,2.0749438,2.3126192,2.6634734,3.3727267,4.4101987,3.874486,2.2899833,0.65643674,0.45648763,0.72811663,0.94692886,1.0487897,0.98465514,0.7167987,0.3772625,0.22258487,0.3734899,0.7997965,1.3430545,1.6071383,1.9542197,2.795515,3.682082,3.2935016,5.409944,5.775889,6.2399216,6.405917,3.6669915,2.4484336,1.931584,1.8863125,2.1353056,2.5616124,2.8332415,2.6974268,1.8334957,0.63002837,0.16222288,0.29049212,1.6109109,2.5276587,2.6898816,3.0218725,1.8561316,2.625747,4.3611546,5.7381625,5.089271,3.4368613,2.7804246,2.7728794,2.897376,2.4522061,2.263575,1.2298758,0.3961256,0.116951376,0.041498873,0.026408374,0.018863125,0.011317875,0.00754525,0.00754525,0.06413463,0.033953626,0.00754525,0.003772625,0.0,0.211267,0.6752999,1.750498,3.6330378,6.3531003,9.899368,12.826925,15.120681,16.856089,18.199142,18.776354,18.549997,17.037174,14.354838,11.208468,10.427535,9.631512,9.156161,9.114662,9.4013815,8.809079,7.9753294,7.145352,6.405917,5.6815734,4.8138695,3.821669,2.886058,2.142851,1.6637276,1.3619176,1.0978339,0.8526133,0.62248313,0.42630664,0.38480774,0.482896,0.6451189,0.8111144,0.9205205,1.0940613,1.086516,0.9997456,0.8903395,0.7507524,0.573439,0.392353,0.27917424,0.28294688,0.40367088,0.5017591,0.3734899,0.33576363,0.392353,0.23013012,0.24522063,0.3772625,0.4979865,0.5055317,0.32444575,0.10940613,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.00754525,0.00754525,0.003772625,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.07922512,0.08677038,0.03772625,0.018863125,0.00754525,0.00754525,0.003772625,0.003772625,0.003772625,0.018863125,0.026408374,0.018863125,0.003772625,0.003772625,0.003772625,0.011317875,0.049044125,0.1056335,0.1659955,0.090543,0.0452715,0.018863125,0.00754525,0.0150905,0.003772625,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.02263575,0.030181,0.10940613,0.362172,0.91297525,1.4335974,1.5015048,1.1657411,0.7432071,0.8186596,1.0638802,1.2261031,1.4675511,1.8938577,2.5804756,2.8634224,2.8294687,2.7992878,3.1237335,4.195159,4.459243,4.1989317,3.9310753,3.8405323,3.7914882,5.0439997,6.6360474,8.246958,9.601331,10.469034,10.751981,10.352083,9.710737,9.318384,9.7296,10.121953,12.261031,15.505488,18.206688,17.708702,16.999449,16.143063,15.577168,15.23386,14.517061,11.529142,7.9413757,4.859141,2.8219235,1.8070874,1.5845025,2.052308,3.138824,4.640329,6.221059,7.779153,8.084735,7.6622014,6.56814,4.376245,3.451952,3.2482302,2.9011486,2.2748928,1.9768555,2.4522061,1.599593,0.66020936,0.18485862,0.071679875,0.049044125,0.018863125,0.0,0.003772625,0.003772625,0.05281675,0.090543,0.08677038,0.06413463,0.06790725,0.05281675,0.056589376,0.124496624,0.17354076,0.0150905,0.018863125,0.05281675,0.10186087,0.17731337,0.3169005,0.48666862,0.7394345,1.0751982,1.4449154,1.7580433,1.9127209,1.9957186,2.1466236,2.4672968,3.0143273,3.2067313,3.4594972,3.5953116,3.6292653,3.7537618,4.146115,4.425289,4.8025517,5.406172,6.2889657,7.541477,8.677037,9.2995205,9.390063,9.337247,9.688101,10.570895,11.121698,11.295239,11.876224,13.026875,12.249713,11.02361,10.155907,9.767326,10.314357,10.8576145,11.140562,11.404645,12.408164,13.313594,14.1926155,14.34352,14.000212,14.335975,16.686321,19.655376,21.647322,21.647322,19.225298,18.957441,20.802254,23.84299,27.136492,29.709421,29.615107,28.509727,28.434275,30.305496,33.90835,35.08164,33.161373,31.524054,31.456148,32.15031,32.116356,32.26726,32.43703,32.72375,33.50091,35.458904,36.402058,36.33038,35.870117,36.281334,37.518757,37.526302,37.375397,37.809246,39.257935,40.67267,42.170403,43.38896,44.415115,45.78835,47.791615,49.534565,51.31902,53.6505,57.211857,61.444744,63.025475,63.23674,62.655758,61.146706,58.717136,55.257637,52.360264,50.183456,47.429443,45.452587,44.76974,43.55118,41.438515,39.53711,38.635452,36.941544,34.542156,31.893772,29.833918,0.0,0.0,0.00754525,0.0150905,0.011317875,0.011317875,0.003772625,0.00754525,0.00754525,0.0,0.0,0.00754525,0.018863125,0.1358145,0.35839936,0.6111652,0.5772116,0.59230214,0.8903395,1.2940104,1.2223305,0.94692886,0.9808825,1.1053791,1.1581959,1.026154,1.0412445,1.2147852,1.327964,1.2638294,1.026154,0.97333723,0.7432071,0.70170826,0.88279426,1.0148361,0.9318384,0.7809334,0.69039035,0.7394345,0.9507015,0.97710985,1.0336993,1.0676528,1.1317875,1.358145,1.9089483,2.2220762,2.2673476,2.142851,2.093807,2.1768045,2.3314822,2.4710693,2.5389767,2.5125682,1.8787673,1.5015048,1.3091009,1.1695137,0.91297525,0.7205714,0.56589377,0.47912338,0.44516975,0.3772625,0.21503963,0.19994913,0.24899325,0.29426476,0.3055826,0.271629,0.45648763,0.7054809,0.84129536,0.6790725,0.5055317,0.35462674,0.24522063,0.18485862,0.1358145,0.1056335,0.11317875,0.17354076,0.26031113,0.31312788,0.4640329,0.47535074,0.362172,0.22258487,0.211267,0.116951376,0.049044125,0.011317875,0.0,0.00754525,0.018863125,0.09808825,0.271629,0.58098423,1.0676528,2.161714,3.7348988,4.8402777,5.0741806,4.5497856,3.8292143,3.2105038,2.516341,1.81086,1.3958713,0.9808825,0.76584285,0.7469798,0.95824677,1.4901869,2.516341,2.8445592,2.2711203,1.2110126,0.70170826,1.086516,1.3656902,1.7542707,1.9730829,1.2449663,0.7167987,0.72811663,1.2411937,2.0296721,2.686109,3.150142,4.195159,5.66271,6.79827,6.247467,8.103599,7.1378064,5.994701,5.4250345,4.2894745,3.059599,2.082489,1.539231,1.4713237,1.7580433,2.3390274,2.7653341,2.595566,1.9730829,1.6071383,1.4977322,1.8485862,2.4182527,3.2482302,4.6856003,4.0970707,3.5764484,3.742444,4.2781568,3.9386206,3.2029586,2.5767028,1.7240896,0.8299775,0.6149379,0.87147635,0.44139713,0.071679875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.07922512,0.2867195,0.7054809,1.2411937,1.539231,2.372981,4.0216184,6.2851934,8.99771,11.759273,14.641558,17.810562,21.537916,21.09652,19.534653,17.16167,13.947394,9.525878,7.5490227,6.4210076,5.987156,6.0814714,6.541732,6.368191,5.9305663,5.43258,4.9534564,4.4630156,3.9801195,3.380272,2.7426984,2.1541688,1.6675003,1.3468271,1.1091517,0.9016574,0.7092535,0.5583485,0.5319401,0.633801,0.784706,0.94692886,1.1280149,1.3355093,1.3770081,1.297783,1.1431054,0.95447415,0.7696155,0.56589377,0.38103512,0.271629,0.31312788,0.36594462,0.29803738,0.26031113,0.31312788,0.43007925,0.51684964,1.0186088,1.2562841,0.95824677,0.24899325,0.07922512,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.00754525,0.00754525,0.003772625,0.00754525,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.003772625,0.041498873,0.05281675,0.033953626,0.02263575,0.011317875,0.003772625,0.0,0.00754525,0.0452715,0.056589376,0.049044125,0.030181,0.0150905,0.00754525,0.030181,0.056589376,0.090543,0.13204187,0.17731337,0.12826926,0.10940613,0.07922512,0.033953626,0.0150905,0.003772625,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.018863125,0.05281675,0.07922512,0.094315626,0.27540162,0.6790725,1.3505998,2.3126192,2.8785129,2.2786655,1.358145,0.7507524,0.8865669,0.94692886,1.0902886,1.1808317,1.1619685,1.0676528,0.91674787,0.6488915,0.5470306,0.7582976,1.3166461,1.7014539,2.5917933,3.874486,5.2665844,6.296511,8.345046,9.986138,11.332966,12.2270775,12.279895,10.929295,8.744945,6.719045,5.624984,6.0324273,7.0246277,9.050528,12.1252165,15.682802,18.565088,18.395319,17.150352,16.388283,16.501461,16.720274,15.158407,12.981603,10.461489,7.9338303,5.7909794,4.6818275,4.29702,4.8063245,5.9117036,6.828451,7.9753294,7.164215,5.926794,4.772371,3.1765501,2.7992878,2.71629,2.4861598,2.003264,1.478869,1.4977322,1.0186088,0.5017591,0.19240387,0.116951376,0.08299775,0.030181,0.0,0.0,0.00754525,0.049044125,0.12826926,0.15845025,0.124496624,0.08299775,0.090543,0.10940613,0.15467763,0.18863125,0.116951376,0.15845025,0.1659955,0.1659955,0.181086,0.241448,0.35462674,0.5319401,0.8111144,1.146878,1.4411428,1.5769572,1.659955,1.7919968,2.052308,2.5012503,2.8634224,3.2444575,3.4670424,3.5651307,3.7763977,4.055572,4.236658,4.4894238,4.949684,5.6891184,6.911449,8.197914,9.163706,9.623966,9.608876,9.378746,9.590013,9.574923,9.363655,9.703192,10.133271,9.899368,9.691874,9.6201935,9.171251,9.310839,9.680555,10.091772,10.597303,11.491416,12.178034,12.46098,12.604341,12.872196,13.513543,15.214996,16.614641,17.263533,16.94286,15.679029,16.029884,18.255732,21.681276,25.374676,28.158873,27.110083,25.450129,24.963459,26.547962,30.181,31.10152,30.12441,29.833918,30.69785,31.078884,30.78462,30.44131,30.286634,30.735577,32.346485,34.77606,35.12691,34.46293,33.851765,34.342205,36.530327,36.685005,36.35679,36.47374,37.375397,38.974987,40.634945,41.95159,42.906063,43.883175,44.773514,45.2715,46.497604,48.659317,51.08134,55.095417,57.50235,59.54711,61.376835,62.052135,60.916576,58.671864,56.04989,53.29587,50.17214,47.633163,46.24484,44.39248,41.646008,38.756176,38.50341,36.945316,34.383705,31.44483,29.04544,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.0150905,0.026408374,0.033953626,0.060362,0.1659955,0.18485862,0.32821837,0.6451189,0.9695646,0.9205205,0.9695646,1.2298758,1.3996439,1.3241913,0.995973,0.965792,1.1657411,1.3468271,1.3656902,1.20724,1.2562841,1.0638802,1.0110635,1.1996948,1.4147344,1.297783,0.995973,0.91297525,1.086516,1.20724,1.0751982,1.0487897,1.0186088,0.9997456,1.1317875,1.6071383,1.9957186,2.3314822,2.546522,2.4710693,2.3692086,2.5087957,2.7879698,2.938875,2.5616124,1.8825399,1.388326,1.1204696,1.0110635,0.8865669,0.77338815,0.5998474,0.41498876,0.271629,0.18863125,0.271629,0.331991,0.3734899,0.36594462,0.24899325,0.20749438,0.21881226,0.241448,0.26031113,0.27917424,0.331991,0.26031113,0.1659955,0.11317875,0.10186087,0.124496624,0.10186087,0.08299775,0.116951376,0.2263575,0.27540162,0.19240387,0.07922512,0.0150905,0.033953626,0.03772625,0.02263575,0.0150905,0.03772625,0.116951376,0.041498873,0.041498873,0.090543,0.20372175,0.42630664,1.3204187,2.8332415,4.1989317,4.8440504,4.3800178,3.5953116,2.9652832,2.293756,1.6373192,1.297783,0.90543,0.63002837,0.48666862,0.482896,0.6413463,1.0751982,1.9353566,2.5578396,2.595566,2.0183544,2.3314822,2.5578396,2.8709676,2.8747404,1.6033657,1.0789708,1.4147344,2.0636258,2.6408374,2.916239,3.7537618,5.0741806,6.221059,6.609639,5.73439,6.462507,5.4174895,4.006528,3.1312788,3.199186,2.6332922,2.0070364,1.6939086,1.7391801,1.8599042,2.2258487,2.565385,2.806833,3.0331905,3.4896781,3.772625,3.2331395,2.8445592,3.1463692,4.2630663,3.9876647,2.8219235,1.9391292,1.690136,1.6071383,1.6939086,1.4675511,0.8601585,0.16976812,0.056589376,0.026408374,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.08677038,0.34330887,0.91297525,2.0145817,3.1539145,4.2027044,5.3910813,7.2698483,8.171506,10.77839,13.3626375,15.562078,18.384,17.904879,16.097792,13.845533,11.465008,8.718536,6.7567716,5.1232247,4.036709,3.5764484,3.7047176,3.7801702,3.6896272,3.4972234,3.2482302,2.9615107,2.704972,2.425798,2.1164427,1.7731338,1.3996439,1.1619685,0.995973,0.87147635,0.7696155,0.694163,0.7205714,0.80734175,0.9280658,1.0676528,1.2449663,1.3732355,1.3770081,1.2638294,1.0714256,0.87147635,0.724344,0.55080324,0.38480774,0.27917424,0.2867195,0.3470815,0.3470815,0.43385187,0.5772116,0.55080324,0.6375736,1.0374719,1.1544232,0.77716076,0.10940613,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.003772625,0.011317875,0.0150905,0.011317875,0.00754525,0.00754525,0.0150905,0.018863125,0.003772625,0.0,0.003772625,0.00754525,0.00754525,0.0,0.003772625,0.0150905,0.02263575,0.02263575,0.018863125,0.011317875,0.00754525,0.02263575,0.06413463,0.06790725,0.049044125,0.033953626,0.026408374,0.041498873,0.06790725,0.08677038,0.09808825,0.11317875,0.1659955,0.14713238,0.14335975,0.10940613,0.056589376,0.0452715,0.030181,0.0150905,0.0150905,0.03772625,0.056589376,0.030181,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.00754525,0.026408374,0.06790725,0.1056335,0.44894236,1.2487389,2.3918443,3.5953116,4.425289,4.08198,2.8596497,1.720317,1.1506506,1.177059,0.9393836,0.8941121,0.77716076,0.52439487,0.24899325,0.08299775,0.026408374,0.011317875,0.011317875,0.026408374,0.663982,2.071171,3.7877154,5.413717,6.6020937,8.605357,10.223814,11.246195,11.559323,11.121698,10.227587,8.6581745,6.964266,5.7683434,5.753253,6.579458,7.24344,8.518587,10.929295,14.762281,16.022339,16.290195,16.59955,17.240896,17.784155,17.154125,16.950403,16.558052,15.596032,13.913441,10.834979,8.137552,6.5040054,5.9003854,5.5985756,5.8211603,4.8440504,3.8895764,3.3048196,2.5540671,2.2598023,2.1088974,1.961765,1.7014539,1.237421,0.9507015,0.69793564,0.46026024,0.3055826,0.392353,0.43385187,0.211267,0.041498873,0.018863125,0.02263575,0.060362,0.15845025,0.20749438,0.18485862,0.150905,0.150905,0.14713238,0.14335975,0.13958712,0.150905,0.21503963,0.24522063,0.26408374,0.28294688,0.28294688,0.29049212,0.39989826,0.62248313,0.9016574,1.1431054,1.2525115,1.3619176,1.50905,1.7467253,2.1088974,2.6106565,3.0822346,3.440634,3.7009451,3.9688015,4.1574326,4.2706113,4.508287,4.98741,5.7607985,6.900131,8.314865,9.714509,10.733118,10.929295,10.197406,9.778644,9.371201,8.967529,8.854351,8.514814,8.52236,8.835487,9.178797,9.024119,9.110889,9.337247,9.778644,10.465261,11.393328,12.208215,12.204442,12.362892,13.030646,13.902123,14.547242,14.807553,14.520834,13.841762,13.249459,13.788944,15.543215,18.546225,22.31885,25.865116,25.733074,24.12971,22.711203,22.643295,24.60506,25.276588,26.623415,28.445593,30.090458,30.433765,29.984823,29.40384,29.24539,29.916916,31.686277,33.474503,33.074604,32.229534,31.878681,32.16163,34.01399,34.859055,35.349495,35.94557,36.930225,38.552456,40.36709,41.672417,42.374123,42.95511,42.838158,42.91361,43.77377,45.309227,46.69378,49.964645,52.899746,55.80844,58.40778,59.811195,59.97342,59.51316,58.30592,56.24984,53.280785,50.624855,47.855747,44.607517,41.121613,38.254417,37.330124,35.91539,33.93476,31.641006,29.584925,0.003772625,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0150905,0.018863125,0.018863125,0.0150905,0.0150905,0.011317875,0.018863125,0.026408374,0.030181,0.049044125,0.094315626,0.28294688,0.3772625,0.39989826,0.6526641,1.1846043,1.5769572,1.6939086,1.5203679,1.1695137,1.0299267,1.0751982,1.2411937,1.388326,1.2940104,1.1619685,1.0148361,0.87147635,0.83752275,1.0940613,1.327964,1.1204696,1.0902886,1.3317367,1.4298248,1.2713746,1.1242423,1.0035182,0.9318384,0.9393836,1.2336484,1.8146327,2.5502944,3.0558262,2.6898816,2.4823873,2.5540671,2.7238352,2.757789,2.372981,1.9730829,1.5920477,1.2261031,0.9205205,0.80356914,0.65643674,0.47912338,0.32444575,0.21881226,0.18485862,0.4074435,0.47535074,0.5055317,0.5055317,0.3961256,0.31312788,0.22258487,0.181086,0.19240387,0.23767537,0.33953625,0.24522063,0.1358145,0.10940613,0.1659955,0.2565385,0.17354076,0.06790725,0.05281675,0.19994913,0.36594462,0.3169005,0.181086,0.06413463,0.0754525,0.090543,0.056589376,0.03772625,0.08299775,0.23390275,0.06790725,0.011317875,0.003772625,0.02263575,0.08677038,0.5885295,1.8448136,3.2142766,4.0970707,3.9348478,3.3010468,2.7087448,2.11267,1.5543215,1.1619685,0.9280658,0.7054809,0.5319401,0.47535074,0.62248313,0.6828451,1.5769572,2.7540162,3.62172,3.5575855,3.8141239,4.006528,4.0178456,3.5651307,2.2069857,2.1051247,2.9313297,3.399135,3.1765501,2.8747404,4.044254,4.825187,4.678055,3.6368105,2.3013012,1.9202662,1.841041,1.4864142,0.9280658,0.86770374,1.5203679,1.8938577,2.2560298,2.5993385,2.6219745,2.5540671,2.3993895,2.4333432,2.9200118,4.08198,4.9949555,4.485651,3.3123648,2.1805773,1.7316349,1.2562841,0.66020936,0.23767537,0.07922512,0.060362,0.060362,0.0452715,0.026408374,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.11317875,0.41498876,1.7391801,3.904667,5.406172,6.198423,7.6697464,6.952948,8.903395,10.103089,9.529651,8.548768,8.918486,8.89585,8.654402,8.45068,8.66572,7.496206,5.5080323,3.7877154,2.837014,2.5578396,2.565385,2.4861598,2.335255,2.1353056,1.9278114,1.659955,1.4901869,1.3656902,1.237421,1.0412445,0.935611,0.8601585,0.814887,0.79602385,0.7997965,0.87902164,0.95447415,1.0299267,1.1129243,1.20724,1.2261031,1.1393328,0.97333723,0.77338815,0.5885295,0.47535074,0.3470815,0.27540162,0.2678564,0.2678564,0.29426476,0.33576363,0.5093044,0.6752999,0.44139713,0.4678055,0.38858038,0.25276586,0.1056335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.003772625,0.011317875,0.02263575,0.02263575,0.02263575,0.026408374,0.041498873,0.011317875,0.00754525,0.003772625,0.003772625,0.0150905,0.003772625,0.00754525,0.0150905,0.018863125,0.0150905,0.011317875,0.018863125,0.033953626,0.049044125,0.049044125,0.03772625,0.033953626,0.030181,0.033953626,0.071679875,0.07922512,0.07922512,0.0754525,0.08677038,0.1659955,0.13958712,0.11317875,0.07922512,0.060362,0.0754525,0.056589376,0.026408374,0.033953626,0.071679875,0.10940613,0.05281675,0.026408374,0.0150905,0.003772625,0.003772625,0.003772625,0.00754525,0.00754525,0.003772625,0.0,0.02263575,0.026408374,0.06790725,0.22258487,0.58098423,2.0485353,4.06689,6.0022464,7.0963078,6.432326,4.425289,2.8747404,1.9391292,1.5241405,1.3204187,0.94692886,0.754525,0.5394854,0.28294688,0.16976812,0.0452715,0.018863125,0.02263575,0.07922512,0.29049212,1.6033657,3.3274553,4.859141,5.80607,6.013564,6.8171334,8.069645,8.850578,8.812852,8.20546,9.009028,9.533423,9.431562,8.782671,8.096053,7.3151197,6.175787,5.674028,6.349328,8.2507305,10.661438,13.343775,15.47908,16.731592,17.225805,17.093763,18.523588,20.711712,22.654613,23.12242,18.87067,14.068119,10.087999,7.4169807,5.66271,4.4743333,3.7575345,3.4368613,3.2369123,2.674791,1.9655377,1.5845025,1.358145,1.1581959,0.90543,0.7205714,0.5885295,0.4640329,0.41498876,0.6187105,0.77338815,0.41498876,0.124496624,0.0754525,0.060362,0.090543,0.15845025,0.1961765,0.1961765,0.23013012,0.24899325,0.21881226,0.1659955,0.124496624,0.124496624,0.1659955,0.23767537,0.32067314,0.38480774,0.3772625,0.2565385,0.27917424,0.41498876,0.6073926,0.79602385,0.8978847,1.0223814,1.2034674,1.4675511,1.841041,2.3277097,2.8181508,3.3274553,3.7877154,4.074435,4.2819295,4.357382,4.5837393,5.093044,5.885295,6.9491754,8.394091,9.967276,11.257513,11.725319,10.978339,10.47658,10.167224,9.899368,9.446653,9.009028,8.646856,8.503497,8.635539,9.027891,9.484379,9.676784,10.038955,10.729345,11.638548,12.445889,12.577931,12.943876,13.7851715,14.667966,14.852824,14.607604,14.056801,13.373956,12.800517,12.679792,13.29473,15.218769,18.474545,22.53389,24.110846,22.933788,20.821117,19.183798,19.021576,19.923233,23.171463,26.40083,28.479546,29.479292,29.192572,28.837946,29.13221,30.158363,31.376923,32.12013,31.422194,30.822346,30.773302,30.645033,31.184519,32.47098,33.753677,34.817554,36.00593,37.680977,39.74838,41.20838,41.830868,42.177948,41.913864,42.249626,42.645752,43.026787,43.766224,46.467422,49.734516,52.779022,55.114277,56.56674,57.566486,58.260647,58.49078,57.649483,54.665337,52.077316,48.16133,43.634182,39.672924,37.948833,35.911617,34.395023,32.840702,31.195837,29.954643,0.0150905,0.003772625,0.00754525,0.0150905,0.011317875,0.0,0.011317875,0.060362,0.060362,0.0150905,0.0150905,0.003772625,0.03772625,0.06790725,0.071679875,0.060362,0.23013012,0.513077,0.73188925,0.8601585,1.0072908,1.4109617,1.750498,1.7731338,1.6448646,1.9391292,1.5354583,1.1695137,1.0525624,1.146878,1.1581959,0.8903395,0.724344,0.62625575,0.63002837,0.8224323,1.2638294,1.3996439,1.2487389,1.0751982,1.4034165,1.6976813,1.448688,1.0902886,0.8526133,0.7922512,0.7582976,1.0035182,1.5052774,2.1315331,2.655928,2.4823873,2.6710186,2.444661,1.7014539,0.9922004,0.8563859,0.814887,0.8262049,0.8262049,0.7167987,0.47157812,0.30181,0.19994913,0.14713238,0.120724,0.21881226,0.49044126,0.8262049,1.0940613,1.1280149,1.1544232,0.8111144,0.47157812,0.2867195,0.21503963,0.13958712,0.1056335,0.14713238,0.31312788,0.6413463,0.95824677,0.6073926,0.20372175,0.026408374,0.0150905,0.26031113,0.32067314,0.26408374,0.17354076,0.1358145,0.11317875,0.071679875,0.041498873,0.026408374,0.0150905,0.003772625,0.00754525,0.02263575,0.060362,0.18485862,0.20749438,0.95447415,2.04099,2.9954643,3.2520027,3.0181,2.7313805,2.3088465,1.7957695,1.358145,0.965792,0.63002837,0.3734899,0.21881226,0.18485862,0.3772625,1.20724,2.1805773,3.059599,3.8141239,4.4630156,4.7874613,4.9345937,4.927048,4.6856003,5.5495315,6.937857,7.0849895,6.085244,5.8890676,7.194396,6.952948,5.342037,3.059599,1.3128735,1.2147852,1.2638294,0.9393836,0.452715,0.73188925,1.9051756,2.142851,1.8146327,1.2789198,0.9016574,1.1581959,1.1732863,1.0336993,0.8601585,0.8224323,0.7884786,0.5319401,0.2867195,0.1358145,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.120724,0.5017591,1.20724,1.991946,2.2748928,1.9202662,1.8146327,2.1503963,2.9200118,3.92353,4.9345937,5.764571,6.1305156,5.9796104,5.4778514,5.062863,3.9801195,3.0520537,2.5691576,2.2899833,2.5201135,2.1843498,1.7693611,1.4901869,1.2826926,1.1091517,0.995973,0.91674787,0.8563859,0.80734175,0.77338815,0.8526133,0.84129536,0.7507524,0.8224323,0.87147635,0.9507015,0.94315624,0.87902164,0.91674787,0.9507015,0.87147635,0.7054809,0.51684964,0.38103512,0.24899325,0.1659955,0.124496624,0.10940613,0.120724,0.10940613,0.09808825,0.10940613,0.124496624,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.030181,0.033953626,0.0452715,0.033953626,0.02263575,0.00754525,0.0,0.0,0.011317875,0.02263575,0.018863125,0.003772625,0.0150905,0.026408374,0.030181,0.02263575,0.0150905,0.0150905,0.0150905,0.033953626,0.0452715,0.041498873,0.0150905,0.003772625,0.03772625,0.08677038,0.10940613,0.060362,0.049044125,0.056589376,0.060362,0.056589376,0.0452715,0.0452715,0.071679875,0.116951376,0.17731337,0.27540162,0.19994913,0.10940613,0.049044125,0.026408374,0.0150905,0.0150905,0.00754525,0.00754525,0.02263575,0.060362,0.060362,0.05281675,0.033953626,0.0150905,0.0150905,0.0150905,0.033953626,0.041498873,0.02263575,0.0,0.060362,0.0754525,0.26031113,0.9507015,2.6106565,6.6247296,10.457717,12.355347,11.216014,6.590776,3.138824,1.4034165,0.7130261,0.5017591,0.32067314,0.150905,0.16976812,0.1659955,0.071679875,0.0,0.0,0.026408374,0.08299775,0.362172,1.267602,3.682082,6.511551,8.66572,9.431562,8.469543,8.175279,8.137552,8.420499,8.537451,7.462252,7.2283497,7.6848373,8.831716,9.842778,9.046755,5.824933,3.7763977,2.8181508,2.9652832,4.3347464,6.3229194,9.337247,12.385528,14.871688,16.618414,18.006739,19.80251,22.254715,24.955914,26.808273,25.721758,22.235851,18.440592,15.086727,11.59705,8.873214,6.9755836,5.7117543,4.727099,3.4934506,2.8219235,2.1881225,1.539231,0.965792,0.68661773,0.6375736,0.46026024,0.27917424,0.19240387,0.29049212,0.27917424,0.23767537,0.21503963,0.20749438,0.18485862,0.23013012,0.33576363,0.3169005,0.21881226,0.3055826,0.4376245,0.44516975,0.35839936,0.24899325,0.19994913,0.211267,0.22258487,0.24899325,0.2678564,0.24522063,0.16976812,0.1358145,0.16976812,0.28294688,0.44139713,0.56589377,0.6790725,0.8224323,1.0450171,1.388326,1.8146327,2.2786655,2.7917426,3.3312278,3.8292143,4.085753,4.168751,4.2894745,4.6252384,5.311856,6.3342376,7.4811153,8.597813,9.552286,10.223814,10.344538,10.201178,9.861642,9.495697,9.397609,9.740918,9.74469,9.488152,9.186342,9.186342,9.673011,10.035183,10.49167,10.993429,11.200924,11.46878,12.396846,13.185325,13.630494,14.143571,14.7170105,14.441608,14.019074,13.739901,13.456953,13.151371,13.517315,14.792462,16.905132,19.470518,20.081682,19.153618,17.701157,16.641048,16.7995,18.033148,19.787418,22.058538,24.63524,27.098766,27.966469,28.411638,29.437794,30.924208,31.629688,31.837183,31.459919,31.1732,30.977024,30.181,30.181,30.531855,31.05625,31.671186,32.38044,34.843964,36.83591,38.635452,40.23882,41.33665,42.80043,43.294643,43.381416,43.67945,44.875374,46.37688,48.025517,49.715652,51.684963,54.503113,55.152004,55.076553,54.820015,53.93345,50.97948,49.22144,47.12386,43.958626,40.11055,37.09245,35.689034,33.94608,31.554235,29.21898,28.67195,0.003772625,0.0,0.0,0.041498873,0.07922512,0.0,0.003772625,0.011317875,0.018863125,0.0150905,0.0150905,0.011317875,0.018863125,0.033953626,0.06413463,0.120724,0.25276586,0.44516975,0.60362,0.7507524,0.995973,1.5920477,1.8863125,1.8448136,1.7429527,2.1315331,2.493705,2.0070364,1.659955,1.750498,1.9278114,1.5241405,1.3430545,1.2261031,1.1506506,1.237421,1.3543724,1.418507,1.599593,1.9164935,2.2447119,2.4899325,2.4069347,2.0070364,1.4826416,1.20724,1.3656902,1.6637276,2.1051247,2.6898816,3.410453,3.4179983,2.8407867,2.0296721,1.2298758,0.5885295,0.45648763,0.5357128,0.6187105,0.6073926,0.5470306,0.35085413,0.20749438,0.124496624,0.08677038,0.060362,0.090543,0.19240387,0.38858038,0.633801,0.7884786,0.8526133,0.80356914,0.7507524,0.6790725,0.45648763,0.4640329,0.4678055,0.5357128,0.8978847,1.9579924,3.078462,2.7125173,2.0975795,2.0183544,2.848332,1.0487897,0.331991,0.17354076,0.27540162,0.55080324,0.51684964,0.3470815,0.17731337,0.06790725,0.026408374,0.033953626,0.030181,0.03772625,0.05281675,0.03772625,0.041498873,0.35839936,1.1091517,2.022127,2.444661,2.3767538,2.3805263,2.4333432,2.474842,2.4069347,2.0862615,1.3920987,1.20724,1.3015556,0.36594462,0.40367088,1.2940104,3.3274553,5.5759397,5.9003854,5.1232247,4.9157305,5.036454,5.191132,5.0741806,5.824933,6.670001,6.273875,5.1760416,5.7909794,5.2250857,4.0593443,2.7087448,1.629774,1.3505998,2.7540162,3.7650797,4.032936,3.832987,4.063117,3.4481792,2.384299,1.3128735,0.5394854,0.23013012,0.32821837,0.30935526,0.241448,0.18485862,0.17731337,0.15845025,0.1056335,0.056589376,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.10186087,0.241448,0.39989826,0.45648763,0.38480774,0.48666862,0.8903395,1.6939086,2.969056,4.1083884,4.9345937,5.43258,5.6476197,5.674028,5.541986,4.8365054,3.8593953,2.886058,2.1541688,1.9164935,1.6561824,1.4147344,1.2223305,1.0638802,0.88279426,0.754525,0.6828451,0.663982,0.724344,0.5998474,0.5998474,0.62248313,0.6451189,0.72811663,0.754525,0.8186596,0.80734175,0.72811663,0.7092535,0.6187105,0.47535074,0.34330887,0.25276586,0.18485862,0.10940613,0.05281675,0.026408374,0.02263575,0.02263575,0.02263575,0.018863125,0.02263575,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.02263575,0.033953626,0.041498873,0.0452715,0.033953626,0.041498873,0.041498873,0.02263575,0.011317875,0.02263575,0.03772625,0.0452715,0.049044125,0.05281675,0.0452715,0.049044125,0.060362,0.06413463,0.06413463,0.0452715,0.03772625,0.03772625,0.041498873,0.026408374,0.033953626,0.05281675,0.060362,0.060362,0.060362,0.07922512,0.08299775,0.08677038,0.071679875,0.02263575,0.041498873,0.071679875,0.08677038,0.10186087,0.18863125,0.15467763,0.116951376,0.11317875,0.15467763,0.211267,0.19994913,0.15845025,0.090543,0.030181,0.03772625,0.03772625,0.056589376,0.06413463,0.041498873,0.003772625,0.05281675,0.060362,0.056589376,0.06413463,0.09808825,0.17731337,0.5281675,1.3166461,2.7011995,4.817642,7.956466,11.231105,11.332966,8.028146,4.1762958,2.2711203,1.3656902,0.9507015,0.70170826,0.47912338,0.41498876,0.2678564,0.14335975,0.14713238,0.3772625,1.3355093,1.9844007,2.5276587,3.5424948,5.9796104,8.356364,9.027891,8.718536,8.167733,8.152642,8.669493,8.627994,8.782671,9.046755,8.511042,7.809334,8.009283,8.835487,9.774872,10.084227,7.7112455,4.8138695,2.9501927,2.6332922,3.2972744,5.5985756,6.530414,8.29223,11.227332,13.822898,15.614895,18.12369,21.051247,24.122164,27.09122,29.090712,28.588953,26.249926,23.062057,20.323132,17.572887,14.086982,10.899114,8.29223,5.7872066,4.1197066,2.8634224,1.9089483,1.2298758,0.87147635,0.76207024,0.70170826,0.5696664,0.3961256,0.3734899,0.754525,0.7809334,0.6149379,0.4376245,0.4640329,0.8337501,0.72811663,0.46026024,0.3055826,0.48666862,0.91674787,1.3619176,1.1431054,0.452715,0.34330887,0.3470815,0.34330887,0.30935526,0.24899325,0.1961765,0.16222288,0.12826926,0.10940613,0.120724,0.16222288,0.23390275,0.3734899,0.5394854,0.724344,0.9507015,1.2600567,1.6260014,2.0900342,2.625747,3.1350515,3.4481792,3.6330378,3.8178966,4.104616,4.5535583,5.1798143,5.8626595,6.590776,7.3415284,8.099826,8.288457,8.443134,8.461998,8.60913,9.495697,9.827688,10.340765,11.057564,11.785681,12.128989,12.393073,11.751727,10.86516,10.352083,10.785934,11.951676,13.124963,13.717264,13.754991,13.875714,14.577423,14.683057,14.422746,14.053028,13.860624,13.788944,14.366156,15.086727,15.716756,16.29774,16.70141,16.229834,15.645076,15.584714,16.55428,18.13878,19.417702,20.662666,22.039675,23.597769,24.412657,26.883726,29.351023,31.214699,32.950108,33.255688,32.301216,31.139246,30.22627,29.411385,28.962442,29.037895,29.724512,31.003431,32.7577,33.73104,35.345722,36.87364,38.08842,39.284344,40.408585,42.060997,43.279552,43.841675,44.26421,44.916874,46.17693,47.60298,48.776268,49.2818,50.534313,50.247593,49.621338,48.8819,47.304943,45.51672,43.82281,42.09118,40.04264,37.239582,34.428974,32.357803,30.777075,29.471746,28.26828,0.0,0.0,0.0,0.02263575,0.049044125,0.00754525,0.0,0.0,0.003772625,0.00754525,0.0150905,0.03772625,0.041498873,0.041498873,0.0452715,0.071679875,0.1358145,0.21881226,0.27540162,0.38103512,0.7167987,0.814887,0.84884065,0.8639311,1.0487897,1.7429527,1.991946,1.6524098,1.5316857,1.961765,2.7879698,3.0218725,2.305074,1.478869,1.1016065,1.4335974,1.4637785,1.6825907,1.991946,2.4823873,3.4255435,3.8858037,3.5160866,2.746471,1.9655377,1.5052774,1.5882751,1.4524606,1.3543724,1.4222796,1.6788181,1.6335466,1.2751472,0.87147635,0.55080324,0.32444575,0.31312788,0.40367088,0.47157812,0.4640329,0.392353,0.29803738,0.32444575,0.41876137,0.51684964,0.55080324,0.49421388,0.43385187,0.3734899,0.32821837,0.29803738,0.35085413,0.3961256,0.41876137,0.44139713,0.49044126,0.331991,0.3169005,0.35085413,0.49421388,0.9620194,1.5052774,1.4977322,1.4109617,1.5467763,2.0372176,1.0978339,0.7130261,0.41498876,0.16976812,0.362172,0.41498876,0.32821837,0.211267,0.14713238,0.17731337,0.20372175,0.150905,0.090543,0.05281675,0.026408374,0.07922512,0.362172,0.7696155,1.2336484,1.750498,1.8334957,2.0485353,2.305074,2.505023,2.516341,2.2447119,1.7278622,1.4034165,1.2034674,0.5394854,0.68661773,2.0673985,4.2291126,6.0248823,5.6363015,4.949684,4.67051,4.5309224,4.293247,3.7537618,3.5424948,3.6669915,3.4783602,3.0181,2.9841464,2.2560298,2.2560298,1.9240388,1.2562841,1.3128735,2.04099,2.3390274,2.2371666,1.9730829,2.033445,1.5656394,0.98465514,0.47535074,0.14335975,0.02263575,0.049044125,0.03772625,0.018863125,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.124496624,0.15467763,0.030181,0.06413463,0.29049212,0.76584285,1.5580941,2.6936543,3.8292143,4.7421894,5.304311,5.455216,5.2552667,4.8138695,4.104616,3.2142766,2.3503454,1.8334957,1.4826416,1.3770081,1.3958713,1.237421,0.8903395,0.6526641,0.59230214,0.63002837,0.5093044,0.47157812,0.44894236,0.4640329,0.52062225,0.59230214,0.6073926,0.65643674,0.6790725,0.6488915,0.58475685,0.452715,0.29803738,0.181086,0.10940613,0.056589376,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.0150905,0.026408374,0.049044125,0.090543,0.07922512,0.071679875,0.071679875,0.071679875,0.05281675,0.056589376,0.094315626,0.1056335,0.08677038,0.08677038,0.08299775,0.09808825,0.1056335,0.10186087,0.08677038,0.0754525,0.06413463,0.0452715,0.026408374,0.02263575,0.041498873,0.049044125,0.0452715,0.03772625,0.041498873,0.10940613,0.1056335,0.071679875,0.041498873,0.0150905,0.033953626,0.049044125,0.071679875,0.10940613,0.15845025,0.14713238,0.150905,0.16222288,0.21503963,0.35839936,0.3772625,0.47912338,0.45648763,0.271629,0.06790725,0.1056335,0.150905,0.12826926,0.041498873,0.0,0.030181,0.030181,0.07922512,0.20372175,0.36971724,0.42630664,0.87902164,1.6637276,2.7313805,4.032936,6.1041074,7.9451485,6.832224,3.500996,2.1503963,1.7882242,2.1390784,2.3993895,2.0900342,1.0601076,0.5093044,0.26031113,0.124496624,0.16222288,0.663982,2.5125682,4.3196554,5.6023483,6.5040054,7.7678347,8.782671,8.763808,8.560086,8.707218,9.454198,9.955957,9.548513,8.91094,8.544995,8.756263,8.590267,7.967784,7.907422,9.114662,11.98563,10.906659,7.8508325,5.0439997,3.531177,3.1916409,3.8669407,3.85185,4.447925,5.9418845,7.6207023,10.521852,13.909668,17.595524,21.402102,25.148317,27.479801,27.743885,26.61587,24.842735,23.265778,21.202152,18.795218,16.11288,13.536179,11.717773,8.001738,5.451443,3.6858547,2.4220252,1.4637785,1.0714256,0.9280658,0.8337501,0.73188925,0.72811663,0.87902164,0.73188925,0.5696664,0.58098423,0.845068,1.2298758,0.8601585,0.59607476,0.73188925,0.9922004,0.98842776,1.0110635,0.7997965,0.45648763,0.4376245,0.452715,0.44516975,0.4376245,0.4074435,0.31312788,0.24899325,0.181086,0.11317875,0.06413463,0.0452715,0.08299775,0.18485862,0.31312788,0.452715,0.6187105,0.8337501,1.146878,1.569412,2.0749438,2.6031113,2.9464202,3.1765501,3.361409,3.561358,3.832987,4.195159,4.568649,4.961002,5.406172,5.9305663,6.4738245,6.692637,6.779407,7.039718,7.8734684,8.137552,8.903395,10.178542,11.517824,12.038446,11.359374,11.521597,11.838497,11.763044,10.872705,11.329193,12.279895,13.053283,13.4644985,13.819125,14.388792,14.600059,14.407655,13.88326,13.230596,13.313594,13.694629,14.056801,14.2077055,14.102073,14.48688,14.879233,15.203679,15.592259,16.41092,17.471025,17.953922,18.199142,18.742401,20.323132,23.499681,25.966978,27.932516,29.716967,31.712687,32.440804,31.822092,30.607307,29.264252,28.030603,27.543936,27.917425,28.709677,29.777328,31.286379,31.972998,34.244118,35.61735,35.821075,36.775547,37.696068,39.10326,40.5444,41.781822,42.777794,42.864567,43.09847,44.0454,45.577084,46.874866,47.187992,47.221947,46.644737,45.5054,44.245346,43.023014,41.604507,40.148273,38.537365,36.398285,33.251915,31.512737,30.105547,28.754948,27.958923,0.0,0.003772625,0.003772625,0.00754525,0.02263575,0.0452715,0.049044125,0.02263575,0.00754525,0.00754525,0.0150905,0.03772625,0.041498873,0.0452715,0.049044125,0.049044125,0.049044125,0.06790725,0.08299775,0.14335975,0.38103512,0.27917424,0.24899325,0.29049212,0.5281675,1.1808317,1.3619176,1.6146835,1.7165444,1.7919968,2.3390274,2.9539654,2.4182527,1.6448646,1.237421,1.4713237,1.3732355,1.5279131,1.7014539,2.022127,2.9803739,3.4444065,3.240685,2.7653341,2.2484846,1.780679,1.6184561,1.2336484,0.8337501,0.5319401,0.35839936,0.30935526,0.26031113,0.21881226,0.18485862,0.15845025,0.19240387,0.2565385,0.30935526,0.3169005,0.241448,0.18485862,0.2565385,0.38103512,0.49421388,0.543258,0.49044126,0.42630664,0.331991,0.241448,0.23767537,0.331991,0.40367088,0.47157812,0.5998474,0.875249,0.6451189,0.5319401,0.5093044,0.5319401,0.52062225,0.43385187,0.41498876,0.47912338,0.6073926,0.7582976,1.1695137,1.7052265,1.8938577,1.6637276,1.3656902,1.6071383,1.418507,1.2751472,1.2487389,1.0072908,1.3656902,1.5316857,1.3166461,0.7809334,0.24899325,0.24522063,0.4376245,0.6187105,0.84884065,1.4600059,2.0485353,2.1051247,2.3616633,2.8521044,2.9049213,3.0256453,2.848332,2.4069347,1.8938577,1.6260014,1.9202662,3.1463692,4.6742826,5.523123,4.398881,3.9876647,3.7952607,3.5500402,3.0935526,2.372981,1.6825907,1.5015048,1.539231,1.50905,1.1280149,0.7696155,2.3390274,2.9954643,2.1277604,1.3430545,1.3053282,0.91297525,0.4376245,0.10186087,0.071679875,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.124496624,0.15467763,0.030181,0.0,0.06790725,0.28294688,0.724344,1.5845025,2.7389257,3.874486,4.7346444,5.1156793,4.938366,4.6742826,4.191386,3.4557245,2.5389767,1.8863125,1.4562333,1.3053282,1.3053282,1.1506506,0.8299775,0.59607476,0.5357128,0.55457586,0.38858038,0.39989826,0.36971724,0.36594462,0.40367088,0.452715,0.47912338,0.5319401,0.6073926,0.6451189,0.5357128,0.36594462,0.21503963,0.11317875,0.056589376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.003772625,0.00754525,0.00754525,0.00754525,0.003772625,0.003772625,0.00754525,0.00754525,0.00754525,0.00754525,0.011317875,0.0150905,0.011317875,0.003772625,0.003772625,0.0150905,0.03772625,0.090543,0.08299775,0.0754525,0.08299775,0.10186087,0.1056335,0.10186087,0.124496624,0.13958712,0.1358145,0.15467763,0.18863125,0.2263575,0.2565385,0.24522063,0.120724,0.10186087,0.0754525,0.03772625,0.00754525,0.00754525,0.030181,0.05281675,0.06413463,0.060362,0.049044125,0.11317875,0.094315626,0.049044125,0.0150905,0.0150905,0.026408374,0.026408374,0.05281675,0.09808825,0.12826926,0.116951376,0.124496624,0.1358145,0.181086,0.32444575,0.43007925,0.5583485,0.663982,0.60362,0.1659955,0.12826926,0.150905,0.124496624,0.0452715,0.011317875,0.018863125,0.0150905,0.0754525,0.21503963,0.39989826,0.45648763,0.935611,1.6486372,2.444661,3.2218218,4.640329,5.323174,4.0178456,1.7165444,1.6448646,2.0900342,2.6483827,2.969056,2.7125173,1.5656394,0.6488915,0.29803738,0.21881226,0.36594462,0.94692886,3.0709167,5.587258,7.5829763,8.597813,8.616675,8.6581745,8.703445,8.944894,9.4127,9.986138,10.042727,9.612649,8.8618965,8.269594,8.627994,9.099571,8.661947,8.831716,10.559577,14.203933,13.788944,10.521852,7.0812173,4.798779,3.6745367,3.0822346,2.6446102,2.4597516,2.6031113,3.138824,5.492942,8.401636,12.083718,16.788181,22.831926,25.487854,26.32915,25.476536,23.360094,20.69662,18.546225,17.263533,16.475054,16.252468,17.093763,15.011275,12.185578,9.163706,6.5568223,5.028909,3.7877154,2.8106055,2.052308,1.5354583,1.3317367,1.267602,0.97333723,0.77716076,0.7809334,0.8639311,1.1317875,0.9242931,1.0374719,1.478869,1.4449154,0.935611,0.60362,0.46026024,0.44139713,0.44139713,0.46026024,0.4678055,0.5093044,0.56212115,0.5357128,0.392353,0.30181,0.23013012,0.15467763,0.071679875,0.060362,0.124496624,0.21503963,0.29803738,0.362172,0.49421388,0.73188925,1.1016065,1.5920477,2.1466236,2.5087957,2.7426984,2.9237845,3.1161883,3.3576362,3.6443558,3.8820312,4.08198,4.2819295,4.538468,5.142088,5.6287565,6.0739264,6.40969,6.4210076,6.5228686,7.1038527,8.190369,9.431562,10.11818,9.7220545,10.555805,11.6008215,11.947904,10.774617,10.325675,11.046246,11.879996,12.377983,12.683565,13.13628,13.758763,14.068119,13.766309,12.709973,12.577931,12.615658,12.698656,12.740154,12.668475,13.2607765,14.181297,14.871688,15.1395445,15.143317,15.497944,15.69412,15.897841,16.716501,19.206434,23.72981,25.310541,25.736847,26.351786,28.05324,29.524563,30.181,29.80751,28.58518,27.072357,26.691322,27.287397,28.113602,28.913399,29.913143,30.407358,32.259716,33.34246,33.448093,34.2743,35.028824,35.9418,37.23581,38.79013,40.114323,40.12187,40.106777,40.87262,42.38544,43.803947,43.283325,42.99661,42.362804,41.33665,40.41613,39.793648,38.767494,37.55648,36.34547,35.274044,32.659615,31.199608,29.841463,28.468227,27.921198,0.003772625,0.0150905,0.00754525,0.00754525,0.026408374,0.0754525,0.094315626,0.049044125,0.0150905,0.0150905,0.0150905,0.0150905,0.018863125,0.041498873,0.0754525,0.0754525,0.03772625,0.0452715,0.07922512,0.11317875,0.12826926,0.29049212,0.44139713,0.5017591,0.55080324,0.8224323,1.0902886,1.841041,1.9730829,1.4109617,1.1053791,1.5203679,1.6750455,1.6260014,1.4713237,1.3053282,1.0789708,0.98465514,0.9242931,0.9507015,1.2449663,1.4147344,1.7278622,1.9844007,2.022127,1.7165444,1.3770081,1.1242423,0.86770374,0.59607476,0.3470815,0.362172,0.35085413,0.29426476,0.20372175,0.1056335,0.07922512,0.12826926,0.17354076,0.17354076,0.116951376,0.049044125,0.02263575,0.018863125,0.026408374,0.041498873,0.049044125,0.08677038,0.14713238,0.26408374,0.5319401,0.66775465,0.73566186,0.84129536,1.0374719,1.3091009,1.2185578,1.0525624,0.9997456,1.0638802,1.0751982,0.84884065,0.5470306,0.38858038,0.452715,0.69039035,1.690136,2.9766011,3.942393,4.13857,3.2784111,3.5160866,3.2859564,3.059599,2.8332415,2.1315331,2.8936033,3.4594972,3.0520537,1.7919968,0.694163,0.9997456,1.358145,1.5958204,1.780679,2.191895,3.1652324,2.7125173,2.6898816,3.4368613,3.772625,4.398881,4.402653,4.0291634,3.572676,3.3953626,3.6254926,4.044254,4.436607,4.29702,2.8294687,2.4710693,2.3578906,2.233394,1.9542197,1.5128226,1.1544232,1.2110126,1.327964,1.3770081,1.4298248,1.4298248,3.3651814,4.1536603,2.969056,1.2336484,1.1091517,0.69039035,0.2565385,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.06413463,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.14713238,0.5470306,1.0110635,1.8259505,2.8558772,3.8971217,4.6856003,4.776143,4.5799665,4.123479,3.4368613,2.5427492,1.8749946,1.4373702,1.1544232,0.9695646,0.814887,0.694163,0.58475685,0.5093044,0.45648763,0.392353,0.36971724,0.33576363,0.32444575,0.32821837,0.34330887,0.392353,0.47535074,0.5885295,0.66020936,0.55080324,0.35839936,0.211267,0.11317875,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.06413463,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.0150905,0.018863125,0.02263575,0.02263575,0.026408374,0.026408374,0.026408374,0.02263575,0.02263575,0.011317875,0.00754525,0.0150905,0.033953626,0.056589376,0.049044125,0.049044125,0.06413463,0.094315626,0.1358145,0.12826926,0.116951376,0.12826926,0.16976812,0.20372175,0.271629,0.331991,0.392353,0.3961256,0.18863125,0.150905,0.07922512,0.030181,0.0150905,0.011317875,0.02263575,0.06790725,0.09808825,0.10186087,0.08677038,0.08677038,0.060362,0.033953626,0.02263575,0.02263575,0.030181,0.026408374,0.03772625,0.071679875,0.11317875,0.090543,0.06790725,0.06790725,0.10186087,0.15845025,0.32821837,0.3734899,0.60362,0.8337501,0.38103512,0.15845025,0.12826926,0.116951376,0.06790725,0.041498873,0.041498873,0.033953626,0.0452715,0.08677038,0.16222288,0.28294688,0.7582976,1.4071891,2.1692593,3.0897799,4.1008434,4.406426,3.9197574,3.0218725,2.5314314,2.7992878,2.5238862,2.2748928,2.1390784,1.7467253,1.026154,0.73188925,0.95824677,1.5958204,2.3277097,4.146115,6.5756855,8.748717,9.895596,9.344792,9.125979,9.439108,9.699419,9.654147,9.386291,8.944894,8.873214,8.809079,8.729855,8.937348,9.97482,10.718028,12.004493,13.890805,15.679029,14.8339615,11.45369,8.080963,5.8702044,4.5837393,3.8103511,3.048281,2.41448,2.022127,1.961765,2.4182527,3.772625,6.6058664,11.608367,19.583696,23.1526,25.02382,24.031622,20.36463,15.558306,12.849561,11.740409,12.3893,14.667966,18.153872,20.904116,20.085455,17.108854,13.687083,11.815862,9.665465,7.4396167,5.379763,3.731126,2.757789,2.3428001,1.8448136,1.4750963,1.2261031,0.8639311,0.8941121,1.0412445,1.5882751,2.161714,1.7429527,1.0299267,0.7205714,0.5998474,0.51684964,0.39989826,0.44516975,0.48666862,0.5885295,0.73566186,0.8299775,0.56212115,0.45648763,0.4074435,0.33953625,0.18863125,0.116951376,0.15845025,0.23013012,0.2678564,0.23013012,0.28294688,0.39989826,0.66775465,1.1053791,1.6486372,2.0372176,2.2748928,2.4899325,2.757789,3.0746894,3.4142256,3.6594462,3.821669,3.9310753,4.0593443,4.402653,5.27413,6.2135134,6.7077274,6.1531515,6.2851934,6.3229194,6.549277,7.0849895,7.9262853,8.8769865,9.616421,10.212496,10.597303,10.559577,9.703192,10.065364,10.529396,10.646348,10.608622,11.00852,12.2119875,13.3626375,13.72481,12.664702,12.136535,11.808316,11.61214,11.566868,11.808316,12.400619,13.132507,13.619176,13.555041,12.728837,12.581704,13.113645,14.249205,16.263786,19.798737,23.458181,23.990122,22.982832,22.239624,23.805264,26.034885,28.007969,28.611588,27.789156,26.547962,26.449873,27.011995,27.73634,28.415411,29.139755,29.298206,29.716967,30.335678,31.082657,31.844728,32.59171,33.549953,34.760967,36.092705,37.23581,37.53762,37.9262,38.51473,39.144756,39.37866,38.61659,37.579117,36.74537,36.224747,35.753166,35.466446,34.843964,34.229027,33.840446,33.75745,32.26726,30.844982,29.558517,28.5135,27.834427,0.0150905,0.026408374,0.011317875,0.00754525,0.0150905,0.0150905,0.0150905,0.00754525,0.00754525,0.0150905,0.0150905,0.0150905,0.033953626,0.056589376,0.0754525,0.0754525,0.026408374,0.033953626,0.05281675,0.056589376,0.030181,0.26408374,0.5319401,0.76207024,0.91674787,0.9922004,0.8337501,0.6828451,0.7809334,1.1431054,1.5580941,1.5920477,1.2525115,0.97333723,0.87902164,0.7922512,0.7809334,0.7696155,0.7922512,0.84129536,0.8563859,0.7205714,0.79602385,0.814887,0.7054809,0.59607476,0.4979865,0.47157812,0.4979865,0.5319401,0.52062225,0.44516975,0.392353,0.3055826,0.21503963,0.23013012,0.181086,0.23013012,0.2263575,0.13958712,0.090543,0.1056335,0.08677038,0.071679875,0.06790725,0.090543,0.07922512,0.041498873,0.0150905,0.1056335,0.45648763,0.4074435,0.3772625,0.40367088,0.49044126,0.62625575,0.80734175,0.9016574,0.875249,0.7582976,0.6111652,0.513077,0.6149379,1.0148361,1.5807298,1.9844007,2.7389257,3.5990841,4.323428,4.5460134,3.7537618,3.180323,3.8593953,3.8292143,2.8181508,2.2447119,2.6710186,3.3350005,2.8407867,1.4901869,1.2826926,3.3463185,5.1873593,5.975838,5.6325293,4.851596,4.7912335,3.8141239,3.0445085,3.138824,4.2706113,4.7233267,4.478106,4.436607,4.6742826,4.45547,4.1498876,4.1574326,3.2821836,1.6825907,0.83752275,0.80356914,0.7582976,0.7394345,0.73188925,0.67152727,0.8299775,1.2638294,1.7391801,2.1768045,2.6408374,3.0671442,2.6446102,1.8561316,1.0487897,0.42630664,0.34330887,0.17354076,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28294688,0.32067314,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.1659955,0.5357128,1.1280149,1.9542197,2.938875,3.953711,4.4177437,4.08198,3.4859054,2.897376,2.335255,1.7844516,1.3807807,1.1996948,1.1317875,0.9016574,0.77716076,0.694163,0.62625575,0.5394854,0.38103512,0.35839936,0.331991,0.331991,0.34330887,0.3055826,0.36594462,0.4640329,0.543258,0.58475685,0.6111652,0.5357128,0.392353,0.21503963,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.0754525,0.0754525,0.026408374,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.041498873,0.060362,0.060362,0.060362,0.071679875,0.0754525,0.06413463,0.03772625,0.0,0.02263575,0.041498873,0.056589376,0.08299775,0.1056335,0.056589376,0.026408374,0.026408374,0.05281675,0.0754525,0.08677038,0.10186087,0.120724,0.13204187,0.1056335,0.1056335,0.124496624,0.17354076,0.23767537,0.27540162,0.27540162,0.15467763,0.0754525,0.071679875,0.060362,0.060362,0.08677038,0.10186087,0.09808825,0.120724,0.071679875,0.041498873,0.041498873,0.056589376,0.0452715,0.033953626,0.049044125,0.08677038,0.1358145,0.19994913,0.18485862,0.12826926,0.07922512,0.071679875,0.120724,0.1358145,0.27540162,0.5017591,0.724344,0.80734175,0.43007925,0.41876137,0.331991,0.116951376,0.090543,0.090543,0.056589376,0.030181,0.026408374,0.0150905,0.271629,0.663982,0.8903395,1.1355602,2.0749438,1.9542197,2.5540671,3.4330888,3.983892,3.4330888,2.7238352,2.0900342,1.6373192,1.4524606,1.5882751,1.8070874,2.1277604,3.3312278,5.281675,6.94163,8.4544525,10.299266,11.404645,11.200924,9.612649,8.771353,9.1825695,9.725827,9.80128,9.337247,8.692128,8.677037,9.024119,9.695646,10.880251,12.928786,14.302021,15.426264,15.961976,14.800008,12.626976,10.26154,8.073418,6.477597,5.9494295,5.2062225,3.9688015,2.8634224,2.2296214,2.1202152,2.3390274,3.108643,5.168496,8.511042,12.404391,15.946886,18.568861,18.715992,16.448645,13.456953,11.834724,10.585986,9.578695,9.439108,11.551778,16.607096,20.915434,22.748928,21.911406,19.7761,18.002966,15.354584,12.1252165,8.82417,6.1644692,4.3196554,3.1010978,2.4333432,2.1579416,1.9994912,1.5241405,1.2940104,1.5505489,2.0485353,2.0598533,1.5241405,1.2864652,1.0450171,0.7054809,0.41121614,0.59607476,0.7130261,0.9280658,1.1732863,1.1581959,0.7582976,0.56589377,0.49044126,0.44516975,0.33576363,0.2263575,0.18863125,0.2263575,0.3055826,0.36594462,0.32821837,0.28294688,0.33953625,0.56212115,0.97710985,1.4147344,1.7354075,2.0183544,2.3201644,2.686109,3.0520537,3.3350005,3.5538127,3.742444,3.9386206,4.2404304,4.9760923,5.66271,6.2625575,7.201941,8.152642,7.6584287,6.8246784,6.5228686,7.4018903,8.488406,9.042982,9.616421,10.3634,11.046246,10.227587,9.431562,8.9788475,8.948667,9.156161,9.4013815,10.502988,12.091263,13.275867,12.664702,12.2119875,11.532914,10.982111,10.853842,11.3669195,10.819888,10.672756,10.880251,11.031156,10.359629,9.95973,10.846297,12.97783,16.003475,19.28566,20.873934,20.500444,19.579924,19.678013,22.522572,24.891779,26.44233,26.498919,25.58217,25.435038,26.121656,26.70264,27.068584,27.370394,28.030603,28.336185,28.539907,28.709677,28.90208,29.158619,30.403585,32.33517,33.855537,34.87792,36.33038,36.918907,36.688778,36.024796,35.458904,35.689034,34.617607,34.010216,33.282097,32.323853,31.493874,31.226017,30.599762,30.558262,31.022295,30.897799,30.788393,29.49061,28.14001,27.287397,26.872408,0.003772625,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.0,0.003772625,0.003772625,0.02263575,0.030181,0.03772625,0.03772625,0.026408374,0.03772625,0.116951376,0.23390275,0.35462674,0.45648763,0.41498876,0.47912338,0.62248313,0.7997965,0.94315624,1.146878,1.1657411,1.0676528,0.8903395,0.6413463,0.5885295,0.66020936,0.7469798,0.77716076,0.7205714,0.6111652,0.47912338,0.36971724,0.32067314,0.35462674,0.3961256,0.47157812,0.49044126,0.43385187,0.362172,0.27540162,0.22258487,0.20372175,0.211267,0.23767537,0.32067314,0.34330887,0.29426476,0.21881226,0.19240387,0.14335975,0.12826926,0.10940613,0.07922512,0.07922512,0.10186087,0.10940613,0.1056335,0.09808825,0.090543,0.07922512,0.0754525,0.060362,0.05281675,0.1056335,0.094315626,0.08677038,0.09808825,0.124496624,0.150905,0.20749438,0.271629,0.38480774,0.51684964,0.58475685,0.6752999,1.2185578,2.335255,3.31991,2.6672459,1.9579924,1.4675511,1.3317367,1.4750963,1.629774,2.4031622,3.289729,3.5802212,3.31991,3.2935016,4.255521,4.515832,3.3010468,1.4222796,1.2449663,1.7165444,2.3616633,2.6974268,2.6106565,2.372981,2.5880208,2.5427492,2.5502944,2.6483827,2.5993385,3.3463185,3.893349,4.5724216,5.3609,5.885295,4.6214657,3.0558262,1.6637276,0.77338815,0.5470306,0.5772116,0.46026024,0.44139713,0.5998474,0.8299775,1.1544232,1.5505489,1.931584,2.1768045,2.1013522,1.5618668,0.91297525,0.49044126,0.32821837,0.1358145,0.07922512,0.116951376,0.09808825,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.06413463,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.071679875,0.32821837,0.77338815,1.4147344,2.252257,3.2557755,3.9725742,3.9989824,3.561358,2.8898308,2.2107582,1.5958204,1.2789198,1.0978339,0.9695646,0.875249,0.80356914,0.7432071,0.69793564,0.633801,0.5017591,0.44894236,0.35085413,0.29426476,0.29803738,0.32821837,0.4678055,0.62248313,0.66775465,0.59230214,0.48666862,0.3772625,0.20372175,0.071679875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.041498873,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.00754525,0.02263575,0.05281675,0.10186087,0.1056335,0.1056335,0.10940613,0.060362,0.05281675,0.05281675,0.0452715,0.030181,0.011317875,0.0452715,0.07922512,0.08677038,0.07922512,0.094315626,0.14335975,0.1659955,0.14713238,0.10940613,0.124496624,0.116951376,0.094315626,0.07922512,0.0754525,0.071679875,0.071679875,0.060362,0.08677038,0.18863125,0.3734899,0.422534,0.35839936,0.29049212,0.2867195,0.392353,0.5281675,0.41876137,0.25276586,0.12826926,0.08677038,0.0754525,0.06790725,0.049044125,0.026408374,0.033953626,0.011317875,0.030181,0.08299775,0.14335975,0.17354076,0.150905,0.09808825,0.0754525,0.12826926,0.3055826,0.36594462,0.38103512,0.44894236,0.573439,0.6375736,0.4640329,0.452715,0.41121614,0.28294688,0.150905,0.124496624,0.094315626,0.060362,0.033953626,0.041498873,0.120724,0.24899325,0.51684964,1.0336993,1.9655377,3.289729,4.183841,4.274384,3.6745367,3.0181,2.6634734,2.305074,2.0258996,1.871222,1.8787673,3.1916409,4.1612053,5.4476705,7.4018903,10.069136,13.015556,14.57365,14.852824,13.909668,11.736636,11.068882,11.359374,11.740409,12.098808,13.04951,12.294985,11.2801485,10.589758,10.95193,13.200415,14.0983,14.11339,13.404137,12.053536,10.065364,8.5563135,7.175533,6.149379,5.5570765,5.3646727,5.100589,4.4931965,3.7348988,2.9954643,2.425798,2.8898308,3.6179473,4.7648253,6.3153744,8.073418,10.585986,13.174006,14.11339,13.35132,12.51757,13.306048,13.151371,12.47607,11.570641,10.585986,11.763044,14.690601,17.765291,19.934551,20.677757,20.255224,19.11589,17.365393,15.113135,12.449662,9.846551,7.673519,6.017337,4.7836885,3.7084904,3.0671442,2.7728794,2.8407867,3.0407357,2.916239,2.2786655,1.8070874,1.5165952,1.2751472,0.8262049,0.66020936,1.0940613,1.3996439,1.2713746,0.8186596,0.66775465,0.77338815,0.87147635,0.7809334,0.4074435,0.33953625,0.3169005,0.35462674,0.4376245,0.5357128,0.55080324,0.5017591,0.4640329,0.4979865,0.66020936,0.9242931,1.1996948,1.478869,1.7580433,2.0258996,2.2862108,2.4974778,2.6974268,2.9351022,3.2670932,3.7575345,4.5460134,5.3344917,5.885295,6.006019,6.360646,6.398372,6.9227667,7.594294,6.960493,7.911195,8.469543,9.22784,10.227587,10.963248,10.34831,9.49947,8.89585,8.677037,8.631766,8.650629,9.348565,10.582213,11.672502,11.3971,10.982111,10.480352,9.922004,9.450426,9.318384,9.325929,9.748463,10.20495,10.137043,8.809079,8.601585,9.963503,12.46098,15.226315,16.969267,16.62973,15.739391,15.611122,17.278622,21.507734,25.789665,27.310032,26.412148,24.537153,24.205162,25.58217,26.585688,27.302486,27.830654,28.275824,28.502182,28.057013,27.476028,27.155355,27.351532,27.027086,27.928743,29.64906,31.663641,33.34246,34.523293,35.08541,34.72324,33.448093,31.599506,31.044931,30.705395,29.984823,29.007713,28.637997,28.898308,28.724768,28.290915,27.85329,27.762747,27.34776,26.845999,26.51778,26.302742,25.808527,0.0,0.003772625,0.011317875,0.018863125,0.02263575,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.011317875,0.011317875,0.03772625,0.0754525,0.07922512,0.0754525,0.120724,0.18863125,0.24899325,0.29049212,0.35462674,0.62248313,0.9808825,1.3204187,1.5430037,1.5656394,1.3920987,1.20724,1.026154,0.7054809,0.60362,0.5998474,0.59607476,0.60362,0.7394345,0.6488915,0.513077,0.33953625,0.18485862,0.15467763,0.18863125,0.23013012,0.271629,0.29803738,0.29426476,0.24899325,0.2263575,0.1961765,0.1659955,0.20372175,0.25276586,0.27917424,0.271629,0.241448,0.21881226,0.19994913,0.181086,0.16222288,0.13958712,0.120724,0.124496624,0.1056335,0.09808825,0.10186087,0.08299775,0.071679875,0.06413463,0.056589376,0.041498873,0.02263575,0.02263575,0.030181,0.033953626,0.030181,0.02263575,0.02263575,0.06413463,0.1659955,0.31312788,0.44139713,0.59230214,0.87147635,1.3468271,1.7354075,1.4298248,1.2751472,1.7014539,2.1692593,2.5767028,3.2670932,4.8327327,5.6853456,5.666483,5.111907,4.8629136,8.197914,11.981857,9.307066,2.0598533,0.90543,0.88279426,1.2261031,1.4864142,1.5580941,1.6825907,2.1013522,2.3428001,2.4182527,2.3692086,2.2560298,2.5389767,3.451952,4.878004,6.4134626,7.394345,4.9044123,2.6634734,1.2034674,0.58475685,0.39989826,0.3772625,0.40367088,0.46026024,0.58098423,0.87147635,1.1695137,1.4901869,1.6976813,1.7278622,1.5656394,1.0902886,0.56589377,0.39989826,0.5093044,0.30935526,0.29049212,0.21503963,0.120724,0.03772625,0.0,0.0,0.10940613,0.124496624,0.030181,0.0,0.18485862,0.150905,0.14713238,0.17731337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.13958712,0.4074435,0.8526133,1.50905,2.41448,3.3840446,3.9084394,3.832987,3.1840954,2.1466236,1.5543215,1.2298758,1.0902886,1.0638802,1.0902886,1.0374719,0.8941121,0.7696155,0.6488915,0.38858038,0.32821837,0.2867195,0.27917424,0.3055826,0.35462674,0.6451189,0.68661773,0.67152727,0.67152727,0.6413463,0.38103512,0.30935526,0.2565385,0.14713238,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.124496624,0.19994913,0.18485862,0.094315626,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.0150905,0.003772625,0.0,0.00754525,0.026408374,0.071679875,0.124496624,0.120724,0.10186087,0.08677038,0.071679875,0.056589376,0.049044125,0.041498873,0.033953626,0.041498873,0.071679875,0.0754525,0.06413463,0.06790725,0.10186087,0.116951376,0.124496624,0.11317875,0.08299775,0.071679875,0.060362,0.056589376,0.06790725,0.07922512,0.071679875,0.049044125,0.030181,0.041498873,0.090543,0.18485862,0.25276586,0.35462674,0.47535074,0.60362,0.7394345,0.97710985,0.68661773,0.362172,0.1961765,0.08677038,0.056589376,0.041498873,0.030181,0.026408374,0.06790725,0.07922512,0.09808825,0.1358145,0.15845025,0.1056335,0.10940613,0.10186087,0.11317875,0.181086,0.35839936,0.482896,0.5281675,0.5772116,0.66775465,0.77716076,0.67152727,0.58098423,0.47912338,0.35839936,0.21503963,0.23013012,0.18485862,0.10940613,0.049044125,0.08299775,0.14713238,0.18863125,0.45648763,1.4637785,3.953711,6.156924,8.699674,8.6732645,5.9532022,3.2255943,2.335255,2.1768045,2.2975287,2.372981,2.1994405,2.9803739,4.825187,6.9869013,9.242931,11.910177,15.101818,15.860115,15.501716,14.886778,14.418973,14.132254,13.781399,14.169979,15.316857,16.448645,14.377474,11.415963,9.805053,10.589758,13.622949,14.437836,13.675766,12.027128,9.955957,7.707473,6.270103,5.5985756,5.1081343,4.798779,5.247721,4.8742313,4.647874,4.236658,3.610402,3.0520537,3.7009451,4.1762958,4.538468,4.983638,5.8173876,6.8661776,7.7150183,7.9036493,7.6508837,7.8696957,10.816116,12.921241,13.600313,13.075918,12.396846,11.6008215,11.891314,12.909923,14.358611,16.007248,17.180534,17.96524,18.225552,17.867151,16.833452,15.158407,13.192869,11.34051,9.710737,8.118689,6.802043,5.9909286,5.4703064,5.0175915,4.38379,3.6066296,2.969056,2.4408884,1.9391292,1.3317367,1.1808317,1.6637276,1.9994912,1.8297231,1.2185578,1.2185578,1.2525115,1.177059,0.95447415,0.6451189,0.5696664,0.47912338,0.44516975,0.47912338,0.56212115,0.63002837,0.63002837,0.59607476,0.56212115,0.5696664,0.66020936,0.8186596,1.0336993,1.2713746,1.4864142,1.7052265,1.9353566,2.161714,2.4182527,2.7879698,3.361409,4.06689,4.7535076,5.2665844,5.451443,5.7004366,6.058836,6.6586833,7.1981683,6.934085,7.0585814,7.175533,7.748972,8.797762,9.914458,10.035183,9.601331,9.024119,8.586494,8.416726,8.4544525,8.60913,9.129752,9.955957,10.748209,11.189606,10.744436,10.03141,9.454198,9.190115,8.850578,8.782671,8.684583,8.318638,7.488661,7.594294,9.242931,11.431054,13.174006,13.539951,12.702429,12.479843,13.649357,16.550507,21.088974,24.767282,25.170954,23.907125,22.571615,22.741383,23.846762,24.854053,25.79721,26.649822,27.355305,27.849518,27.770292,27.445847,27.14781,27.064812,26.374422,25.933023,26.40083,27.80802,29.56229,30.863846,31.350513,31.097748,30.26777,29.113348,28.1966,28.215462,27.434528,25.944342,25.642532,25.72553,25.72553,25.51049,25.19359,25.091728,25.012505,25.02382,25.07664,24.986095,24.442837,0.0,0.0,0.003772625,0.011317875,0.0150905,0.00754525,0.0150905,0.00754525,0.003772625,0.00754525,0.00754525,0.00754525,0.003772625,0.030181,0.07922512,0.090543,0.08299775,0.090543,0.09808825,0.10186087,0.11317875,0.20749438,0.4678055,0.7809334,1.0638802,1.2638294,1.2525115,1.1355602,1.0940613,1.0978339,0.9016574,0.79602385,0.7997965,0.88279426,1.0487897,1.3166461,1.1431054,0.8903395,0.6187105,0.3734899,0.181086,0.13204187,0.1659955,0.23013012,0.27917424,0.29049212,0.241448,0.25276586,0.271629,0.27540162,0.27917424,0.21881226,0.23767537,0.2678564,0.27540162,0.24522063,0.26031113,0.23767537,0.20749438,0.17731337,0.1659955,0.15845025,0.11317875,0.08299775,0.07922512,0.056589376,0.049044125,0.05281675,0.056589376,0.049044125,0.030181,0.026408374,0.030181,0.026408374,0.018863125,0.0150905,0.003772625,0.0150905,0.06413463,0.14335975,0.24899325,0.392353,0.47157812,0.46026024,0.40367088,0.43385187,0.845068,1.7919968,2.493705,2.8596497,3.5123138,4.6327834,5.240176,5.4174895,5.304311,5.089271,8.043237,11.729091,9.359882,2.493705,1.0223814,0.845068,1.1657411,1.4901869,1.7354075,2.2447119,3.6745367,4.29702,4.187614,3.5538127,2.7502437,2.1579416,2.8445592,4.274384,5.9003854,7.164215,4.7836885,3.2218218,2.0145817,1.1129243,0.845068,0.77338815,0.9205205,1.0714256,1.0827434,0.9016574,1.0336993,1.0676528,1.1053791,1.1317875,0.9997456,0.8262049,0.6451189,0.6187105,0.6790725,0.4979865,0.41121614,0.24522063,0.1358145,0.09808825,0.030181,0.00754525,0.10940613,0.181086,0.14335975,0.0,0.18485862,0.150905,0.14713238,0.17731337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.18863125,0.5055317,1.026154,1.7919968,2.795515,3.6481283,3.92353,3.470815,2.384299,1.7618159,1.358145,1.1732863,1.1581959,1.2185578,1.20724,1.0789708,0.9205205,0.72811663,0.41876137,0.3772625,0.33576363,0.31312788,0.32821837,0.3961256,0.5696664,0.4640329,0.392353,0.46026024,0.58098423,0.271629,0.24899325,0.24522063,0.14713238,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.011317875,0.011317875,0.018863125,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.033953626,0.071679875,0.06790725,0.041498873,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.06790725,0.116951376,0.08677038,0.049044125,0.030181,0.026408374,0.0,0.0,0.0,0.049044125,0.18485862,0.44516975,0.5885295,0.4678055,0.26031113,0.08677038,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.0150905,0.011317875,0.018863125,0.030181,0.0452715,0.06413463,0.11317875,0.13958712,0.13204187,0.10186087,0.06413463,0.056589376,0.041498873,0.026408374,0.02263575,0.049044125,0.060362,0.041498873,0.033953626,0.049044125,0.08677038,0.06790725,0.06413463,0.06413463,0.060362,0.03772625,0.033953626,0.049044125,0.06790725,0.08299775,0.0754525,0.05281675,0.041498873,0.049044125,0.06790725,0.0754525,0.12826926,0.26408374,0.44139713,0.59607476,0.6488915,0.8601585,0.6790725,0.44894236,0.30935526,0.16976812,0.1056335,0.06790725,0.0452715,0.060362,0.14713238,0.15467763,0.14713238,0.14713238,0.14713238,0.090543,0.150905,0.19994913,0.20372175,0.1961765,0.31312788,0.4376245,0.47535074,0.5017591,0.5470306,0.6187105,0.59607476,0.52062225,0.44139713,0.3772625,0.3055826,0.452715,0.44139713,0.27917424,0.0754525,0.06413463,0.116951376,0.15467763,0.7092535,2.1805773,4.8553686,6.6586833,11.076427,12.958967,11.004747,7.7301087,4.274384,3.640583,3.7537618,3.451952,2.505023,2.8143783,5.247721,8.028146,10.321902,12.2270775,14.517061,15.592259,15.856343,15.784663,15.916705,16.4411,16.361876,16.505234,16.878725,16.65614,14.11339,11.317875,10.303039,11.578186,14.136025,13.600313,12.253486,10.487898,8.669493,7.145352,6.3455553,5.904158,5.3646727,4.878004,5.2099953,5.2854476,5.251494,4.961002,4.4101987,3.7613072,4.3422914,4.4931965,4.104616,3.4783602,3.3312278,3.410453,3.229367,3.1124156,3.270866,3.7952607,6.5002327,8.82417,10.284176,11.050018,11.951676,11.638548,11.400873,11.159425,11.208468,12.215759,13.177779,14.618922,16.014793,17.052265,17.652113,17.384256,16.414692,15.331948,14.385019,13.4644985,12.483616,10.997202,9.703192,8.677037,7.352846,6.089017,4.991183,3.9801195,3.078462,2.3880715,2.3314822,2.5012503,2.6408374,2.5880208,2.2673476,2.1579416,1.9051756,1.569412,1.2336484,1.026154,0.8601585,0.66775465,0.5583485,0.5470306,0.55457586,0.5998474,0.62248313,0.6149379,0.5772116,0.52062225,0.51684964,0.58475685,0.72811663,0.9205205,1.1317875,1.3505998,1.599593,1.8599042,2.1466236,2.4861598,3.0331905,3.6028569,4.142342,4.5950575,4.930821,5.198677,5.73439,6.2663302,6.6813188,7.0548086,6.63982,6.4210076,6.6360474,7.322665,8.296002,9.22784,9.533423,9.22784,8.646856,8.439363,8.692128,8.27714,8.054554,8.465771,9.559832,10.465261,10.287949,9.756008,9.318384,9.159933,8.846806,8.511042,7.9300575,7.277394,7.111398,7.99042,9.408927,10.736891,11.400873,10.872705,10.20495,10.861387,12.917468,16.033657,19.48561,21.205925,20.873934,20.232588,20.334448,21.553007,22.326395,22.90738,23.533634,24.307022,25.189817,25.951887,26.310287,26.563053,26.736593,26.600779,26.136745,24.963459,24.265524,24.556017,25.661396,26.695095,27.04972,26.981813,26.729048,26.506464,25.63876,25.58217,24.97855,23.778856,23.220507,22.92247,22.89606,22.95265,22.967741,22.862108,22.95265,23.186554,23.280869,23.099783,22.68102,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.00754525,0.0150905,0.0150905,0.011317875,0.003772625,0.011317875,0.030181,0.041498873,0.049044125,0.05281675,0.05281675,0.056589376,0.1056335,0.07922512,0.071679875,0.090543,0.14713238,0.25276586,0.4376245,0.6187105,0.8111144,0.95824677,0.8865669,0.8563859,1.0450171,1.4298248,1.8825399,2.2069857,1.8146327,1.4449154,1.1544232,0.9016574,0.5281675,0.39989826,0.44516975,0.5093044,0.5093044,0.452715,0.29426476,0.2565385,0.29803738,0.35085413,0.31312788,0.20372175,0.211267,0.25276586,0.2565385,0.20372175,0.23767537,0.20372175,0.15845025,0.1358145,0.150905,0.15467763,0.10940613,0.06413463,0.03772625,0.026408374,0.033953626,0.056589376,0.06413463,0.05281675,0.03772625,0.026408374,0.02263575,0.0150905,0.00754525,0.0150905,0.003772625,0.0,0.00754525,0.026408374,0.071679875,0.17354076,0.32067314,0.422534,0.4376245,0.35462674,0.62625575,1.0789708,1.3920987,1.5731846,1.9429018,1.9994912,2.3088465,2.938875,3.5953116,3.6368105,3.7763977,3.772625,3.2746384,2.3465726,1.4449154,1.2940104,1.8184053,2.2899833,2.4823873,2.674791,5.010046,6.3455553,6.3908267,5.2137675,3.2670932,2.0258996,2.1881225,3.0331905,4.1310244,5.3759904,4.4516973,4.376245,3.6971724,2.4182527,1.9957186,1.7429527,1.8221779,1.9693103,1.841041,1.0072908,0.8978847,0.58475685,0.513077,0.6526641,0.5319401,0.5017591,0.62625575,0.6413463,0.52439487,0.482896,0.30181,0.181086,0.14713238,0.15467763,0.06413463,0.011317875,0.0,0.11317875,0.2263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.120724,0.38858038,0.8299775,1.4524606,2.3201644,3.289729,3.8593953,3.772625,3.0369632,2.2711203,1.750498,1.4562333,1.3355093,1.3015556,1.3505998,1.3543724,1.2449663,1.0450171,0.8526133,0.88279426,0.67152727,0.482896,0.43385187,0.5017591,0.3734899,0.24899325,0.18485862,0.211267,0.32444575,0.17354076,0.12826926,0.124496624,0.10940613,0.07922512,0.041498873,0.05281675,0.090543,0.124496624,0.116951376,0.08677038,0.07922512,0.10186087,0.12826926,0.10186087,0.09808825,0.090543,0.06413463,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.00754525,0.026408374,0.071679875,0.1659955,0.14713238,0.07922512,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.1358145,0.28294688,0.3734899,0.21881226,0.08677038,0.018863125,0.011317875,0.0,0.0,0.0,0.09808825,0.3734899,0.8941121,0.9318384,0.5394854,0.16222288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.041498873,0.0754525,0.090543,0.08299775,0.05281675,0.094315626,0.15467763,0.17731337,0.13958712,0.05281675,0.049044125,0.030181,0.011317875,0.011317875,0.03772625,0.026408374,0.0150905,0.018863125,0.0452715,0.071679875,0.06790725,0.06413463,0.071679875,0.07922512,0.060362,0.071679875,0.090543,0.10186087,0.1056335,0.094315626,0.08677038,0.08299775,0.09808825,0.12826926,0.1358145,0.15845025,0.1961765,0.26408374,0.31312788,0.2565385,0.36971724,0.49044126,0.5583485,0.543258,0.43385187,0.31312788,0.20749438,0.14713238,0.14713238,0.23767537,0.181086,0.150905,0.124496624,0.1056335,0.120724,0.2263575,0.31312788,0.29426476,0.211267,0.26031113,0.3055826,0.26408374,0.2263575,0.21503963,0.18485862,0.2678564,0.29049212,0.31312788,0.35462674,0.392353,0.6111652,0.6488915,0.44139713,0.120724,0.00754525,0.003772625,0.056589376,0.9016574,2.493705,4.032936,4.538468,9.684328,14.25675,15.633758,13.773854,7.2094865,5.455216,5.0213637,4.08198,2.474842,3.108643,5.938112,9.076936,11.348056,12.298758,12.996693,14.894323,16.52787,17.120173,16.588232,17.912424,18.715992,18.421728,16.980585,14.86037,12.996693,12.185578,12.611885,13.864397,14.920732,12.321393,10.502988,8.971302,7.7942433,7.605612,7.745199,7.2057137,6.349328,5.50426,4.991183,5.824933,5.904158,5.6778007,5.2892203,4.557331,4.749735,4.504514,3.4934506,1.991946,0.87147635,0.69039035,0.6752999,0.95447415,1.4147344,1.7391801,2.372981,2.9124665,4.0480266,5.8626595,7.8206515,9.239159,10.555805,11.125471,11.057564,11.219787,10.838752,11.5857315,12.7477,13.932304,15.101818,15.920478,16.131744,16.290195,16.667458,17.278622,17.663431,16.177015,14.618922,13.3626375,11.348056,9.344792,7.6584287,6.1833324,4.9685473,4.195159,4.014073,3.6179473,3.3689542,3.3651814,3.451952,3.1124156,2.5993385,2.1013522,1.720317,1.4675511,1.1695137,0.90543,0.76207024,0.7167987,0.63002837,0.573439,0.5583485,0.55080324,0.52062225,0.44894236,0.43385187,0.47157812,0.5696664,0.73566186,0.9507015,1.1657411,1.3845534,1.6448646,1.931584,2.2183034,2.637065,3.0633714,3.4972234,3.9008942,4.2064767,4.4705606,5.010046,5.6400743,6.2927384,7.009537,6.8397694,6.7152724,6.7077274,6.8359966,7.069899,8.36391,9.35611,9.4127,8.737399,8.360137,8.710991,8.0206,7.4811153,7.5490227,7.9451485,8.7600355,8.948667,8.782671,8.552541,8.529905,8.858124,9.020347,8.635539,7.9791017,7.9715567,9.378746,10.072908,10.401127,10.33322,9.450426,9.027891,10.099318,12.223305,14.664193,16.407146,16.263786,16.075155,16.74291,18.470772,20.768301,21.371922,21.258741,21.11161,21.353058,22.130219,23.077147,23.75622,24.582424,25.385994,25.412401,24.963459,23.72981,22.571615,21.956678,21.952906,22.56407,22.93756,23.126192,23.19787,23.243143,23.035648,22.696112,22.488617,22.266033,21.477554,20.89657,20.700394,20.787165,20.92675,20.772074,20.745665,21.017294,21.081429,20.858843,20.692848,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.02263575,0.03772625,0.0452715,0.0452715,0.056589376,0.05281675,0.10186087,0.21503963,0.35085413,0.44894236,0.5093044,0.6073926,0.7432071,0.83752275,0.97333723,1.1544232,1.5015048,1.9881734,2.425798,1.8297231,1.8259505,1.9240388,1.8334957,1.478869,1.3317367,1.3166461,1.3317367,1.2940104,1.0978339,0.66020936,0.3734899,0.21503963,0.15467763,0.1659955,0.19240387,0.16976812,0.120724,0.071679875,0.0452715,0.056589376,0.041498873,0.03772625,0.041498873,0.030181,0.041498873,0.03772625,0.02263575,0.0150905,0.0150905,0.041498873,0.056589376,0.049044125,0.03772625,0.060362,0.060362,0.05281675,0.041498873,0.026408374,0.0150905,0.003772625,0.0,0.00754525,0.011317875,0.0,0.011317875,0.1056335,0.31312788,0.5017591,0.36594462,0.41498876,0.72811663,1.3694628,2.1994405,2.8822856,3.1539145,3.429316,3.1124156,2.282438,1.7089992,1.8184053,2.1579416,2.1956677,1.7731338,1.1129243,1.6373192,3.0331905,3.874486,3.2482302,0.7469798,1.1883769,3.2670932,4.5535583,4.146115,2.6710186,1.9240388,2.022127,2.7426984,3.6783094,4.22534,4.496969,5.194905,5.3156285,4.6214657,3.6330378,2.655928,2.3918443,2.2598023,1.9089483,1.2525115,0.8978847,0.67152727,0.56589377,0.5319401,0.45648763,0.4074435,0.422534,0.41121614,0.3470815,0.27540162,0.24899325,0.18863125,0.12826926,0.0754525,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.27540162,0.633801,1.1581959,2.0372176,3.1652324,4.074435,4.4403796,4.074435,3.0746894,2.4672968,2.173032,2.022127,1.7542707,1.7919968,1.8749946,1.8749946,1.8070874,1.8297231,2.0258996,1.4524606,0.94692886,0.79602385,0.7469798,0.62625575,0.79602385,0.9242931,0.8111144,0.3961256,0.63002837,0.6488915,0.6149379,0.55457586,0.3961256,0.19994913,0.271629,0.46026024,0.6149379,0.58098423,0.43385187,0.38858038,0.38103512,0.38103512,0.38103512,0.36971724,0.26408374,0.14335975,0.05281675,0.0150905,0.003772625,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.00754525,0.033953626,0.1056335,0.20372175,0.14713238,0.056589376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.17354076,0.45648763,0.7394345,0.70170826,0.2263575,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.1056335,0.17731337,0.18485862,0.124496624,0.0754525,0.08677038,0.090543,0.08677038,0.0754525,0.0754525,0.06413463,0.033953626,0.02263575,0.03772625,0.060362,0.060362,0.05281675,0.05281675,0.071679875,0.120724,0.14713238,0.14335975,0.13204187,0.120724,0.120724,0.120724,0.1659955,0.211267,0.21503963,0.1659955,0.13204187,0.1056335,0.116951376,0.15845025,0.18485862,0.20749438,0.2678564,0.3055826,0.3055826,0.3055826,0.4376245,0.52062225,0.76207024,1.0676528,1.0072908,0.7394345,0.4979865,0.35085413,0.29803738,0.27540162,0.13958712,0.16222288,0.150905,0.071679875,0.060362,0.1358145,0.21503963,0.28294688,0.331991,0.38103512,0.32067314,0.21503963,0.14713238,0.1358145,0.1358145,0.19994913,0.18485862,0.20372175,0.27917424,0.36594462,0.29426476,0.26408374,0.26031113,0.21503963,0.030181,0.018863125,0.033953626,0.31312788,1.2525115,3.3878171,3.180323,6.3153744,10.484125,13.272095,12.162943,6.058836,3.1954134,2.071171,1.6825907,1.50905,3.059599,6.8171334,11.053791,14.215251,14.924504,14.215251,14.603831,16.222288,18.248188,18.919714,19.923233,20.19109,19.798737,18.617905,16.31283,14.86037,14.1926155,14.132254,14.347293,14.358611,12.453435,10.495442,8.669493,7.5565677,8.118689,7.8508325,7.360391,6.507778,5.406172,4.45547,4.7120085,4.9685473,5.3344917,5.692891,5.692891,5.251494,4.353609,3.1539145,1.9579924,1.2525115,1.0186088,0.94315624,0.80734175,0.56589377,0.33576363,0.32444575,0.36594462,0.60362,1.1695137,2.1805773,3.5990841,5.142088,7.039718,9.035437,10.38981,10.963248,11.155652,11.140562,11.11038,11.231105,12.449662,13.196642,13.856852,14.800008,16.388283,17.731337,18.278368,18.131235,17.063583,14.509516,12.0082655,10.321902,8.98262,7.7716074,6.700182,5.832478,4.9647746,4.3800178,4.085753,3.8292143,3.5990841,3.1539145,2.7238352,2.335255,1.8448136,1.478869,1.2411937,1.1129243,1.0336993,0.9016574,0.754525,0.6451189,0.5772116,0.52062225,0.41121614,0.38858038,0.4376245,0.5470306,0.694163,0.8563859,0.98842776,1.1317875,1.297783,1.4864142,1.6939086,1.9391292,2.1994405,2.584248,3.0445085,3.3878171,3.731126,3.953711,4.3800178,5.191132,6.4247804,7.326438,7.835742,8.118689,8.156415,7.7678347,8.375228,9.371201,9.510788,8.616675,7.5527954,7.3075747,7.201941,7.3377557,7.5301595,7.3075747,8.322411,8.409182,8.058327,7.699928,7.7376537,8.552541,9.737145,10.574668,10.668983,9.948412,9.850324,9.74469,9.608876,9.26934,8.379,7.816879,8.43559,9.948412,11.778135,13.060828,12.89106,13.241914,14.894323,17.618158,20.157135,20.243906,19.53088,18.731083,18.406637,18.983849,20.202406,21.617142,23.088465,24.167437,24.091984,22.496162,21.051247,19.798737,18.85558,18.402864,18.817854,18.968758,19.191343,19.579924,19.957186,20.153362,20.29295,20.349539,20.258997,19.927006,19.255478,18.776354,18.62545,18.614132,18.233097,18.391546,18.72731,18.919714,18.923487,18.934805,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.011317875,0.011317875,0.00754525,0.00754525,0.026408374,0.03772625,0.049044125,0.060362,0.06413463,0.0452715,0.049044125,0.05281675,0.06413463,0.090543,0.1659955,0.44139713,0.95824677,1.4750963,1.7580433,1.5845025,1.5920477,1.8485862,2.2258487,2.5201135,2.463524,2.0975795,2.425798,2.5578396,2.0862615,1.0789708,0.9695646,1.2751472,1.388326,1.1959221,1.0978339,1.0186088,0.965792,0.7394345,0.38858038,0.21503963,0.19240387,0.23013012,0.29426476,0.33953625,0.32821837,0.22258487,0.19240387,0.18863125,0.16976812,0.07922512,0.071679875,0.08299775,0.0754525,0.049044125,0.041498873,0.026408374,0.02263575,0.030181,0.05281675,0.08677038,0.06413463,0.08677038,0.08677038,0.05281675,0.041498873,0.018863125,0.011317875,0.00754525,0.003772625,0.0,0.011317875,0.08299775,0.362172,0.60362,0.1961765,0.41121614,0.663982,1.3619176,2.4974778,3.640583,4.436607,6.1342883,8.235641,9.65792,8.75249,8.695901,7.8810134,6.1531515,4.4630156,4.847823,5.8702044,6.33801,6.296511,5.7872066,4.8365054,3.0897799,2.8030603,2.8407867,2.5540671,1.7919968,1.5543215,1.7354075,2.3578906,3.338773,4.4818783,5.270357,5.8400235,6.247467,6.1833324,4.9987283,4.647874,3.953711,3.097325,2.2371666,1.5203679,1.2336484,0.784706,0.59607476,0.724344,0.83752275,0.8563859,0.86770374,0.77716076,0.58098423,0.3734899,0.29049212,0.18485862,0.09808825,0.0452715,0.0150905,0.003772625,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.030181,0.018863125,0.018863125,0.02263575,0.011317875,0.003772625,0.0,0.0,0.003772625,0.011317875,0.02263575,0.0754525,0.23013012,0.52062225,0.97710985,1.7467253,2.7653341,3.8556228,4.659192,4.636556,3.9159849,3.308592,2.9766011,2.8596497,2.6597006,3.2331395,4.5761943,5.798525,6.417235,6.3832817,5.6325293,3.9499383,2.4484336,1.5845025,1.1732863,1.3543724,1.6033657,1.6863633,1.5316857,1.2147852,1.3958713,1.4147344,1.4562333,1.4411428,1.0186088,0.814887,0.9242931,1.177059,1.3543724,1.2034674,0.9393836,0.8111144,0.724344,0.633801,0.56589377,0.58098423,0.4979865,0.35839936,0.19994913,0.06413463,0.041498873,0.05281675,0.03772625,0.0,0.003772625,0.0,0.0,0.0,0.00754525,0.02263575,0.041498873,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.071679875,0.094315626,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.090543,0.14713238,0.13958712,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.011317875,0.026408374,0.05281675,0.056589376,0.07922512,0.06790725,0.0452715,0.026408374,0.026408374,0.030181,0.03772625,0.0452715,0.049044125,0.041498873,0.03772625,0.030181,0.033953626,0.05281675,0.08677038,0.08677038,0.11317875,0.150905,0.20372175,0.29426476,0.3961256,0.362172,0.27917424,0.22258487,0.23013012,0.271629,0.28294688,0.27540162,0.2565385,0.23013012,0.13204187,0.09808825,0.120724,0.18485862,0.2565385,0.27917424,0.25276586,0.27917424,0.41876137,0.6828451,0.7394345,0.6752999,0.694163,0.8903395,1.237421,1.0186088,0.7922512,0.6187105,0.482896,0.26408374,0.14713238,0.12826926,0.14335975,0.14713238,0.14713238,0.24899325,0.26408374,0.23013012,0.1961765,0.23390275,0.35085413,0.271629,0.18485862,0.17731337,0.23390275,0.20749438,0.2263575,0.362172,0.55080324,0.58475685,0.40367088,0.31312788,0.29426476,0.27917424,0.1659955,0.124496624,0.15467763,0.40367088,1.0525624,2.2899833,2.5616124,2.9049213,4.768598,7.3075747,7.3868,4.466788,2.8709676,1.8749946,1.177059,0.8865669,3.0256453,7.665974,12.826925,16.520325,16.776863,14.392565,14.690601,16.720274,19.032892,19.715738,18.1086,16.516552,14.879233,13.2607765,11.830952,11.423509,10.785934,10.812344,11.389555,11.393328,10.212496,8.695901,7.6282477,7.3490734,7.7640624,8.160188,7.383027,6.1531515,4.8629136,3.5877664,3.874486,3.9612563,3.7763977,3.3915899,3.029418,2.757789,2.3993895,2.1088974,1.8825399,1.5580941,1.3619176,1.2147852,1.0072908,0.72811663,0.45648763,0.23013012,0.17731337,0.21881226,0.3734899,0.7432071,1.4335974,2.293756,3.6556737,5.3910813,6.911449,8.099826,9.578695,10.834979,11.465008,11.155652,11.849815,11.46878,11.329193,11.657412,11.555551,12.47607,13.913441,14.916959,14.841507,13.377728,11.578186,10.20495,9.065618,8.096053,7.3453007,6.458734,5.5797124,4.9647746,4.636556,4.3913355,3.983892,3.4745877,2.969056,2.5087957,2.0787163,1.7014539,1.4335974,1.2902378,1.2336484,1.1581959,1.0110635,0.87147635,0.7582976,0.66775465,0.5470306,0.40367088,0.36594462,0.42630664,0.5470306,0.6451189,0.6828451,0.72811663,0.7997965,0.90543,1.0336993,1.1996948,1.3770081,1.5618668,1.7580433,1.9730829,2.3616633,2.6182017,3.0331905,3.7273536,4.678055,6.039973,7.5527954,8.677037,9.193887,9.1825695,8.669493,9.009028,9.14107,8.699674,8.028146,7.5716586,7.5490227,7.454707,7.1793056,7.0284004,7.964011,8.661947,8.903395,8.650629,8.054554,7.835742,8.511042,9.280658,9.756008,9.97482,9.7296,9.797507,10.457717,11.083972,10.121953,8.729855,8.043237,8.29223,9.288202,10.423763,11.219787,12.434572,14.11339,15.954432,17.301258,17.346529,16.874952,16.588232,16.678776,16.822134,18.666948,20.066593,20.685303,20.52308,19.942095,18.851807,17.520071,16.490145,15.954432,15.7657995,16.101564,16.320375,16.497688,16.705183,17.01831,17.112627,17.222033,17.210714,17.063583,16.90136,16.807045,16.882498,16.810818,16.59955,16.573141,16.87118,17.120173,17.452164,17.761518,17.716248,0.00754525,0.00754525,0.003772625,0.00754525,0.0150905,0.00754525,0.00754525,0.00754525,0.011317875,0.0150905,0.0150905,0.02263575,0.02263575,0.02263575,0.02263575,0.030181,0.049044125,0.08677038,0.16222288,0.2565385,0.31312788,0.26031113,0.19994913,0.18863125,0.24522063,0.38858038,0.6828451,1.1204696,1.5845025,1.9504471,2.082489,2.3428001,2.6295197,2.625747,2.305074,1.9240388,1.901403,2.2786655,2.8521044,2.8898308,1.1242423,0.70170826,1.0487897,1.1204696,0.7469798,0.6149379,0.7884786,0.94692886,0.8903395,0.62625575,0.3470815,0.35462674,0.35462674,0.331991,0.28294688,0.20372175,0.12826926,0.13204187,0.1659955,0.18863125,0.17354076,0.21881226,0.3055826,0.36594462,0.35462674,0.24899325,0.19994913,0.12826926,0.06790725,0.03772625,0.03772625,0.033953626,0.049044125,0.049044125,0.030181,0.018863125,0.00754525,0.00754525,0.00754525,0.011317875,0.018863125,0.030181,0.14335975,0.39989826,0.5885295,0.20749438,0.22258487,0.32444575,0.63002837,1.1355602,1.6976813,2.1202152,2.957738,4.0517993,4.8742313,4.5460134,4.534695,5.27413,5.7079816,5.2137675,3.6028569,4.6554193,6.809588,8.461998,8.692128,7.250985,5.1156793,4.002755,3.8669407,4.7535076,6.790725,7.3981175,5.311856,3.9386206,4.7421894,7.2283497,8.937348,9.439108,9.537196,9.363655,8.371455,7.9262853,6.6247296,4.991183,3.440634,2.282438,1.8221779,1.2411937,1.0186088,1.2487389,1.6260014,2.0145817,2.3578906,2.0598533,1.2411937,0.76207024,0.5055317,0.3055826,0.16222288,0.071679875,0.02263575,0.003772625,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.018863125,0.02263575,0.033953626,0.05281675,0.06413463,0.05281675,0.026408374,0.00754525,0.0,0.00754525,0.033953626,0.06790725,0.12826926,0.22258487,0.392353,0.6828451,1.2298758,2.04099,3.0633714,4.06689,4.640329,4.3422914,3.821669,3.4859054,3.4859054,3.6896272,4.7421894,6.1795597,7.383027,7.8810134,7.356619,6.4210076,4.719554,3.0746894,1.9127209,1.2713746,1.237421,1.388326,1.5845025,1.7165444,1.7316349,1.690136,1.5958204,1.5543215,1.4750963,1.0751982,0.8903395,1.116697,1.4260522,1.5543215,1.2864652,0.9393836,0.79602385,0.6828451,0.56212115,0.52062225,0.5055317,0.4640329,0.38103512,0.2565385,0.1056335,0.06413463,0.071679875,0.056589376,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.07922512,0.10186087,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.03772625,0.06413463,0.090543,0.120724,0.16976812,0.15467763,0.10186087,0.05281675,0.026408374,0.02263575,0.018863125,0.0150905,0.026408374,0.041498873,0.030181,0.0150905,0.018863125,0.026408374,0.049044125,0.090543,0.12826926,0.15845025,0.20372175,0.27917424,0.39989826,0.5885295,0.62625575,0.62625575,0.6111652,0.5357128,0.5319401,0.58098423,0.66020936,0.68661773,0.5470306,0.2678564,0.1659955,0.19240387,0.29426476,0.4376245,0.38480774,0.271629,0.3169005,0.5696664,0.90543,0.724344,0.7167987,0.98465514,1.327964,1.2600567,0.8337501,0.58098423,0.45648763,0.38480774,0.23013012,0.150905,0.1358145,0.17731337,0.23013012,0.23013012,0.36971724,0.3772625,0.3055826,0.21503963,0.181086,0.23013012,0.1961765,0.17731337,0.1961765,0.20372175,0.30181,0.47912338,0.58098423,0.5885295,0.60362,0.4640329,0.28294688,0.1961765,0.21503963,0.2263575,0.17731337,0.15467763,0.2867195,0.6149379,1.116697,2.3805263,2.9426475,3.31991,3.7877154,4.3913355,4.67051,3.3576362,2.1390784,1.6033657,1.2261031,3.4217708,8.028146,12.543978,15.124454,14.607604,13.275867,14.898096,18.334957,20.832436,17.999193,13.434318,10.502988,8.805306,7.99042,7.756517,8.069645,8.382772,9.088254,9.7069645,8.903395,8.831716,7.2358947,5.9117036,5.59103,5.9532022,6.7077274,6.673774,5.704209,4.123479,2.7313805,2.5767028,2.9011486,2.8521044,2.3956168,2.3013012,2.3390274,2.4710693,2.6031113,2.6332922,2.4295704,2.2183034,1.8523588,1.4562333,1.0676528,0.62625575,0.32444575,0.18863125,0.1358145,0.13204187,0.21503963,0.452715,0.9016574,1.8334957,3.1840954,4.5761943,6.258785,7.635793,8.782671,9.627739,9.95973,10.321902,9.789962,9.163706,8.801534,8.605357,8.639311,10.001229,11.159425,11.227332,9.944639,8.83926,8.114917,7.5716586,7.145352,6.911449,6.270103,5.492942,4.889322,4.52715,4.247976,3.8971217,3.4368613,2.9049213,2.3692086,1.9240388,1.5845025,1.3430545,1.237421,1.2487389,1.3204187,1.1808317,1.0148361,0.875249,0.77338815,0.69039035,0.49044126,0.33953625,0.29803738,0.35839936,0.43007925,0.42630664,0.41121614,0.41876137,0.45648763,0.5319401,0.62625575,0.724344,0.8262049,0.94315624,1.0940613,1.3430545,1.599593,1.9579924,2.4484336,3.0445085,3.8820312,5.692891,7.564113,8.963757,9.737145,9.163706,8.858124,8.756263,8.703445,8.45068,8.729855,8.639311,8.431817,8.303548,8.405409,8.477088,8.503497,8.91094,9.450426,9.186342,8.959985,9.020347,9.092027,9.114662,9.265567,9.7296,10.49167,11.45369,12.061082,11.317875,10.246449,8.948667,8.345046,8.639311,9.2995205,10.299266,11.646093,12.917468,13.79649,14.079436,14.173752,14.5132885,14.939595,15.279131,15.328176,16.116653,16.803272,17.078674,16.852316,16.260014,15.471535,14.7321005,14.162435,13.856852,13.8870325,13.992666,13.88326,13.819125,13.913441,14.147344,14.2077055,14.249205,14.302021,14.468017,14.924504,14.667966,14.649103,14.652876,14.694374,15.041456,15.592259,16.06761,16.505234,16.795727,16.712729,0.00754525,0.00754525,0.003772625,0.00754525,0.0150905,0.011317875,0.00754525,0.00754525,0.00754525,0.011317875,0.0150905,0.03772625,0.03772625,0.03772625,0.033953626,0.030181,0.041498873,0.071679875,0.14335975,0.24522063,0.32821837,0.331991,0.241448,0.22258487,0.3169005,0.44894236,0.59230214,0.935611,1.4109617,1.9089483,2.2748928,2.4974778,2.4522061,2.203213,1.8825399,1.6976813,1.599593,1.6448646,2.0258996,2.1692593,0.7432071,0.4074435,0.70170826,0.7997965,0.52062225,0.32067314,0.5093044,0.694163,0.7922512,0.7809334,0.7130261,0.935611,0.9997456,0.77338815,0.35839936,0.08677038,0.08299775,0.0754525,0.08677038,0.116951376,0.16222288,0.23767537,0.331991,0.41121614,0.4376245,0.36971724,0.30935526,0.211267,0.14335975,0.10940613,0.060362,0.03772625,0.02263575,0.018863125,0.018863125,0.00754525,0.00754525,0.00754525,0.00754525,0.011317875,0.018863125,0.026408374,0.116951376,0.271629,0.36594462,0.18863125,0.10940613,0.116951376,0.13204187,0.14713238,0.19994913,0.5055317,0.7507524,1.0412445,1.297783,1.2411937,0.98842776,2.2560298,3.5764484,3.6858547,1.5580941,1.991946,4.1612053,6.089017,6.779407,6.2399216,5.8664317,5.6551647,5.994701,7.2585306,9.81637,9.756008,7.24344,5.583485,6.2361493,8.82417,10.910432,12.027128,13.072145,14.109617,14.369928,9.922004,7.7225633,5.994701,4.2291126,3.2105038,2.8143783,2.505023,2.5087957,2.8294687,3.2369123,3.5424948,3.651901,3.0860074,2.04099,1.3732355,0.875249,0.5357128,0.3055826,0.150905,0.060362,0.06413463,0.1358145,0.10940613,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.02263575,0.0452715,0.07922512,0.1056335,0.11317875,0.094315626,0.05281675,0.018863125,0.0,0.0150905,0.0754525,0.12826926,0.20372175,0.35839936,0.543258,0.56212115,0.77716076,1.2487389,1.961765,2.8634224,3.863168,4.168751,3.9499383,3.783943,3.942393,4.38379,5.3986263,6.462507,7.2660756,7.4773426,6.749226,5.8588867,4.4516973,3.0671442,2.0070364,1.3015556,1.0336993,1.0978339,1.3656902,1.690136,1.9127209,1.6561824,1.4222796,1.3241913,1.2826926,1.0148361,0.8563859,1.0638802,1.3053282,1.3468271,1.0525624,0.724344,0.60362,0.5055317,0.392353,0.35839936,0.32821837,0.32067314,0.29803738,0.2263575,0.1056335,0.060362,0.06790725,0.05281675,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.003772625,0.0,0.00754525,0.018863125,0.03772625,0.05281675,0.056589376,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.06413463,0.07922512,0.090543,0.10940613,0.17731337,0.15467763,0.10940613,0.0754525,0.06790725,0.07922512,0.05281675,0.030181,0.033953626,0.056589376,0.049044125,0.02263575,0.018863125,0.026408374,0.0452715,0.071679875,0.14713238,0.17731337,0.22258487,0.32444575,0.4979865,0.754525,0.9393836,1.1544232,1.2864652,1.0110635,0.9205205,1.0638802,1.2261031,1.2449663,1.0110635,0.60362,0.3470815,0.24899325,0.28294688,0.3734899,0.2867195,0.211267,0.27540162,0.47535074,0.6790725,0.49421388,0.66775465,1.1431054,1.5165952,1.0450171,0.47912338,0.30181,0.32821837,0.38103512,0.2867195,0.18863125,0.14713238,0.17731337,0.241448,0.2867195,0.46026024,0.44139713,0.32821837,0.1961765,0.124496624,0.14335975,0.15467763,0.18485862,0.26031113,0.38103512,0.69793564,0.8903395,0.7884786,0.4979865,0.38480774,0.31312788,0.20372175,0.14713238,0.150905,0.18863125,0.16976812,0.14335975,0.17354076,0.271629,0.40367088,1.50905,3.500996,4.134797,3.3350005,3.2067313,4.564876,3.8480775,2.5616124,1.6712729,1.6109109,3.5689032,6.752999,9.933322,12.095036,12.457208,13.124963,15.150862,17.40312,17.614386,12.385528,8.00551,5.413717,4.2102494,4.195159,5.3684454,5.994701,6.9755836,8.054554,8.541223,7.3151197,7.062354,5.666483,4.5988297,4.2894745,4.115934,4.689373,5.885295,6.149379,5.142088,3.7499893,3.289729,3.5877664,3.561358,3.078462,2.9652832,3.2670932,3.500996,3.4557245,3.1048703,2.6068838,2.323937,2.0485353,1.7995421,1.539231,1.1732863,0.7205714,0.392353,0.20749438,0.14713238,0.13204187,0.15467763,0.38480774,0.9393836,1.780679,2.7238352,4.1574326,5.119452,6.0248823,6.9755836,7.7904706,8.446907,8.552541,8.156415,7.54525,7.232122,6.8359966,7.5905213,8.182823,7.9413757,6.8473144,6.300284,5.96452,5.7419353,5.643847,5.7909794,5.6023483,4.9760923,4.221567,3.610402,3.399135,3.3915899,2.9728284,2.3956168,1.8636768,1.5354583,1.3392819,1.1657411,1.056335,1.0714256,1.2713746,1.2713746,1.1883769,1.0940613,1.0148361,0.9280658,0.694163,0.47535074,0.35839936,0.3470815,0.3734899,0.35462674,0.31312788,0.27540162,0.2678564,0.2867195,0.32444575,0.362172,0.422534,0.5093044,0.6149379,0.7582976,0.97710985,1.2713746,1.5958204,1.8448136,2.2371666,3.6028569,5.3156285,6.9265394,8.171506,8.3525915,8.518587,8.582722,8.526133,8.394091,9.190115,9.390063,9.435335,9.6201935,10.069136,10.3634,10.303039,10.220041,10.235131,10.223814,10.521852,10.069136,9.348565,8.782671,8.733627,9.367428,10.163452,11.234878,12.30253,12.679792,11.646093,10.325675,9.4013815,9.129752,9.34102,9.857869,10.631257,11.374464,11.827179,11.747954,11.68382,12.536433,13.441863,13.970031,14.139798,14.128481,14.128481,14.053028,13.826671,13.377728,12.936331,12.740154,12.581704,12.494934,12.7477,12.37421,11.868678,11.536687,11.46878,11.536687,11.608367,11.676274,11.849815,12.253486,13.023102,12.781653,12.743927,12.830698,13.053283,13.528633,14.132254,14.679284,15.252723,15.697892,15.629986,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.02263575,0.026408374,0.02263575,0.0150905,0.018863125,0.0452715,0.0452715,0.0452715,0.0452715,0.026408374,0.018863125,0.030181,0.0452715,0.07922512,0.150905,0.27540162,0.20749438,0.17354076,0.23013012,0.27917424,0.28294688,0.633801,1.1506506,1.6486372,1.9504471,1.9466745,1.6373192,1.5807298,1.8221779,1.9051756,1.3656902,1.0223814,0.69039035,0.33953625,0.056589376,0.29049212,0.5055317,0.6111652,0.5583485,0.35839936,0.38103512,0.43385187,0.5772116,0.79602385,1.026154,1.3996439,1.599593,1.3091009,0.66775465,0.27540162,0.25276586,0.15467763,0.060362,0.018863125,0.049044125,0.10186087,0.14335975,0.181086,0.23390275,0.3055826,0.26408374,0.21503963,0.211267,0.2263575,0.16222288,0.124496624,0.071679875,0.0452715,0.049044125,0.033953626,0.026408374,0.02263575,0.02263575,0.026408374,0.02263575,0.018863125,0.02263575,0.03772625,0.056589376,0.090543,0.10940613,0.1056335,0.09808825,0.09808825,0.090543,0.59607476,1.0676528,1.6637276,2.1390784,1.8749946,1.3204187,1.5128226,1.5430037,1.1355602,0.60362,0.3470815,0.56589377,0.8563859,1.3468271,2.7087448,4.4931965,5.7607985,6.617184,7.232122,7.8319697,6.7114997,6.832224,7.2660756,7.8017883,8.948667,11.099063,12.872196,14.849052,16.848543,17.938831,9.461743,6.8699503,5.7683434,4.5007415,4.1574326,4.0970707,4.2291126,4.5120597,4.8553686,5.1043615,5.138315,4.659192,3.7047176,2.6144292,2.0183544,1.2713746,0.8224323,0.51684964,0.27917424,0.12826926,0.15467763,0.2867195,0.22258487,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.09808825,0.1056335,0.13958712,0.15845025,0.15467763,0.120724,0.071679875,0.02263575,0.0,0.018863125,0.09808825,0.181086,0.27917424,0.52439487,0.7582976,0.5470306,0.47535074,0.6073926,0.9393836,1.5467763,2.5767028,3.4594972,3.7009451,3.8141239,4.036709,4.323428,4.82896,5.451443,5.9003854,5.956975,5.458988,4.7233267,3.6745367,2.7200627,1.9994912,1.3732355,1.0374719,1.0374719,1.2411937,1.5241405,1.750498,1.4600059,1.1393328,1.0412445,1.1204696,1.0450171,0.9507015,1.0299267,1.1053791,1.0450171,0.7507524,0.49044126,0.39989826,0.3470815,0.27917424,0.2263575,0.19994913,0.20749438,0.211267,0.17731337,0.10186087,0.06413463,0.0754525,0.056589376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.00754525,0.003772625,0.011317875,0.041498873,0.041498873,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.00754525,0.003772625,0.00754525,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.003772625,0.011317875,0.02263575,0.03772625,0.05281675,0.060362,0.041498873,0.026408374,0.033953626,0.06790725,0.06790725,0.049044125,0.05281675,0.08677038,0.12826926,0.09808825,0.07922512,0.0754525,0.08299775,0.07922512,0.05281675,0.03772625,0.041498873,0.05281675,0.056589376,0.1358145,0.16976812,0.21503963,0.32444575,0.5394854,0.875249,1.20724,1.659955,2.0145817,1.7014539,1.5203679,1.6373192,1.6863633,1.5543215,1.3958713,1.0374719,0.6187105,0.3169005,0.17354076,0.120724,0.07922512,0.1056335,0.15845025,0.19994913,0.20749438,0.22258487,0.5319401,0.95824677,1.1732863,0.694163,0.21503963,0.17731337,0.34330887,0.4979865,0.45648763,0.41121614,0.29426476,0.21503963,0.23390275,0.362172,0.47157812,0.3961256,0.24522063,0.116951376,0.06413463,0.13958712,0.18863125,0.25276586,0.41498876,0.7997965,1.1619685,1.1204696,0.79602385,0.38480774,0.1358145,0.071679875,0.1358145,0.181086,0.15845025,0.13204187,0.14713238,0.16222288,0.16222288,0.18485862,0.31312788,0.39989826,3.0822346,5.032682,4.8553686,3.0897799,3.6858547,4.2102494,3.3840446,1.8523588,2.1881225,3.8443048,5.3269467,7.7414265,10.8576145,13.094781,14.6302395,15.663939,14.777372,11.491416,6.258785,4.2291126,3.180323,2.8256962,3.2633207,4.98741,5.481624,6.560595,7.3377557,7.3075747,6.3417826,5.251494,4.466788,4.142342,3.9499383,3.0671442,2.927557,5.160951,7.2396674,7.8432875,6.881268,6.4021444,6.2021956,5.7381625,4.983638,4.432834,4.7572803,4.776143,4.3422914,3.5500402,2.7540162,2.4786146,2.4559789,2.4559789,2.372981,2.214531,1.5354583,0.8639311,0.41876137,0.23767537,0.19994913,0.181086,0.27917424,0.52439487,0.8978847,1.3166461,2.022127,2.7389257,3.6254926,4.5837393,5.2628117,6.477597,7.567886,8.001738,7.699928,7.0057645,6.881268,7.183078,7.201941,6.651138,5.674028,5.5004873,5.089271,4.6327834,4.3800178,4.606375,4.817642,4.425289,3.5990841,2.7426984,2.4974778,2.7238352,2.3201644,1.7655885,1.3543724,1.2223305,1.1921495,1.0714256,0.91674787,0.8526133,1.0751982,1.297783,1.4298248,1.4939595,1.4826416,1.3656902,1.1016065,0.86770374,0.724344,0.6752999,0.66020936,0.59607476,0.5394854,0.4640329,0.38480774,0.32821837,0.3055826,0.29803738,0.30935526,0.35085413,0.4074435,0.5470306,0.7092535,0.9393836,1.1732863,1.2411937,1.5430037,2.082489,2.8898308,3.9197574,5.081726,6.085244,7.333983,8.009283,7.997965,7.8810134,8.560086,9.476834,10.344538,11.080199,11.827179,12.996693,13.373956,12.294985,10.544487,10.31813,10.967021,10.257768,9.21275,8.499724,8.428044,8.529905,8.76758,9.846551,11.646093,13.200415,12.147853,11.378237,10.70671,10.170997,10.005001,9.714509,9.6201935,9.884277,10.344538,10.49167,10.227587,10.970794,11.876224,12.506252,12.823153,12.81938,12.577931,12.189351,11.759273,11.389555,11.370691,11.498961,11.608367,11.7026825,11.970539,11.223559,10.533169,9.997457,9.654147,9.488152,9.556059,9.7069645,9.978593,10.446399,11.208468,11.351829,11.544232,11.710228,11.876224,12.151625,12.566614,12.921241,13.532406,14.203933,14.222796,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.06413463,0.071679875,0.056589376,0.030181,0.018863125,0.02263575,0.041498873,0.05281675,0.0150905,0.026408374,0.08677038,0.14713238,0.2263575,0.3961256,0.482896,0.41121614,0.28294688,0.20749438,0.3055826,0.56212115,0.73566186,0.724344,0.6187105,0.7167987,1.1808317,1.8938577,2.5314314,2.6974268,1.8938577,1.20724,1.146878,0.87147635,0.31312788,0.1659955,0.8865669,0.9393836,0.66020936,0.35839936,0.32067314,0.24899325,0.24899325,0.41121614,0.62248313,0.55080324,0.41498876,0.5470306,0.77716076,0.95824677,0.94692886,0.69039035,0.41498876,0.1659955,0.0,0.0,0.02263575,0.049044125,0.07922512,0.10940613,0.120724,0.15845025,0.20372175,0.20372175,0.17354076,0.19994913,0.29426476,0.21881226,0.14713238,0.13204187,0.1056335,0.071679875,0.05281675,0.08299775,0.1358145,0.120724,0.08677038,0.049044125,0.018863125,0.00754525,0.030181,0.030181,0.02263575,0.033953626,0.06790725,0.090543,0.06790725,0.18863125,0.35462674,0.44516975,0.33576363,0.4074435,0.49044126,0.48666862,0.3961256,0.33576363,0.663982,0.663982,0.42630664,0.16976812,0.24522063,0.7092535,1.4939595,2.1390784,2.4710693,2.595566,4.1310244,8.20546,10.853842,11.034928,10.61994,13.902123,14.468017,12.966512,10.442626,8.333729,6.7680893,5.994701,5.583485,5.3156285,5.1571784,5.304311,5.2665844,5.243949,5.3609,5.692891,6.5455046,6.4738245,4.7836885,2.5087957,2.4107075,1.4600059,1.0751982,0.7809334,0.43385187,0.21503963,0.150905,0.071679875,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.060362,0.24522063,0.14713238,0.15845025,0.18863125,0.181086,0.1056335,0.056589376,0.018863125,0.0,0.0,0.0,0.16976812,0.35085413,0.39989826,0.31312788,0.23013012,0.21503963,0.29426476,0.4979865,0.87902164,1.5241405,2.5276587,3.1425967,3.3953626,3.3463185,3.127506,3.2142766,3.4368613,3.5839937,3.5424948,3.3123648,3.0897799,2.7804246,2.3880715,1.9353566,1.4335974,1.0676528,0.8865669,0.8903395,1.0450171,1.2525115,1.2525115,1.0148361,0.83752275,0.87147635,1.1280149,1.2034674,1.2864652,1.297783,1.1280149,0.6413463,0.35839936,0.271629,0.27917424,0.29803738,0.27540162,0.23767537,0.23767537,0.24522063,0.23390275,0.19994913,0.16222288,0.18863125,0.12826926,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.02263575,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.056589376,0.041498873,0.018863125,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.056589376,0.08677038,0.08677038,0.0150905,0.003772625,0.00754525,0.0150905,0.018863125,0.030181,0.030181,0.02263575,0.0150905,0.018863125,0.030181,0.06790725,0.13958712,0.150905,0.1056335,0.090543,0.056589376,0.0452715,0.056589376,0.07922512,0.090543,0.1056335,0.1358145,0.1659955,0.22258487,0.38103512,0.8941121,1.2713746,1.7467253,2.3126192,2.71629,2.4974778,2.11267,1.5618668,1.1280149,1.3732355,1.2864652,0.9016574,0.5017591,0.25276586,0.1659955,0.15467763,0.124496624,0.120724,0.14713238,0.18485862,0.15845025,0.29049212,0.4979865,0.6187105,0.41121614,0.26408374,0.19994913,0.24899325,0.41876137,0.68661773,1.1016065,0.86770374,0.52062225,0.38858038,0.59607476,0.362172,0.21503963,0.150905,0.1358145,0.0754525,0.11317875,0.241448,0.41121614,0.6790725,1.1883769,0.995973,0.543258,0.29803738,0.331991,0.32067314,0.1358145,0.1659955,0.21503963,0.21503963,0.23013012,0.20372175,0.18863125,0.21881226,0.35085413,0.65643674,1.0827434,1.6109109,3.651901,5.534441,2.516341,3.187868,4.98741,5.4212623,4.38379,4.164978,5.715527,7.8508325,11.721546,16.218515,17.987877,16.927769,16.935314,15.848798,12.717519,7.798016,4.82896,4.4177437,5.4703064,6.560595,5.9494295,5.8890676,7.1302614,7.0849895,5.6098933,4.9760923,5.3269467,5.05909,4.3686996,3.5538127,3.006782,1.871222,4.142342,7.492433,10.11818,10.725573,10.227587,9.303293,8.065872,6.809588,6.043745,5.956975,5.926794,5.772116,5.534441,5.462761,5.511805,5.1647234,4.6290107,4.0706625,3.6330378,2.8747404,1.7882242,0.86770374,0.36971724,0.32067314,0.28294688,0.26408374,0.35085413,0.58475685,0.9620194,1.5731846,2.1164427,2.686109,3.199186,3.4179983,4.3196554,6.058836,7.2924843,7.5792036,7.3868,7.786698,8.710991,9.333474,8.944894,6.94163,7.0170827,6.2361493,5.0854983,4.168751,4.2404304,4.315883,4.3800178,4.2517486,3.7763977,2.837014,2.3616633,2.033445,1.81086,1.6486372,1.4637785,1.3656902,1.2223305,1.0638802,0.9507015,0.97710985,1.3053282,1.7089992,2.0560806,2.233394,2.1353056,1.8297231,1.5807298,1.4524606,1.4411428,1.4637785,1.2940104,1.1883769,1.0223814,0.7922512,0.59607476,0.4979865,0.4074435,0.35462674,0.3470815,0.3961256,0.5055317,0.62625575,0.77338815,0.9620194,1.20724,1.3015556,1.4109617,1.6712729,2.1768045,2.9464202,3.5689032,4.3913355,5.5985756,6.8661776,7.356619,7.624475,9.348565,11.751727,13.890805,14.649103,14.637785,13.981348,11.921495,9.318384,8.68081,8.560086,7.9715567,7.654656,7.696155,7.537705,7.515069,7.8923316,8.703445,9.65792,10.148361,10.902886,11.332966,11.472552,11.2650585,10.544487,9.774872,9.318384,9.175024,9.273112,9.431562,9.525878,9.752235,10.155907,10.627484,10.895341,10.834979,10.929295,10.868933,10.559577,10.133271,10.423763,10.884023,11.204697,11.212241,10.834979,10.627484,10.170997,9.488152,8.778898,8.439363,8.341274,8.43559,8.722309,9.329701,10.514306,10.842525,11.144334,11.348056,11.3971,11.261286,11.480098,11.619685,11.84227,12.147853,12.3289385,0.011317875,0.02263575,0.02263575,0.018863125,0.011317875,0.011317875,0.030181,0.06790725,0.08299775,0.0754525,0.090543,0.15845025,0.14713238,0.120724,0.124496624,0.18485862,0.392353,0.59607476,0.76584285,0.8186596,0.63002837,0.5093044,0.3961256,0.29049212,0.211267,0.18485862,0.271629,0.392353,0.5017591,0.68661773,1.1581959,1.3958713,1.4147344,1.3619176,1.2147852,0.7809334,0.6149379,0.5281675,0.41498876,0.36971724,0.6790725,0.9016574,0.95447415,1.0110635,1.1355602,1.2864652,1.0450171,0.9016574,0.8941121,0.95824677,0.91674787,0.5470306,0.49421388,0.60362,0.7696155,0.9205205,0.9205205,0.8601585,0.7092535,0.47912338,0.2565385,0.1056335,0.06413463,0.060362,0.056589376,0.049044125,0.06413463,0.07922512,0.090543,0.116951376,0.150905,0.13958712,0.094315626,0.08677038,0.116951376,0.13204187,0.11317875,0.07922512,0.06413463,0.08299775,0.10940613,0.094315626,0.0452715,0.0150905,0.011317875,0.00754525,0.00754525,0.003772625,0.011317875,0.026408374,0.041498873,0.018863125,0.060362,0.13204187,0.19240387,0.18863125,0.76207024,0.8299775,0.59607476,0.2867195,0.12826926,0.26408374,0.3169005,0.271629,0.1659955,0.071679875,0.271629,1.6071383,3.0143273,3.983892,4.5460134,5.353355,7.001992,8.66572,9.631512,9.314611,9.95973,10.18986,9.408927,7.907422,6.8435416,6.5002327,6.7114997,7.3415284,7.888559,7.466025,7.0246277,6.439871,5.832478,5.4250345,5.5193505,6.0814714,6.085244,5.198677,3.904667,3.4859054,1.7731338,1.0487897,0.694163,0.4074435,0.2263575,0.1358145,0.07922512,0.0754525,0.11317875,0.1358145,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.06790725,0.18485862,0.17354076,0.18485862,0.181086,0.14713238,0.08299775,0.033953626,0.00754525,0.0,0.0,0.0,0.033953626,0.4074435,0.6790725,0.6451189,0.32821837,0.2565385,0.32821837,0.47157812,0.62625575,0.7432071,1.3355093,2.0108092,2.5012503,2.6785638,2.565385,2.6031113,2.8143783,3.0331905,3.2218218,3.4594972,3.4632697,2.9011486,2.293756,1.8674494,1.5430037,1.2562841,1.0714256,1.0072908,1.0638802,1.2147852,1.2826926,1.1581959,1.0186088,1.0110635,1.2261031,1.5165952,1.7542707,1.7957695,1.5354583,0.90920264,0.58098423,0.47912338,0.49044126,0.5281675,0.543258,0.5470306,0.5696664,0.58098423,0.55080324,0.4678055,0.38103512,0.29426476,0.15845025,0.02263575,0.011317875,0.02263575,0.02263575,0.018863125,0.011317875,0.011317875,0.030181,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.09808825,0.049044125,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.003772625,0.018863125,0.0150905,0.018863125,0.026408374,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.049044125,0.06413463,0.08677038,0.07922512,0.041498873,0.0150905,0.003772625,0.00754525,0.018863125,0.026408374,0.030181,0.060362,0.041498873,0.03772625,0.05281675,0.056589376,0.033953626,0.049044125,0.06790725,0.07922512,0.06790725,0.030181,0.041498873,0.056589376,0.056589376,0.07922512,0.120724,0.23013012,0.41498876,0.65643674,0.94315624,0.95824677,1.0638802,1.3392819,1.7957695,2.372981,2.4295704,2.0598533,1.931584,2.1315331,2.191895,1.6561824,1.1431054,0.69793564,0.392353,0.32821837,0.26408374,0.23767537,0.24899325,0.29426476,0.32821837,0.3055826,0.25276586,0.23013012,0.23767537,0.20372175,0.51684964,0.7884786,0.935611,1.0638802,1.478869,1.7882242,1.6637276,1.2487389,0.754525,0.47157812,0.3772625,0.35085413,0.41498876,0.5319401,0.5772116,0.67152727,0.784706,0.9922004,1.3204187,1.7655885,1.2449663,0.7054809,0.56212115,0.7205714,0.5998474,0.4074435,0.42630664,0.52062225,0.573439,0.4979865,0.5998474,0.58098423,0.4979865,0.45648763,0.59607476,0.60362,0.98842776,2.686109,4.8025517,4.6290107,2.957738,4.1762958,5.511805,5.855114,5.753253,8.201687,12.853333,15.882751,15.924251,14.071891,14.883006,15.814844,15.988385,14.784918,11.838497,7.356619,7.2924843,8.948667,10.231359,9.650374,7.907422,7.3453007,7.2585306,7.043491,6.19465,6.7039547,5.451443,4.08198,3.3764994,3.2255943,3.7009451,5.040227,6.719045,8.578949,10.850069,11.785681,11.41219,10.20495,9.073163,9.348565,9.752235,8.782671,7.6584287,6.8246784,5.9494295,5.764571,5.2099953,4.7233267,4.5196047,4.561104,4.104616,3.0520537,1.8372684,0.90543,0.69793564,0.52439487,0.422534,0.38858038,0.41876137,0.48666862,0.87147635,1.478869,2.1881225,2.806833,3.0633714,3.1576872,4.191386,6.2663302,8.722309,10.155907,11.661184,13.340002,13.947394,13.034419,10.933067,9.87296,8.499724,7.435844,7.009537,7.220804,8.484633,8.575176,8.043237,7.284939,6.549277,5.281675,4.666737,3.9348478,3.0143273,2.5389767,2.372981,2.3956168,2.3880715,2.2862108,2.173032,2.1692593,2.505023,2.7841973,2.806833,2.5502944,2.1768045,1.9164935,1.7957695,1.780679,1.7957695,1.8184053,1.8334957,1.7316349,1.4939595,1.1808317,0.87902164,0.663982,0.5357128,0.48666862,0.5055317,0.6375736,0.7809334,0.87902164,0.91674787,0.9242931,0.9922004,1.086516,1.2638294,1.569412,2.0183544,2.5502944,3.1765501,4.0216184,5.0553174,6.1078796,6.485142,7.9791017,9.786189,11.000975,10.646348,10.38981,9.344792,8.09228,7.115171,6.802043,6.85486,6.63982,6.590776,6.8473144,7.24344,7.435844,7.6697464,7.779153,7.835742,8.156415,9.099571,10.057818,10.842525,11.249968,11.057564,10.227587,9.49947,9.291975,9.7220545,10.612394,10.740664,10.235131,9.616421,9.239159,9.2844305,9.318384,9.359882,9.276885,9.171251,9.337247,10.344538,10.914205,11.102836,10.933067,10.419991,9.929549,9.393836,8.809079,8.254503,7.914967,7.8432875,8.0206,8.239413,8.548768,9.242931,10.1294985,10.763299,10.914205,10.718028,10.650121,10.487898,10.627484,10.827434,10.978339,11.072655,0.1358145,0.07922512,0.049044125,0.030181,0.07922512,0.33576363,0.19240387,0.12826926,0.12826926,0.15467763,0.14335975,0.15467763,0.15467763,0.13958712,0.16976812,0.36594462,0.754525,1.026154,1.1053791,0.9620194,0.62248313,0.5998474,0.5772116,0.452715,0.29049212,0.30935526,0.35839936,0.41121614,0.52062225,0.7432071,1.1280149,1.2826926,1.2789198,1.3053282,1.2902378,0.8865669,0.97710985,0.90920264,0.7469798,0.62248313,0.73566186,0.7582976,0.694163,0.9205205,1.3505998,1.4449154,1.237421,1.086516,0.95824677,0.8337501,0.694163,0.5017591,0.43007925,0.39989826,0.39989826,0.48666862,0.62625575,0.7696155,0.7922512,0.663982,0.44894236,0.24522063,0.14713238,0.08677038,0.041498873,0.02263575,0.026408374,0.026408374,0.033953626,0.049044125,0.06413463,0.041498873,0.041498873,0.06790725,0.120724,0.21881226,0.29426476,0.24522063,0.16976812,0.124496624,0.116951376,0.1056335,0.06413463,0.033953626,0.018863125,0.0,0.0,0.0,0.003772625,0.011317875,0.030181,0.026408374,0.056589376,0.1056335,0.15467763,0.1358145,0.6111652,0.663982,0.49044126,0.2565385,0.094315626,0.090543,0.116951376,0.13958712,0.13958712,0.094315626,0.120724,0.8224323,1.7240896,2.5389767,3.169005,3.3727267,3.9159849,5.100589,7.073672,9.820143,14.588741,12.344029,8.903395,6.9982195,6.25124,6.462507,7.250985,8.262049,8.899622,8.326183,7.5112963,7.1868505,6.749226,6.039973,5.349582,4.847823,4.436607,3.9197574,3.3123648,2.8558772,1.5543215,1.0525624,0.76207024,0.452715,0.23013012,0.211267,0.14713238,0.094315626,0.0754525,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.06790725,0.120724,0.29426476,0.27540162,0.1961765,0.124496624,0.0754525,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.211267,0.40367088,0.452715,0.35085413,0.30935526,0.31312788,0.331991,0.362172,0.4376245,0.724344,1.2940104,1.931584,2.4182527,2.546522,2.3956168,2.305074,2.372981,2.674791,3.2482302,3.169005,2.71629,2.2786655,1.9881734,1.7467253,1.5052774,1.3505998,1.2826926,1.297783,1.3807807,1.4147344,1.358145,1.2902378,1.3015556,1.478869,1.8863125,2.2711203,2.41448,2.1692593,1.4449154,0.9695646,0.784706,0.7507524,0.80734175,0.9393836,1.0487897,1.1016065,1.0789708,0.9620194,0.754525,0.60362,0.392353,0.18863125,0.05281675,0.02263575,0.030181,0.026408374,0.0150905,0.00754525,0.00754525,0.030181,0.03772625,0.026408374,0.00754525,0.0,0.0150905,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.049044125,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.00754525,0.011317875,0.018863125,0.030181,0.018863125,0.011317875,0.011317875,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.041498873,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.030181,0.0150905,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.05281675,0.08677038,0.049044125,0.05281675,0.05281675,0.03772625,0.02263575,0.011317875,0.018863125,0.026408374,0.049044125,0.120724,0.150905,0.1659955,0.15467763,0.124496624,0.08677038,0.03772625,0.02263575,0.030181,0.041498873,0.041498873,0.049044125,0.0754525,0.090543,0.094315626,0.11317875,0.211267,0.41121614,0.69039035,1.0638802,1.5882751,1.1695137,1.116697,1.2789198,1.5241405,1.7655885,1.780679,1.7957695,1.9881734,2.2069857,1.991946,1.5505489,1.237421,0.9507015,0.6752999,0.47535074,0.36594462,0.33576363,0.35085413,0.40367088,0.52062225,0.40367088,0.25276586,0.150905,0.17354076,0.39989826,0.9205205,1.3996439,1.5731846,1.5656394,1.871222,2.5616124,2.493705,2.0145817,1.4335974,0.9997456,0.88279426,0.8186596,0.7997965,0.8186596,0.875249,1.0751982,1.2751472,1.6448646,2.0183544,1.9240388,1.3920987,0.88279426,0.6149379,0.58098423,0.5055317,0.5093044,0.52062225,0.5998474,0.68661773,0.573439,0.5319401,0.51684964,0.573439,0.6828451,0.73566186,0.513077,0.83752275,1.6071383,3.1840954,6.4021444,5.8513412,6.858632,8.303548,9.397609,9.691874,9.178797,11.431054,13.641812,14.302021,13.185325,15.396083,16.252468,16.026112,14.758509,12.261031,9.540969,9.676784,10.967021,12.14408,12.377983,11.555551,11.216014,11.374464,11.491416,10.465261,8.605357,6.368191,4.5196047,3.640583,4.1310244,5.3759904,6.643593,7.5527954,8.529905,10.797253,13.577678,14.84528,14.226569,12.649611,12.3289385,9.725827,8.167733,7.3679366,6.9227667,6.3116016,5.8098426,5.062863,4.4516973,4.1008434,3.8858037,3.3463185,2.7238352,2.052308,1.4222796,1.0035182,0.8111144,0.69039035,0.6111652,0.55080324,0.49421388,0.573439,0.80734175,1.2826926,1.8938577,2.3088465,2.1692593,2.4182527,3.6669915,5.726845,7.598067,9.016574,11.442371,13.358865,13.792717,12.325166,10.9594755,9.665465,8.507269,7.8017883,8.122461,9.529651,10.095545,10.163452,9.793735,8.7600355,7.5565677,6.6549106,5.8890676,5.172269,4.5196047,4.0517993,3.8895764,3.99521,4.183841,4.1197066,3.821669,3.7990334,3.7801702,3.5764484,3.0935526,2.5502944,2.1503963,1.9806281,2.0145817,2.1051247,2.2899833,2.4559789,2.4899325,2.3314822,1.9693103,1.5543215,1.2638294,1.0601076,0.9205205,0.83752275,0.86770374,0.97333723,1.0902886,1.146878,1.0450171,0.9695646,0.995973,1.1204696,1.3355093,1.629774,2.0900342,2.6182017,3.2670932,4.063117,4.9760923,5.515578,6.1908774,7.2057137,8.216777,8.345046,7.7904706,7.273621,6.670001,6.013564,5.4891696,5.5382137,5.7079816,6.085244,6.8171334,8.114917,8.6581745,8.299775,7.654656,7.2585306,7.5792036,8.311093,9.258021,10.103089,10.801025,11.604594,10.940613,9.891823,9.4127,9.680555,10.103089,10.691619,10.412445,9.522105,8.495952,8.039464,8.07719,8.141325,8.137552,8.118689,8.262049,8.89585,9.439108,9.725827,9.74469,9.627739,9.461743,9.167479,8.756263,8.303548,7.9451485,7.752744,7.779153,7.888559,8.088508,8.52236,9.25425,9.989911,10.344538,10.280403,10.114408,9.782416,9.7069645,9.737145,9.846551,10.125726,0.34330887,0.25276586,0.181086,0.120724,0.14335975,0.40367088,0.2867195,0.24522063,0.3055826,0.38858038,0.30935526,0.19240387,0.16222288,0.181086,0.29426476,0.62248313,0.9922004,1.2600567,1.3091009,1.116697,0.7582976,0.8337501,1.0978339,1.2713746,1.2147852,0.9318384,1.1695137,1.2336484,1.1280149,0.94692886,0.8978847,0.8601585,0.8526133,0.9620194,1.0978339,0.9808825,1.3166461,1.4335974,1.3694628,1.177059,0.935611,0.8526133,0.845068,1.0638802,1.3845534,1.4147344,1.1280149,0.9695646,0.97710985,1.0186088,0.77338815,0.5281675,0.35839936,0.24899325,0.20372175,0.25276586,0.35085413,0.4640329,0.55080324,0.55457586,0.41121614,0.26408374,0.17731337,0.120724,0.07922512,0.071679875,0.030181,0.0150905,0.0150905,0.02263575,0.026408374,0.011317875,0.018863125,0.041498873,0.094315626,0.19994913,0.33953625,0.32821837,0.271629,0.22258487,0.16976812,0.124496624,0.08677038,0.056589376,0.033953626,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.026408374,0.0452715,0.0754525,0.10186087,0.071679875,0.27540162,0.30181,0.2867195,0.2867195,0.271629,0.13204187,0.06413463,0.07922512,0.14335975,0.17354076,0.094315626,0.23390275,0.7092535,1.629774,3.0746894,3.0746894,2.727608,2.7125173,3.712263,6.417235,11.385782,9.2995205,6.470052,5.587258,5.7004366,6.617184,7.594294,8.29223,8.446907,7.9036493,7.5792036,7.786698,7.4697976,6.3531003,4.9421387,4.2781568,3.2935016,2.7238352,2.6144292,2.3201644,1.2713746,0.9507015,0.7809334,0.52439487,0.30935526,0.29049212,0.1659955,0.056589376,0.0150905,0.00754525,0.056589376,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.090543,0.181086,0.19994913,0.30181,0.25276586,0.1659955,0.094315626,0.056589376,0.033953626,0.011317875,0.0,0.0,0.0,0.0,0.0452715,0.23013012,0.47912338,0.51684964,0.392353,0.35085413,0.35462674,0.38480774,0.4376245,0.4376245,0.80734175,1.3204187,1.7844516,2.022127,1.9240388,1.8070874,1.8749946,2.2673476,3.0709167,3.0218725,2.7728794,2.5087957,2.2899833,2.0749438,1.8976303,1.8070874,1.7580433,1.750498,1.7995421,1.7919968,1.7165444,1.6335466,1.6222287,1.7844516,2.2598023,2.7804246,3.0897799,2.9539654,2.1692593,1.5430037,1.2751472,1.2298758,1.3241913,1.5241405,1.6675003,1.6976813,1.6071383,1.3770081,0.98465514,0.724344,0.422534,0.18863125,0.06413463,0.03772625,0.03772625,0.02263575,0.00754525,0.0,0.0,0.0150905,0.02263575,0.026408374,0.018863125,0.00754525,0.041498873,0.05281675,0.033953626,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.018863125,0.011317875,0.02263575,0.18485862,0.21881226,0.15845025,0.056589376,0.00754525,0.00754525,0.0150905,0.026408374,0.033953626,0.018863125,0.0150905,0.02263575,0.041498873,0.05281675,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.030181,0.0150905,0.0150905,0.011317875,0.02263575,0.026408374,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.056589376,0.00754525,0.00754525,0.02263575,0.049044125,0.0754525,0.08677038,0.026408374,0.0150905,0.030181,0.049044125,0.056589376,0.049044125,0.03772625,0.030181,0.05281675,0.13958712,0.19994913,0.26408374,0.2678564,0.21881226,0.18485862,0.13958712,0.08677038,0.049044125,0.041498873,0.056589376,0.0754525,0.08677038,0.10940613,0.15467763,0.20372175,0.4074435,0.5772116,0.875249,1.3204187,1.7882242,1.327964,1.1921495,1.2600567,1.4600059,1.7618159,1.569412,2.052308,2.3918443,2.2560298,1.7919968,1.4864142,1.2789198,1.0902886,0.87902164,0.6413463,0.573439,0.44139713,0.35462674,0.3734899,0.47912338,0.33953625,0.18863125,0.09808825,0.1358145,0.38103512,0.8903395,1.297783,1.4600059,1.5731846,2.1768045,2.848332,2.6182017,2.1315331,1.7580433,1.6033657,1.539231,1.3505998,1.177059,1.1204696,1.2487389,1.4750963,1.7127718,2.0673985,2.335255,1.9730829,1.2487389,0.91674787,0.694163,0.56212115,0.76207024,0.91297525,0.8639311,0.8224323,0.8262049,0.73188925,0.5017591,0.43007925,0.62248313,0.9242931,0.9242931,0.79602385,1.1883769,1.4411428,2.1202152,5.010046,7.5263867,9.922004,11.532914,12.140307,11.974312,11.23865,11.879996,13.004238,14.011529,14.588741,18.157644,18.225552,17.274849,15.671484,11.676274,9.435335,8.654402,8.835487,9.654147,10.974566,11.276376,13.355092,14.690601,14.354838,13.015556,9.612649,7.2358947,5.8173876,5.300538,5.6287565,6.3417826,7.7187905,9.21275,10.61994,12.064855,15.24895,17.369165,17.338985,15.46399,13.472044,9.333474,7.8508325,7.3981175,7.01331,6.360646,5.4967146,4.617693,3.874486,3.2670932,2.6521554,1.961765,1.7429527,1.6675003,1.4637785,0.94315624,0.80734175,0.7696155,0.76207024,0.754525,0.73188925,0.6526641,0.58098423,0.694163,1.0412445,1.5430037,1.5430037,1.4147344,1.7655885,2.8445592,4.5422406,5.987156,8.201687,10.510533,11.936585,11.216014,10.54826,9.699419,8.782671,8.231868,8.790216,9.767326,9.982366,9.789962,9.650374,10.155907,9.144843,8.088508,7.333983,6.8661776,6.277648,5.6778007,5.383536,5.4363527,5.6400743,5.583485,5.379763,5.2590394,5.0741806,4.7233267,4.1498876,3.5990841,3.2105038,3.1425967,3.2520027,3.1010978,3.0633714,3.1425967,3.150142,2.9841464,2.6219745,2.233394,1.8674494,1.5505489,1.3015556,1.1355602,1.0827434,1.1581959,1.2864652,1.3770081,1.2902378,1.1544232,1.1242423,1.1996948,1.3656902,1.599593,1.9391292,2.3767538,2.9086938,3.5462675,4.3083377,5.0666356,5.3759904,5.7796617,6.330465,6.579458,6.398372,6.3908267,6.138061,5.587258,5.040227,4.8930945,5.0062733,5.5004873,6.6134114,8.68081,9.027891,8.533678,7.7678347,7.232122,7.364164,7.575431,7.937603,8.541223,9.563604,11.287694,11.246195,10.201178,9.593785,9.676784,9.525878,10.050273,10.020092,9.110889,7.7301087,7.0246277,7.986647,8.43559,8.428044,8.156415,7.9300575,7.99042,8.299775,8.560086,8.684583,8.809079,8.903395,8.8769865,8.692128,8.420499,8.231868,7.907422,7.624475,7.5037513,7.586749,7.8206515,8.262049,8.869441,9.378746,9.623966,9.544742,9.152389,8.801534,8.5563135,8.511042,8.782671,0.59230214,0.52439487,0.422534,0.31312788,0.23013012,0.23013012,0.3169005,0.362172,0.46026024,0.5583485,0.4678055,0.26408374,0.241448,0.32444575,0.4979865,0.8224323,0.9997456,1.1996948,1.3166461,1.2902378,1.1242423,1.5467763,2.1202152,2.584248,2.625747,1.8938577,2.323937,2.4107075,1.9806281,1.2411937,0.7696155,0.47912338,0.27540162,0.29049212,0.5281675,0.87147635,1.2864652,1.5279131,1.6524098,1.5882751,1.1732863,1.0676528,1.2110126,1.2940104,1.2638294,1.3166461,0.97333723,0.77338815,0.9620194,1.2864652,1.0072908,0.5583485,0.29426476,0.19994913,0.23013012,0.32821837,0.29803738,0.24522063,0.27917424,0.35085413,0.2565385,0.23013012,0.19240387,0.16222288,0.15467763,0.1659955,0.08677038,0.049044125,0.049044125,0.060362,0.056589376,0.026408374,0.00754525,0.0150905,0.0452715,0.08677038,0.1961765,0.24522063,0.271629,0.271629,0.20749438,0.13204187,0.090543,0.06790725,0.0452715,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0150905,0.0150905,0.10940613,0.2867195,0.41876137,0.24899325,0.1056335,0.0754525,0.14713238,0.21503963,0.13958712,0.2263575,0.7130261,1.9202662,4.2328854,4.244203,3.169005,1.8033148,0.7507524,0.422534,0.965792,1.991946,3.4444065,4.8440504,5.2892203,6.971811,7.6207023,7.605612,7.281166,6.9869013,7.4396167,7.9225125,7.6395655,6.379509,4.52715,4.4818783,3.1124156,2.2409391,2.252257,2.0862615,1.0412445,0.7582976,0.69039035,0.5583485,0.392353,0.4074435,0.22258487,0.090543,0.071679875,0.03772625,0.11317875,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.150905,0.29803738,0.31312788,0.20749438,0.33953625,0.35839936,0.18863125,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.28294688,0.724344,0.7809334,0.58475685,0.51684964,0.5470306,0.5885295,0.52062225,0.362172,0.47157812,0.65643674,0.8337501,1.0035182,1.1619685,1.3166461,1.5656394,2.0296721,2.8596497,3.0256453,2.969056,2.8030603,2.6068838,2.4333432,2.3465726,2.335255,2.3314822,2.3314822,2.4031622,2.41448,2.323937,2.1805773,2.093807,2.2107582,2.674791,3.289729,3.7914882,3.863168,3.1237335,2.3918443,2.0447628,1.9768555,2.071171,2.2069857,2.2598023,2.2107582,2.033445,1.6939086,1.1204696,0.7092535,0.36594462,0.14335975,0.0452715,0.03772625,0.03772625,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.011317875,0.05281675,0.06790725,0.049044125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.018863125,0.02263575,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.003772625,0.03772625,0.06413463,0.056589376,0.02263575,0.033953626,0.35462674,0.44894236,0.35462674,0.23390275,0.362172,0.124496624,0.05281675,0.06413463,0.090543,0.09808825,0.1056335,0.090543,0.06790725,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.02263575,0.041498873,0.033953626,0.041498873,0.0452715,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.071679875,0.124496624,0.026408374,0.026408374,0.0452715,0.06790725,0.07922512,0.056589376,0.018863125,0.00754525,0.026408374,0.060362,0.090543,0.090543,0.05281675,0.030181,0.049044125,0.120724,0.20372175,0.29803738,0.32444575,0.2867195,0.29049212,0.26408374,0.17731337,0.10940613,0.090543,0.090543,0.116951376,0.11317875,0.150905,0.23390275,0.331991,0.6111652,0.70170826,0.94315624,1.3166461,1.448688,1.2713746,1.177059,1.1921495,1.4222796,2.0447628,1.7995421,2.516341,2.8143783,2.3314822,1.7316349,1.5015048,1.2600567,1.0827434,0.9922004,0.935611,0.9205205,0.5696664,0.29426476,0.22258487,0.21503963,0.15467763,0.071679875,0.030181,0.056589376,0.15467763,0.5055317,0.65643674,0.76207024,1.1204696,2.173032,2.4220252,2.1503963,1.8825399,1.8787673,2.1390784,2.2069857,1.9202662,1.6222287,1.5430037,1.7769064,1.8938577,2.071171,2.203213,2.1881225,1.9164935,1.0487897,0.9808825,0.94692886,0.84884065,1.237421,1.4524606,1.4147344,1.3204187,1.2487389,1.20724,0.80356914,0.5394854,0.65643674,0.98842776,0.965792,1.1619685,1.7919968,2.1202152,1.9655377,1.7127718,6.587003,10.834979,12.830698,12.649611,12.076173,13.151371,14.283158,14.551015,14.426518,15.769572,20.175999,20.353312,20.055275,18.889534,12.3289385,7.9451485,5.572167,4.6327834,4.8855495,6.4247804,7.2057137,11.69891,14.286931,13.483362,11.955449,9.273112,7.7640624,7.3113475,7.3377557,6.79827,6.5228686,8.0206,10.812344,13.604086,14.317112,16.331694,17.946377,17.96524,16.0827,12.879742,10.582213,9.74469,8.937348,7.7225633,6.6586833,5.1798143,4.0178456,3.127506,2.3956168,1.6524098,0.9922004,0.8978847,1.0148361,1.0299267,0.6790725,0.6526641,0.6828451,0.7432071,0.8224323,0.91674787,0.90920264,0.8186596,0.67152727,0.62625575,0.97710985,1.1959221,1.1657411,1.2336484,1.750498,3.0746894,4.9157305,6.33801,7.8961043,9.25425,9.190115,9.537196,9.039209,8.552541,8.582722,9.25425,9.5032425,8.703445,7.4584794,7.1076255,9.737145,9.265567,8.3525915,7.673519,7.3868,7.1340337,6.620957,6.387054,6.368191,6.3531003,5.987156,6.228604,6.3644185,6.2663302,5.9494295,5.587258,5.353355,5.2137675,5.3269467,5.4476705,4.8968673,4.293247,3.9461658,3.6481283,3.3048196,2.9313297,2.6408374,2.2409391,1.8297231,1.4826416,1.2525115,1.1695137,1.2185578,1.3355093,1.448688,1.478869,1.4298248,1.3958713,1.4298248,1.5543215,1.7580433,1.9730829,2.323937,2.7502437,3.289729,4.06689,5.036454,5.6023483,5.723072,5.4967146,5.172269,5.6589375,5.753253,5.613666,5.3609,5.0968165,4.7572803,4.5309224,4.772371,5.7909794,7.8319697,8.024373,7.8923316,7.4207535,6.85486,6.7152724,6.5040054,6.1908774,6.4436436,7.6018395,9.654147,10.487898,9.899368,9.465516,9.537196,9.273112,9.469289,9.593785,8.7600355,7.2623034,6.5832305,8.835487,10.095545,10.34831,9.903141,9.371201,8.763808,8.345046,8.175279,8.167733,8.107371,8.126234,8.209232,8.235641,8.194141,8.197914,7.7942433,7.273621,6.94163,6.8774953,6.9265394,7.1906233,7.5603404,8.047009,8.52236,8.729855,8.409182,7.937603,7.4697976,7.17176,7.213259,0.8224323,0.77338815,0.6790725,0.56589377,0.4640329,0.42630664,0.56212115,0.38480774,0.18863125,0.1358145,0.26031113,0.17354076,0.44516975,0.66020936,0.6752999,0.62625575,0.68661773,0.7582976,0.84129536,1.0374719,1.5241405,3.308592,3.8178966,3.5689032,3.0256453,2.625747,2.686109,2.5917933,2.082489,1.3656902,1.0978339,0.8299775,0.47157812,0.6111652,1.177059,1.4335974,1.1544232,0.90920264,0.8601585,0.8941121,0.62625575,0.77338815,0.7092535,0.633801,0.66020936,0.7922512,0.965792,0.77716076,0.5696664,0.43385187,0.21503963,0.21503963,0.26031113,0.271629,0.25276586,0.29049212,0.33953625,0.38858038,0.4376245,0.452715,0.36594462,0.48666862,0.38103512,0.26031113,0.21503963,0.23013012,0.21503963,0.20372175,0.19240387,0.1659955,0.090543,0.041498873,0.02263575,0.033953626,0.060362,0.060362,0.03772625,0.056589376,0.08677038,0.09808825,0.060362,0.071679875,0.0754525,0.056589376,0.02263575,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.011317875,0.033953626,0.0452715,0.033953626,0.049044125,0.07922512,0.08677038,0.0150905,0.18485862,0.1358145,0.06413463,0.071679875,0.1659955,0.27917424,0.452715,0.76207024,1.2525115,1.9391292,1.5580941,0.94315624,0.46026024,0.25276586,0.23013012,0.98465514,3.9386206,7.466025,9.205205,6.058836,7.5829763,7.1038527,6.63982,6.8435416,6.9869013,6.696409,6.696409,7.062354,6.990674,4.8063245,4.244203,3.0256453,1.9127209,1.2223305,0.7922512,0.633801,0.6149379,0.5772116,0.45648763,0.26031113,0.724344,0.63002837,0.452715,0.35462674,0.18485862,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.049044125,0.07922512,0.090543,0.26408374,1.1581959,1.3694628,0.67152727,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.120724,0.41498876,0.8526133,1.0374719,0.8903395,0.67152727,0.5093044,0.41121614,0.4979865,0.33576363,0.29426476,0.44139713,0.56589377,0.7092535,0.9393836,1.2562841,1.6524098,2.0900342,2.384299,2.5578396,2.6295197,2.625747,2.5804756,2.5917933,2.6483827,2.727608,2.8294687,2.9766011,3.1463692,3.2520027,3.229367,3.1010978,2.9916916,3.259548,3.8480775,4.538468,4.927048,4.4403796,3.6707642,3.169005,2.916239,2.8294687,2.7313805,2.6106565,2.4786146,2.214531,1.7655885,1.1431054,0.6073926,0.25276586,0.06413463,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.026408374,0.08677038,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.018863125,0.003772625,0.0150905,0.1358145,0.1961765,0.16976812,0.1056335,0.1056335,0.19240387,0.21503963,0.26408374,0.63002837,1.8146327,0.63002837,0.16222288,0.056589376,0.120724,0.3055826,0.392353,0.29426476,0.17731337,0.09808825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.05281675,0.1358145,0.05281675,0.041498873,0.06413463,0.08299775,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.06413463,0.0754525,0.06413463,0.060362,0.056589376,0.0452715,0.0452715,0.0452715,0.0452715,0.056589376,0.07922512,0.090543,0.07922512,0.049044125,0.03772625,0.094315626,0.29049212,0.27917424,0.31312788,0.31312788,0.26408374,0.23013012,0.20372175,0.150905,0.1358145,0.13958712,0.090543,0.21503963,0.27917424,0.33576363,0.392353,0.44139713,0.6149379,0.83752275,0.965792,0.9620194,0.9016574,0.8865669,1.1129243,1.1921495,1.0940613,1.1280149,1.4600059,1.8070874,1.9051756,1.6486372,1.0978339,1.1581959,1.056335,1.0374719,1.2185578,1.5731846,1.3505998,0.72811663,0.271629,0.13204187,0.0452715,0.02263575,0.0150905,0.026408374,0.1056335,0.35085413,0.5470306,0.56589377,0.5319401,0.62248313,1.0978339,1.4147344,2.0258996,2.516341,2.7502437,2.8822856,2.9313297,2.7691069,2.4333432,2.1541688,2.3503454,2.214531,2.3201644,2.2296214,1.8561316,1.4637785,1.4637785,1.5580941,1.4449154,1.1431054,0.94692886,1.3241913,1.6750455,1.991946,2.2107582,2.1956677,1.539231,0.8526133,0.5281675,0.5772116,0.62625575,1.0638802,2.1466236,2.4861598,1.991946,1.8448136,4.5950575,7.643338,9.703192,10.940613,12.955194,9.891823,10.506761,11.427281,11.631002,12.434572,15.769572,19.896824,23.707176,24.122164,16.11288,8.83926,6.0211096,5.2099953,4.7648253,3.8593953,5.1798143,7.5226145,9.0807085,9.171251,8.254503,8.084735,7.9413757,7.5075235,6.749226,5.9192486,6.3342376,8.288457,11.351829,14.354838,15.380992,16.271332,16.731592,15.75071,13.687083,12.283667,14.015302,13.909668,11.853588,9.148616,8.514814,5.7079816,3.6858547,2.4295704,1.7769064,1.4335974,1.1544232,0.8563859,0.63002837,0.58098423,0.8224323,0.94692886,0.7922512,0.6111652,0.56589377,0.7469798,0.9922004,1.0601076,0.9808825,0.80734175,0.6111652,0.7809334,0.9507015,1.1431054,1.5467763,2.546522,4.3309736,6.1229706,7.564113,8.567632,9.337247,9.461743,8.601585,7.914967,7.752744,7.6923823,7.032173,6.1078796,5.0553174,4.353609,4.7912335,6.4021444,6.156924,6.0286546,6.560595,6.8661776,6.3531003,6.2436943,6.587003,6.7454534,5.402399,6.0248823,6.40969,6.519096,6.515323,6.760544,7.1981683,7.4471617,7.515069,7.3868,7.0359454,5.9117036,4.870459,3.9989824,3.31991,2.806833,2.5276587,2.2560298,1.9127209,1.50905,1.1431054,1.0223814,0.97333723,1.0902886,1.3317367,1.5430037,1.6260014,1.6561824,1.7052265,1.8070874,1.9542197,2.1956677,2.5314314,2.8634224,3.2255943,3.7990334,4.8742313,5.6363015,5.696664,5.221313,4.927048,4.9157305,4.859141,4.8402777,4.82896,4.67051,4.485651,4.459243,4.432834,4.4630156,4.7912335,6.7944975,6.6813188,5.772116,5.028909,5.0666356,5.2854476,5.20245,5.1043615,5.4212623,6.7152724,7.9828744,8.216777,8.235641,8.379,8.514814,9.601331,10.47658,9.989911,8.424272,7.5226145,9.303293,11.664956,13.328684,13.853079,13.59654,11.581959,9.4127,8.239413,8.009283,7.4471617,7.201941,7.1793056,7.281166,7.3188925,6.9869013,6.537959,6.270103,6.096562,5.987156,5.9494295,6.085244,6.330465,6.63982,6.983129,7.322665,7.3868,7.1981683,6.8397694,6.4926877,6.470052,1.7995421,1.6750455,1.5958204,1.3770081,1.0601076,0.91674787,1.0487897,1.0186088,0.8865669,0.7469798,0.7092535,0.8299775,1.2713746,1.3656902,1.0940613,1.0638802,1.056335,0.9507015,0.94315624,1.1091517,1.3920987,2.2183034,3.0671442,2.8747404,2.003264,2.2447119,2.11267,1.8674494,1.6712729,1.6033657,1.6486372,1.2223305,0.86770374,0.6413463,0.6451189,1.0186088,0.95447415,1.0035182,1.0186088,0.84884065,0.35839936,0.5319401,0.724344,0.875249,0.9695646,1.026154,1.0110635,1.4977322,1.7052265,1.4335974,1.056335,0.7809334,0.62248313,0.5394854,0.48666862,0.3734899,0.3470815,0.41121614,0.5281675,0.6451189,0.694163,0.67152727,0.5998474,0.4678055,0.3055826,0.19240387,0.13204187,0.14335975,0.18863125,0.23013012,0.2263575,0.26408374,0.23013012,0.16222288,0.09808825,0.049044125,0.02263575,0.02263575,0.041498873,0.06413463,0.09808825,0.060362,0.0452715,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.018863125,0.00754525,0.00754525,0.026408374,0.033953626,0.033953626,0.049044125,0.11317875,0.39989826,0.36594462,0.21881226,0.14713238,0.30181,0.331991,0.35462674,0.43007925,0.5696664,0.754525,0.72811663,0.55080324,0.331991,0.18863125,0.25276586,0.6375736,1.6825907,3.1916409,4.7610526,5.802297,6.300284,6.488915,6.7039547,6.971811,7.001992,6.436098,5.764571,5.20245,4.7044635,3.9650288,3.138824,2.6144292,2.1277604,1.6071383,1.1581959,1.0186088,0.965792,0.8865669,0.66775465,0.211267,0.24522063,0.5055317,0.513077,0.2263575,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.0754525,0.21503963,0.52062225,1.0186088,1.146878,0.7432071,0.02263575,0.003772625,0.0,0.1056335,0.36971724,0.7809334,0.392353,0.116951376,0.06413463,0.271629,0.7205714,1.0110635,0.9507015,0.875249,0.875249,0.76584285,0.8224323,0.513077,0.2565385,0.20749438,0.26031113,0.3169005,0.452715,0.66020936,0.9393836,1.2600567,1.6410918,1.9768555,2.214531,2.3503454,2.4069347,2.5389767,2.776652,3.0520537,3.2746384,3.3425457,3.7763977,4.191386,4.395108,4.3347464,4.0782075,4.112161,4.6327834,5.4250345,6.047518,5.832478,4.927048,4.1310244,3.4972234,3.0143273,2.6332922,2.354118,2.1353056,1.8674494,1.4901869,0.97333723,0.5055317,0.1659955,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.00754525,0.018863125,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.003772625,0.011317875,0.02263575,0.018863125,0.02263575,0.03772625,0.03772625,0.030181,0.0150905,0.0150905,0.026408374,0.041498873,0.13204187,0.3734899,0.5885295,0.633801,0.39989826,0.27917424,0.15467763,0.150905,0.3772625,0.935611,0.573439,0.27917424,0.120724,0.1056335,0.16976812,0.15845025,0.13204187,0.14713238,0.16976812,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.030181,0.0452715,0.0452715,0.03772625,0.049044125,0.049044125,0.049044125,0.03772625,0.02263575,0.011317875,0.011317875,0.011317875,0.00754525,0.0,0.0,0.011317875,0.011317875,0.02263575,0.05281675,0.10186087,0.11317875,0.08677038,0.06413463,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.033953626,0.0150905,0.011317875,0.018863125,0.018863125,0.011317875,0.02263575,0.030181,0.041498873,0.049044125,0.049044125,0.041498873,0.030181,0.060362,0.14335975,0.271629,0.38858038,0.38480774,0.3470815,0.32821837,0.32444575,0.27917424,0.15467763,0.27540162,0.42630664,0.5017591,0.5319401,0.59607476,0.633801,0.6828451,0.7167987,0.6488915,0.56589377,0.62625575,0.69793564,0.72811663,0.76584285,0.80356914,0.7394345,0.76207024,0.8941121,1.0186088,1.056335,1.20724,1.0940613,0.73188925,0.513077,0.56212115,0.5885295,0.60362,0.62248313,0.6451189,0.5998474,0.47535074,0.32067314,0.17731337,0.08299775,0.056589376,0.030181,0.018863125,0.033953626,0.08299775,0.21881226,0.33576363,0.4074435,0.4678055,0.6111652,0.86770374,1.4637785,2.2183034,2.8634224,3.0671442,2.8219235,2.4107075,2.2975287,2.4522061,2.372981,2.0636258,2.1390784,2.1692593,2.1202152,2.3428001,2.9766011,2.957738,2.5691576,2.0900342,1.7882242,1.4260522,1.2525115,1.4637785,2.0560806,2.8445592,2.282438,1.5920477,1.0638802,0.7884786,0.6488915,1.0789708,1.8787673,2.493705,3.4745877,6.4738245,7.1000805,7.6207023,7.9300575,8.114917,8.439363,7.1906233,6.9152217,8.065872,10.246449,12.204442,13.162688,14.984866,16.576914,17.010767,15.528125,13.132507,10.578441,8.650629,7.4282985,6.2889657,7.111398,8.179051,8.446907,7.914967,7.643338,8.91094,10.023865,10.38981,9.9257765,9.107117,11.3971,13.494679,15.343266,16.682549,17.052265,17.123945,17.916197,16.618414,13.622949,12.50248,13.034419,12.73261,11.3669195,9.450426,8.22055,6.587003,4.8666863,3.519859,2.6295197,1.8976303,1.6071383,1.3430545,1.0978339,0.87147635,0.6790725,0.7130261,0.77716076,0.77716076,0.724344,0.7582976,0.91674787,1.0223814,1.1053791,1.1581959,1.146878,1.1053791,0.9808825,0.91297525,1.0072908,1.3166461,2.1315331,3.6368105,5.4250345,7.009537,7.835742,8.07719,7.6282477,7.0963078,6.7944975,6.7643166,6.2021956,5.300538,4.3196554,3.5575855,3.350091,3.8895764,4.5460134,5.2250857,5.8513412,6.3417826,5.1345425,4.919503,5.251494,5.4174895,4.436607,5.100589,5.6400743,5.9117036,5.9796104,6.138061,6.6058664,6.903904,7.0548086,7.0887623,7.0585814,6.326692,5.4288073,4.644101,4.0706625,3.6368105,3.4255435,3.1840954,2.795515,2.263575,1.7316349,1.267602,1.0223814,0.95824677,1.0487897,1.297783,1.5580941,1.7429527,1.9051756,2.082489,2.3088465,2.5993385,2.8596497,3.1350515,3.4972234,4.044254,4.4931965,4.798779,4.991183,5.20245,5.66271,5.111907,4.538468,4.074435,3.742444,3.4368613,3.3123648,3.4179983,3.4557245,3.4029078,3.4972234,4.08198,4.247976,4.2630663,4.2819295,4.3083377,4.4403796,4.4403796,4.406426,4.508287,4.979865,5.613666,5.934339,6.2135134,6.620957,7.183078,7.8508325,8.36391,8.526133,8.499724,8.827943,10.182315,11.680047,12.540206,12.506252,11.838497,10.665211,9.522105,8.537451,7.748972,7.1302614,6.5832305,6.3342376,6.2625575,6.228604,6.085244,5.798525,5.5495315,5.3684454,5.2590394,5.194905,5.2326307,5.3759904,5.621211,5.9494295,6.360646,6.4511886,6.5002327,6.4511886,6.258785,5.885295,3.289729,2.8785129,2.6672459,2.463524,2.203213,1.9542197,1.9844007,1.7618159,1.5467763,1.3807807,1.0902886,1.4222796,1.7580433,1.8787673,1.81086,1.8146327,1.5807298,1.3166461,1.3958713,1.81086,2.2183034,2.3503454,2.565385,2.444661,2.123988,2.3088465,1.991946,1.4335974,1.2411937,1.5052774,1.7957695,1.6222287,1.4411428,1.1808317,0.9808825,1.20724,1.116697,1.1204696,1.1280149,0.9922004,0.5357128,0.5583485,0.56589377,0.58098423,0.6375736,0.7922512,0.76584285,0.9507015,1.3053282,1.5618668,1.2110126,0.8186596,0.59230214,0.5017591,0.482896,0.422534,0.45648763,0.48666862,0.6111652,0.8337501,1.0450171,1.2034674,1.3128735,1.267602,1.0487897,0.694163,0.4678055,0.41121614,0.41876137,0.4678055,0.5885295,0.6488915,0.513077,0.32821837,0.211267,0.23767537,0.10940613,0.090543,0.14713238,0.21503963,0.18863125,0.08299775,0.041498873,0.02263575,0.0150905,0.00754525,0.00754525,0.00754525,0.026408374,0.06413463,0.10186087,0.08299775,0.056589376,0.0452715,0.05281675,0.03772625,0.060362,0.06790725,0.056589376,0.0452715,0.06413463,0.19240387,0.17731337,0.13204187,0.120724,0.181086,0.30181,0.392353,0.44516975,0.452715,0.40367088,0.44894236,0.60362,0.5055317,0.2565385,0.41498876,0.48666862,0.84884065,1.8033148,3.5424948,6.1116524,6.5530496,6.722818,7.0359454,7.364164,7.001992,6.4511886,5.7306175,4.930821,4.104616,3.2972744,2.252257,1.6524098,1.2751472,0.9997456,0.8111144,0.76584285,0.7582976,0.7054809,0.55080324,0.29049212,0.32067314,0.30935526,0.21503963,0.07922512,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.181086,0.4640329,1.0827434,1.1808317,0.6413463,0.08677038,0.060362,0.02263575,0.05281675,0.18485862,0.392353,0.1961765,0.12826926,0.150905,0.25276586,0.47535074,0.66020936,0.66775465,0.60362,0.6451189,1.0186088,0.77338815,0.56589377,0.3772625,0.2263575,0.1358145,0.12826926,0.14713238,0.23767537,0.44894236,0.814887,1.4298248,1.659955,1.8297231,2.071171,2.3465726,2.7087448,3.2784111,3.7990334,4.0706625,3.9273026,4.3385186,4.870459,5.2288585,5.2967653,5.1269975,5.160951,5.594803,6.3116016,6.934085,6.828451,5.772116,4.727099,3.7952607,3.0256453,2.425798,2.071171,1.9504471,1.9504471,1.7693611,0.9318384,0.44139713,0.20372175,0.16222288,0.17354076,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.00754525,0.00754525,0.003772625,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.018863125,0.00754525,0.011317875,0.02263575,0.06413463,0.090543,0.08299775,0.060362,0.0452715,0.08299775,0.120724,0.16222288,0.18485862,0.1358145,0.1358145,0.35462674,0.6451189,0.784706,0.5017591,0.36594462,0.18485862,0.120724,0.241448,0.5357128,0.5017591,0.31312788,0.15845025,0.10940613,0.14713238,0.07922512,0.0754525,0.10940613,0.13958712,0.1056335,0.056589376,0.033953626,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.033953626,0.056589376,0.060362,0.0452715,0.05281675,0.0754525,0.0754525,0.056589376,0.033953626,0.0150905,0.00754525,0.00754525,0.003772625,0.0,0.0,0.011317875,0.030181,0.06413463,0.1056335,0.120724,0.14713238,0.12826926,0.090543,0.0452715,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.011317875,0.011317875,0.0,0.0,0.003772625,0.003772625,0.0,0.00754525,0.041498873,0.041498873,0.03772625,0.049044125,0.094315626,0.120724,0.271629,0.52062225,0.7469798,0.7432071,0.48666862,0.3734899,0.32444575,0.31312788,0.33576363,0.36594462,0.55080324,0.7469798,0.90543,1.0714256,1.3241913,1.2600567,1.0299267,0.7884786,0.6828451,0.55080324,0.55080324,0.6451189,0.7884786,0.90543,0.7582976,0.67152727,0.663982,0.68661773,0.6451189,0.5470306,0.543258,0.46026024,0.3055826,0.23013012,0.271629,0.29426476,0.30181,0.30935526,0.32821837,0.35839936,0.35462674,0.30181,0.211267,0.1358145,0.090543,0.0452715,0.02263575,0.0150905,0.0150905,0.08677038,0.21503963,0.35085413,0.4376245,0.38858038,0.49421388,0.8563859,1.599593,2.4710693,2.867195,2.3805263,2.0447628,2.082489,2.3390274,2.2899833,2.1692593,2.161714,2.173032,2.2409391,2.5540671,3.5689032,4.002755,3.6481283,2.8558772,2.5578396,1.9278114,1.6222287,1.5580941,1.7240896,2.1654868,2.1164427,1.7467253,1.267602,0.875249,0.72811663,0.9507015,1.629774,2.5238862,4.1008434,7.5188417,9.563604,8.971302,8.296002,8.273367,7.8395147,7.8961043,7.6207023,8.024373,9.224068,10.416218,10.27663,9.797507,9.933322,10.7557535,11.434827,12.6345215,11.69891,10.238904,9.1825695,8.790216,8.99771,8.624221,7.828197,7.24344,8.00551,8.948667,10.054046,10.70671,10.570895,9.601331,11.465008,14.109617,16.580687,18.044466,17.7917,17.591751,18.376457,17.761518,15.282904,12.400619,13.087236,13.045737,11.608367,9.465516,8.643084,7.364164,5.6551647,4.115934,3.0181,2.2975287,1.8070874,1.3543724,0.95447415,0.633801,0.4376245,0.52439487,0.7582976,0.8941121,0.8865669,0.90920264,0.8601585,0.84129536,0.8903395,1.0035182,1.1355602,1.2147852,1.2223305,1.20724,1.1921495,1.20724,1.3807807,2.033445,3.2444575,4.640329,5.402399,6.1305156,6.677546,6.9982195,6.8850408,5.945657,5.270357,4.8553686,4.349837,3.7047176,3.1840954,3.048281,3.4330888,4.0291634,4.504514,4.496969,3.6745367,3.5274043,3.6745367,3.8480775,3.904667,4.5460134,5.0138187,5.311856,5.4967146,5.6891184,5.753253,5.907931,6.013564,6.017337,5.956975,5.7192993,5.342037,4.9987283,4.7346444,4.496969,4.3724723,4.4215164,4.2630663,3.7198083,2.848332,2.2258487,1.7278622,1.3732355,1.2034674,1.2638294,1.4600059,1.7052265,1.9957186,2.3428001,2.7615614,3.138824,3.2859564,3.4481792,3.7575345,4.214022,4.647874,4.745962,4.8968673,5.2665844,5.824933,5.7796617,5.3194013,4.564876,3.7348988,3.127506,2.8558772,2.71629,2.595566,2.4974778,2.5314314,2.757789,3.0633714,3.3727267,3.6292653,3.7990334,3.893349,3.8480775,3.7650797,3.7499893,3.9159849,4.195159,4.395108,4.6554193,5.0062733,5.3759904,5.9305663,6.4474163,7.1793056,8.394091,10.344538,11.766817,12.30253,12.215759,11.800771,11.351829,10.695392,9.808825,8.7751255,7.7150183,6.7567716,6.187105,5.87775,5.572167,5.323174,5.511805,5.2665844,4.957229,4.7233267,4.6026025,4.538468,4.534695,4.6252384,4.8138695,5.093044,5.4703064,6.013564,6.1833324,6.1418333,5.9796104,5.692891,4.3347464,3.7952607,4.0404816,4.002755,3.4029078,2.746471,2.776652,2.625747,2.4220252,2.1805773,1.7919968,2.474842,2.7653341,2.8407867,2.8030603,2.7011995,2.2447119,1.7769064,1.8448136,2.463524,3.1350515,3.2821836,2.9766011,2.7502437,2.7540162,2.7691069,2.3616633,1.6825907,1.388326,1.6033657,1.8938577,1.5467763,1.3430545,1.2336484,1.2562841,1.5241405,1.5241405,1.4562333,1.5279131,1.6410918,1.3958713,1.4298248,1.20724,0.8865669,0.6111652,0.5394854,0.46026024,0.44894236,0.9695646,1.6976813,1.4977322,1.1242423,0.8978847,0.72811663,0.573439,0.43007925,0.6488915,0.8526133,1.0902886,1.3770081,1.6788181,1.8900851,2.0560806,2.1051247,1.9655377,1.5731846,1.1280149,0.9242931,0.7582976,0.6526641,0.8337501,0.7884786,0.58475685,0.38480774,0.29049212,0.33576363,0.16976812,0.211267,0.271629,0.26031113,0.18485862,0.0754525,0.030181,0.0150905,0.011317875,0.02263575,0.026408374,0.049044125,0.06790725,0.08299775,0.13204187,0.10940613,0.06790725,0.05281675,0.06790725,0.07922512,0.07922512,0.071679875,0.056589376,0.03772625,0.02263575,0.0150905,0.018863125,0.041498873,0.071679875,0.06413463,0.2263575,0.3169005,0.36971724,0.3772625,0.29803738,0.38858038,0.6752999,0.6526641,0.362172,0.38480774,0.36594462,0.7167987,1.6825907,3.31991,5.4967146,6.3153744,6.5002327,6.628502,6.8359966,6.790725,6.304056,5.666483,4.8742313,3.942393,2.9237845,1.9164935,1.2034674,0.7507524,0.55457586,0.63002837,0.754525,0.77338815,0.68661773,0.5394854,0.4376245,0.62248313,0.6752999,0.41876137,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.10186087,0.33576363,0.9242931,0.965792,0.41876137,0.09808825,0.08677038,0.033953626,0.0,0.02263575,0.10940613,0.22258487,0.26031113,0.21881226,0.17354076,0.2867195,0.38103512,0.4074435,0.33576363,0.31312788,0.6790725,0.41498876,0.34330887,0.29803738,0.21881226,0.1358145,0.10186087,0.056589376,0.05281675,0.15467763,0.41876137,0.98465514,1.1091517,1.2298758,1.5505489,2.04099,2.7615614,3.7537618,4.606375,4.957229,4.4894238,4.719554,5.2099953,5.643847,5.8702044,5.8966126,6.0286546,6.3719635,6.8737226,7.273621,7.092535,5.9909286,4.8025517,3.6896272,2.7691069,2.1202152,1.9579924,2.2409391,2.2862108,1.8070874,0.935611,0.4640329,0.2678564,0.23767537,0.23390275,0.06413463,0.06790725,0.0452715,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.018863125,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0150905,0.026408374,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.0452715,0.033953626,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.071679875,0.08299775,0.08677038,0.10186087,0.120724,0.17354076,0.18863125,0.14335975,0.09808825,0.211267,0.19240387,0.181086,0.18863125,0.20749438,0.22258487,0.27917424,0.3470815,0.482896,0.6149379,0.52439487,0.42630664,0.30181,0.27540162,0.38103512,0.58098423,0.5772116,0.35462674,0.17354076,0.1358145,0.18485862,0.09808825,0.06790725,0.071679875,0.08677038,0.1056335,0.056589376,0.03772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.003772625,0.0,0.0,0.00754525,0.0150905,0.033953626,0.03772625,0.030181,0.033953626,0.056589376,0.060362,0.049044125,0.033953626,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.018863125,0.049044125,0.08677038,0.12826926,0.1659955,0.15467763,0.14713238,0.13204187,0.10940613,0.08299775,0.06413463,0.026408374,0.02263575,0.030181,0.033953626,0.033953626,0.03772625,0.033953626,0.0150905,0.0,0.00754525,0.0,0.0,0.00754525,0.02263575,0.049044125,0.06790725,0.05281675,0.030181,0.041498873,0.10186087,0.1659955,0.3734899,0.69793564,0.95824677,0.7922512,0.5055317,0.422534,0.3961256,0.35839936,0.35839936,0.452715,0.663982,0.8865669,1.0940613,1.3317367,1.7580433,1.629774,1.2110126,0.7884786,0.663982,0.6488915,0.663982,0.9318384,1.2826926,1.1581959,0.8526133,0.83752275,0.8262049,0.6828451,0.41876137,0.3772625,0.35462674,0.31312788,0.24899325,0.18485862,0.18485862,0.16222288,0.15845025,0.18485862,0.23013012,0.27917424,0.2565385,0.2263575,0.20749438,0.19240387,0.13958712,0.07922512,0.03772625,0.02263575,0.026408374,0.06413463,0.14713238,0.24899325,0.32444575,0.29426476,0.32821837,0.46026024,0.95447415,1.6750455,2.1164427,1.6637276,1.5807298,1.8636768,2.2598023,2.2598023,2.2296214,2.1654868,2.1466236,2.2371666,2.4861598,3.150142,3.640583,3.5160866,2.938875,2.686109,2.1541688,1.9089483,1.8863125,1.961765,1.9391292,2.0145817,1.8938577,1.599593,1.2449663,1.0525624,1.237421,1.5958204,3.2935016,5.643847,6.1229706,8.710991,8.809079,8.439363,8.20546,7.2924843,7.284939,7.7942433,8.650629,9.382519,9.208978,8.443134,7.032173,6.3832817,6.85486,7.7301087,10.005001,10.533169,10.099318,9.567377,9.884277,9.944639,9.137298,7.960239,7.1566696,7.699928,8.793989,9.329701,9.680555,9.676784,8.612903,9.759781,13.268322,17.195625,19.640285,18.742401,17.595524,18.018057,17.863379,16.014793,12.377983,12.37421,12.219532,10.914205,8.865668,7.8998766,7.115171,5.594803,4.123479,3.1161883,2.6408374,2.093807,1.478869,0.88279426,0.4376245,0.29803738,0.3470815,0.55080324,0.7130261,0.7997965,0.9280658,0.9318384,0.9205205,0.8941121,0.87147635,0.8978847,1.0676528,1.2261031,1.3166461,1.3468271,1.3807807,1.3958713,1.50905,2.003264,2.806833,3.4783602,4.244203,5.1043615,5.7683434,5.8437963,4.847823,4.4139714,4.504514,4.6516466,4.515832,3.8782585,3.350091,3.2331395,3.31991,3.3689542,3.1010978,2.806833,2.8106055,2.9011486,3.0935526,3.6481283,4.195159,4.6856003,5.089271,5.3458095,5.353355,5.119452,5.1043615,5.0062733,4.779916,4.6252384,4.6516466,4.6818275,4.7535076,4.8553686,4.927048,5.0025005,5.1873593,5.451443,5.4288073,4.432834,3.6066296,2.987919,2.474842,2.0560806,1.8070874,1.7278622,1.8599042,2.1164427,2.493705,3.0746894,3.6254926,3.8405323,3.9499383,4.1197066,4.432834,4.7308717,4.7874613,4.919503,5.270357,5.8136153,6.3644185,6.3644185,5.7796617,4.7535076,3.5839937,2.9501927,2.4861598,2.1503963,1.9240388,1.8372684,1.9240388,2.1692593,2.4786146,2.8030603,3.138824,3.2935016,3.270866,3.2067313,3.199186,3.3161373,3.4632697,3.5349495,3.62172,3.7688525,3.942393,4.606375,5.311856,6.2814207,7.7150183,9.789962,11.117926,11.498961,11.419736,11.276376,11.370691,10.993429,10.099318,8.98262,7.835742,6.7869525,6.221059,5.6891184,5.1345425,4.772371,5.0666356,4.8553686,4.515832,4.236658,4.0895257,4.0178456,4.002755,4.055572,4.187614,4.4101987,4.749735,5.594803,5.9984736,6.1041074,6.0248823,5.824933,4.878004,4.515832,5.402399,5.8400235,5.05909,3.2255943,3.4217708,3.5236318,3.3953626,3.1312788,3.0709167,4.014073,4.1574326,3.9763467,3.7348988,3.4934506,2.776652,2.2107582,2.1768045,2.6597006,3.2670932,3.7877154,3.640583,3.2784111,3.0030096,2.957738,2.6521554,2.191895,1.931584,1.9542197,2.0673985,1.1657411,0.7167987,0.7884786,1.2411937,1.6976813,1.7542707,1.6448646,1.8372684,2.263575,2.3314822,2.4069347,2.1202152,1.6071383,1.0676528,0.77338815,0.48666862,0.482896,1.0035182,1.6976813,1.659955,1.4147344,1.4222796,1.2789198,0.90543,0.5772116,0.7997965,1.2147852,1.6373192,2.0296721,2.4861598,2.4710693,2.584248,2.7238352,2.746471,2.4672968,1.7769064,1.4147344,1.0601076,0.72811663,0.77338815,0.56212115,0.38480774,0.29803738,0.32067314,0.41498876,0.2678564,0.3055826,0.27917424,0.14335975,0.071679875,0.033953626,0.011317875,0.0,0.003772625,0.02263575,0.033953626,0.07922512,0.07922512,0.041498873,0.060362,0.06413463,0.049044125,0.033953626,0.03772625,0.08677038,0.056589376,0.033953626,0.02263575,0.018863125,0.02263575,0.0150905,0.02263575,0.033953626,0.041498873,0.05281675,0.17731337,0.16976812,0.17731337,0.22258487,0.19994913,0.33576363,0.5885295,0.6790725,0.5319401,0.27917424,0.45648763,0.8563859,1.6863633,2.848332,3.9461658,5.0854983,5.613666,5.775889,5.904158,6.432326,6.0022464,5.3948536,4.6026025,3.6858547,2.757789,2.0108092,1.4373702,0.98465514,0.7582976,0.98842776,1.1053791,1.086516,0.965792,0.7884786,0.6375736,0.8639311,1.2902378,0.9620194,0.090543,0.056589376,0.05281675,0.056589376,0.06790725,0.07922512,0.056589376,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.049044125,0.2678564,0.5055317,0.45648763,0.16976812,0.049044125,0.060362,0.0754525,0.10186087,0.181086,0.3734899,0.56212115,0.44516975,0.22258487,0.08677038,0.21503963,0.26408374,0.271629,0.21503963,0.1056335,0.0,0.0,0.0,0.041498873,0.10940613,0.150905,0.124496624,0.08299775,0.049044125,0.041498873,0.1056335,0.331991,0.422534,0.573439,0.90920264,1.4939595,2.505023,3.7877154,4.889322,5.342037,4.6856003,4.749735,5.142088,5.6098933,6.0022464,6.25124,6.4511886,6.6549106,6.8850408,6.9755836,6.571913,5.541986,4.327201,3.1916409,2.3428001,1.9579924,2.1277604,2.7011995,2.4522061,1.4222796,0.91674787,0.66775465,0.52062225,0.38103512,0.241448,0.19994913,0.21881226,0.150905,0.071679875,0.02263575,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.018863125,0.02263575,0.02263575,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.030181,0.05281675,0.0452715,0.018863125,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.003772625,0.05281675,0.08299775,0.071679875,0.041498873,0.026408374,0.026408374,0.018863125,0.003772625,0.003772625,0.10940613,0.150905,0.16976812,0.18863125,0.21503963,0.24899325,0.2263575,0.14335975,0.13958712,0.4640329,0.36594462,0.23767537,0.124496624,0.11317875,0.32821837,0.8601585,0.6451189,0.36594462,0.32821837,0.47157812,0.43007925,0.43385187,0.5093044,0.66020936,0.8526133,0.6790725,0.35839936,0.15845025,0.14335975,0.1961765,0.120724,0.06413463,0.03772625,0.041498873,0.06413463,0.011317875,0.00754525,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.041498873,0.03772625,0.026408374,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.02263575,0.030181,0.033953626,0.02263575,0.026408374,0.026408374,0.033953626,0.041498873,0.041498873,0.10186087,0.13958712,0.1659955,0.181086,0.15845025,0.120724,0.13204187,0.16976812,0.21881226,0.28294688,0.12826926,0.08299775,0.08299775,0.090543,0.09808825,0.11317875,0.08677038,0.0452715,0.011317875,0.02263575,0.00754525,0.003772625,0.026408374,0.071679875,0.120724,0.08677038,0.056589376,0.033953626,0.030181,0.056589376,0.16222288,0.33576363,0.6111652,0.8224323,0.6149379,0.543258,0.5093044,0.49044126,0.44894236,0.32821837,0.33953625,0.56212115,0.8186596,1.0374719,1.237421,1.6524098,1.4901869,1.1317875,0.83752275,0.73566186,0.91297525,1.056335,1.5543215,2.0787163,1.6184561,1.1393328,1.0940613,1.086516,0.91674787,0.55457586,0.58098423,0.6073926,0.543258,0.39989826,0.26408374,0.181086,0.1358145,0.12826926,0.14713238,0.15467763,0.18863125,0.13958712,0.116951376,0.150905,0.19994913,0.16976812,0.1056335,0.056589376,0.041498873,0.071679875,0.12826926,0.18863125,0.2678564,0.32821837,0.27917424,0.31312788,0.35085413,0.55080324,0.90920264,1.2298758,1.1053791,1.2826926,1.7278622,2.1881225,2.1805773,2.203213,2.2183034,2.2371666,2.293756,2.444661,2.4182527,2.5314314,2.565385,2.4974778,2.5087957,2.2673476,2.1013522,2.3163917,2.727608,2.6295197,2.233394,1.991946,1.8297231,1.690136,1.539231,1.8259505,1.7731338,4.134797,7.3490734,5.5382137,6.19465,7.4169807,7.907422,7.2396674,5.847569,5.1232247,6.651138,8.959985,10.555805,9.9257765,8.484633,7.17176,6.2361493,5.9532022,6.609639,7.9225125,8.990166,9.442881,9.397609,9.461743,9.533423,9.533423,9.039209,8.130007,7.394345,8.75249,8.703445,8.4544525,8.231868,7.3000293,8.431817,12.566614,17.384256,20.458946,19.270569,16.890041,16.516552,16.260014,14.890551,11.846043,10.661438,10.099318,9.21275,7.748972,6.126743,6.085244,5.036454,3.9008942,3.1727777,2.9200118,2.4522061,1.8033148,1.116697,0.56212115,0.35462674,0.2263575,0.23013012,0.30935526,0.44894236,0.70170826,0.935611,1.0601076,1.0336993,0.8903395,0.73566186,0.845068,0.98465514,1.1204696,1.2600567,1.4411428,1.6033657,1.6825907,1.7655885,1.991946,2.5427492,2.8294687,3.1916409,3.5387223,3.7650797,3.7613072,3.863168,4.115934,4.5912848,4.930821,4.3385186,3.9197574,3.6783094,3.3727267,3.0181,2.867195,2.6785638,2.6785638,2.8294687,3.127506,3.591539,4.002755,4.5422406,5.040227,5.292993,5.062863,4.8402777,4.745962,4.4177437,3.9159849,3.7047176,3.6594462,3.7499893,4.002755,4.3875628,4.8100967,5.1043615,5.194905,5.7494807,6.511551,6.300284,5.3986263,4.7346444,4.13857,3.5462675,3.029418,2.6672459,2.4559789,2.4031622,2.5804756,3.1237335,3.8065786,4.274384,4.5196047,4.6214657,4.7535076,4.689373,4.7421894,4.927048,5.2665844,5.80607,6.5945487,7.0963078,6.9869013,6.0776987,4.3121104,3.3689542,2.727608,2.2560298,1.8863125,1.599593,1.4373702,1.4411428,1.6260014,1.9655377,2.3880715,2.637065,2.7125173,2.7502437,2.8294687,2.9841464,3.150142,3.187868,3.1425967,3.138824,3.3576362,4.285702,5.149633,5.907931,6.590776,7.3000293,8.194141,9.061845,9.808825,10.461489,11.155652,11.072655,10.340765,9.258021,8.111144,7.1566696,6.4964604,5.66271,4.9421387,4.5422406,4.640329,4.5309224,4.2781568,4.025391,3.8405323,3.712263,3.6783094,3.7084904,3.7990334,3.9801195,4.3121104,5.119452,5.8098426,6.2625575,6.4210076,6.307829,5.7683434,5.8173876,5.994701,7.496206,8.473316,4.044254,4.4818783,4.2706113,3.9688015,4.0706625,5.036454,5.5495315,4.7874613,4.0970707,3.9461658,3.9197574,2.625747,2.4672968,2.5125682,2.2748928,1.7391801,1.8599042,2.5880208,2.5314314,1.7127718,1.5430037,1.6750455,1.7278622,1.8938577,2.1390784,2.2107582,1.3317367,0.7092535,0.80734175,1.4147344,1.6486372,1.0638802,0.7696155,0.9393836,1.4524606,1.8938577,1.4411428,1.2638294,1.2336484,1.4071891,2.0296721,1.3807807,0.72811663,0.4074435,0.41498876,0.36594462,0.3055826,1.1959221,1.690136,1.4675511,1.237421,0.69793564,0.7394345,1.1883769,1.9504471,2.9766011,2.595566,2.8332415,3.169005,3.2331395,2.806833,1.8561316,1.4335974,1.146878,0.7997965,0.3961256,0.1659955,0.071679875,0.13204187,0.392353,0.91674787,0.67152727,0.25276586,0.00754525,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.00754525,0.0150905,0.026408374,0.0754525,0.26031113,0.26031113,0.24899325,0.26408374,0.21503963,0.19994913,0.4074435,0.7130261,0.9016574,0.65643674,1.3015556,1.1242423,1.1732863,1.8599042,2.9464202,3.8971217,4.961002,6.0626082,6.7756343,6.2851934,5.9796104,5.492942,4.640329,3.5160866,2.5012503,1.9278114,1.6109109,1.4411428,1.4411428,1.7693611,1.1732863,1.0601076,1.1242423,1.1393328,0.9318384,0.79602385,0.8903395,0.69039035,0.26408374,0.27540162,0.26408374,0.27917424,0.34330887,0.3961256,0.27540162,0.056589376,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.060362,0.27917424,0.181086,0.05281675,0.011317875,0.0,0.0,0.2565385,0.52062225,0.6790725,0.76207024,0.59230214,0.3470815,0.23767537,0.26408374,0.21503963,0.116951376,0.071679875,0.03772625,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.030181,0.02263575,0.033953626,0.1056335,0.27540162,0.2867195,0.3169005,0.4074435,0.63002837,1.0676528,1.9089483,2.9615107,3.8480775,4.2819295,4.074435,4.2102494,4.606375,5.149633,5.7117543,6.1644692,6.2851934,6.1795597,6.187105,6.168242,5.5080323,4.557331,3.3840446,2.4371157,2.04099,2.3956168,2.6144292,2.3956168,1.7844516,1.0751982,0.7922512,1.20724,1.4147344,1.1242423,0.56589377,0.44139713,0.44139713,0.3055826,0.150905,0.056589376,0.030181,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.0,0.011317875,0.0150905,0.0452715,0.1056335,0.150905,0.12826926,0.13204187,0.08677038,0.0150905,0.0150905,0.05281675,0.071679875,0.071679875,0.056589376,0.0452715,0.071679875,0.049044125,0.03772625,0.1358145,0.48666862,0.633801,0.52439487,0.29803738,0.20372175,0.59607476,2.3277097,1.6524098,0.67152727,0.2867195,0.21503963,0.3470815,0.45648763,0.52062225,0.62248313,0.91674787,0.3772625,0.150905,0.071679875,0.049044125,0.060362,0.03772625,0.02263575,0.00754525,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.041498873,0.0754525,0.11317875,0.11317875,0.08299775,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.033953626,0.071679875,0.120724,0.08677038,0.0754525,0.10186087,0.11317875,0.0150905,0.0754525,0.10186087,0.094315626,0.071679875,0.060362,0.120724,0.23767537,0.3961256,0.5998474,0.87147635,0.38103512,0.22258487,0.19994913,0.20749438,0.24522063,0.2678564,0.211267,0.120724,0.0452715,0.0452715,0.02263575,0.0150905,0.05281675,0.10940613,0.120724,0.03772625,0.02263575,0.041498873,0.071679875,0.1056335,0.27917424,0.41121614,0.5696664,0.76207024,0.94692886,0.87147635,0.5998474,0.43385187,0.39989826,0.23013012,0.25276586,0.46026024,0.7167987,0.91674787,0.9922004,1.1619685,0.86770374,0.7696155,0.9808825,1.0525624,1.3468271,1.8599042,2.4069347,2.7653341,2.655928,1.629774,1.2261031,1.2034674,1.2638294,1.0676528,0.7997965,0.68661773,0.6488915,0.56589377,0.27540162,0.1056335,0.08677038,0.1056335,0.1056335,0.1056335,0.08299775,0.041498873,0.0150905,0.026408374,0.0754525,0.0754525,0.056589376,0.0452715,0.071679875,0.1659955,0.31312788,0.5055317,0.84884065,1.0374719,0.36594462,0.29426476,0.40367088,0.63002837,0.91297525,1.20724,1.50905,1.780679,1.7919968,1.6335466,1.6939086,2.293756,2.7087448,2.848332,2.7615614,2.6408374,2.8596497,3.0331905,2.727608,2.372981,3.2670932,3.2784111,3.0407357,2.9803739,3.180323,3.3878171,2.323937,1.3543724,1.0638802,1.4298248,1.8297231,1.9542197,1.9466745,3.0105548,5.9418845,11.151879,8.627994,8.262049,8.152642,7.273621,5.492942,5.6891184,7.466025,9.654147,11.5857315,13.13628,10.70671,8.488406,7.5075235,7.8319697,8.575176,9.076936,9.748463,10.574668,10.770844,8.805306,7.828197,9.186342,10.691619,11.091517,10.054046,8.835487,8.575176,8.099826,7.2283497,6.7756343,8.567632,12.064855,15.399856,17.271078,16.954176,15.049001,13.343775,12.943876,12.702429,9.246704,9.2844305,9.016574,8.058327,6.6134114,5.4778514,5.723072,5.1345425,4.266839,3.519859,3.127506,2.493705,1.9127209,1.4298248,1.026154,0.6111652,0.3169005,0.1358145,0.056589376,0.090543,0.27540162,0.3734899,0.47157812,0.6111652,0.784706,0.9318384,0.94315624,0.95447415,1.0525624,1.2449663,1.4637785,1.5505489,1.5731846,1.6524098,1.8334957,2.0900342,2.1013522,2.1315331,2.425798,3.0030096,3.663219,3.893349,3.6858547,3.3764994,3.0897799,2.7615614,3.5689032,3.832987,3.8443048,3.731126,3.4632697,2.7691069,2.2107582,2.214531,2.8332415,3.7386713,4.032936,4.195159,4.3724723,4.587512,4.745962,4.708236,4.689373,4.398881,3.8895764,3.5689032,3.2520027,3.0897799,3.2331395,3.6858547,4.3347464,4.640329,4.640329,4.776143,5.66271,8.118689,7.8621507,6.9265394,5.987156,5.311856,4.776143,4.4705606,3.6443558,2.9954643,2.8030603,2.916239,3.3538637,4.0404816,4.749735,5.2175403,5.1571784,5.0213637,4.9421387,5.1345425,5.5268955,5.783434,6.4926877,7.2094865,7.250985,6.3153744,4.4705606,3.8593953,3.3123648,2.9124665,2.6106565,2.2598023,1.8787673,1.6222287,1.5467763,1.690136,2.0447628,2.263575,2.3654358,2.4333432,2.5314314,2.71629,2.9615107,3.1048703,3.2029586,3.3576362,3.7235808,5.040227,5.745708,5.873977,5.6400743,5.43258,5.847569,6.609639,7.665974,8.873214,9.993684,10.665211,10.567122,9.797507,8.586494,7.277394,6.4134626,5.726845,5.040227,4.4215164,4.22534,4.3121104,4.3422914,4.2517486,4.0291634,3.7235808,3.6481283,3.6783094,3.7688525,3.9461658,4.2894745,4.9119577,5.6061206,6.277648,6.8435416,7.2472124,5.80607,5.832478,6.043745,6.7379084,7.3905725,6.6322746,6.387054,6.79827,7.17176,7.250985,7.2094865,6.470052,5.66271,5.1081343,4.8402777,4.5912848,3.8065786,3.108643,2.727608,2.674791,2.7540162,2.5804756,2.7011995,2.6710186,2.3805263,2.052308,2.022127,1.7391801,1.9466745,2.4522061,2.1164427,1.478869,1.086516,1.0148361,1.2751472,1.8297231,2.3767538,2.354118,2.123988,1.8636768,1.5618668,1.5505489,1.841041,2.444661,2.9766011,2.6521554,1.780679,1.931584,2.0183544,1.6033657,0.87902164,0.48666862,0.56212115,0.9695646,1.3317367,1.0525624,0.58475685,0.573439,0.7809334,1.026154,1.1808317,0.84129536,0.88279426,1.1129243,1.297783,1.1355602,1.0336993,0.8299775,0.66775465,0.58475685,0.543258,0.43007925,0.31312788,0.17731337,0.094315626,0.20749438,0.14713238,0.056589376,0.03772625,0.124496624,0.27917424,0.36971724,0.41498876,0.30181,0.1056335,0.08677038,0.06413463,0.02263575,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.011317875,0.011317875,0.0150905,0.011317875,0.0,0.0,0.00754525,0.0150905,0.018863125,0.041498873,0.116951376,0.271629,0.5394854,0.77716076,0.69039035,0.4640329,0.66775465,0.8941121,0.9280658,0.7432071,0.84129536,1.0714256,1.4373702,2.1843498,3.7877154,4.534695,4.957229,5.2628117,5.5004873,5.5797124,5.564622,5.1156793,4.349837,3.4217708,2.5276587,1.991946,1.4713237,1.0412445,0.87902164,1.2562841,0.91297525,1.0110635,1.0525624,0.8903395,0.724344,0.8224323,0.8941121,0.663982,0.2867195,0.3470815,0.16976812,0.09808825,0.73188925,1.7769064,2.0447628,1.267602,0.7167987,0.5281675,0.5281675,0.1961765,0.1358145,0.071679875,0.02263575,0.003772625,0.011317875,0.030181,0.060362,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.29426476,1.20724,0.6488915,0.0754525,0.003772625,0.0,0.0,0.05281675,0.35839936,0.7205714,0.5319401,0.48666862,0.573439,0.5055317,0.29049212,0.24899325,0.23013012,0.09808825,0.00754525,0.0,0.0,0.0,0.0,0.033953626,0.09808825,0.13958712,0.10940613,0.071679875,0.090543,0.18863125,0.35839936,0.5583485,0.7092535,0.77338815,0.8111144,0.94692886,1.4260522,1.9730829,2.7540162,3.482133,3.3915899,3.3576362,3.5689032,4.0216184,4.587512,5.028909,4.6252384,4.3800178,4.221567,4.0404816,3.6669915,3.4934506,3.2633207,3.138824,3.2859564,3.874486,3.8367596,3.3274553,2.6672459,1.9806281,1.1732863,1.0110635,1.116697,1.0827434,0.77338815,0.30935526,0.13204187,0.060362,0.06413463,0.1056335,0.13958712,0.13958712,0.1056335,0.05281675,0.0,0.0,0.011317875,0.003772625,0.003772625,0.0150905,0.02263575,0.033953626,0.0150905,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0150905,0.02263575,0.018863125,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.011317875,0.00754525,0.0150905,0.03772625,0.06790725,0.041498873,0.0452715,0.056589376,0.0754525,0.11317875,0.10940613,0.08299775,0.041498873,0.0150905,0.02263575,0.03772625,0.026408374,0.094315626,0.452715,1.4524606,1.9127209,1.0978339,0.3734899,0.24522063,0.362172,0.98465514,1.0638802,1.1242423,1.3015556,1.3241913,0.88279426,0.62625575,0.41498876,0.27540162,0.40367088,0.1961765,0.09808825,0.06413463,0.060362,0.060362,0.0452715,0.026408374,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.026408374,0.06413463,0.056589376,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.011317875,0.026408374,0.03772625,0.03772625,0.05281675,0.06790725,0.0754525,0.06413463,0.23390275,0.38480774,0.51684964,0.66020936,0.8903395,1.3430545,1.1016065,0.76207024,0.56589377,0.4074435,0.24899325,0.20372175,0.2263575,0.27917424,0.3169005,0.20372175,0.150905,0.13958712,0.16222288,0.181086,0.14713238,0.1358145,0.18863125,0.2263575,0.071679875,0.018863125,0.049044125,0.120724,0.20372175,0.29049212,0.3055826,0.26031113,0.2565385,0.41498876,0.8601585,1.0601076,1.0374719,0.95447415,0.8639311,0.694163,0.66020936,0.86770374,1.1091517,1.2940104,1.4562333,1.1657411,0.845068,0.694163,0.784706,1.0525624,1.267602,1.7618159,1.9768555,1.8070874,1.569412,1.5203679,1.5505489,1.5580941,1.3845534,0.83752275,0.6149379,0.49421388,0.5017591,0.52439487,0.29803738,0.15845025,0.11317875,0.10186087,0.08677038,0.056589376,0.033953626,0.026408374,0.041498873,0.06790725,0.08677038,0.08677038,0.08299775,0.08299775,0.13204187,0.33953625,0.3772625,0.41876137,0.5017591,0.5696664,0.4640329,0.5583485,0.76584285,0.995973,1.1506506,1.1317875,1.2110126,1.5203679,1.8599042,2.1164427,2.2560298,2.2673476,2.1277604,2.0258996,2.142851,2.625747,3.1312788,3.3538637,3.3161373,3.31991,3.9499383,4.0970707,3.6330378,3.5462675,3.9574835,4.0970707,3.4330888,2.8709676,2.372981,1.9202662,1.5128226,1.871222,1.8485862,2.0372176,3.2029586,6.296511,6.7756343,7.0963078,8.099826,9.156161,8.152642,8.710991,10.352083,11.830952,12.472299,12.185578,10.303039,8.684583,8.477088,9.763554,11.54046,12.147853,12.566614,12.989148,12.83447,10.733118,10.20495,11.133017,12.079946,12.083718,10.653893,9.627739,9.235386,8.926031,8.503497,8.130007,9.846551,11.117926,12.038446,12.355347,11.472552,10.446399,10.257768,10.506761,10.585986,9.710737,8.575176,8.016829,7.484888,6.7567716,5.9532022,5.541986,5.349582,5.142088,4.7308717,3.9574835,2.7653341,2.0258996,1.6184561,1.3355093,0.8903395,0.40367088,0.1358145,0.026408374,0.02263575,0.06790725,0.1056335,0.26408374,0.41876137,0.56589377,0.8224323,1.1053791,1.4637785,1.5958204,1.5015048,1.478869,1.5731846,1.6033657,1.5958204,1.5618668,1.5052774,1.7014539,2.0070364,2.4710693,3.0445085,3.5764484,3.1840954,2.6521554,2.2862108,2.2183034,2.3956168,2.9954643,3.8103511,4.5007415,4.8138695,4.5761943,3.8782585,3.3350005,3.1425967,3.5123138,4.678055,5.643847,5.3910813,5.1232247,5.160951,4.927048,4.0706625,3.893349,4.0480266,4.3385186,4.6931453,3.9461658,3.3915899,3.2935016,3.7575345,4.7346444,5.9494295,6.749226,7.4282985,8.409182,10.27663,10.325675,9.627739,8.541223,7.2396674,5.715527,5.05909,4.561104,3.9159849,3.2067313,2.927557,3.0822346,3.4859054,3.983892,4.4743333,4.90064,5.6551647,5.938112,5.828706,5.5570765,5.4891696,5.7683434,6.304056,6.4738245,5.9720654,4.8138695,4.191386,3.7009451,3.3764994,3.2520027,3.3576362,3.1727777,2.7200627,2.4484336,2.493705,2.6898816,3.059599,3.150142,3.180323,3.2935016,3.5953116,3.983892,4.22534,4.3083377,4.266839,4.1762958,4.1762958,4.3875628,4.466788,4.346064,4.236658,4.7874613,5.3571277,6.0814714,7.1038527,8.578949,10.461489,11.631002,11.747954,10.7218,8.729855,7.3453007,6.356873,5.5759397,4.9647746,4.6554193,4.5233774,4.5837393,4.6554193,4.6026025,4.29702,3.9989824,3.904667,4.0593443,4.376245,4.640329,5.0213637,5.5759397,6.304056,6.907676,6.7831798,6.620957,6.8133607,7.4207535,8.031919,8.243186,7.6886096,7.575431,8.07719,8.394091,8.194141,7.624475,7.805561,7.4169807,6.900131,6.488915,6.205968,5.4174895,4.5950575,4.0782075,3.9159849,3.874486,3.6443558,3.3048196,3.097325,3.0407357,2.9237845,2.938875,2.8747404,2.9539654,2.9426475,2.1466236,1.7995421,1.3204187,0.9808825,0.9507015,1.2902378,1.9240388,2.1692593,2.1277604,1.9806281,1.9730829,2.2560298,2.7879698,3.4330888,3.9763467,4.115934,3.802806,2.7011995,1.6976813,1.1280149,0.7884786,1.1846043,1.3091009,1.2789198,1.1091517,0.7432071,0.4376245,0.8299775,1.1732863,1.1695137,0.9620194,0.86770374,1.0299267,1.267602,1.358145,1.0450171,1.2147852,1.4449154,1.4260522,1.1280149,0.8262049,0.7432071,0.72811663,0.573439,0.29426476,0.15845025,0.2263575,0.15845025,0.094315626,0.10940613,0.18485862,0.24522063,0.31312788,0.24522063,0.08677038,0.09808825,0.07922512,0.030181,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.011317875,0.0,0.00754525,0.011317875,0.0452715,0.090543,0.094315626,0.29049212,0.52062225,0.6375736,0.59607476,0.46026024,0.9922004,1.146878,1.2147852,1.237421,0.9997456,0.7809334,1.0978339,1.690136,2.4974778,3.6594462,3.92353,4.3347464,4.821415,5.300538,5.6589375,5.564622,4.919503,4.1989317,3.5538127,2.7879698,2.2296214,1.6222287,1.146878,0.9808825,1.2751472,1.3920987,1.1619685,0.8299775,0.6073926,0.663982,0.573439,0.5055317,0.4074435,0.27540162,0.17354076,0.1358145,0.3055826,0.965792,1.8976303,2.3503454,1.720317,1.0978339,0.8563859,0.965792,0.97710985,0.56589377,0.30181,0.1358145,0.056589376,0.071679875,0.10186087,0.08299775,0.03772625,0.0,0.0,0.0,0.0,0.116951376,0.24899325,0.08299775,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.09808825,0.46026024,1.6146835,0.875249,0.120724,0.00754525,0.0,0.071679875,0.181086,0.41121614,0.60362,0.3169005,0.5093044,0.59607476,0.5017591,0.35462674,0.47157812,0.43385187,0.16976812,0.0,0.0,0.0,0.0,0.049044125,0.11317875,0.181086,0.26031113,0.30181,0.3055826,0.41121614,0.56212115,0.49044126,0.56589377,0.59607476,0.6073926,0.69039035,0.9695646,1.5958204,1.9693103,2.214531,2.3578906,2.305074,2.4522061,2.5880208,2.7389257,2.9049213,3.0445085,2.7389257,2.6068838,2.6408374,2.8030603,3.0030096,3.31991,3.6858547,4.0970707,4.4705606,4.636556,4.274384,3.5424948,2.7313805,1.9466745,1.1091517,0.8563859,0.8563859,0.8903395,0.724344,0.10940613,0.0452715,0.056589376,0.120724,0.211267,0.3055826,0.32821837,0.27540162,0.17731337,0.08677038,0.06413463,0.06790725,0.0452715,0.02263575,0.018863125,0.041498873,0.094315626,0.056589376,0.011317875,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.011317875,0.03772625,0.011317875,0.011317875,0.018863125,0.03772625,0.071679875,0.0754525,0.0452715,0.018863125,0.011317875,0.0150905,0.026408374,0.033953626,0.10186087,0.41498876,1.237421,1.9768555,1.2525115,0.5093044,0.32821837,0.4074435,0.66020936,0.7582976,0.9016574,1.1732863,1.5279131,0.62625575,0.392353,0.28294688,0.120724,0.120724,0.07922512,0.056589376,0.05281675,0.049044125,0.041498873,0.0452715,0.026408374,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.03772625,0.033953626,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.033953626,0.033953626,0.060362,0.116951376,0.1961765,0.23767537,0.25276586,0.29426476,0.3772625,0.5017591,0.79602385,0.69793564,0.5055317,0.35462674,0.2263575,0.18863125,0.211267,0.30181,0.4376245,0.58098423,0.52439487,0.3961256,0.331991,0.33953625,0.31312788,0.241448,0.21881226,0.24522063,0.2678564,0.16222288,0.09808825,0.1056335,0.16222288,0.2263575,0.23390275,0.24899325,0.24522063,0.271629,0.3734899,0.59230214,0.7130261,0.7997965,0.90920264,1.0186088,0.9997456,0.8865669,1.0940613,1.3505998,1.4977322,1.4901869,1.3505998,1.3053282,1.1581959,0.965792,1.026154,1.0978339,1.2525115,1.2789198,1.1619685,1.0676528,1.116697,1.1996948,1.1695137,0.97710985,0.6488915,0.60362,0.6488915,0.6413463,0.5055317,0.2678564,0.15467763,0.08299775,0.056589376,0.06413463,0.071679875,0.07922512,0.094315626,0.1056335,0.1056335,0.120724,0.09808825,0.090543,0.14713238,0.26031113,0.392353,0.41121614,0.46026024,0.51684964,0.6111652,0.8186596,1.1506506,1.4298248,1.5882751,1.5958204,1.4524606,1.388326,1.50905,1.6712729,1.8561316,2.1654868,2.282438,2.463524,2.516341,2.4710693,2.5691576,3.0256453,3.6783094,4.0291634,4.1083884,4.447925,4.515832,4.266839,4.1008434,4.104616,4.032936,4.0517993,3.500996,2.7502437,2.0787163,1.6373192,1.780679,1.7429527,1.7882242,2.505023,4.798779,4.425289,4.6856003,5.9494295,7.7829256,8.948667,10.759526,11.521597,10.95193,9.842778,10.080454,10.061591,9.880505,10.642575,12.219532,13.253232,13.12119,13.404137,13.898351,14.04171,12.917468,11.295239,10.774617,10.797253,10.823661,10.344538,10.072908,10.299266,10.763299,11.155652,11.133017,12.491161,13.283413,13.196642,12.057309,9.846551,9.061845,8.963757,9.220296,9.525878,9.590013,8.66572,7.8432875,7.1679873,6.719045,6.587003,6.8963585,7.3415284,7.352846,6.598321,4.961002,3.3840446,2.2711203,1.6561824,1.3505998,0.94315624,0.41876137,0.12826926,0.0150905,0.00754525,0.00754525,0.0150905,0.094315626,0.181086,0.30181,0.573439,0.79602385,1.1544232,1.4600059,1.6825907,1.9466745,1.9994912,2.0070364,1.9806281,1.901403,1.7240896,1.6750455,1.8749946,2.2183034,2.5578396,2.7238352,2.3767538,1.9089483,1.6750455,1.7995421,2.1956677,2.7011995,3.0709167,3.610402,4.3649273,5.1081343,4.821415,4.4177437,4.3422914,4.719554,5.353355,6.006019,5.885295,5.8211603,6.149379,6.7152724,6.156924,5.59103,5.560849,6.085244,6.6662283,6.617184,6.2436943,6.138061,6.579458,7.537705,8.443134,8.744945,9.193887,10.005001,10.846297,11.268831,10.695392,9.371201,7.726336,6.3719635,5.745708,5.243949,4.640329,3.953711,3.451952,3.259548,3.308592,3.5802212,4.093298,4.881777,6.19465,6.4549613,6.149379,5.726845,5.572167,5.692891,5.983383,6.1078796,5.87775,5.2628117,4.7233267,4.247976,3.874486,3.6368105,3.5764484,3.3915899,3.1237335,2.9351022,2.8936033,2.9728284,3.259548,3.5839937,3.7990334,3.8858037,3.953711,4.006528,3.9989824,3.9084394,3.742444,3.5274043,3.3161373,3.3274553,3.429316,3.5274043,3.5424948,3.85185,4.2706113,5.032682,6.2021956,7.6848373,9.688101,11.680047,13.068373,13.340002,12.042219,9.714509,7.8923316,6.590776,5.8136153,5.5382137,5.1873593,5.0553174,5.0062733,4.961002,4.8968673,4.821415,4.5912848,4.4894238,4.5988297,4.776143,5.0553174,5.572167,6.2399216,6.8397694,7.0057645,8.29223,8.586494,9.280658,9.895596,10.069136,9.552286,8.952439,9.039209,9.175024,8.963757,8.228095,8.941121,9.050528,8.75249,8.307321,8.031919,6.952948,6.2361493,5.666483,5.168496,4.779916,4.7044635,4.255521,4.0593443,4.2102494,4.247976,3.6481283,3.2935016,3.059599,2.7389257,2.052308,1.8146327,1.6260014,1.3807807,1.116697,1.0035182,1.1808317,1.4260522,1.6410918,1.8334957,2.1013522,2.2673476,2.8445592,3.7499893,4.7950063,5.696664,5.8702044,4.5837393,3.048281,1.9994912,1.690136,2.4371157,2.293756,1.8636768,1.4939595,1.2789198,0.9280658,1.0525624,1.2223305,1.20724,0.9808825,1.1280149,1.5430037,1.901403,1.9504471,1.5165952,1.50905,1.6071383,1.6260014,1.4600059,1.0789708,1.0751982,1.0638802,0.84129536,0.4640329,0.26408374,0.35839936,0.27540162,0.18863125,0.16222288,0.1659955,0.14335975,0.15467763,0.14713238,0.17731337,0.43385187,0.3470815,0.24899325,0.16222288,0.11317875,0.120724,0.1358145,0.1358145,0.12826926,0.10940613,0.060362,0.02263575,0.011317875,0.00754525,0.00754525,0.00754525,0.0150905,0.011317875,0.03772625,0.08299775,0.08677038,0.36594462,0.5998474,0.6413463,0.5394854,0.5583485,1.4713237,1.6863633,1.720317,1.720317,1.4637785,1.1808317,1.4335974,2.0636258,2.806833,3.2972744,3.651901,4.2630663,4.938366,5.5268955,5.915476,5.692891,4.9760923,4.353609,3.904667,3.199186,2.4107075,1.7995421,1.4298248,1.297783,1.3241913,1.3355093,1.0412445,0.65643674,0.40367088,0.48666862,0.3055826,0.25276586,0.27540162,0.28294688,0.10186087,0.30935526,0.6073926,0.97710985,1.358145,1.6524098,1.3920987,1.0035182,0.79602385,0.845068,1.0072908,0.6149379,0.36594462,0.19994913,0.1056335,0.120724,0.17354076,0.1659955,0.124496624,0.090543,0.10940613,0.071679875,0.041498873,0.13958712,0.26031113,0.08299775,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.16976812,0.4979865,1.2110126,0.6375736,0.08677038,0.00754525,0.0,0.071679875,0.181086,0.35462674,0.4979865,0.35839936,0.42630664,0.52439487,0.55457586,0.543258,0.6413463,0.5357128,0.271629,0.06413463,0.0,0.0,0.0,0.09808825,0.17731337,0.21503963,0.29049212,0.3961256,0.46026024,0.59607476,0.7130261,0.49044126,0.49044126,0.45648763,0.4979865,0.7054809,1.1657411,1.7957695,1.8599042,1.6524098,1.4222796,1.3958713,1.5958204,1.6825907,1.659955,1.5807298,1.5543215,1.629774,2.1088974,2.493705,2.7087448,3.0897799,3.380272,3.6745367,4.0291634,4.29702,4.1310244,3.470815,2.6219745,1.8259505,1.2034674,0.72811663,0.8299775,0.84129536,0.7432071,0.49421388,0.0,0.05281675,0.11317875,0.211267,0.34330887,0.48666862,0.51684964,0.44516975,0.32067314,0.19994913,0.17354076,0.12826926,0.0754525,0.030181,0.011317875,0.026408374,0.07922512,0.049044125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.003772625,0.0,0.0,0.003772625,0.0150905,0.030181,0.049044125,0.02263575,0.00754525,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.003772625,0.018863125,0.003772625,0.0,0.0,0.003772625,0.018863125,0.033953626,0.018863125,0.0150905,0.033953626,0.056589376,0.071679875,0.07922512,0.15467763,0.3961256,0.935611,1.5279131,1.1808317,0.6828451,0.46026024,0.58098423,0.8224323,0.8526133,0.80356914,0.8941121,1.4373702,0.5470306,0.29426476,0.20749438,0.090543,0.033953626,0.02263575,0.02263575,0.026408374,0.026408374,0.018863125,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.018863125,0.02263575,0.02263575,0.02263575,0.02263575,0.0150905,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.060362,0.03772625,0.030181,0.071679875,0.15845025,0.26408374,0.181086,0.094315626,0.056589376,0.071679875,0.08677038,0.18485862,0.24522063,0.23767537,0.18863125,0.16976812,0.17354076,0.2263575,0.362172,0.5772116,0.8224323,0.965792,0.8601585,0.6752999,0.5319401,0.48666862,0.3772625,0.30935526,0.28294688,0.28294688,0.24899325,0.241448,0.29049212,0.3470815,0.36594462,0.30181,0.32067314,0.38858038,0.52062225,0.62625575,0.52062225,0.52439487,0.59607476,0.7922512,1.0412445,1.1091517,0.965792,1.146878,1.3694628,1.5279131,1.6788181,1.7655885,1.7014539,1.4449154,1.1393328,1.116697,1.1959221,1.0940613,1.0186088,0.995973,0.8601585,0.7469798,0.7582976,0.72811663,0.62248313,0.5017591,0.52439487,0.573439,0.5394854,0.3961256,0.19994913,0.11317875,0.05281675,0.030181,0.03772625,0.060362,0.07922512,0.10186087,0.10186087,0.094315626,0.10186087,0.09808825,0.1358145,0.23767537,0.362172,0.38480774,0.422534,0.52062225,0.70170826,0.97710985,1.3355093,1.659955,1.9353566,1.9994912,1.8674494,1.7278622,1.629774,1.6184561,1.6335466,1.7165444,2.033445,2.2296214,2.6182017,2.9351022,3.0558262,2.9615107,3.2520027,3.85185,4.2592936,4.436607,4.82896,5.4250345,5.7306175,5.828706,5.6513925,4.9987283,5.0741806,4.927048,4.2404304,3.2029586,2.5201135,2.2220762,2.0070364,1.9353566,2.516341,4.7044635,5.1647234,4.8666863,5.409944,7.213259,9.540969,14.162435,14.939595,12.713746,9.669238,9.333474,9.371201,9.507015,10.416218,11.608367,11.442371,10.668983,10.812344,11.551778,12.3893,12.649611,10.744436,9.7220545,9.4013815,9.559832,9.929549,10.740664,11.834724,12.970284,13.913441,14.434063,14.890551,15.313085,14.996184,13.58145,11.072655,9.857869,9.107117,8.892077,9.178797,9.812597,9.042982,8.084735,7.2924843,6.888813,6.964266,7.877241,8.956212,9.092027,7.877241,5.6287565,3.9612563,2.8747404,2.173032,1.6222287,0.935611,0.44516975,0.14335975,0.02263575,0.011317875,0.0,0.003772625,0.02263575,0.049044125,0.116951376,0.29426476,0.38480774,0.6073926,0.935611,1.3128735,1.6976813,1.7693611,1.8334957,1.8938577,1.9466745,1.961765,1.9127209,2.082489,2.3465726,2.5502944,2.4823873,2.233394,1.81086,1.5618668,1.6222287,1.8825399,2.0749438,1.9730829,2.1390784,2.8256962,3.953711,4.45547,4.9685473,5.2552667,5.342037,5.50426,5.8928404,6.270103,6.820906,7.443389,7.745199,7.77538,7.3905725,7.635793,8.654402,9.699419,10.103089,9.955957,9.793735,9.793735,9.789962,10.144588,10.137043,10.287949,10.653893,10.797253,11.091517,10.521852,9.261794,7.805561,6.952948,6.485142,6.039973,5.583485,5.089271,4.5422406,4.093298,3.8367596,3.8782585,4.3083377,5.2288585,6.549277,6.85486,6.6549106,6.307829,6.0286546,5.7872066,5.9984736,6.1795597,6.085244,5.704209,5.191132,4.738417,4.3385186,3.9876647,3.6745367,3.3651814,3.229367,3.1765501,3.150142,3.1237335,3.2218218,3.5651307,3.7763977,3.731126,3.5500402,3.3651814,3.1916409,3.0633714,2.987919,2.9351022,2.9539654,2.9766011,3.0633714,3.199186,3.3312278,3.4029078,3.6179473,4.2630663,5.3873086,6.8133607,8.262049,10.367173,12.694883,14.558559,15.015047,13.030646,10.540714,8.341274,6.858632,6.1606965,5.87775,5.670255,5.50426,5.3910813,5.3873086,5.5268955,5.3269467,5.0854983,5.0062733,5.2099953,5.383536,5.692891,6.277648,7.020855,7.5301595,11.431054,11.800771,12.08749,12.468526,12.936331,13.290957,11.879996,11.242422,11.216014,11.193378,10.152134,10.559577,10.653893,10.246449,9.5032425,8.922258,7.598067,7.092535,6.628502,5.956975,5.349582,5.5004873,5.2137675,5.093044,5.1835866,5.0138187,3.640583,2.7351532,2.214531,1.9579924,1.8033148,1.5731846,1.9164935,2.0673985,1.780679,1.3505998,1.0902886,1.0751982,1.3091009,1.6448646,1.7769064,1.7240896,2.3390274,3.500996,4.8553686,5.847569,6.651138,6.8397694,5.975838,4.5309224,3.874486,4.195159,3.270866,2.5389767,2.463524,2.5201135,1.9504471,1.2864652,1.0072908,1.1355602,1.2223305,1.7957695,2.2183034,2.5427492,2.6408374,2.2107582,1.9240388,1.5203679,1.3845534,1.5128226,1.5052774,1.5769572,1.4864142,1.1506506,0.69039035,0.42630664,0.41121614,0.32821837,0.27917424,0.2867195,0.30181,0.3169005,0.23767537,0.18863125,0.3169005,0.7809334,0.6488915,0.5998474,0.4678055,0.29803738,0.35085413,0.41121614,0.44516975,0.4678055,0.4376245,0.27917424,0.094315626,0.030181,0.018863125,0.026408374,0.026408374,0.0150905,0.011317875,0.018863125,0.030181,0.018863125,0.25276586,0.49044126,0.66020936,0.79602385,1.0374719,1.6712729,2.0749438,2.3805263,2.5389767,2.323937,2.033445,2.1164427,2.535204,3.0105548,3.0256453,3.783943,4.478106,5.111907,5.6551647,6.039973,5.80607,5.221313,4.7006907,4.255521,3.5123138,2.5767028,1.9655377,1.6637276,1.5543215,1.4109617,1.0299267,0.97333723,0.8186596,0.4979865,0.3169005,0.211267,0.2565385,0.30181,0.271629,0.19240387,0.543258,0.72811663,0.7469798,0.6752999,0.66020936,0.8865669,0.9808825,0.9280658,0.7922512,0.7167987,0.72811663,0.6752999,0.6526641,0.69793564,0.8111144,0.88279426,0.8299775,0.6413463,0.41121614,0.3169005,0.32821837,0.20372175,0.08299775,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11317875,0.331991,0.5583485,0.45648763,0.17731337,0.003772625,0.003772625,0.0150905,0.018863125,0.026408374,0.181086,0.4376245,0.5470306,0.23767537,0.40367088,0.6375736,0.7167987,0.62248313,0.51684964,0.41121614,0.33576363,0.2678564,0.11317875,0.10186087,0.150905,0.18485862,0.18485862,0.21503963,0.32067314,0.42630664,0.52062225,0.5357128,0.35462674,0.38480774,0.42630664,0.573439,0.87902164,1.3355093,1.6373192,1.3543724,1.0223814,0.88279426,0.8941121,0.9695646,1.0110635,1.0035182,0.98842776,1.0789708,1.5656394,2.4861598,2.9124665,2.7917426,2.938875,2.9200118,2.7426984,2.6634734,2.6710186,2.505023,1.8636768,1.1996948,0.7092535,0.46026024,0.3772625,0.7922512,0.8262049,0.573439,0.22258487,0.041498873,0.120724,0.20372175,0.331991,0.5055317,0.6790725,0.6790725,0.58475685,0.44139713,0.3055826,0.271629,0.15845025,0.0754525,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.018863125,0.030181,0.026408374,0.011317875,0.0,0.0,0.0,0.0,0.018863125,0.09808825,0.049044125,0.0150905,0.00754525,0.0150905,0.030181,0.041498873,0.02263575,0.003772625,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.003772625,0.02263575,0.049044125,0.10186087,0.181086,0.26408374,0.27917424,0.28294688,0.32821837,0.55080324,1.1619685,1.2600567,1.2034674,0.9922004,0.76584285,0.8224323,0.9620194,1.1355602,1.0299267,0.8186596,1.1506506,0.66775465,0.35085413,0.18485862,0.116951376,0.06790725,0.018863125,0.003772625,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.060362,0.07922512,0.06790725,0.030181,0.018863125,0.00754525,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.011317875,0.03772625,0.056589376,0.030181,0.033953626,0.10186087,0.19994913,0.23390275,0.116951376,0.049044125,0.02263575,0.030181,0.05281675,0.10940613,0.16222288,0.1659955,0.1358145,0.150905,0.1659955,0.211267,0.35462674,0.58098423,0.80734175,1.1129243,1.1242423,0.8978847,0.62625575,0.60362,0.5281675,0.41121614,0.31312788,0.26408374,0.24899325,0.35462674,0.55457586,0.7092535,0.7469798,0.6375736,0.5583485,0.663982,0.88279426,1.0148361,0.73566186,0.6828451,0.6790725,0.84129536,1.1091517,1.2487389,1.0714256,1.2826926,1.4675511,1.5845025,1.961765,2.0862615,1.7580433,1.3732355,1.1959221,1.3958713,1.4977322,1.3128735,1.1959221,1.1544232,0.8601585,0.6526641,0.5998474,0.5696664,0.48666862,0.35839936,0.3169005,0.21881226,0.181086,0.19994913,0.12826926,0.06790725,0.05281675,0.03772625,0.018863125,0.018863125,0.030181,0.03772625,0.041498873,0.041498873,0.0452715,0.11317875,0.211267,0.3169005,0.39989826,0.38480774,0.44139713,0.56212115,0.87147635,1.327964,1.7240896,1.8599042,2.0749438,2.0862615,1.8976303,1.7957695,1.7429527,1.7580433,1.8184053,1.9164935,2.0560806,2.1541688,2.3692086,2.776652,3.2331395,3.3576362,3.4066803,3.6254926,3.9310753,4.3309736,4.889322,6.066381,6.8171334,7.4169807,7.6508837,6.8171334,6.587003,7.33021,7.0774446,5.4778514,3.8103511,2.8407867,2.3277097,2.1805773,2.6634734,4.3875628,7.3717093,6.8058157,6.319147,7.443389,9.635284,17.056038,19.089483,17.1164,13.445636,11.314102,9.325929,8.20546,8.22055,8.624221,7.6395655,6.692637,6.673774,7.5603404,8.959985,10.114408,9.163706,8.9788475,9.246704,9.612649,9.680555,11.129244,12.672247,14.011529,15.135772,16.335466,16.414692,16.320375,15.920478,14.969776,13.098554,11.197151,9.756008,8.993938,9.092027,10.182315,9.307066,8.337502,7.6018395,7.194396,6.990674,7.7678347,9.099571,9.442881,8.239413,5.934339,4.38379,3.6745367,3.0671442,2.1881225,1.0072908,0.44894236,0.14713238,0.030181,0.011317875,0.0,0.011317875,0.018863125,0.030181,0.0452715,0.0754525,0.10186087,0.211267,0.3772625,0.573439,0.76207024,0.91297525,1.0902886,1.2826926,1.4977322,1.7919968,2.1202152,2.474842,2.8898308,3.240685,3.2255943,2.8709676,2.3918443,2.0447628,1.8900851,1.780679,1.4750963,1.2562841,1.1657411,1.3053282,1.8334957,2.9426475,4.515832,5.2779026,5.191132,5.4703064,5.945657,6.851087,8.039464,8.888305,8.265821,8.741172,9.329701,10.393582,11.830952,13.072145,13.27964,13.223051,12.947649,12.400619,11.41219,11.947904,11.691365,11.32542,11.125471,10.955703,10.506761,9.827688,8.922258,8.013056,7.541477,7.2472124,7.020855,6.790725,6.48137,6.0286546,5.4740787,5.028909,4.8365054,5.040227,5.772116,6.6360474,7.1340337,7.2962565,7.1566696,6.752999,6.013564,6.1305156,6.3417826,6.258785,5.8513412,5.3382645,4.957229,4.636556,4.3007927,3.8895764,3.470815,3.2972744,3.289729,3.3161373,3.2105038,3.1463692,3.2972744,3.3727267,3.289729,3.169005,2.8445592,2.686109,2.776652,3.0633714,3.3878171,3.6292653,3.5575855,3.4255435,3.380272,3.4896781,3.4481792,3.4481792,3.7650797,4.5422406,5.802297,6.462507,8.080963,10.574668,13.460726,15.856343,15.818617,13.702174,10.872705,8.299775,6.571913,6.356873,6.156924,5.983383,5.8400235,5.723072,5.885295,5.9192486,5.7909794,5.6778007,5.983383,5.926794,5.8928404,6.356873,7.2170315,7.805561,17.180534,17.912424,17.629477,17.482344,17.927513,18.723537,18.161417,16.905132,16.365646,16.086473,13.717264,14.618922,13.419228,11.299012,9.103344,7.3075747,6.221059,5.987156,6.1078796,6.1418333,5.692891,5.8513412,5.643847,5.0025005,4.0480266,3.097325,2.6710186,2.5012503,2.1768045,1.7165444,1.5731846,1.6448646,1.8372684,2.093807,2.2673476,2.1202152,2.0372176,1.8221779,1.750498,1.7995421,1.6788181,2.191895,3.169005,3.3312278,2.6106565,2.1956677,5.089271,6.4436436,6.677546,6.379509,6.3153744,6.304056,4.90064,3.6934,3.2670932,3.2029586,2.595566,2.0673985,1.8523588,2.123988,2.9916916,4.7346444,4.376245,3.9688015,4.0178456,3.4934506,3.3727267,3.259548,2.727608,2.1503963,2.7011995,2.565385,2.5804756,2.2975287,1.659955,0.97710985,0.6451189,0.4376245,0.30935526,0.25276586,0.29049212,0.754525,0.7054809,0.41876137,0.14713238,0.120724,0.24522063,0.694163,0.7205714,0.3734899,0.5357128,0.6790725,0.8639311,1.0412445,1.0827434,0.77716076,0.25276586,0.094315626,0.10186087,0.124496624,0.0754525,0.0150905,0.03772625,0.1056335,0.13958712,0.030181,0.17731337,0.56212115,0.8224323,0.8903395,0.97710985,1.4524606,2.0749438,3.1124156,4.115934,3.9197574,3.2482302,2.9916916,2.9426475,2.916239,2.7313805,2.867195,3.2557755,4.134797,5.281675,6.0286546,5.8928404,5.455216,4.870459,4.183841,3.3425457,3.0105548,2.2786655,1.7240896,1.6410918,2.0447628,2.2899833,2.0749438,1.6863633,1.2336484,0.67152727,0.3772625,0.23013012,0.15845025,0.14335975,0.23013012,0.422534,0.39989826,0.32067314,0.27917424,0.3055826,1.4411428,2.282438,2.6295197,2.535204,2.305074,2.4522061,2.3578906,2.5125682,2.9954643,3.5085413,3.519859,3.0218725,2.142851,1.1581959,0.48666862,0.9280658,0.5885295,0.181086,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.24899325,0.6790725,1.0223814,0.5583485,0.1961765,0.02263575,0.026408374,0.0754525,0.10186087,0.124496624,0.19240387,0.30181,0.41121614,0.181086,0.21503963,0.3772625,0.5017591,0.36594462,0.513077,0.63002837,1.0299267,1.3468271,0.56589377,0.5017591,0.2867195,0.12826926,0.094315626,0.1056335,0.14335975,0.25276586,0.331991,0.32821837,0.24522063,0.1961765,0.28294688,0.51684964,0.8224323,1.0676528,0.95824677,0.9393836,0.8111144,0.62625575,0.68661773,0.8224323,0.8639311,0.87147635,0.95447415,1.297783,2.0787163,1.6976813,1.116697,0.8639311,1.0223814,1.0714256,0.88279426,0.7469798,0.724344,0.62625575,0.784706,0.9808825,1.0450171,0.9280658,0.67152727,0.392353,0.12826926,0.041498873,0.12826926,0.21503963,0.31312788,0.4376245,0.59607476,0.76207024,0.8865669,0.83752275,0.694163,0.5319401,0.38103512,0.26031113,0.1358145,0.05281675,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.07922512,0.150905,0.1659955,0.08677038,0.018863125,0.003772625,0.0150905,0.0150905,0.0150905,0.00754525,0.003772625,0.0150905,0.0150905,0.16222288,0.39989826,0.65643674,0.83752275,0.8639311,0.87147635,0.7054809,0.77338815,2.0296721,1.8825399,1.7731338,1.6637276,1.478869,1.1129243,0.5998474,1.086516,1.1959221,0.6488915,0.26031113,0.08677038,0.06413463,0.11317875,0.150905,0.090543,0.056589376,0.026408374,0.02263575,0.030181,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.060362,0.120724,0.19240387,0.19240387,0.116951376,0.030181,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.0452715,0.00754525,0.018863125,0.15845025,0.32067314,0.19994913,0.05281675,0.00754525,0.0,0.003772625,0.0150905,0.05281675,0.07922512,0.1056335,0.124496624,0.1358145,0.124496624,0.150905,0.22258487,0.3055826,0.3055826,0.3772625,0.46026024,0.49044126,0.47157812,0.45648763,0.56589377,0.4678055,0.30181,0.17731337,0.150905,0.2867195,0.66775465,1.1129243,1.3807807,1.1732863,0.8224323,0.9997456,1.2110126,1.2223305,1.0525624,0.88279426,0.8563859,1.0336993,1.4071891,1.9089483,1.5165952,2.022127,2.3163917,2.0485353,1.6335466,1.6071383,1.4750963,1.297783,1.3015556,1.8599042,1.4826416,1.1883769,1.0902886,1.1544232,1.1883769,0.9808825,0.8941121,0.6790725,0.3470815,0.150905,0.090543,0.06790725,0.056589376,0.056589376,0.090543,0.090543,0.071679875,0.049044125,0.030181,0.030181,0.041498873,0.03772625,0.030181,0.033953626,0.0452715,0.19240387,0.2565385,0.31312788,0.38480774,0.45648763,0.5055317,0.6111652,0.8601585,1.2110126,1.478869,1.7240896,1.8749946,1.931584,1.8938577,1.7693611,1.7580433,1.8561316,1.9579924,2.022127,2.0447628,2.2409391,2.3880715,2.41448,2.3578906,2.3805263,2.003264,2.6295197,3.5085413,4.1197066,4.1800685,4.0103,4.304565,5.0553174,6.145606,7.352846,7.854605,9.363655,9.703192,7.960239,4.4705606,2.4069347,1.7014539,2.2598023,3.1425967,2.5314314,4.217795,5.0062733,4.6554193,4.4101987,6.971811,13.370183,16.954176,18.43682,18.184053,16.218515,12.740154,9.839006,8.495952,8.2507305,7.1868505,6.319147,6.2399216,6.930312,7.9413757,8.394091,8.137552,8.952439,10.484125,11.389555,9.337247,9.654147,10.4049,11.45369,12.845788,14.784918,17.421982,17.769064,16.7995,15.086727,12.815607,10.838752,9.382519,8.677037,8.729855,9.337247,9.167479,8.201687,7.4169807,7.115171,6.881268,7.0510364,7.7376537,8.394091,8.265821,6.3644185,4.8138695,4.123479,3.5047686,2.5578396,1.2525115,0.30935526,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.05281675,0.124496624,0.20372175,0.2867195,0.3961256,0.55457586,0.7582976,0.9507015,1.0827434,1.1431054,1.8033148,2.4182527,3.2331395,4.06689,4.2894745,3.7763977,3.380272,3.2670932,3.2482302,2.806833,2.1956677,2.0258996,1.8674494,1.5769572,1.297783,1.7618159,2.6106565,3.7499893,5.0213637,6.1795597,6.643593,7.6093845,8.929804,10.265312,11.106608,11.891314,13.879487,15.362129,15.660167,15.135772,15.101818,15.128226,14.950912,14.758509,15.196134,17.625704,15.433809,13.309821,12.736382,11.993175,10.529396,9.676784,8.98262,8.360137,8.103599,8.00551,7.9791017,7.9451485,7.809334,7.492433,6.9680386,6.4436436,6.043745,5.881522,6.0286546,6.3945994,6.9152217,7.435844,7.7301087,7.5226145,6.752999,6.19465,5.8966126,5.704209,5.2628117,4.8968673,4.7233267,4.5761943,4.3422914,3.953711,3.610402,3.4330888,3.3425457,3.259548,3.1124156,3.0746894,3.2972744,3.6254926,4.036709,4.6214657,3.6707642,3.4972234,3.9914372,4.878004,5.7079816,5.938112,5.089271,4.3385186,4.063117,3.8443048,3.6368105,3.5953116,3.783943,4.214022,4.8365054,4.9119577,5.945657,7.7037,10.095545,13.185325,15.626213,15.9695215,14.045483,10.661438,7.5829763,6.5568223,6.043745,5.885295,5.915476,5.96452,6.0512905,6.4134626,6.4964604,6.3644185,6.6662283,6.1908774,6.009792,6.1418333,6.549277,7.111398,18.621677,18.289686,18.23687,18.565088,18.964987,18.723537,18.297232,17.067356,16.075155,15.565851,14.973549,14.188843,12.140307,10.367173,9.378746,8.639311,7.6697464,6.8058157,6.156924,5.7683434,5.6287565,4.938366,4.738417,4.2064767,3.308592,2.8030603,2.9426475,3.229367,3.380272,3.3123648,3.1463692,3.893349,4.1574326,3.942393,3.429316,2.9992368,3.0407357,2.9313297,2.6974268,2.5880208,3.0822346,3.2821836,3.350091,3.2633207,3.187868,3.4670424,4.123479,4.647874,5.0553174,5.4401255,5.96452,6.6624556,5.9230213,4.191386,2.3805263,1.8485862,1.991946,2.0447628,1.9881734,1.8863125,1.9051756,2.516341,3.097325,3.7952607,4.4215164,4.432834,4.195159,4.4931965,4.587512,4.22534,3.651901,3.3236825,3.6292653,4.1008434,4.085753,2.757789,2.1277604,1.6410918,1.1544232,0.7092535,0.5696664,0.73188925,0.9280658,0.91674787,0.7884786,0.98842776,1.1016065,1.0072908,0.7922512,0.5319401,0.29049212,0.543258,0.59230214,0.5583485,0.513077,0.47157812,0.3961256,0.36594462,0.29049212,0.181086,0.16222288,0.08299775,0.03772625,0.03772625,0.06413463,0.07922512,0.26408374,0.5772116,0.84129536,1.2411937,2.3314822,2.916239,3.2142766,3.6971724,4.247976,4.1272516,2.7540162,2.8030603,3.1199608,3.108643,2.7200627,2.7087448,3.5387223,4.8930945,6.3229194,7.224577,6.7379084,6.1833324,5.6476197,5.1571784,4.696918,4.745962,4.5422406,3.5764484,2.1843498,1.5316857,1.297783,1.2562841,1.3845534,1.4713237,1.1242423,0.43007925,0.14713238,0.071679875,0.08299775,0.13204187,0.16976812,0.14335975,0.181086,0.5093044,1.4411428,1.569412,3.3463185,5.251494,6.3417826,6.247467,6.9491754,9.650374,7.809334,2.3088465,1.4335974,1.750498,1.6976813,1.3128735,0.76584285,0.3772625,0.35839936,0.21881226,0.090543,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.482896,1.1204696,1.3656902,0.422534,0.07922512,0.003772625,0.00754525,0.026408374,0.071679875,0.07922512,0.07922512,0.07922512,0.08299775,0.211267,0.14713238,0.23767537,0.482896,0.52439487,0.7997965,0.9280658,0.814887,0.63002837,0.79602385,1.6637276,1.2034674,0.5357128,0.2565385,0.422534,0.65643674,0.69793564,0.4979865,0.20749438,0.16976812,0.19994913,0.331991,0.482896,0.60362,0.6526641,0.66020936,0.5017591,0.36971724,0.35085413,0.44139713,0.58475685,0.73566186,0.87147635,0.965792,0.965792,1.0072908,0.69039035,0.38858038,0.271629,0.30181,0.55457586,0.8865669,0.84884065,0.5394854,0.5885295,0.9808825,1.4034165,1.6335466,1.5505489,1.146878,0.7507524,0.5885295,0.56589377,0.59230214,0.58098423,0.69793564,0.84884065,0.98465514,1.0638802,1.0676528,0.9507015,0.7582976,0.5885295,0.4074435,0.05281675,0.026408374,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.056589376,0.049044125,0.030181,0.0452715,0.08677038,0.10186087,0.041498873,0.018863125,0.03772625,0.10186087,0.211267,0.10186087,0.06790725,0.33576363,0.8865669,1.448688,0.694163,0.38480774,0.40367088,0.70170826,1.3355093,1.3241913,1.1242423,0.9318384,0.7922512,0.5998474,0.28294688,0.3772625,0.56589377,0.633801,0.4678055,0.12826926,0.026408374,0.03772625,0.06413463,0.030181,0.02263575,0.011317875,0.00754525,0.02263575,0.030181,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.1056335,0.18485862,0.07922512,0.056589376,0.060362,0.060362,0.041498873,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.056589376,0.02263575,0.071679875,0.16976812,0.26031113,0.28294688,0.150905,0.033953626,0.0,0.0,0.0,0.003772625,0.018863125,0.026408374,0.049044125,0.06790725,0.05281675,0.049044125,0.05281675,0.09808825,0.16222288,0.16976812,0.17731337,0.24899325,0.33576363,0.3734899,0.26408374,0.28294688,0.40367088,0.513077,0.5394854,0.44516975,0.38480774,0.6375736,1.0412445,1.3468271,1.1883769,1.8863125,2.7841973,3.2369123,3.0709167,2.5804756,1.7542707,1.6033657,1.8749946,2.2598023,2.3578906,2.282438,2.6219745,2.867195,2.7615614,2.3163917,2.565385,2.6521554,2.6068838,2.4786146,2.323937,1.7240896,1.3694628,1.1204696,0.87902164,0.59230214,0.3961256,0.271629,0.17354076,0.090543,0.030181,0.018863125,0.0150905,0.030181,0.071679875,0.12826926,0.10940613,0.06413463,0.030181,0.018863125,0.018863125,0.02263575,0.026408374,0.030181,0.03772625,0.071679875,0.14713238,0.26031113,0.38103512,0.45648763,0.43385187,0.6073926,0.84129536,1.0714256,1.2600567,1.3807807,1.4524606,1.50905,1.5241405,1.5015048,1.478869,1.5052774,1.6486372,1.8825399,2.1315331,2.263575,2.293756,2.4899325,2.6446102,2.6672459,2.5767028,2.4031622,2.7238352,3.6066296,4.5724216,4.5950575,4.979865,5.511805,6.126743,7.039718,8.744945,11.18206,11.566868,11.747954,11.634775,9.205205,6.8133607,5.462761,4.930821,4.908185,5.010046,7.0849895,8.382772,7.2924843,4.957229,5.2779026,10.344538,15.728074,19.723284,20.043957,13.837989,8.729855,6.541732,6.126743,6.2135134,5.4174895,4.851596,5.0553174,5.8211603,6.964266,8.296002,7.665974,8.009283,9.148616,10.250222,9.789962,8.809079,9.291975,10.265312,11.249968,12.234623,14.079436,15.294222,15.241405,13.890805,11.815862,10.016319,8.360137,7.1981683,6.677546,6.749226,7.4396167,8.224322,9.092027,9.684328,9.288202,8.160188,7.4396167,6.8397694,6.0550632,4.776143,4.2706113,3.9159849,3.4783602,2.7389257,1.4713237,0.5394854,0.13958712,0.02263575,0.011317875,0.0,0.0,0.0,0.011317875,0.026408374,0.041498873,0.06790725,0.116951376,0.18863125,0.271629,0.32444575,0.452715,0.62625575,0.80356914,0.9695646,1.1581959,1.4939595,1.8787673,2.3503454,2.8407867,3.1765501,3.1539145,3.0709167,2.9841464,2.9086938,2.8332415,2.5917933,2.776652,2.8936033,2.746471,2.444661,2.5087957,2.8030603,3.2444575,3.832987,4.6290107,6.673774,9.092027,11.876224,14.973549,18.297232,21.65864,23.654358,22.813063,19.783646,17.346529,16.52787,16.146835,16.158154,16.761772,18.421728,19.979822,18.293459,15.55076,13.000465,10.967021,9.895596,9.163706,8.624221,8.243186,8.103599,8.190369,8.314865,8.416726,8.428044,8.284684,7.9451485,7.4584794,6.952948,6.511551,6.2097406,6.2361493,6.56814,7.149124,7.8017883,8.216777,7.635793,7.020855,6.436098,5.904158,5.3873086,5.0213637,4.847823,4.7572803,4.5799665,4.063117,3.7990334,3.8820312,3.8895764,3.7009451,3.5160866,3.6745367,3.8103511,4.08198,4.429062,4.5761943,4.315883,4.353609,4.606375,4.9534564,5.2175403,5.2250857,4.659192,4.164978,3.9801195,3.9197574,3.8367596,3.7613072,3.7273536,3.783943,4.006528,4.4139714,5.3382645,7.066127,9.386291,11.59705,13.607859,15.324403,15.414946,13.517315,10.246449,8.360137,6.9227667,6.221059,6.1342883,6.126743,6.228604,6.571913,6.937857,7.194396,7.303802,7.284939,7.0472636,6.6850915,6.432326,6.670001,12.37421,12.257258,12.291212,12.411936,12.46098,12.185578,12.064855,11.487643,11.106608,11.144334,11.3820095,10.895341,10.0465,9.431562,9.092027,8.503497,7.624475,6.7039547,5.904158,5.3986263,5.3684454,5.2854476,5.617439,5.7192993,5.492942,5.3684454,5.243949,4.678055,4.146115,3.8178966,3.519859,3.2784111,3.0671442,2.9652832,2.9766011,3.0181,3.2746384,3.3689542,3.3123648,3.2255943,3.361409,3.108643,2.8521044,2.8936033,3.3274553,4.0593443,4.8100967,5.6287565,6.458734,7.488661,9.178797,8.27714,6.802043,4.9232755,3.127506,2.1805773,1.7919968,1.8297231,2.1843498,2.7691069,3.5274043,3.059599,2.9652832,3.5575855,4.817642,6.398372,6.696409,7.069899,7.5112963,7.5527954,6.2889657,4.930821,4.4403796,4.557331,4.666737,3.7990334,3.7273536,3.6707642,3.3312278,2.6332922,1.7014539,0.98842776,1.2147852,1.2826926,1.0110635,1.1129243,0.98842776,0.77716076,0.66775465,0.6828451,0.68661773,0.543258,0.76584285,0.83752275,0.66775465,0.5885295,0.543258,0.4640329,0.362172,0.29049212,0.33953625,0.32067314,0.36971724,0.41121614,0.3961256,0.32067314,0.58098423,1.5354583,2.384299,2.8332415,3.0897799,5.160951,6.6624556,7.3075747,7.1038527,6.368191,4.8553686,3.99521,3.6028569,3.4745877,3.3953626,3.5877664,4.323428,5.4740787,6.888813,8.394091,7.2698483,7.911195,8.416726,8.062099,7.322665,7.281166,6.1418333,4.1498876,2.0787163,1.267602,2.0560806,2.2673476,1.9466745,1.4373702,1.3732355,0.3734899,0.08299775,0.049044125,0.060362,0.124496624,0.14713238,0.15845025,0.2678564,0.633801,1.448688,5.6400743,6.617184,6.1229706,5.451443,5.409944,7.152897,8.182823,5.802297,1.418507,0.55080324,0.6752999,0.68661773,0.55457586,0.32821837,0.15845025,0.09808825,0.056589376,0.026408374,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20372175,0.49421388,0.7054809,0.62625575,0.1659955,0.030181,0.06413463,0.124496624,0.116951376,0.0754525,0.0452715,0.041498873,0.071679875,0.12826926,0.29803738,0.2678564,0.43385187,0.7432071,0.7092535,0.88279426,1.026154,0.90920264,0.814887,1.539231,2.2598023,1.7391801,1.0374719,0.6828451,0.6790725,0.68661773,0.6375736,0.4376245,0.17354076,0.1056335,0.22258487,0.35462674,0.43385187,0.42630664,0.3772625,0.5055317,0.36594462,0.21881226,0.16976812,0.16976812,0.23013012,0.33576363,0.46026024,0.5319401,0.45648763,0.44894236,0.271629,0.11317875,0.090543,0.26031113,0.5998474,0.784706,0.8186596,0.7809334,0.83752275,1.0601076,1.3166461,1.4562333,1.3958713,1.1393328,1.056335,0.8601585,0.7205714,0.70170826,0.754525,1.0072908,1.2826926,1.4562333,1.4298248,1.1053791,0.9205205,0.694163,0.5017591,0.32444575,0.06413463,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.00754525,0.011317875,0.05281675,0.116951376,0.15845025,0.071679875,0.030181,0.0452715,0.1358145,0.31312788,0.21503963,0.10186087,0.19994913,0.543258,0.9620194,0.38858038,0.28294688,0.47535074,0.88279426,1.4977322,1.5241405,0.8337501,0.35462674,0.32067314,0.25276586,0.13204187,0.116951376,0.18863125,0.271629,0.2263575,0.060362,0.011317875,0.02263575,0.041498873,0.02263575,0.011317875,0.003772625,0.003772625,0.00754525,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.041498873,0.056589376,0.06413463,0.0754525,0.1056335,0.03772625,0.018863125,0.018863125,0.030181,0.03772625,0.026408374,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.049044125,0.13204187,0.20749438,0.29426476,0.39989826,0.362172,0.19240387,0.06413463,0.011317875,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.033953626,0.049044125,0.030181,0.030181,0.030181,0.056589376,0.09808825,0.120724,0.11317875,0.1358145,0.16976812,0.18485862,0.13204187,0.13958712,0.27540162,0.5998474,0.9808825,1.1053791,1.0751982,1.1016065,1.1619685,1.267602,1.4750963,2.6068838,3.361409,3.4368613,2.9841464,2.584248,2.7011995,3.0935526,3.3953626,3.4217708,3.150142,2.9011486,2.9313297,3.0105548,2.969056,2.71629,2.746471,2.8709676,3.029418,3.029418,2.5314314,1.5656394,1.0035182,0.66775465,0.43385187,0.21503963,0.11317875,0.056589376,0.026408374,0.011317875,0.0,0.0150905,0.030181,0.041498873,0.056589376,0.08299775,0.06413463,0.05281675,0.05281675,0.060362,0.060362,0.030181,0.03772625,0.06790725,0.11317875,0.1961765,0.1961765,0.3470815,0.482896,0.543258,0.5357128,0.8186596,1.1053791,1.2826926,1.3430545,1.3845534,1.3807807,1.3091009,1.2034674,1.1242423,1.1393328,1.0072908,1.0601076,1.3015556,1.6675003,2.0183544,2.1956677,2.384299,2.5427492,2.6521554,2.7087448,2.8332415,3.4142256,4.6516466,5.994701,6.145606,6.379509,7.537705,8.492179,8.990166,9.64283,11.317875,12.189351,12.925014,13.174006,11.555551,9.590013,8.20546,7.537705,7.6584287,8.567632,10.148361,10.329447,8.7600355,6.221059,4.6252384,6.2399216,9.623966,12.985375,14.037937,10.005001,5.2326307,3.229367,2.9992368,3.4179983,3.199186,3.180323,3.682082,4.6327834,5.832478,6.9869013,7.0812173,7.360391,8.179051,9.21275,9.435335,9.190115,10.238904,11.140562,11.227332,10.627484,11.034928,12.261031,12.838243,12.242168,10.853842,10.001229,8.620448,7.0812173,5.9532022,5.994701,6.990674,8.6732645,10.604849,12.140307,12.4307995,9.529651,7.364164,5.836251,4.7610526,3.8669407,3.4594972,3.1048703,2.8936033,2.5691576,1.5165952,0.7432071,0.30935526,0.116951376,0.06790725,0.06413463,0.049044125,0.02263575,0.018863125,0.033953626,0.0452715,0.071679875,0.11317875,0.17731337,0.271629,0.38858038,0.5017591,0.6187105,0.76207024,0.95824677,1.2525115,1.7052265,2.2862108,2.9954643,3.6330378,3.8141239,3.5160866,3.4632697,3.5953116,3.783943,3.8556228,3.5387223,3.3274553,3.229367,3.2670932,3.482133,3.9273026,4.376245,4.402653,3.9763467,3.4557245,4.8327327,7.183078,9.982366,13.083464,16.716501,20.787165,23.258234,22.797974,19.90437,16.927769,15.181043,14.045483,13.890805,14.532151,15.207452,15.516807,15.445127,14.826416,13.502225,11.344283,9.759781,8.643084,7.9753294,7.673519,7.564113,7.586749,7.726336,7.877241,7.9753294,8.009283,7.964011,7.835742,7.6131573,7.333983,7.069899,7.062354,7.326438,7.805561,8.367682,8.82417,8.518587,7.914967,7.224577,6.56814,5.994701,5.481624,5.089271,4.7950063,4.5120597,4.08198,3.7990334,3.7462165,3.8405323,3.953711,3.9273026,4.1574326,4.3347464,4.696918,5.138315,5.2137675,4.949684,4.870459,4.919503,5.032682,5.1232247,5.2665844,5.160951,4.9534564,4.798779,4.870459,4.402653,3.99521,3.7386713,3.6971724,3.9008942,4.45547,5.3759904,6.651138,8.182823,9.789962,11.593277,13.845533,15.467763,15.543215,13.328684,10.925522,9.035437,7.6508837,6.85486,6.7869525,6.72659,6.809588,6.9944468,7.2057137,7.322665,7.3490734,6.990674,6.579458,6.247467,5.938112,6.7379084,6.7454534,6.8058157,6.700182,6.462507,6.387054,6.349328,6.307829,6.5530496,6.9944468,7.149124,7.145352,7.2698483,7.5905213,7.888559,7.6622014,6.7831798,5.753253,4.98741,4.689373,4.8365054,5.330719,5.8588867,6.119198,6.0324273,5.7570257,5.534441,4.5535583,3.651901,3.1199608,2.727608,2.1466236,1.8599042,1.931584,2.2598023,2.5804756,3.0105548,3.2029586,3.2369123,3.1916409,3.1237335,2.9086938,2.5880208,2.5993385,3.0746894,3.8405323,4.949684,6.2323766,7.5037513,8.718536,9.948412,8.258276,6.2097406,4.7836885,4.074435,3.2784111,2.463524,2.3616633,2.987919,4.22534,5.8098426,3.9499383,2.957738,3.1312788,4.4931965,6.752999,7.7716074,8.09228,8.744945,9.49947,8.8769865,7.4207535,6.0512905,5.1458607,4.696918,4.3121104,4.425289,4.398881,4.0216184,3.2520027,2.2107582,1.3204187,1.3392819,1.4034165,1.2147852,1.0299267,0.8639311,0.8111144,0.90920264,1.0902886,1.1883769,0.7394345,1.0072908,1.1506506,0.965792,0.8941121,0.7884786,0.6073926,0.452715,0.40367088,0.5017591,0.46026024,0.55080324,0.6413463,0.7167987,0.875249,1.4449154,2.625747,3.7235808,4.5761943,5.5797124,7.54525,8.741172,9.06939,8.843033,8.7751255,8.016829,5.885295,4.323428,3.8971217,3.802806,4.0103,4.429062,5.093044,6.092789,7.5565677,7.2623034,8.356364,9.250477,9.148616,8.058327,6.964266,5.221313,3.3727267,1.8674494,1.0902886,1.9164935,2.0070364,1.4901869,0.8526133,0.9205205,0.27540162,0.19994913,0.33576363,0.43007925,0.32821837,0.23767537,0.18863125,0.2565385,0.49044126,0.9318384,5.119452,5.247721,3.8292143,2.6483827,2.7389257,4.168751,3.7386713,2.2673476,0.72811663,0.24522063,0.18485862,0.15467763,0.116951376,0.06413463,0.018863125,0.0150905,0.02263575,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.26031113,0.392353,0.27917424,0.05281675,0.018863125,0.033953626,0.094315626,0.15845025,0.1358145,0.07922512,0.0452715,0.049044125,0.08677038,0.15845025,0.271629,0.3772625,0.5470306,0.7432071,0.80356914,1.1016065,1.3920987,1.4600059,1.4977322,2.1277604,1.9089483,1.4222796,1.0638802,0.95824677,0.965792,0.80734175,0.6111652,0.482896,0.422534,0.32821837,0.47157812,0.5583485,0.55457586,0.482896,0.4376245,0.543258,0.35462674,0.15845025,0.06413463,0.02263575,0.018863125,0.056589376,0.11317875,0.14713238,0.120724,0.15467763,0.09808825,0.041498873,0.0754525,0.271629,0.5394854,0.5998474,0.6526641,0.7507524,0.7922512,0.9016574,0.9808825,0.98465514,0.935611,0.9016574,1.116697,0.94315624,0.7997965,0.875249,1.1091517,1.327964,1.4260522,1.4864142,1.4449154,1.0940613,0.8111144,0.56212115,0.36594462,0.20749438,0.06413463,0.033953626,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.07922512,0.16976812,0.21881226,0.14713238,0.060362,0.030181,0.06413463,0.1358145,0.20749438,0.1961765,0.18485862,0.211267,0.27540162,0.35839936,0.26031113,0.17354076,0.19994913,0.32821837,0.44139713,0.21881226,0.23390275,0.4376245,0.8299775,1.4750963,1.4826416,0.63002837,0.0754525,0.11317875,0.14335975,0.10940613,0.06413463,0.03772625,0.033953626,0.02263575,0.003772625,0.003772625,0.0150905,0.026408374,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.030181,0.124496624,0.27540162,0.19240387,0.08299775,0.049044125,0.060362,0.05281675,0.03772625,0.033953626,0.05281675,0.07922512,0.12826926,0.116951376,0.08299775,0.0452715,0.02263575,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.033953626,0.10940613,0.2263575,0.35839936,0.5281675,0.47912338,0.21881226,0.06413463,0.033953626,0.018863125,0.00754525,0.0,0.0,0.00754525,0.0150905,0.02263575,0.030181,0.02263575,0.018863125,0.018863125,0.033953626,0.06790725,0.1056335,0.1659955,0.18863125,0.15467763,0.090543,0.08299775,0.090543,0.18485862,0.62248313,1.267602,1.5920477,1.7165444,1.8334957,1.8448136,1.8599042,2.2107582,2.9011486,3.029418,2.7804246,2.425798,2.335255,3.0331905,3.6028569,3.953711,4.06689,3.9688015,3.9273026,3.9461658,3.8669407,3.6443558,3.338773,3.380272,3.2218218,3.0369632,2.7728794,2.1353056,1.2147852,0.663982,0.35462674,0.181086,0.07922512,0.041498873,0.030181,0.02263575,0.0150905,0.018863125,0.033953626,0.041498873,0.03772625,0.030181,0.033953626,0.026408374,0.033953626,0.049044125,0.060362,0.056589376,0.124496624,0.3961256,0.55457586,0.513077,0.43385187,0.49421388,0.5772116,0.6111652,0.6073926,0.663982,0.965792,1.2261031,1.3845534,1.4562333,1.5241405,1.4562333,1.2751472,1.0978339,1.0072908,1.0223814,0.83752275,0.845068,1.0525624,1.3807807,1.6524098,1.8334957,1.9768555,2.123988,2.3126192,2.584248,3.108643,4.123479,5.553304,6.8963585,7.24344,7.164215,8.235641,9.337247,9.914458,10.005001,10.321902,11.080199,11.857361,12.181807,11.52537,10.831206,10.208723,9.737145,9.514561,9.661693,10.250222,9.993684,9.1825695,7.8734684,5.873977,4.640329,5.3684454,7.533932,9.235386,7.194396,3.8669407,2.1088974,1.7429527,2.1541688,2.293756,2.5012503,2.7879698,3.482133,4.5233774,5.4703064,5.8513412,6.247467,7.164215,8.333729,8.703445,8.763808,10.56335,12.019584,12.045992,10.559577,9.495697,10.465261,11.581959,11.936585,11.6008215,11.638548,10.872705,9.590013,8.360137,8.043237,8.567632,9.7220545,11.502733,13.400364,14.4114275,11.487643,8.394091,6.145606,4.949684,4.191386,3.3953626,2.6597006,2.305074,2.1805773,1.6825907,1.1091517,0.66775465,0.41121614,0.29803738,0.20372175,0.1358145,0.09808825,0.08677038,0.08677038,0.0754525,0.094315626,0.14335975,0.2263575,0.3470815,0.4979865,0.5885295,0.66020936,0.7582976,0.90543,1.1280149,1.539231,2.0636258,2.7351532,3.3463185,3.4670424,3.1727777,3.2935016,3.8556228,4.61392,5.070408,4.779916,4.2027044,3.7688525,3.712263,4.06689,5.7494807,7.394345,7.828197,6.7077274,4.5422406,3.9914372,4.8742313,6.3455553,8.0206,9.986138,12.562841,14.7170105,15.569623,15.060319,13.962485,12.58925,11.551778,11.170743,11.065109,10.182315,10.050273,10.876478,11.6008215,11.574413,10.544487,9.261794,8.209232,7.5716586,7.326438,7.24344,7.0548086,6.9793563,6.9869013,7.0963078,7.3717093,7.4018903,7.533932,7.6697464,7.77538,7.865923,8.024373,8.296002,8.6732645,9.103344,9.457971,9.261794,8.6732645,7.8923316,7.073672,6.3342376,5.753253,5.2779026,4.9119577,4.5950575,4.2027044,3.8858037,3.7688525,3.9914372,4.406426,4.5799665,4.8063245,5.0515447,5.4476705,5.9003854,6.0739264,5.881522,5.783434,5.8664317,6.043745,6.0701537,6.2323766,6.149379,5.9494295,5.7419353,5.6287565,4.7346444,4.006528,3.5953116,3.572676,3.9310753,4.4743333,5.0666356,5.7607985,6.628502,7.7338815,9.2995205,11.551778,13.981348,15.671484,15.267814,13.249459,11.472552,9.865415,8.518587,7.6848373,7.356619,7.0510364,6.8737226,6.851087,6.9152217,6.85486,6.488915,6.1078796,5.764571,5.27413,4.7950063,4.496969,4.4403796,4.2102494,3.874486,3.9574835,3.8254418,3.9989824,4.4630156,4.881777,4.5912848,4.5988297,4.8327327,5.458988,6.277648,6.7152724,5.764571,4.647874,4.0291634,4.044254,4.2630663,4.5799665,4.7648253,4.6629643,4.247976,3.610402,3.7084904,3.2859564,2.727608,2.2484846,1.9127209,2.2447119,2.5993385,2.7992878,2.8219235,2.8181508,3.059599,2.9237845,2.7200627,2.674791,2.9086938,3.187868,2.9615107,2.757789,2.8596497,3.3010468,4.1800685,5.666483,7.073672,7.779153,7.1981683,6.1229706,4.244203,3.4934506,3.942393,3.8103511,3.2218218,3.2746384,4.074435,5.4778514,7.069899,4.3309736,3.1124156,2.9803739,3.7537618,5.485397,6.749226,6.888813,7.4999785,8.835487,9.812597,9.461743,7.8244243,5.983383,4.659192,4.236658,4.0782075,3.8707132,3.361409,2.6219745,2.0258996,1.6939086,1.5052774,1.5618668,1.6373192,1.1996948,1.1581959,1.2411937,1.448688,1.6184561,1.4600059,1.0374719,1.1581959,1.2298758,1.1242423,1.1431054,0.95447415,0.7205714,0.5281675,0.44894236,0.5394854,0.44516975,0.52439487,0.6752999,0.94315624,1.5241405,2.6031113,3.4896781,4.3913355,5.9192486,9.099571,8.59404,7.8244243,7.254758,7.326438,8.465771,8.858124,6.609639,4.7346444,4.1008434,3.4179983,3.5236318,3.6707642,3.9310753,4.4516973,5.4665337,7.020855,7.224577,7.352846,7.432071,6.255012,4.1536603,2.7804246,2.071171,1.690136,1.0186088,0.8224323,0.5055317,0.24522063,0.13204187,0.18485862,0.46026024,1.0751982,1.418507,1.2261031,0.59230214,0.2867195,0.12826926,0.094315626,0.1659955,0.34330887,0.23390275,0.14713238,0.13958712,0.23390275,0.4376245,0.48666862,0.2867195,0.23767537,0.32821837,0.120724,0.06413463,0.026408374,0.00754525,0.0,0.003772625,0.011317875,0.041498873,0.0452715,0.018863125,0.0,0.0,0.0,0.0,0.0,0.00754525,0.033953626,0.211267,0.2678564,0.150905,0.018863125,0.030181,0.060362,0.08299775,0.09808825,0.090543,0.09808825,0.08677038,0.0754525,0.0754525,0.090543,0.16222288,0.41121614,0.52062225,0.5394854,0.87147635,1.4411428,1.9466745,2.263575,2.384299,2.4371157,1.2940104,0.7884786,0.73188925,0.9205205,1.1393328,1.0789708,0.77338815,0.6828451,0.8563859,0.90543,0.91297525,0.8526133,0.76207024,0.6790725,0.6451189,0.5696664,0.3055826,0.094315626,0.02263575,0.011317875,0.003772625,0.0,0.0,0.00754525,0.03772625,0.011317875,0.003772625,0.02263575,0.06413463,0.120724,0.21881226,0.33953625,0.3734899,0.33953625,0.3772625,0.52062225,0.58475685,0.5998474,0.62248313,0.72811663,1.026154,0.91297525,0.8903395,1.1355602,1.50905,1.5015048,1.2336484,1.0827434,1.1129243,1.0450171,0.6752999,0.41498876,0.23767537,0.11317875,0.0,0.03772625,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.1659955,0.35085413,0.482896,0.4074435,0.24522063,0.14335975,0.17731337,0.30181,0.32821837,0.3734899,0.4074435,0.46026024,0.49421388,0.392353,0.23013012,0.24899325,0.32821837,0.38103512,0.35085413,0.2678564,0.16222288,0.21503963,0.5357128,1.1317875,0.94315624,0.3734899,0.03772625,0.07922512,0.15845025,0.120724,0.060362,0.030181,0.03772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.06413463,0.20372175,0.47912338,0.29426476,0.094315626,0.060362,0.094315626,0.09808825,0.0754525,0.1056335,0.19994913,0.32444575,0.42630664,0.36971724,0.23390275,0.1056335,0.06790725,0.030181,0.018863125,0.00754525,0.0,0.0,0.003772625,0.0,0.0,0.011317875,0.049044125,0.21503963,0.4678055,0.5394854,0.39989826,0.2678564,0.120724,0.06413463,0.060362,0.06790725,0.06790725,0.041498873,0.0150905,0.00754525,0.0150905,0.02263575,0.0150905,0.00754525,0.0150905,0.03772625,0.094315626,0.23767537,0.32444575,0.28294688,0.16222288,0.120724,0.1056335,0.16976812,0.5885295,1.237421,1.6109109,2.0636258,2.516341,2.7841973,2.8785129,2.9841464,2.7540162,2.4107075,2.3277097,2.505023,2.5540671,2.987919,3.187868,3.4594972,3.8593953,4.2064767,4.9685473,5.1647234,4.889322,4.3649273,3.92353,4.2291126,3.7386713,2.927557,2.0862615,1.3543724,0.9016574,0.5885295,0.362172,0.19994913,0.13204187,0.094315626,0.0754525,0.06413463,0.05281675,0.056589376,0.049044125,0.026408374,0.011317875,0.011317875,0.02263575,0.018863125,0.0150905,0.0150905,0.011317875,0.003772625,0.211267,0.80734175,1.2034674,1.2110126,1.056335,1.0978339,0.94692886,0.7582976,0.6526641,0.7432071,0.9808825,1.1544232,1.2826926,1.388326,1.50905,1.418507,1.2525115,1.146878,1.1544232,1.2147852,1.1204696,1.177059,1.3355093,1.4826416,1.4449154,1.4524606,1.5279131,1.6712729,1.9127209,2.293756,3.1199608,4.3611546,5.66271,6.7077274,7.24344,7.009537,7.3792543,8.22055,9.242931,10.012547,9.884277,9.733373,9.88805,10.295494,10.502988,10.79348,10.967021,10.627484,9.65792,8.213005,7.9791017,7.986647,8.412953,8.733627,7.7112455,5.696664,4.749735,5.8588867,7.5829763,6.047518,4.689373,3.4632697,2.7917426,2.6483827,2.5578396,2.6483827,2.4559789,2.6031113,3.229367,3.983892,3.983892,4.5460134,5.832478,7.3075747,7.7338815,7.232122,9.261794,11.472552,12.351574,11.231105,9.87296,11.027383,12.777881,14.056801,14.618922,14.7321005,14.339747,13.562587,12.54775,11.476325,10.9594755,10.797253,11.717773,13.50977,15.01882,13.50977,10.352083,7.7640624,6.4549613,5.6023483,4.2819295,3.0860074,2.3503454,2.123988,2.1466236,1.7240896,1.2902378,0.9507015,0.69793564,0.392353,0.26031113,0.21881226,0.21881226,0.22258487,0.19994913,0.211267,0.24899325,0.33953625,0.4678055,0.5772116,0.6149379,0.65643674,0.7092535,0.7696155,0.8337501,0.97333723,1.177059,1.4260522,1.6788181,1.8448136,2.003264,2.4786146,3.591539,5.0854983,6.126743,5.994701,5.221313,4.4705606,4.1197066,4.293247,6.983129,9.97482,11.514051,10.759526,7.7678347,5.20245,4.0517993,3.783943,3.8405323,3.6594462,3.6783094,4.5422406,6.0701537,7.91874,9.574923,9.752235,9.786189,9.454198,8.511042,6.7077274,6.6549106,7.122716,7.533932,7.7678347,8.167733,8.114917,7.779153,7.541477,7.492433,7.4509344,7.2057137,6.960493,6.752999,6.7039547,7.001992,6.900131,7.118943,7.4773426,7.865923,8.22055,8.586494,8.89585,9.288202,9.733373,10.072908,9.87296,9.34102,8.518587,7.5263867,6.560595,5.956975,5.560849,5.3759904,5.2552667,4.9119577,4.557331,4.4705606,4.727099,5.172269,5.409944,5.5382137,5.798525,6.168242,6.598321,7.009537,7.2623034,7.250985,7.4471617,7.77538,7.6584287,7.432071,6.964266,6.571913,6.3153744,6.013564,4.768598,3.8782585,3.4255435,3.4368613,3.8820312,4.1989317,4.236658,4.4743333,5.0439997,5.7494807,7.0548086,9.073163,11.581959,13.970031,15.203679,14.377474,13.12119,11.695138,10.137043,8.235641,7.7301087,7.1604424,6.7114997,6.4511886,6.3229194,6.205968,5.9418845,5.553304,5.138315,4.859141,4.3800178,4.063117,3.4783602,2.8256962,2.4559789,2.8822856,2.9464202,3.3350005,3.8367596,4.187614,4.0895257,4.187614,4.678055,5.198677,5.6287565,6.119198,5.119452,4.7120085,4.6629643,4.6290107,4.164978,3.591539,3.31991,3.308592,3.3764994,3.218049,3.610402,4.0103,3.8707132,3.3538637,3.3425457,4.745962,6.1041074,6.7077274,6.40969,5.613666,4.772371,3.4557245,2.5880208,2.5540671,3.187868,3.712263,3.8895764,3.7499893,3.5085413,3.5689032,3.9612563,5.515578,6.307829,5.794752,4.8063245,3.8178966,2.444661,1.6222287,1.6109109,2.0145817,2.0145817,2.8936033,4.2592936,5.5457587,5.9984736,4.8855495,4.5422406,4.142342,3.92353,5.2175403,5.3759904,5.0138187,4.9647746,5.7607985,7.6131573,8.360137,7.4282985,5.80607,4.236658,3.2331395,3.429316,4.3121104,4.4818783,3.6254926,2.5012503,2.2598023,2.323937,2.4295704,2.372981,2.0296721,1.7731338,1.5241405,1.5731846,1.7391801,1.3732355,1.177059,1.2562841,1.2562841,1.1204696,1.0827434,0.6187105,0.45648763,0.40367088,0.35839936,0.32067314,0.43007925,0.6790725,0.98842776,1.3317367,1.7089992,3.2331395,4.2102494,5.198677,6.85486,9.918231,5.96452,4.3611546,3.2670932,2.1051247,1.5580941,2.142851,3.1237335,3.8178966,3.6481283,2.1353056,2.7238352,2.8785129,3.1237335,3.904667,5.5985756,7.3717093,6.1908774,5.0439997,4.715781,3.7990334,3.2142766,2.674791,1.9655377,1.2864652,1.2525115,1.2864652,0.91297525,0.5583485,0.43007925,0.5017591,1.5279131,3.7160356,4.014073,2.1315331,0.52062225,0.116951376,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.120724,0.21881226,0.21503963,0.1056335,0.030181,0.041498873,0.06413463,0.094315626,0.13958712,0.21503963,0.19994913,0.16222288,0.124496624,0.116951376,0.150905,0.1659955,0.44139713,0.65643674,0.79602385,1.1732863,1.5430037,2.0636258,2.757789,3.2784111,2.897376,2.1654868,1.4071891,0.8563859,0.6488915,0.80734175,1.0525624,0.8941121,0.8224323,1.0902886,1.7240896,1.2713746,0.8865669,0.694163,0.633801,0.42630664,0.1358145,0.041498873,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.26408374,0.5696664,0.87147635,0.94692886,1.177059,0.91674787,0.84884065,1.1204696,1.327964,1.1431054,0.9242931,0.814887,0.83752275,0.8865669,0.55457586,0.29803738,0.14713238,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.0754525,0.211267,0.56589377,0.6375736,0.45648763,0.56589377,0.87902164,0.67152727,0.40367088,0.3734899,0.47535074,0.573439,0.48666862,0.21881226,0.33576363,0.36594462,0.29049212,0.5357128,0.46026024,0.23013012,0.1659955,0.47157812,1.267602,0.362172,0.056589376,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.071679875,0.0452715,0.0452715,0.06413463,0.0754525,0.071679875,0.0452715,0.071679875,0.1056335,0.2678564,0.59230214,1.0072908,1.0299267,0.73566186,0.35085413,0.07922512,0.090543,0.056589376,0.026408374,0.00754525,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.09808825,0.22258487,0.4074435,0.62248313,0.7922512,0.3055826,0.15467763,0.22258487,0.3470815,0.33576363,0.19994913,0.0754525,0.0150905,0.02263575,0.0452715,0.056589376,0.041498873,0.018863125,0.00754525,0.0452715,0.1659955,0.3169005,0.38480774,0.34330887,0.24522063,0.16976812,0.23390275,0.46026024,0.7922512,1.0978339,2.293756,2.7389257,2.9841464,3.1199608,2.776652,2.203213,2.425798,3.2444575,3.9688015,3.4330888,3.7386713,3.7047176,3.350091,2.9351022,2.9615107,4.67051,4.5761943,3.8405323,3.3010468,3.4481792,3.5953116,3.3764994,2.8030603,1.9542197,0.97710985,0.9016574,0.663982,0.42630664,0.27917424,0.23013012,0.19240387,0.17354076,0.15467763,0.12826926,0.090543,0.056589376,0.026408374,0.026408374,0.049044125,0.060362,0.03772625,0.02263575,0.00754525,0.003772625,0.0150905,0.0754525,0.35839936,1.0148361,1.9089483,2.595566,1.9730829,1.3845534,0.9393836,0.7054809,0.7167987,0.8865669,0.9507015,0.875249,0.7394345,0.70170826,0.7997965,0.935611,1.0978339,1.3128735,1.6184561,1.5430037,1.6637276,1.7165444,1.6524098,1.6184561,1.6524098,1.6524098,1.7655885,1.9881734,2.1956677,2.8558772,3.7348988,4.7610526,5.7570257,6.439871,6.2814207,6.643593,7.115171,7.9489207,10.084227,11.295239,11.257513,11.091517,11.200924,11.261286,9.869187,9.156161,8.7600355,8.345046,7.6131573,7.6622014,6.4021444,6.047518,6.760544,6.6360474,6.1229706,4.6327834,3.6368105,3.874486,5.342037,6.205968,5.6287565,4.395108,3.059599,1.9240388,2.082489,2.1768045,2.305074,2.3616633,2.0447628,2.033445,2.7540162,4.0404816,5.4740787,6.379509,6.0739264,7.032173,8.68081,10.182315,10.438853,11.8045435,14.369928,17.056038,18.949896,19.31584,18.085964,16.731592,15.384765,14.015302,12.449662,10.997202,10.570895,11.566868,13.649357,15.762027,14.222796,11.981857,9.918231,8.397863,7.2623034,5.541986,4.4441524,3.7763977,3.3538637,2.9766011,2.584248,2.1843498,1.7165444,1.1619685,0.56589377,0.44139713,0.36594462,0.36594462,0.43007925,0.5017591,0.51684964,0.47157812,0.46026024,0.5017591,0.56589377,0.5017591,0.47912338,0.52062225,0.62625575,0.7469798,0.87147635,1.146878,1.2261031,1.1016065,1.1129243,1.4675511,2.123988,3.7047176,5.836251,7.141579,6.809588,5.492942,4.3385186,4.014073,4.6856003,5.9305663,8.273367,10.850069,12.344029,11.000975,7.7037,5.5080323,4.8365054,5.2099953,5.2326307,4.255521,3.7198083,3.9159849,4.7874613,5.934339,7.1679873,8.235641,8.639311,8.160188,6.8661776,5.6815734,5.2967653,5.4665337,5.847569,5.983383,6.6058664,7.0887623,7.624475,8.084735,8.009283,8.401636,8.6732645,8.518587,7.9791017,7.432071,7.3453007,7.745199,8.111144,8.22055,8.14887,8.503497,8.892077,9.424017,10.023865,10.453944,10.514306,10.216269,9.6051035,8.744945,7.7225633,6.8435416,6.3945994,6.4964604,6.900131,6.971811,6.5228686,6.1720147,6.043745,6.0814714,6.058836,5.9117036,6.0776987,6.5341864,7.254758,8.194141,9.110889,8.869441,8.710991,8.843033,8.4544525,7.3075747,6.7341356,6.405917,6.304056,6.7454534,4.961002,4.0480266,3.7198083,3.7348988,3.904667,3.6368105,3.5538127,3.6330378,3.9197574,4.515832,5.775889,7.654656,9.737145,11.627231,12.970284,13.422999,12.645839,11.121698,9.288202,7.5527954,7.273621,6.9567204,6.5945487,6.2135134,5.8588867,5.7117543,5.485397,5.20245,4.919503,4.7006907,6.5643673,6.3342376,5.4967146,4.13857,2.7917426,2.4182527,3.1539145,3.9348478,4.032936,3.4217708,2.746471,3.85185,4.4101987,4.919503,5.643847,6.620957,4.9345937,4.4516973,4.9987283,5.775889,5.349582,4.5233774,4.3196554,4.678055,4.8855495,3.5839937,4.123479,4.063117,3.5953116,3.0445085,2.8785129,3.5990841,4.640329,5.7796617,6.507778,6.006019,5.828706,5.270357,4.515832,3.9348478,4.08198,3.7952607,3.8141239,3.783943,3.6858547,3.8141239,4.187614,5.05909,6.8774953,8.382772,6.6134114,5.409944,4.164978,3.0860074,2.323937,1.9655377,2.2296214,3.0143273,3.5651307,3.640583,3.5047686,3.5462675,4.08198,4.6252384,5.010046,5.3759904,5.534441,5.0025005,4.3347464,4.104616,4.9157305,6.7152724,7.0963078,5.96452,4.0970707,3.1237335,2.957738,3.361409,3.7952607,3.802806,2.9916916,2.5804756,2.2975287,2.1881225,2.1579416,1.991946,1.8146327,1.8938577,2.0900342,2.1768045,1.8485862,1.3996439,1.1732863,1.1053791,1.1317875,1.1921495,1.0336993,1.0336993,0.9393836,0.69039035,0.41876137,0.46026024,0.7205714,1.0412445,1.448688,2.161714,2.757789,4.587512,6.4738245,7.7678347,8.329956,6.6322746,3.7914882,1.7278622,1.0299267,0.95824677,1.2298758,1.6712729,2.191895,2.5502944,2.3428001,1.8749946,1.9730829,2.3465726,2.8785129,3.5990841,4.244203,4.1498876,4.1762958,4.3422914,3.7990334,3.2821836,3.0671442,2.7879698,2.1843498,1.0940613,0.543258,0.35839936,0.26408374,0.16222288,0.1358145,0.38103512,0.845068,0.875249,0.4376245,0.1056335,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.090543,0.094315626,0.071679875,0.06413463,0.07922512,0.10940613,0.150905,0.1961765,0.24899325,0.31312788,0.4376245,0.44516975,0.3772625,0.29803738,0.2867195,0.38858038,0.33576363,0.4074435,0.7997965,1.6373192,1.9164935,1.780679,1.5920477,1.569412,1.7882242,2.8332415,2.5616124,1.7957695,1.1355602,0.94315624,1.0978339,0.814887,0.7884786,1.0676528,1.0789708,0.84884065,0.8186596,0.86770374,0.79602385,0.3055826,0.090543,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.018863125,0.08677038,0.07922512,0.033953626,0.0,0.0,0.0,0.0,0.071679875,0.14713238,0.14713238,0.0,0.0150905,0.05281675,0.27917424,0.62248313,0.77338815,1.1921495,1.2411937,1.0450171,0.7582976,0.5470306,0.68661773,0.77338815,0.7130261,0.55457586,0.5055317,0.34330887,0.19994913,0.08677038,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.00754525,0.00754525,0.03772625,0.43007925,0.47912338,0.35839936,0.21503963,0.19994913,0.26031113,0.26031113,0.26031113,0.29426476,0.34330887,0.3470815,0.6111652,0.965792,1.0714256,0.4376245,0.2867195,0.47912338,0.68661773,0.7809334,0.7922512,0.5319401,0.20372175,0.060362,0.28294688,0.9997456,0.4640329,0.13204187,0.003772625,0.0150905,0.02263575,0.003772625,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.041498873,0.0452715,0.071679875,0.09808825,0.10186087,0.090543,0.07922512,0.08299775,0.06790725,0.06790725,0.13204187,0.27540162,0.49421388,0.5885295,0.3734899,0.16222288,0.0754525,0.06790725,0.049044125,0.041498873,0.030181,0.018863125,0.03772625,0.07922512,0.049044125,0.0150905,0.0,0.0,0.06790725,0.26031113,0.6187105,0.98465514,0.98842776,0.68661773,0.5017591,0.45648763,0.513077,0.58098423,0.24899325,0.1056335,0.05281675,0.041498873,0.056589376,0.060362,0.041498873,0.026408374,0.026408374,0.033953626,0.06790725,0.150905,0.28294688,0.422534,0.5017591,0.33953625,0.513077,0.7092535,0.8299775,0.98842776,1.6486372,2.1881225,2.6068838,3.0746894,3.92353,3.5462675,3.7160356,4.22534,4.776143,4.9723196,4.817642,4.0480266,2.9992368,2.655928,4.644101,4.82896,4.2592936,3.742444,3.5689032,3.5085413,3.1576872,2.3805263,1.6939086,1.2638294,0.8903395,0.83752275,0.86770374,0.70170826,0.38858038,0.29049212,0.25276586,0.241448,0.24522063,0.241448,0.21503963,0.12826926,0.094315626,0.090543,0.08677038,0.060362,0.03772625,0.02263575,0.0150905,0.011317875,0.003772625,0.06413463,0.18485862,0.4979865,0.9695646,1.3996439,1.418507,1.267602,1.0072908,0.784706,0.8262049,0.9393836,0.9922004,0.9393836,0.77338815,0.543258,0.4074435,0.44516975,0.6187105,0.9205205,1.3732355,1.7580433,1.9994912,2.071171,2.0673985,2.2296214,2.263575,2.2786655,2.4069347,2.7125173,3.1727777,3.6292653,4.214022,4.82896,5.5004873,6.379509,7.24344,8.016829,8.507269,9.001483,10.269085,14.388792,16.248695,15.901614,13.841762,11.042474,9.416472,9.088254,8.8618965,8.175279,7.1000805,6.5945487,6.439871,6.7831798,7.0849895,6.1116524,6.7831798,6.888813,6.466279,5.994701,6.4134626,6.537959,4.7421894,2.848332,1.7165444,1.2261031,1.6410918,1.7919968,1.8749946,1.9957186,2.1654868,1.6260014,1.6675003,2.3578906,3.4594972,4.4139714,5.572167,7.3075747,8.98262,9.842778,8.98262,10.506761,14.6151495,18.61036,20.643805,19.719511,16.893814,15.422491,13.788944,11.695138,10.095545,9.559832,9.9257765,11.050018,12.619431,14.162435,13.52486,12.494934,11.529142,10.729345,9.839006,8.243186,6.5756855,5.4288073,4.8100967,4.146115,3.6896272,3.0218725,2.142851,1.1846043,0.43007925,0.6488915,0.784706,0.80356914,0.7394345,0.68661773,0.56212115,0.41876137,0.38858038,0.44894236,0.44139713,0.362172,0.38480774,0.4640329,0.573439,0.68661773,0.86770374,1.1016065,1.267602,1.3694628,1.5279131,1.6863633,2.0673985,2.9124665,4.036709,4.8327327,4.376245,3.5462675,3.0143273,3.0897799,3.731126,4.938366,6.8925858,9.156161,10.846297,10.63503,8.405409,6.7379084,6.205968,6.820906,8.016829,8.409182,7.567886,6.628502,6.006019,5.3873086,5.20245,5.674028,6.511551,7.194396,6.9755836,6.25124,5.6853456,5.4703064,5.613666,5.934339,6.047518,6.0701537,6.2625575,6.8058157,7.779153,8.695901,9.276885,9.669238,10.065364,10.676529,9.861642,9.2844305,9.009028,9.099571,9.661693,10.238904,9.7296,9.601331,10.20495,10.7557535,11.11038,11.219787,11.106608,10.812344,10.382264,9.650374,9.114662,8.729855,8.439363,8.167733,7.726336,7.2396674,6.862405,6.620957,6.4134626,6.3153744,6.9152217,7.6508837,8.186596,8.412953,9.193887,9.103344,8.601585,7.9338303,7.122716,6.33801,6.2021956,6.5040054,6.7944975,6.3644185,5.6853456,4.961002,4.3800178,4.104616,4.29702,4.6252384,4.557331,4.3800178,4.432834,5.0779533,6.5228686,8.058327,9.344792,10.220041,10.710483,11.740409,12.162943,11.676274,10.355856,8.650629,7.6395655,6.779407,6.2399216,5.9796104,5.7607985,5.624984,5.485397,5.2779026,4.9723196,4.564876,7.4773426,7.0774446,6.1720147,4.7233267,3.1765501,2.4522061,2.848332,3.3274553,3.519859,3.3953626,3.270866,4.0706625,4.0404816,4.3007927,5.138315,6.0022464,5.2892203,5.142088,5.7004366,6.379509,5.847569,4.8100967,4.8930945,5.3156285,5.304311,4.0895257,4.0404816,3.8895764,3.712263,3.5953116,3.6141748,4.3309736,4.938366,5.323174,5.4967146,5.59103,6.466279,6.7114997,6.417235,5.7683434,5.0439997,3.8178966,3.1199608,2.9237845,2.9916916,2.9049213,3.4557245,3.821669,4.8138695,6.349328,7.466025,7.8961043,6.379509,4.5422406,3.2255943,2.5012503,2.9200118,4.425289,6.5040054,7.665974,5.4665337,4.485651,4.436607,4.7950063,5.311856,6.013564,6.771862,6.330465,5.342037,4.406426,4.0782075,4.659192,4.768598,4.2102494,3.4066803,3.3727267,3.31991,3.2482302,3.240685,3.2255943,2.9841464,2.927557,3.1916409,3.0935526,2.5012503,1.8372684,1.7014539,2.1692593,2.8030603,2.9766011,1.8674494,1.3920987,1.2147852,1.1883769,1.20724,1.2110126,1.1544232,1.1996948,1.1317875,0.965792,0.935611,0.7432071,0.86770374,1.3204187,2.0560806,2.9615107,3.3915899,4.093298,5.3458095,6.677546,6.881268,5.50426,3.1350515,1.358145,0.6790725,0.51684964,0.6451189,0.8337501,1.1280149,1.5316857,2.0108092,2.6483827,2.04099,1.7240896,2.1805773,2.8332415,3.1840954,3.2557755,3.3274553,3.31991,2.8106055,2.3465726,2.11267,1.8636768,1.4298248,0.7054809,0.33953625,0.23013012,0.19240387,0.150905,0.14713238,0.06413463,0.049044125,0.033953626,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.120724,0.56212115,0.43007925,0.20372175,0.1056335,0.090543,0.12826926,0.1961765,0.29803738,0.41121614,0.4640329,0.77716076,0.83752275,0.77338815,0.69039035,0.6488915,0.62625575,0.73566186,0.814887,0.9318384,1.3694628,1.4373702,1.2336484,1.0601076,1.1355602,1.6109109,2.0183544,1.9542197,1.6448646,1.3015556,1.1317875,1.1996948,1.0525624,0.814887,0.63002837,0.63002837,0.7922512,0.87147635,0.79602385,0.5583485,0.211267,0.06790725,0.011317875,0.0,0.0,0.0,0.0,0.0,0.00754525,0.056589376,0.20749438,0.14335975,0.06413463,0.011317875,0.0,0.0,0.0,0.03772625,0.071679875,0.071679875,0.0,0.0,0.13204187,0.29426476,0.4979865,0.8601585,1.0902886,1.146878,1.0148361,0.76584285,0.55080324,0.59607476,0.6526641,0.6413463,0.5772116,0.5394854,0.44139713,0.3055826,0.15845025,0.041498873,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.00754525,0.00754525,0.00754525,0.003772625,0.003772625,0.018863125,0.42630664,0.5093044,0.38103512,0.19994913,0.16222288,0.33953625,0.6149379,0.6073926,0.32821837,0.1659955,0.181086,0.34330887,0.52439487,0.5696664,0.26408374,0.3169005,0.5017591,0.66775465,0.7092535,0.58098423,0.29803738,0.09808825,0.033953626,0.16222288,0.573439,0.36971724,0.14335975,0.02263575,0.018863125,0.041498873,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.090543,0.0754525,0.06413463,0.05281675,0.056589376,0.094315626,0.181086,0.3772625,0.452715,0.35839936,0.19994913,0.090543,0.049044125,0.060362,0.124496624,0.26408374,0.30935526,0.21503963,0.271629,0.4979865,0.6451189,0.1961765,0.049044125,0.02263575,0.018863125,0.03772625,0.071679875,0.056589376,0.030181,0.018863125,0.018863125,0.1659955,0.31312788,0.49044126,0.6451189,0.6451189,0.56212115,0.4376245,0.34330887,0.30181,0.29426476,0.18485862,0.17354076,0.20372175,0.23013012,0.24522063,0.09808825,0.049044125,0.05281675,0.07922512,0.08677038,0.090543,0.13204187,0.20749438,0.29803738,0.392353,0.3470815,0.6149379,0.91674787,1.1280149,1.3091009,1.8184053,2.0258996,2.3956168,3.0143273,3.5990841,3.62172,3.9197574,4.0480266,4.014073,4.266839,3.9461658,3.2859564,2.674791,2.6898816,4.112161,4.659192,4.146115,3.5990841,3.3538637,3.0671442,2.4069347,1.5731846,0.9997456,0.77716076,0.66020936,0.7205714,0.69039035,0.543258,0.3470815,0.29426476,0.25276586,0.2263575,0.241448,0.2678564,0.20749438,0.124496624,0.090543,0.071679875,0.060362,0.05281675,0.094315626,0.07922512,0.0452715,0.041498873,0.10186087,0.19240387,0.23767537,0.3169005,0.5583485,1.1355602,1.5543215,1.539231,1.2261031,0.845068,0.72811663,0.8526133,0.8978847,0.814887,0.633801,0.44894236,0.32821837,0.29049212,0.35085413,0.59607476,1.1657411,1.9164935,2.2447119,2.4182527,2.5804756,2.727608,2.6483827,2.8747404,3.2218218,3.5575855,3.7650797,3.983892,4.402653,4.8553686,5.4665337,6.6662283,8.043237,8.790216,9.129752,9.450426,10.33322,13.588995,16.101564,17.022083,16.03743,13.347548,12.3289385,11.378237,9.869187,7.9791017,6.670001,6.089017,6.4247804,7.3075747,8.013056,7.4735703,8.114917,8.941121,8.348819,7.0774446,8.194141,7.5527954,6.058836,4.236658,2.5502944,1.3920987,1.690136,1.8033148,1.750498,1.7089992,1.9881734,1.8485862,1.7354075,2.0145817,2.8521044,4.2328854,5.379763,6.990674,8.465771,9.2995205,9.088254,10.510533,14.045483,17.384256,19.081938,18.53868,16.124199,14.11339,11.974312,9.854096,8.601585,8.850578,9.34102,10.095545,11.004747,11.830952,11.921495,11.98563,11.947904,11.642321,10.812344,9.1825695,7.6282477,6.470052,5.7306175,5.1081343,4.9685473,4.376245,3.3010468,2.0145817,1.0751982,0.8941121,0.7507524,0.7432071,0.84129536,0.87902164,0.73566186,0.6149379,0.56212115,0.513077,0.27540162,0.271629,0.362172,0.47535074,0.573439,0.663982,0.8224323,0.9808825,1.1016065,1.1921495,1.2864652,1.3505998,1.4298248,1.629774,1.961765,2.354118,2.4597516,2.4408884,2.444661,2.5804756,2.9464202,3.6669915,5.138315,7.424526,9.491924,9.208978,8.333729,7.6810646,7.564113,7.986647,8.639311,9.590013,9.65792,9.175024,8.345046,7.24344,6.187105,5.7872066,5.847569,6.0626082,6.013564,6.1305156,6.0512905,5.824933,5.6061206,5.674028,5.9117036,6.5756855,6.8661776,6.7944975,7.2094865,8.243186,9.242931,10.125726,10.853842,11.442371,11.125471,10.725573,10.529396,10.668983,11.102836,11.52537,11.563096,11.993175,12.528888,11.8045435,11.793225,11.898859,11.978085,11.974312,11.925267,11.378237,10.827434,10.34831,9.952185,9.612649,9.2844305,9.012801,8.416726,7.594294,7.1302614,6.7680893,6.8774953,7.1868505,7.4471617,7.4169807,7.6320205,7.6923823,7.816879,7.956466,7.779153,6.9567204,6.1041074,5.8588867,6.1229706,6.0701537,5.594803,5.2779026,5.0779533,5.036454,5.292993,5.028909,4.7836885,4.6327834,4.7421894,5.3571277,6.700182,8.00551,8.937348,9.397609,9.525878,10.850069,11.879996,12.2119875,11.6875925,10.408672,9.009028,7.7376537,6.7039547,6.017337,5.772116,5.6023483,5.492942,5.3684454,5.1458607,4.7610526,7.8961043,7.91874,6.990674,5.59103,4.255521,3.5689032,3.4368613,3.742444,4.036709,4.0895257,3.9008942,4.063117,3.8593953,4.0782075,4.881777,5.8211603,5.745708,5.9192486,6.436098,6.9454026,6.628502,5.9607477,6.115425,6.092789,5.5268955,4.67051,4.2706113,4.2027044,4.3121104,4.4630156,4.5422406,5.0213637,5.2288585,5.062863,4.776143,5.010046,5.987156,6.5266414,6.428553,5.692891,4.508287,3.5387223,3.097325,3.1916409,3.4972234,3.3764994,3.802806,3.832987,3.8669407,4.496969,6.4964604,7.956466,7.0548086,5.6400743,4.4516973,3.1614597,2.9992368,4.4403796,7.250985,9.759781,8.865668,7.356619,6.0739264,5.6363015,6.1116524,7.0057645,7.7678347,7.364164,6.187105,4.817642,4.0291634,3.5538127,3.1425967,2.8143783,2.7087448,3.1161883,3.2067313,3.1048703,2.8407867,2.595566,2.7087448,3.0746894,3.7160356,3.893349,3.380272,2.4522061,1.9278114,2.3993895,3.138824,3.3236825,2.0636258,1.5920477,1.3392819,1.3317367,1.4449154,1.3958713,1.3091009,1.3241913,1.3392819,1.2902378,1.1431054,0.8865669,1.0450171,1.8146327,3.0445085,4.266839,4.3309736,3.6179473,3.6066296,4.406426,4.7535076,3.651901,2.282438,1.1695137,0.5319401,0.29049212,0.29049212,0.3470815,0.46026024,0.7582976,1.4977322,2.7691069,1.8033148,1.1317875,1.5769572,2.252257,2.71629,2.886058,2.957738,3.006782,3.006782,2.1503963,1.6260014,1.2223305,0.84884065,0.5017591,0.27917424,0.18485862,0.14713238,0.12826926,0.1358145,0.030181,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0452715,0.211267,0.8111144,0.58098423,0.26031113,0.14713238,0.120724,0.16222288,0.2678564,0.45648763,0.6828451,0.8186596,1.0487897,1.1016065,1.0601076,0.97710985,0.8865669,0.79602385,1.0072908,1.0751982,0.9695646,1.0789708,1.0374719,1.0186088,1.177059,1.4562333,1.6109109,1.3392819,1.2600567,1.2487389,1.2411937,1.2298758,1.2600567,1.2147852,0.95824677,0.663982,0.80356914,0.94692886,0.8563859,0.58098423,0.26031113,0.10186087,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.0,0.00754525,0.049044125,0.1659955,0.1056335,0.049044125,0.011317875,0.0,0.0,0.0,0.02263575,0.056589376,0.08299775,0.06790725,0.0150905,0.13204187,0.211267,0.30181,0.694163,0.8526133,0.935611,1.0035182,1.0751982,1.1317875,0.9922004,1.0487897,1.1695137,1.2147852,1.0412445,0.73188925,0.47157812,0.2565385,0.1056335,0.049044125,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.026408374,0.026408374,0.0452715,0.041498873,0.030181,0.026408374,0.056589376,0.27540162,0.33576363,0.271629,0.16222288,0.120724,0.2867195,0.65643674,0.7205714,0.42630664,0.16222288,0.14713238,0.12826926,0.124496624,0.14335975,0.150905,0.2565385,0.35085413,0.3961256,0.3734899,0.26408374,0.32067314,0.20749438,0.08677038,0.0754525,0.20749438,0.17731337,0.08299775,0.018863125,0.011317875,0.026408374,0.018863125,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.041498873,0.06790725,0.1358145,0.120724,0.08677038,0.06413463,0.07922512,0.14335975,0.23013012,0.4376245,0.5281675,0.44516975,0.29803738,0.18863125,0.116951376,0.07922512,0.08677038,0.18485862,0.181086,0.15845025,0.29049212,0.55457586,0.7394345,0.23013012,0.05281675,0.018863125,0.018863125,0.03772625,0.071679875,0.10186087,0.12826926,0.1358145,0.10940613,0.19994913,0.26408374,0.29049212,0.2867195,0.27917424,0.40367088,0.32821837,0.20372175,0.11317875,0.071679875,0.17731337,0.331991,0.5394854,0.694163,0.573439,0.4376245,0.3734899,0.32067314,0.26408374,0.23013012,0.24522063,0.271629,0.271629,0.2678564,0.3169005,0.452715,0.80734175,1.1732863,1.4034165,1.4147344,1.9051756,2.0258996,2.3163917,2.8747404,3.3651814,3.6330378,3.7877154,3.482133,2.8936033,2.704972,2.4295704,2.1805773,2.2220762,2.637065,3.3274553,3.7914882,3.259548,2.7502437,2.595566,2.4371157,1.6184561,0.9507015,0.5772116,0.47157812,0.452715,0.51684964,0.42630664,0.32444575,0.271629,0.25276586,0.21881226,0.18863125,0.19994913,0.21881226,0.14713238,0.08299775,0.056589376,0.049044125,0.049044125,0.0452715,0.116951376,0.116951376,0.08299775,0.071679875,0.13204187,0.23767537,0.24899325,0.23013012,0.35085413,0.87902164,1.4071891,1.5015048,1.2713746,0.9242931,0.7432071,0.7696155,0.73566186,0.6111652,0.44139713,0.33953625,0.30935526,0.2678564,0.271629,0.43007925,0.90920264,1.629774,2.0598533,2.354118,2.5691576,2.6785638,2.584248,2.8294687,3.2067313,3.5764484,3.8405323,3.9273026,4.1272516,4.515832,5.2326307,6.507778,7.8621507,8.756263,9.431562,10.03141,10.589758,12.849561,14.84528,16.309057,16.923996,16.320375,16.116653,14.581196,12.272349,9.854096,8.099826,7.6093845,7.6395655,8.065872,8.360137,7.594294,8.91094,10.287949,9.812597,8.035691,7.967784,7.7640624,6.2663302,4.4139714,2.7841973,1.5882751,1.5656394,1.5958204,1.6033657,1.6675003,1.9994912,2.444661,2.5012503,2.6710186,3.3010468,4.606375,5.956975,7.2472124,8.469543,9.65792,10.906659,12.770335,15.486626,17.629477,18.459454,17.923742,16.203424,13.702174,11.1631975,9.22784,8.4544525,8.89585,8.865668,8.748717,8.854351,9.420244,10.159679,10.819888,11.234878,11.223559,10.597303,9.144843,7.9451485,7.043491,6.417235,5.975838,5.987156,5.4891696,4.45547,3.1010978,1.8976303,1.4034165,1.0336993,0.90543,0.9808825,1.0751982,0.97333723,0.88279426,0.7394345,0.5093044,0.18485862,0.2263575,0.36594462,0.48666862,0.55080324,0.5998474,0.7092535,0.80356914,0.84129536,0.84129536,0.8526133,0.86770374,0.7922512,0.7205714,0.7469798,0.9507015,1.3656902,1.7618159,2.0560806,2.2560298,2.474842,2.7992878,3.8103511,5.594803,7.2358947,6.832224,6.881268,7.7301087,8.892077,9.937095,10.506761,11.321648,11.778135,11.54046,10.684074,9.703192,8.809079,8.016829,7.352846,6.828451,6.4474163,6.6662283,6.94163,6.881268,6.507778,6.2663302,6.515323,7.3717093,7.7829256,7.6282477,7.707473,8.356364,9.273112,10.137043,10.79348,11.272603,11.638548,11.6008215,11.532914,11.61214,11.815862,12.272349,12.992921,13.977575,14.739646,14.283158,13.63804,13.347548,13.298503,13.411682,13.660675,12.925014,12.268577,11.853588,11.61214,11.272603,10.831206,10.461489,9.710737,8.6732645,7.960239,7.462252,7.0548086,6.8058157,6.673774,6.519096,6.4134626,6.5643673,7.1566696,7.964011,8.333729,7.5075235,6.360646,5.934339,6.228604,6.1720147,5.704209,5.4401255,5.4665337,5.6363015,5.59103,5.13077,4.979865,4.9534564,5.070408,5.5382137,6.5643673,7.541477,8.213005,8.533678,8.695901,9.955957,11.11038,11.751727,11.68382,10.929295,9.782416,8.650629,7.496206,6.4926877,6.0286546,5.7607985,5.5495315,5.3948536,5.2590394,5.028909,7.9489207,8.541223,7.7150183,6.628502,5.824933,5.2288585,4.7006907,5.036454,5.413717,5.2137675,4.0178456,3.7575345,3.802806,4.1612053,4.889322,6.092789,5.9418845,6.1644692,6.7077274,7.333983,7.6131573,7.8206515,7.865923,7.254758,6.2097406,5.6853456,5.3609,5.2175403,5.2175403,5.2892203,5.3269467,5.3910813,5.281675,5.0741806,4.859141,4.749735,4.772371,4.919503,4.6742826,3.8895764,2.776652,2.9351022,3.8707132,4.7233267,5.0251365,4.7233267,4.772371,4.678055,4.376245,4.1197066,4.45547,5.5759397,5.8890676,5.8588867,5.3948536,3.8480775,2.9011486,3.500996,5.413717,8.039464,10.393582,9.5183325,7.7640624,6.952948,7.484888,8.307321,8.952439,8.499724,6.8850408,4.8629136,4.0103,3.591539,3.187868,2.8709676,2.6936543,2.6974268,2.625747,2.704972,2.5502944,2.2560298,2.3880715,2.9916916,3.6330378,4.2706113,4.587512,4.0178456,2.6634734,2.8030603,3.2067313,3.1652324,2.4710693,1.9881734,1.4977322,1.4600059,1.7618159,1.7240896,1.6184561,1.6071383,1.6825907,1.6373192,1.0827434,0.98465514,1.3392819,2.2899833,3.712263,5.2288585,4.930821,3.5689032,2.463524,2.1805773,2.5238862,2.0145817,1.3920987,0.8224323,0.42630664,0.26408374,0.13958712,0.09808825,0.1056335,0.29803738,0.95824677,1.871222,1.4600059,0.97333723,1.0336993,1.6222287,2.2069857,2.5880208,2.8785129,3.2331395,3.8593953,2.5578396,1.8523588,1.3694628,0.90920264,0.48666862,0.18485862,0.09808825,0.071679875,0.041498873,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.003772625,0.0,0.0,0.0,0.003772625,0.0150905,0.06413463,0.21503963,0.6149379,0.4074435,0.24522063,0.31312788,0.31312788,0.35839936,0.5319401,0.8262049,1.1657411,1.4034165,1.3053282,1.2600567,1.2034674,1.0940613,0.94315624,0.875249,0.98842776,1.0110635,0.9318384,1.0072908,0.9808825,1.1317875,1.5165952,1.8561316,1.5165952,1.2789198,1.0940613,1.0336993,1.086516,1.1921495,1.2185578,1.1581959,1.1506506,1.2562841,1.4524606,1.2147852,0.80356914,0.3734899,0.06790725,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.11317875,0.16222288,0.1358145,0.060362,0.033953626,0.018863125,0.05281675,0.2565385,0.5093044,0.69793564,0.95824677,1.3166461,1.6675003,1.6788181,1.9655377,2.2258487,2.2220762,1.7769064,1.1393328,0.66020936,0.35462674,0.19994913,0.1056335,0.056589376,0.018863125,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.003772625,0.003772625,0.003772625,0.00754525,0.011317875,0.00754525,0.018863125,0.02263575,0.026408374,0.03772625,0.071679875,0.12826926,0.1358145,0.10186087,0.06790725,0.116951376,0.13958712,0.13958712,0.13204187,0.1056335,0.00754525,0.08299775,0.3169005,0.42630664,0.33953625,0.19994913,0.20749438,0.116951376,0.0754525,0.11317875,0.1358145,0.1358145,0.120724,0.08677038,0.056589376,0.056589376,0.5281675,0.4074435,0.15467763,0.0150905,0.02263575,0.03772625,0.07922512,0.07922512,0.03772625,0.0,0.011317875,0.02263575,0.018863125,0.0150905,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.056589376,0.09808825,0.10940613,0.11317875,0.116951376,0.090543,0.06790725,0.08299775,0.181086,0.23013012,0.26031113,0.271629,0.27540162,0.30181,0.3055826,0.26031113,0.19994913,0.16222288,0.19994913,0.18863125,0.18863125,0.211267,0.24899325,0.27917424,0.1358145,0.06790725,0.041498873,0.03772625,0.056589376,0.10940613,0.20749438,0.29426476,0.331991,0.26408374,0.14335975,0.124496624,0.14713238,0.15845025,0.124496624,0.36594462,0.33953625,0.22258487,0.1358145,0.124496624,0.2263575,0.44139713,0.784706,1.056335,0.814887,0.814887,0.77716076,0.6526641,0.49421388,0.46026024,0.49421388,0.52062225,0.5281675,0.5093044,0.49044126,0.6828451,1.0374719,1.3920987,1.5882751,1.4713237,1.8825399,2.11267,2.3314822,2.7200627,3.4557245,3.6141748,3.3463185,2.7200627,1.9202662,1.2487389,1.1280149,1.3128735,1.8070874,2.4710693,3.0030096,2.4597516,1.720317,1.3807807,1.5052774,1.6222287,0.8903395,0.482896,0.31312788,0.28294688,0.30935526,0.27917424,0.23767537,0.2263575,0.23390275,0.21503963,0.19994913,0.17731337,0.16222288,0.1358145,0.08677038,0.05281675,0.0452715,0.05281675,0.06413463,0.0452715,0.09808825,0.124496624,0.13204187,0.13204187,0.15467763,0.2565385,0.2565385,0.23390275,0.2678564,0.45648763,0.7922512,0.94692886,0.94315624,0.8526133,0.80734175,0.7092535,0.5772116,0.42630664,0.2867195,0.22258487,0.2565385,0.2678564,0.29049212,0.38103512,0.6073926,0.9997456,1.5430037,1.9202662,2.071171,2.2183034,2.2862108,2.3277097,2.4786146,2.837014,3.4330888,3.5123138,3.4896781,3.8065786,4.5799665,5.594803,6.7152724,8.065872,9.473062,10.567122,10.789707,12.774108,13.615403,14.5283785,15.965749,17.652113,18.274595,16.961721,14.992412,13.011784,11.042474,10.495442,9.590013,8.699674,7.726336,6.092789,8.703445,11.091517,11.302785,9.193887,6.439871,7.3151197,5.2854476,3.1161883,1.9994912,1.5505489,1.2487389,1.4109617,1.8900851,2.584248,3.4557245,4.274384,4.708236,4.8930945,5.0439997,5.4703064,7.1378064,8.526133,10.061591,12.00072,14.4152,16.807045,19.051756,20.172226,19.825144,18.289686,16.51278,13.747445,11.212241,9.65792,9.344792,9.333474,8.495952,7.394345,6.760544,7.4999785,8.707218,9.49947,9.914458,9.967276,9.623966,8.5563135,7.6093845,6.983129,6.692637,6.537959,6.571913,6.1720147,5.2854476,4.0178456,2.6446102,2.1164427,1.6675003,1.3468271,1.1808317,1.1808317,1.0827434,0.97333723,0.7130261,0.362172,0.16976812,0.211267,0.34330887,0.452715,0.49421388,0.5093044,0.5696664,0.6375736,0.633801,0.56589377,0.5357128,0.51684964,0.44894236,0.46026024,0.5885295,0.784706,1.0412445,1.3355093,1.6788181,2.0296721,2.3163917,2.4522061,3.048281,3.8556228,4.4630156,4.3121104,4.7120085,6.79827,9.457971,11.849815,13.404137,14.215251,14.547242,14.083209,13.015556,12.034674,11.876224,11.336739,10.574668,9.74469,8.990166,8.458225,8.458225,8.461998,8.303548,8.16396,8.088508,8.2507305,8.52236,8.820397,9.125979,9.310839,9.623966,9.914458,10.235131,10.86516,11.725319,11.996947,11.98563,11.940358,12.064855,12.66093,13.619176,14.800008,16.116653,17.527617,16.897587,16.177015,15.656394,15.497944,15.731846,14.815099,14.117163,13.721037,13.472044,12.958967,12.264804,11.574413,10.801025,9.933322,9.046755,8.541223,7.9526935,7.375482,6.900131,6.6058664,6.5832305,6.696409,7.1038527,7.748972,8.329956,7.673519,7.115171,7.2170315,7.6093845,6.983129,6.3417826,5.8400235,5.6589375,5.6363015,5.2665844,5.4250345,5.66271,5.7306175,5.670255,5.836251,6.405917,6.9680386,7.3000293,7.466025,7.7904706,8.805306,9.861642,10.480352,10.510533,10.103089,9.5183325,8.944894,8.20546,7.3679366,6.749226,6.2814207,5.80607,5.4778514,5.3080835,5.1571784,7.0963078,6.6813188,6.3945994,6.6058664,6.8435416,5.7683434,4.779916,4.715781,5.5759397,6.175787,4.1498876,3.783943,3.4444065,3.6481283,4.4215164,5.3269467,5.594803,5.485397,5.836251,6.760544,7.673519,8.567632,8.8618965,8.43559,7.7602897,7.91874,7.515069,6.6662283,6.006019,5.87775,6.3153744,6.8171334,6.4021444,5.80607,5.3873086,5.142088,4.274384,3.591539,3.2935016,3.059599,2.0447628,2.191895,4.4139714,5.764571,5.1647234,3.4179983,3.4179983,3.4632697,3.2369123,3.0256453,3.7235808,4.0517993,4.2894745,4.504514,4.7044635,4.8365054,4.5912848,5.198677,6.0286546,6.571913,6.439871,6.013564,6.571913,7.3679366,8.296002,9.918231,12.51757,12.178034,9.280658,5.451443,3.5689032,3.8141239,4.1498876,4.3196554,4.1762958,3.663219,2.9049213,2.4786146,2.2711203,2.2069857,2.2447119,2.8521044,3.7462165,4.8025517,5.715527,5.994701,3.7613072,3.7537618,3.8254418,3.218049,2.5314314,2.1164427,1.629774,1.5882751,1.9089483,1.9089483,2.0183544,2.082489,2.033445,1.8523588,1.5731846,1.6222287,1.9881734,2.3201644,2.7615614,3.983892,4.7044635,3.893349,2.5389767,1.6335466,2.1805773,1.3996439,0.8865669,0.6526641,0.56589377,0.33576363,0.21503963,0.120724,0.06413463,0.1056335,0.33576363,1.4826416,2.674791,2.1768045,0.7167987,1.50905,1.8523588,2.0862615,2.2371666,2.282438,2.1353056,1.539231,1.478869,1.2713746,0.7432071,0.24522063,0.09808825,0.033953626,0.026408374,0.041498873,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.026408374,0.030181,0.018863125,0.0,0.0,0.0,0.018863125,0.041498873,0.07922512,0.150905,0.26408374,0.271629,0.5394854,0.94692886,0.8865669,0.935611,1.237421,1.6524098,2.0145817,2.1353056,1.8297231,1.5882751,1.3958713,1.2223305,1.0525624,0.90543,0.9808825,1.0638802,1.056335,0.94692886,0.87147635,0.965792,1.20724,1.478869,1.5430037,1.1732863,1.0186088,0.9997456,1.0450171,1.0827434,1.0601076,0.9808825,1.2185578,1.6976813,1.8938577,1.5241405,0.95824677,0.38480774,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16976812,0.17731337,0.090543,0.0,0.0,0.1358145,0.2867195,0.52439487,0.83752275,1.1431054,2.1692593,2.9011486,3.1048703,2.7879698,2.2296214,1.629774,0.9393836,0.5017591,0.3470815,0.21503963,0.116951376,0.0452715,0.00754525,0.0,0.0,0.011317875,0.0150905,0.00754525,0.003772625,0.0150905,0.0150905,0.02263575,0.041498873,0.056589376,0.030181,0.041498873,0.0452715,0.06413463,0.1056335,0.1659955,0.21503963,0.26408374,0.21503963,0.090543,0.030181,0.041498873,0.056589376,0.056589376,0.0452715,0.0452715,0.27917424,0.34330887,0.271629,0.12826926,0.030181,0.056589376,0.041498873,0.03772625,0.049044125,0.060362,0.071679875,0.056589376,0.0452715,0.0452715,0.0452715,0.20372175,0.18863125,0.090543,0.00754525,0.0452715,0.13204187,0.362172,0.392353,0.18485862,0.0,0.011317875,0.041498873,0.06790725,0.071679875,0.0452715,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.06790725,0.1056335,0.124496624,0.1358145,0.16222288,0.1056335,0.056589376,0.056589376,0.1056335,0.20372175,0.24899325,0.23013012,0.181086,0.1659955,0.27917424,0.36971724,0.4074435,0.38480774,0.33576363,0.31312788,0.36971724,0.41121614,0.3772625,0.24522063,0.15845025,0.12826926,0.116951376,0.1056335,0.090543,0.17731337,0.30935526,0.44139713,0.5093044,0.41121614,0.14335975,0.06790725,0.056589376,0.06413463,0.1358145,0.32067314,0.4376245,0.44516975,0.35839936,0.26031113,0.18485862,0.18485862,0.30181,0.47157812,0.5357128,0.4376245,0.47535074,0.48666862,0.4979865,0.7167987,0.72811663,0.80734175,0.9507015,1.0638802,0.9318384,0.8224323,0.9205205,1.2751472,1.8372684,2.4710693,2.6295197,2.3767538,2.4031622,2.7351532,2.746471,2.4182527,1.8938577,1.3505998,0.87147635,0.44139713,0.47912338,1.0751982,1.8938577,2.5502944,2.625747,1.478869,0.7696155,0.5319401,0.5357128,0.3055826,0.14713238,0.09808825,0.09808825,0.11317875,0.1358145,0.1358145,0.15467763,0.211267,0.27917424,0.29049212,0.25276586,0.19994913,0.15467763,0.124496624,0.0754525,0.10186087,0.09808825,0.071679875,0.0452715,0.0452715,0.120724,0.1659955,0.21881226,0.31312788,0.47157812,0.59607476,0.6451189,0.59607476,0.49044126,0.44139713,0.271629,0.14713238,0.14713238,0.271629,0.44139713,0.5885295,0.48666862,0.32821837,0.22258487,0.19994913,0.22258487,0.24899325,0.26408374,0.29049212,0.35085413,0.59607476,1.2147852,1.6222287,1.7542707,2.0598533,2.4031622,2.3390274,2.2786655,2.4182527,2.7615614,2.8709676,2.8634224,3.0331905,3.482133,4.104616,5.4703064,7.24344,8.89585,9.982366,10.11818,10.616167,10.650121,11.370691,12.951422,14.588741,16.28265,16.478827,15.369675,13.751218,13.030646,11.955449,10.005001,8.043237,6.4964604,5.3269467,7.779153,12.193124,13.200415,10.272858,7.7225633,8.001738,6.277648,3.953711,2.123988,1.5882751,1.3920987,2.3578906,3.8405323,5.715527,8.375228,9.329701,10.325675,10.148361,8.888305,7.9489207,8.122461,10.570895,14.056801,17.384256,19.410156,20.715485,22.130219,22.416937,21.073883,18.327412,15.347038,12.442118,10.623712,10.076681,10.163452,9.416472,8.171506,6.7643166,5.885295,6.5455046,7.756517,8.669493,9.001483,8.76758,8.314865,7.4735703,6.4210076,5.847569,5.915476,6.255012,6.828451,6.790725,5.885295,4.447925,3.3878171,2.71629,1.9806281,1.4675511,1.2185578,1.0223814,0.7167987,0.5583485,0.33953625,0.09808825,0.120724,0.16976812,0.2565385,0.35462674,0.4376245,0.47157812,0.48666862,0.6073926,0.65643674,0.58475685,0.48666862,0.4376245,0.44516975,0.55080324,0.73566186,0.9318384,1.0412445,1.2336484,1.5505489,1.9504471,2.305074,2.1466236,2.335255,2.6823363,3.006782,3.127506,3.7613072,5.323174,7.8319697,10.853842,13.487134,15.98084,17.4333,17.538933,16.403374,14.57365,14.32843,14.249205,13.905896,13.249459,12.604341,11.359374,10.242677,9.850324,10.299266,11.216014,10.751981,10.03141,9.718282,9.831461,9.733373,10.321902,10.084227,9.623966,9.473062,10.069136,11.536687,12.525115,12.958967,12.992921,13.015556,13.113645,14.045483,15.580941,17.493662,19.53088,20.960705,20.519308,19.17248,17.784155,17.135263,17.195625,16.984358,16.395828,15.460217,14.313339,13.72481,13.377728,12.781653,11.857361,10.940613,10.121953,9.469289,8.975075,8.571404,8.13378,8.265821,8.118689,7.816879,7.8319697,8.941121,8.477088,8.737399,9.1825695,9.337247,8.790216,7.141579,6.7944975,6.2323766,5.413717,5.7683434,6.609639,7.149124,7.1868505,6.8246784,6.470052,6.541732,6.8171334,6.779407,6.507778,6.670001,7.6810646,8.831716,9.748463,10.103089,9.627739,8.944894,8.646856,8.511042,8.397863,8.239413,7.4094353,6.5530496,5.9117036,5.4740787,4.9760923,6.5945487,6.832224,7.0548086,7.2924843,7.141579,5.7419353,4.979865,4.979865,5.523123,6.085244,5.836251,5.5193505,5.3609,5.300538,5.292993,5.2892203,4.776143,4.3800178,4.7233267,6.2323766,9.14107,9.201432,8.790216,8.031919,7.220804,6.832224,6.8774953,7.1302614,7.413208,7.5301595,7.2585306,6.6134114,5.8928404,5.349582,4.9723196,4.496969,4.889322,4.285702,3.5123138,2.9539654,2.5578396,2.674791,3.8443048,4.187614,3.4255435,2.8822856,2.4899325,2.4371157,2.8143783,3.270866,3.0256453,3.5538127,4.115934,4.5196047,4.749735,4.983638,5.587258,6.319147,7.039718,7.7602897,8.661947,8.684583,8.186596,7.4999785,7.224577,8.22055,12.50248,13.943622,12.574159,9.261794,5.7419353,4.5724216,6.092789,7.009537,6.4436436,5.934339,5.0477724,4.3422914,3.9197574,3.5500402,2.6597006,2.6634734,3.1652324,4.0216184,5.0251365,5.9117036,5.541986,4.3309736,3.5689032,3.4745877,3.180323,2.5201135,1.8976303,1.6410918,1.8070874,2.1881225,2.6408374,2.8030603,2.655928,2.2371666,1.6335466,1.2336484,1.327964,1.871222,2.727608,3.6669915,3.4859054,2.6823363,1.871222,1.5316857,1.9730829,1.3770081,0.814887,0.44139713,0.2867195,0.24899325,0.2263575,0.17731337,0.11317875,0.06790725,0.1056335,0.32444575,0.6752999,0.77716076,0.6375736,0.6790725,1.1016065,1.4562333,1.720317,1.8863125,1.9542197,1.8938577,1.8523588,1.3392819,0.5319401,0.2565385,0.18863125,0.21503963,0.41121614,0.5281675,0.0150905,0.05281675,0.0452715,0.041498873,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.003772625,0.0,0.0,0.0,0.011317875,0.0452715,0.1056335,0.18863125,0.30935526,0.452715,0.7205714,1.1544232,1.7391801,1.6825907,1.4524606,1.3770081,1.5128226,1.6712729,1.4826416,1.5015048,1.5279131,1.4675511,1.297783,1.1204696,1.026154,0.95824677,0.875249,0.72811663,0.6149379,0.56212115,0.58475685,0.69793564,0.94315624,0.94692886,0.9507015,1.0223814,1.1431054,1.2185578,1.086516,0.98842776,1.177059,1.6184561,1.9881734,1.780679,1.2600567,0.6451189,0.15467763,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033953626,0.033953626,0.06790725,0.09808825,0.0,0.026408374,0.056589376,0.16976812,0.3961256,0.72811663,1.3430545,2.0900342,2.6295197,2.8106055,2.6672459,2.1956677,1.237421,0.7582976,0.80734175,0.5055317,0.241448,0.116951376,0.049044125,0.018863125,0.03772625,0.060362,0.094315626,0.11317875,0.1056335,0.08677038,0.07922512,0.120724,0.15467763,0.15845025,0.150905,0.124496624,0.09808825,0.08299775,0.0754525,0.056589376,0.06790725,0.08299775,0.07922512,0.056589376,0.056589376,0.116951376,0.17731337,0.17354076,0.10940613,0.071679875,0.124496624,0.20749438,0.27540162,0.2565385,0.030181,0.033953626,0.026408374,0.0150905,0.011317875,0.011317875,0.0150905,0.011317875,0.00754525,0.00754525,0.00754525,0.041498873,0.06790725,0.10940613,0.16222288,0.181086,0.21503963,0.32067314,0.3169005,0.17354076,0.0,0.003772625,0.00754525,0.0150905,0.0150905,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.026408374,0.026408374,0.041498873,0.033953626,0.026408374,0.0452715,0.094315626,0.16222288,0.18485862,0.21881226,0.271629,0.29049212,0.331991,0.38480774,0.44516975,0.482896,0.44516975,0.5885295,0.77338815,0.95447415,1.0601076,1.0148361,0.724344,0.45648763,0.3055826,0.32067314,0.543258,0.5394854,0.5017591,0.51684964,0.513077,0.27917424,0.1659955,0.09808825,0.071679875,0.094315626,0.18485862,0.4074435,0.77716076,1.3091009,1.6863633,1.297783,0.69793564,0.32444575,0.17354076,0.1659955,0.120724,0.15845025,0.20372175,0.2867195,0.5017591,0.97333723,1.6410918,2.0560806,1.9051756,1.4034165,1.297783,1.0601076,0.9318384,1.1619685,1.8070874,2.71629,3.3048196,3.0407357,2.4786146,1.9202662,1.4147344,1.0676528,0.79602385,0.5885295,0.45648763,0.43007925,0.69039035,1.0336993,1.388326,1.8787673,2.8332415,1.7127718,0.9242931,0.4678055,0.26031113,0.14713238,0.056589376,0.05281675,0.07922512,0.090543,0.0754525,0.15467763,0.22258487,0.23390275,0.1961765,0.181086,0.17354076,0.124496624,0.07922512,0.060362,0.10186087,0.1659955,0.120724,0.090543,0.13958712,0.26408374,0.30935526,0.29803738,0.27917424,0.271629,0.25276586,0.422534,0.86770374,1.1657411,1.1393328,0.8563859,0.5696664,0.25276586,0.094315626,0.10186087,0.1358145,0.1659955,0.14713238,0.10940613,0.08299775,0.0754525,0.20749438,0.2678564,0.27540162,0.27917424,0.35085413,0.5772116,0.9393836,1.2147852,1.4713237,2.1088974,2.3805263,2.282438,2.1051247,2.04099,2.1881225,2.2484846,2.5427492,2.9803739,3.519859,4.1536603,5.089271,6.217286,7.092535,7.6584287,8.262049,8.907167,9.608876,10.646348,12.098808,13.841762,18.13878,17.984104,16.365646,15.049001,14.592513,13.607859,11.623458,10.329447,9.684328,7.937603,9.903141,12.340257,12.687338,11.348056,11.6875925,11.363147,8.2507305,5.0779533,3.308592,3.1124156,2.8596497,4.779916,6.1342883,7.1340337,10.929295,13.766309,14.532151,13.290957,11.00852,9.559832,11.16697,14.6302395,17.512526,18.761265,18.689585,19.723284,20.783392,20.85507,19.628967,17.497435,14.879233,12.6345215,11.234878,10.631257,10.246449,9.454198,8.371455,7.2283497,6.4210076,6.485142,7.4999785,8.182823,7.9941926,7.115171,6.4474163,5.926794,5.5193505,5.323174,5.270357,5.1345425,6.156924,6.7567716,6.6058664,5.7306175,4.5233774,3.3350005,1.9693103,0.9507015,0.44894236,0.30181,0.241448,0.1961765,0.1358145,0.08677038,0.120724,0.150905,0.2263575,0.30935526,0.38858038,0.47157812,0.5357128,0.573439,0.5470306,0.47535074,0.41498876,0.38480774,0.3961256,0.47157812,0.6187105,0.8337501,0.80734175,0.95824677,1.2223305,1.4977322,1.6561824,1.6561824,2.3013012,2.7125173,2.6144292,2.3465726,2.5502944,3.380272,4.82896,6.771862,8.959985,11.400873,14.947141,18.135008,19.927006,19.700647,17.70493,16.056292,15.026365,14.335975,13.151371,12.2119875,11.491416,10.899114,10.484125,10.419991,10.816116,10.533169,10.103089,9.8239155,9.748463,9.989911,9.559832,8.763808,8.2507305,8.98262,10.076681,11.69891,13.290957,14.362384,14.494425,14.4152,14.679284,15.686575,17.56157,20.16468,22.620659,23.812809,23.631723,22.424482,21.017294,20.775846,21.175745,21.379465,20.602304,18.1086,16.82968,15.78089,14.879233,14.083209,13.392818,12.73261,12.015811,11.321648,10.816116,10.7557535,10.159679,9.593785,9.310839,9.26934,9.099571,9.495697,9.099571,8.197914,7.1038527,6.1531515,5.5683947,5.4288073,5.4288073,5.5268955,5.9494295,6.217286,6.2323766,6.096562,5.96452,6.0286546,6.2399216,6.2851934,6.1644692,5.9984736,6.0211096,6.790725,7.8810134,9.0543,10.042727,10.544487,10.495442,10.280403,9.903141,9.310839,8.409182,7.541477,6.477597,5.80607,5.583485,5.3156285,5.372218,4.930821,4.878004,5.111907,5.406172,5.4174895,5.7570257,6.587003,7.2396674,7.183078,6.043745,5.036454,4.534695,4.5497856,5.0213637,5.7909794,4.908185,4.508287,4.8063245,6.0701537,8.627994,9.695646,9.793735,9.318384,8.571404,7.7602897,7.0548086,6.964266,7.24344,7.466025,7.0170827,6.168242,5.515578,5.0025005,4.6516466,4.561104,5.198677,4.859141,4.3309736,3.9348478,3.5274043,3.1312788,3.2029586,3.097325,2.7615614,2.727608,2.8634224,2.8747404,2.8709676,2.7728794,2.3314822,2.6785638,3.531177,4.274384,4.749735,5.2779026,5.772116,6.0248823,6.1342883,6.4134626,7.4018903,8.356364,7.8131065,6.677546,5.7419353,5.6551647,7.564113,10.374719,12.166716,11.955449,9.699419,7.854605,7.7414265,7.707473,6.9869013,5.704209,5.5268955,5.692891,5.9984736,6.1041074,5.5080323,4.606375,3.8443048,3.7160356,4.4516973,6.017337,6.6360474,5.6023483,4.183841,3.218049,3.138824,2.655928,2.7200627,2.987919,3.1463692,2.927557,2.6219745,2.6710186,2.6332922,2.4861598,2.6446102,2.6106565,2.2899833,2.0598533,2.2862108,3.3312278,2.9766011,2.4220252,2.022127,1.9240388,2.0673985,1.1883769,0.68661773,0.43385187,0.34330887,0.3470815,0.331991,0.27540162,0.1659955,0.049044125,0.0452715,0.07922512,0.21503963,0.46026024,0.724344,0.8224323,0.7469798,1.0148361,1.3166461,1.5316857,1.7429527,1.8372684,1.6637276,1.1808317,0.5772116,0.27917424,0.16222288,0.16976812,0.29803738,0.3772625,0.07922512,0.09808825,0.05281675,0.02263575,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.05281675,0.056589376,0.056589376,0.0754525,0.15467763,0.060362,0.033953626,0.071679875,0.16976812,0.33576363,0.60362,0.9280658,1.1581959,1.4524606,2.2560298,2.3088465,1.9844007,1.6260014,1.4260522,1.4373702,1.3732355,1.478869,1.5618668,1.5505489,1.4675511,1.388326,1.2864652,1.1355602,0.9242931,0.663982,0.4979865,0.422534,0.43385187,0.543258,0.784706,0.845068,0.88279426,0.97710985,1.1091517,1.1883769,1.0789708,1.1808317,1.3732355,1.5656394,1.7014539,1.6637276,1.3920987,0.875249,0.29803738,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.049044125,0.0,0.0,0.0,0.041498873,0.16222288,0.38858038,0.87147635,1.4109617,1.8976303,2.2560298,2.4371157,2.0862615,1.2411937,0.69793564,0.59607476,0.422534,0.331991,0.2867195,0.32444575,0.45648763,0.6790725,0.6790725,0.59607476,0.49421388,0.4074435,0.35462674,0.35085413,0.331991,0.28294688,0.211267,0.14713238,0.116951376,0.13204187,0.124496624,0.07922512,0.02263575,0.056589376,0.1358145,0.20749438,0.241448,0.21503963,0.18863125,0.181086,0.13958712,0.07922512,0.056589376,0.11317875,0.21503963,0.2867195,0.26031113,0.0754525,0.05281675,0.049044125,0.049044125,0.041498873,0.026408374,0.033953626,0.018863125,0.011317875,0.06413463,0.23767537,0.362172,0.19994913,0.07922512,0.08677038,0.08677038,0.116951376,0.1659955,0.17354076,0.11317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.0150905,0.0,0.0,0.018863125,0.033953626,0.056589376,0.094315626,0.17354076,0.2867195,0.362172,0.42630664,0.47157812,0.4678055,0.44139713,0.42630664,0.43007925,0.44139713,0.41876137,0.5055317,0.69039035,1.0148361,1.5731846,2.516341,1.8297231,1.297783,1.0751982,1.1619685,1.4071891,1.3241913,1.5316857,1.7278622,1.7467253,1.5543215,1.3128735,0.9808825,0.58475685,0.23767537,0.14335975,0.21503963,0.5319401,1.1808317,1.8825399,1.9693103,1.0223814,0.482896,0.23013012,0.14335975,0.071679875,0.08299775,0.094315626,0.16222288,0.392353,0.935611,1.3128735,1.5731846,1.5279131,1.2789198,1.2223305,1.297783,1.4147344,1.9466745,2.8030603,3.399135,3.5236318,3.1010978,2.4710693,1.7882242,0.9922004,0.8224323,0.7130261,0.6413463,0.6149379,0.7092535,0.97710985,1.1242423,1.1883769,1.3166461,1.7957695,1.2638294,0.7205714,0.331991,0.13958712,0.071679875,0.056589376,0.06790725,0.07922512,0.07922512,0.071679875,0.10186087,0.15845025,0.18485862,0.16976812,0.16222288,0.15467763,0.13958712,0.1056335,0.0754525,0.116951376,0.150905,0.13958712,0.17731337,0.32444575,0.5772116,0.46026024,0.43385187,0.42630664,0.3961256,0.33576363,0.3734899,0.6111652,0.98842776,1.3392819,1.3996439,1.1431054,0.7092535,0.32821837,0.120724,0.14335975,0.09808825,0.08677038,0.094315626,0.10186087,0.10940613,0.17354076,0.22258487,0.24899325,0.3055826,0.48666862,0.7507524,1.1016065,1.4562333,1.7731338,2.0749438,2.0673985,2.052308,2.0258996,2.0296721,2.1353056,2.3163917,2.746471,3.3010468,3.9008942,4.5120597,5.2552667,5.9909286,6.4436436,6.6322746,6.900131,7.4811153,8.348819,9.246704,10.367173,12.366665,16.271332,16.87118,16.376965,15.645076,14.177525,12.687338,11.076427,10.061591,10.26154,12.215759,12.872196,13.570132,12.706201,10.834979,10.665211,13.147598,11.34051,8.397863,6.2625575,5.643847,5.485397,6.760544,8.20546,9.906913,13.29473,15.331948,15.230087,13.849306,12.310076,12.034674,14.841507,19.549744,22.439573,22.541435,21.65864,21.062565,20.168453,19.017803,17.753973,16.618414,14.841507,13.057055,11.668729,10.763299,10.133271,9.590013,8.484633,7.2962565,6.511551,6.617184,7.4697976,7.858378,7.4471617,6.417235,5.4703064,5.2326307,5.240176,5.194905,4.90064,4.255521,4.2781568,5.0477724,5.7192993,5.8966126,5.613666,4.346064,2.4408884,0.91674787,0.1961765,0.120724,0.120724,0.10940613,0.1056335,0.120724,0.150905,0.17354076,0.23390275,0.30181,0.36594462,0.41876137,0.47535074,0.52062225,0.56589377,0.59607476,0.52439487,0.52062225,0.573439,0.6790725,0.8299775,0.9808825,0.9205205,0.9507015,1.0714256,1.2185578,1.2751472,1.2826926,1.690136,2.1051247,2.2484846,1.931584,1.780679,1.9466745,2.5201135,3.5424948,5.0175915,7.145352,10.963248,15.275358,18.908396,20.69662,19.76101,18.372684,17.237123,16.275105,14.588741,13.306048,12.559069,12.155397,11.9064045,11.661184,11.823407,11.234878,10.393582,9.691874,9.393836,9.559832,9.14107,8.213005,7.586749,8.793989,9.767326,11.438599,13.415455,14.856597,14.494425,15.339493,16.003475,17.105082,18.923487,21.405874,23.835445,25.642532,26.90636,26.940315,24.295706,22.975286,22.8357,22.730066,21.967995,20.323132,19.379974,18.23687,17.172989,16.301512,15.573396,14.875461,14.18507,13.434318,12.815607,12.777881,11.966766,11.091517,10.431308,10.035183,9.7069645,9.533423,8.869441,7.7640624,6.477597,5.5004873,5.300538,4.9949555,4.979865,5.251494,5.4212623,5.43258,5.2892203,5.0741806,4.9421387,5.1043615,5.3948536,5.485397,5.6023483,5.7872066,5.915476,6.1305156,6.964266,8.118689,9.318384,10.306811,10.627484,10.555805,10.246449,9.733373,8.91094,7.960239,6.960493,6.2663302,5.9796104,5.9682927,4.6214657,3.6669915,3.180323,3.150142,3.4859054,4.036709,5.330719,6.7831798,7.564113,7.1679873,5.4288073,4.293247,3.7537618,3.7650797,4.2517486,5.119452,4.7610526,5.010046,5.798525,6.952948,8.216777,9.906913,10.540714,10.412445,9.922004,9.590013,8.326183,7.164215,6.6322746,6.6549106,6.5945487,6.255012,5.783434,5.194905,4.719554,4.8327327,5.1873593,5.353355,5.7079816,5.9984736,5.3269467,4.7233267,4.032936,3.5990841,3.5160866,3.5953116,3.4444065,3.270866,3.0860074,2.8445592,2.4597516,2.3314822,2.7728794,3.5424948,4.8553686,7.375482,7.3113475,7.1906233,6.862405,6.560595,6.903904,7.6395655,7.699928,6.7869525,5.3986263,4.82896,5.409944,8.13378,10.827434,11.910177,10.386037,8.733627,8.016829,7.726336,7.201941,5.6363015,5.8664317,6.8058157,7.673519,8.001738,7.6320205,6.688864,5.6513925,4.9421387,4.9534564,6.0776987,6.530414,6.2361493,5.406172,4.4215164,3.8292143,3.169005,3.218049,3.440634,3.4217708,2.8596497,2.0673985,1.841041,2.022127,2.584248,3.6330378,4.0404816,3.6745367,3.0143273,2.655928,3.2935016,2.969056,2.5276587,2.1466236,1.9051756,1.7693611,1.1355602,0.814887,0.6111652,0.45648763,0.3961256,0.362172,0.29803738,0.17731337,0.060362,0.0754525,0.10940613,0.17354076,0.32067314,0.5470306,0.80734175,0.6828451,0.7997965,1.0186088,1.2562841,1.50905,1.629774,1.448688,1.0789708,0.6526641,0.31312788,0.15467763,0.14713238,0.18863125,0.20749438,0.12826926,0.181086,0.07922512,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.094315626,0.14713238,0.14713238,0.15467763,0.23013012,0.41876137,0.7469798,0.4074435,0.2263575,0.21503963,0.35462674,0.59230214,0.84129536,1.0223814,1.1317875,1.3355093,1.961765,2.1315331,2.003264,1.7316349,1.4750963,1.3656902,1.448688,1.5807298,1.6373192,1.6071383,1.6033657,1.6863633,1.6561824,1.4524606,1.1091517,0.7582976,0.55457586,0.48666862,0.5319401,0.6526641,0.7922512,0.7394345,0.7809334,0.8865669,1.0072908,1.0638802,1.0223814,1.1808317,1.3166461,1.3317367,1.2638294,1.3204187,1.2487389,0.86770374,0.32067314,0.056589376,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026408374,0.03772625,0.060362,0.19240387,0.48666862,0.784706,1.1280149,1.5128226,1.871222,1.7354075,1.358145,1.0487897,0.91297525,0.8639311,0.88279426,0.8526133,0.91297525,1.1091517,1.4109617,1.418507,1.2223305,1.0072908,0.8563859,0.7394345,0.7130261,0.62248313,0.47912338,0.32821837,0.23013012,0.241448,0.2867195,0.29803738,0.26031113,0.211267,0.21881226,0.2565385,0.2867195,0.27917424,0.21503963,0.13958712,0.09808825,0.060362,0.030181,0.0452715,0.11317875,0.16976812,0.20749438,0.211267,0.15467763,0.1056335,0.071679875,0.056589376,0.05281675,0.056589376,0.049044125,0.026408374,0.018863125,0.08677038,0.29426476,0.44139713,0.24899325,0.06413463,0.018863125,0.011317875,0.033953626,0.060362,0.07922512,0.06790725,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.049044125,0.03772625,0.03772625,0.05281675,0.06413463,0.08299775,0.120724,0.19994913,0.30935526,0.41121614,0.47535074,0.51684964,0.56589377,0.46026024,0.36971724,0.32067314,0.32067314,0.35085413,0.43385187,0.5885295,0.8526133,1.4260522,2.6672459,2.263575,1.8599042,1.7731338,2.2220762,3.3350005,3.5462675,3.92353,3.9763467,3.5764484,2.9464202,2.5729303,2.2673476,1.6825907,0.8941121,0.422534,0.211267,0.29049212,0.694163,1.2864652,1.750498,1.0676528,0.663982,0.44139713,0.31312788,0.21503963,0.181086,0.23013012,0.35462674,0.58098423,0.9507015,1.0186088,1.1129243,1.0978339,1.0035182,1.0336993,1.3317367,1.8938577,2.6974268,3.4255435,3.4783602,3.4066803,2.8106055,2.142851,1.5920477,1.0601076,1.2110126,1.3015556,1.237421,1.146878,1.3807807,1.3732355,1.1317875,0.86770374,0.7092535,0.7092535,0.62625575,0.392353,0.19240387,0.094315626,0.05281675,0.08299775,0.08677038,0.090543,0.09808825,0.08677038,0.08299775,0.124496624,0.16976812,0.181086,0.14335975,0.16976812,0.20749438,0.19994913,0.15467763,0.13958712,0.14335975,0.1961765,0.29426476,0.452715,0.7167987,0.633801,0.59607476,0.573439,0.543258,0.47535074,0.42630664,0.4074435,0.58475685,0.9205205,1.1808317,1.1242423,0.87902164,0.5470306,0.27540162,0.271629,0.20749438,0.16222288,0.1659955,0.23013012,0.36594462,0.47535074,0.482896,0.45648763,0.482896,0.663982,0.90920264,1.2110126,1.5580941,1.8636768,1.9768555,1.9051756,1.9881734,2.093807,2.1843498,2.2899833,2.6898816,3.1539145,3.6669915,4.172523,4.606375,5.194905,5.802297,6.296511,6.6586833,6.9793563,7.413208,7.779153,8.096053,8.903395,11.283921,14.524607,16.22606,16.97304,16.505234,13.732355,11.69891,10.0465,9.110889,9.714509,13.155144,14.007756,14.241659,12.985375,10.702937,9.201432,11.978085,11.200924,9.2844305,7.7716074,7.33021,6.9454026,7.7640624,9.1825695,10.816116,12.521342,13.057055,12.611885,12.294985,12.872196,14.754736,18.350048,22.371666,24.48811,24.378702,23.726038,22.100037,19.768555,17.64834,16.263786,15.735619,14.939595,13.370183,11.751727,10.570895,10.076681,10.314357,9.891823,8.91094,7.8508325,7.5263867,7.6093845,7.3792543,6.7341356,5.7872066,4.889322,4.9044123,4.983638,4.870459,4.4139714,3.5802212,2.9954643,3.4745877,4.191386,4.7648253,5.251494,4.2328854,2.4408884,0.965792,0.2678564,0.16976812,0.120724,0.11317875,0.12826926,0.15845025,0.19240387,0.2263575,0.271629,0.331991,0.38103512,0.38858038,0.42630664,0.49044126,0.60362,0.7092535,0.67152727,0.66775465,0.7432071,0.91297525,1.1355602,1.2940104,1.2411937,1.2336484,1.2713746,1.3128735,1.2562841,1.1619685,1.3015556,1.7089992,2.082489,1.7957695,1.4147344,1.2185578,1.3015556,1.7240896,2.4823873,3.783943,6.349328,9.982366,14.064346,17.580433,18.534906,18.576405,18.433046,18.03692,16.531643,14.958458,14.128481,13.792717,13.641812,13.328684,13.3626375,12.510024,11.332966,10.370946,10.125726,10.408672,10.597303,10.065364,9.424017,10.510533,11.231105,12.113899,13.249459,14.18507,13.947394,15.328176,16.614641,18.229324,20.19109,22.111355,24.118391,26.046204,28.038149,29.124664,27.200626,25.506718,24.857826,24.250433,23.314823,22.29244,22.10381,21.149336,20.013775,19.021576,18.202915,17.523844,17.037174,16.229834,15.113135,14.241659,13.264549,12.261031,11.23865,10.374719,10.001229,9.461743,8.793989,7.960239,7.01331,6.1003346,5.7494807,5.7306175,5.6023483,5.2854476,5.0477724,5.070408,4.938366,4.715781,4.564876,4.7572803,4.957229,5.1043615,5.3269467,5.5759397,5.6325293,5.873977,6.537959,7.5112963,8.616675,9.6051035,9.827688,9.673011,9.382519,9.039209,8.563859,7.8206515,7.149124,6.677546,6.466279,6.530414,4.357382,3.561358,2.9011486,2.4861598,2.2786655,2.1013522,3.4934506,4.927048,5.7683434,5.6513925,4.478106,3.7348988,3.482133,3.361409,3.2520027,3.2670932,3.904667,5.0025005,6.3945994,7.635793,7.986647,9.710737,10.585986,10.823661,10.895341,11.532914,10.499215,8.616675,7.273621,6.881268,6.8737226,6.983129,6.620957,5.9682927,5.349582,5.247721,5.2175403,5.726845,6.722818,7.496206,6.651138,6.1720147,5.3194013,4.7308717,4.636556,4.847823,3.9159849,3.3350005,3.338773,3.6556737,3.5085413,2.9124665,2.4484336,2.8030603,4.82896,9.548513,10.280403,10.170997,9.58624,8.884532,8.420499,7.9941926,8.688355,8.299775,6.6586833,5.6400743,7.001992,8.707218,9.955957,9.933322,7.8244243,6.8963585,7.0887623,7.4094353,7.201941,6.1418333,6.1833324,7.24344,8.13378,8.36391,8.137552,8.096053,7.9791017,7.4584794,6.647365,6.089017,6.006019,6.579458,7.1793056,7.0963078,5.560849,4.093298,3.187868,2.7389257,2.4823873,2.033445,1.3656902,0.91674787,1.2336484,2.372981,3.863168,4.7836885,5.0515447,4.768598,4.183841,3.682082,3.059599,2.5578396,2.0183544,1.4901869,1.2223305,1.2713746,1.177059,0.8639311,0.4640329,0.30181,0.28294688,0.241448,0.1659955,0.09808825,0.13204187,0.116951376,0.071679875,0.06413463,0.16976812,0.49044126,0.8563859,0.8262049,0.8601585,1.086516,1.297783,1.4562333,1.4109617,1.1091517,0.663982,0.35839936,0.23390275,0.20749438,0.20749438,0.18485862,0.116951376,0.2263575,0.10186087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.011317875,0.06413463,0.18863125,0.32444575,0.33953625,0.29049212,0.38480774,0.62625575,0.98842776,1.3958713,0.91674787,0.5281675,0.38103512,0.5017591,0.76584285,0.9280658,0.8526133,0.83752275,0.9997456,1.3053282,1.5052774,1.6373192,1.6788181,1.6184561,1.4524606,1.6071383,1.6712729,1.6448646,1.6033657,1.6863633,1.9504471,2.052308,1.8334957,1.3619176,0.95447415,0.7205714,0.6413463,0.69039035,0.80734175,0.8865669,0.6413463,0.66020936,0.784706,0.9016574,0.9393836,0.90920264,0.9393836,0.95824677,0.91297525,0.7884786,0.8337501,0.84884065,0.62625575,0.23390275,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.05281675,0.06413463,0.056589376,0.15467763,0.17354076,0.30181,0.573439,0.97710985,1.4600059,1.659955,1.8146327,1.9127209,1.9579924,1.9504471,1.8863125,1.7882242,1.7467253,1.8221779,2.0145817,2.0636258,1.7882242,1.5015048,1.3204187,1.1544232,1.0374719,0.8903395,0.7054809,0.52439487,0.452715,0.4979865,0.52062225,0.52062225,0.5055317,0.46026024,0.38480774,0.31312788,0.22258487,0.116951376,0.049044125,0.011317875,0.0,0.0,0.00754525,0.041498873,0.06790725,0.0452715,0.06413463,0.1358145,0.18485862,0.124496624,0.060362,0.018863125,0.02263575,0.071679875,0.03772625,0.011317875,0.0150905,0.05281675,0.120724,0.19240387,0.150905,0.0754525,0.026408374,0.02263575,0.026408374,0.0452715,0.07922512,0.090543,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.03772625,0.071679875,0.07922512,0.0754525,0.0754525,0.08299775,0.090543,0.11317875,0.17354076,0.24522063,0.29803738,0.32444575,0.362172,0.4979865,0.362172,0.23767537,0.17731337,0.1961765,0.30181,0.4640329,0.5772116,0.63002837,0.80734175,1.4826416,1.9164935,1.8900851,2.2409391,3.5047686,5.915476,6.485142,6.6360474,6.2814207,5.5759397,4.8930945,4.0291634,3.610402,2.938875,1.9693103,1.3166461,0.8337501,0.6413463,0.7092535,0.965792,1.3166461,1.1921495,1.0487897,0.8224323,0.56589377,0.43007925,0.39989826,0.573439,0.8526133,1.1016065,1.1431054,1.3505998,1.3845534,1.177059,0.9016574,0.9808825,1.2449663,2.1843498,3.0860074,3.4481792,2.9954643,3.0897799,2.4484336,1.7391801,1.3317367,1.3166461,1.7278622,2.0636258,2.0183544,1.7655885,1.9730829,1.6109109,0.98465514,0.4678055,0.22258487,0.19994913,0.19240387,0.150905,0.1056335,0.071679875,0.056589376,0.09808825,0.090543,0.09808825,0.120724,0.09808825,0.10186087,0.13958712,0.18485862,0.18863125,0.120724,0.20372175,0.3169005,0.38858038,0.38480774,0.3055826,0.20749438,0.2565385,0.34330887,0.44894236,0.6375736,0.754525,0.7130261,0.6790725,0.6752999,0.6073926,0.513077,0.41121614,0.3055826,0.2565385,0.35839936,0.5017591,0.5885295,0.5319401,0.392353,0.35839936,0.33953625,0.28294688,0.30181,0.4640329,0.7922512,1.0223814,0.9620194,0.8262049,0.7582976,0.8111144,0.965792,1.1393328,1.3543724,1.6071383,1.8749946,2.0296721,2.1654868,2.2673476,2.3616633,2.516341,3.127506,3.5236318,3.8858037,4.244203,4.478106,4.8100967,5.3194013,6.066381,6.9869013,7.8961043,8.311093,8.103599,7.9791017,8.718536,11.204697,14.27184,16.708956,17.904879,17.25976,14.200161,12.00072,10.106862,9.042982,9.273112,11.204697,12.792972,13.52486,13.060828,11.438599,9.103344,9.110889,8.239413,7.405663,7.0812173,7.3075747,6.436098,7.375482,8.669493,9.4013815,9.1976595,8.782671,8.75249,9.971047,12.626976,16.252468,20.089228,22.03213,22.884743,23.1941,23.277096,21.881226,19.508244,17.30503,15.916705,15.467763,15.24895,13.7700815,11.925267,10.521852,10.253995,11.427281,12.185578,11.8045435,10.427535,9.084481,7.914967,6.828451,5.847569,5.028909,4.4743333,4.6026025,4.504514,4.1989317,3.7084904,3.059599,2.9011486,3.0633714,3.2670932,3.5047686,4.0291634,3.270866,1.9202662,0.86770374,0.41121614,0.2565385,0.120724,0.10186087,0.12826926,0.16976812,0.23013012,0.27917424,0.30935526,0.35462674,0.40367088,0.39989826,0.41121614,0.4678055,0.5696664,0.6752999,0.7092535,0.69793564,0.7696155,0.97710985,1.2789198,1.5279131,1.6033657,1.7165444,1.7580433,1.690136,1.5241405,1.3392819,1.4335974,1.7919968,2.11267,1.8184053,1.3468271,1.0940613,1.0487897,1.1846043,1.4449154,1.7618159,2.5804756,4.515832,7.654656,11.559323,13.845533,15.690348,17.354074,18.5085,18.229324,17.150352,16.765545,16.573141,16.286423,15.848798,16.188334,15.422491,14.034165,12.706201,12.291212,12.619431,13.52486,13.664448,13.102326,13.298503,13.58145,13.422999,13.204187,13.196642,13.570132,14.800008,16.275105,18.221779,20.375948,21.983086,23.635496,25.348267,27.283625,29.06053,29.769783,29.06053,28.373913,27.37794,26.076384,24.827644,25.159636,24.371157,23.1526,21.934042,20.904116,20.300495,20.032639,19.161163,17.463482,15.46399,14.305794,13.290957,12.083718,10.838752,10.201178,9.880505,9.390063,8.892077,8.311093,7.3377557,6.670001,7.062354,6.802043,5.723072,5.2062225,5.330719,5.300538,5.1458607,5.0553174,5.372218,5.353355,5.311856,5.330719,5.3759904,5.2779026,5.847569,6.417235,7.1566696,8.035691,8.797762,8.741172,8.371455,7.9451485,7.598067,7.333983,6.9982195,6.7077274,6.5643673,6.537959,6.462507,3.4179983,2.9426475,2.5767028,2.1843498,1.750498,1.358145,1.6146835,2.5012503,3.5651307,4.172523,3.5236318,2.305074,1.8523588,1.81086,1.901403,1.9391292,2.7200627,3.5839937,4.304565,4.9723196,5.9984736,9.012801,10.370946,11.457462,12.608112,13.106099,12.925014,12.079946,11.442371,10.744436,8.620448,7.7904706,7.352846,6.9944468,6.587003,6.2097406,6.0286546,5.8702044,5.583485,5.111907,4.5007415,3.7688525,3.5123138,3.4594972,3.6783094,4.5912848,4.7044635,3.9876647,3.7198083,4.217795,4.851596,4.315883,3.5500402,3.218049,4.0178456,6.670001,12.672247,12.811834,11.476325,10.714255,10.238904,9.763554,10.220041,10.299266,8.922258,5.247721,6.541732,8.424272,9.574923,9.22784,7.141579,6.651138,6.4134626,6.1606965,5.798525,5.372218,5.198677,5.855114,6.590776,7.281166,8.394091,9.224068,9.733373,9.74469,8.82417,6.270103,7.1264887,8.677037,9.639057,9.307066,7.537705,4.8402777,3.1312788,2.5578396,2.546522,1.7995421,1.2034674,0.9507015,1.0374719,1.5807298,2.837014,5.0477724,6.7454534,7.2396674,6.356873,4.4403796,2.6446102,2.214531,2.0070364,1.6260014,1.418507,1.4071891,1.3845534,0.9808825,0.33953625,0.1056335,0.20372175,0.23013012,0.19240387,0.14335975,0.1659955,0.14335975,0.08299775,0.041498873,0.16222288,0.68661773,1.297783,1.0827434,0.91297525,1.0525624,1.1732863,1.4298248,1.4411428,1.1280149,0.6488915,0.38103512,0.392353,0.241448,0.094315626,0.030181,0.030181,0.041498873,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.03772625,0.0,0.0,0.19240387,0.51684964,0.76584285,0.59607476,0.4979865,0.9318384,1.388326,1.50905,1.0676528,1.1053791,0.6828451,0.29803738,0.21503963,0.47157812,0.98465514,1.3505998,1.4147344,1.3430545,1.6486372,1.8070874,1.9730829,2.0900342,2.0636258,1.7693611,1.7089992,1.418507,1.2487389,1.3468271,1.6637276,2.04099,2.4031622,2.2484846,1.6260014,1.1129243,0.8224323,0.7092535,0.76584285,0.9507015,1.20724,0.7054809,0.6149379,0.72811663,0.86770374,0.91674787,0.7582976,0.73566186,0.6790725,0.52062225,0.27540162,0.21503963,0.32821837,0.331991,0.16976812,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14713238,0.071679875,0.0,0.0,0.0,0.0,0.0,0.06790725,0.181086,0.23013012,0.1659955,0.2263575,0.5055317,1.056335,1.8599042,2.4823873,2.674791,2.7804246,2.927557,3.0369632,2.8181508,2.7426984,2.625747,2.4899325,2.5616124,2.6597006,2.2371666,1.81086,1.5920477,1.4939595,1.1544232,0.965792,0.845068,0.7432071,0.67152727,0.66020936,0.59230214,0.5357128,0.47157812,0.29049212,0.20372175,0.21881226,0.14713238,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.02263575,0.00754525,0.0,0.00754525,0.0452715,0.1659955,0.116951376,0.041498873,0.011317875,0.0,0.011317875,0.071679875,0.16222288,0.21503963,0.090543,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.00754525,0.02263575,0.026408374,0.0150905,0.0150905,0.041498873,0.08677038,0.150905,0.26031113,0.36971724,0.35839936,0.2678564,0.181086,0.23013012,0.23013012,0.19240387,0.150905,0.15467763,0.29049212,0.41121614,0.4074435,0.4074435,0.56589377,1.0676528,1.7769064,1.6788181,2.8445592,5.4250345,7.6584287,7.6848373,7.066127,6.8171334,7.567886,9.582467,6.8737226,4.738417,3.4029078,2.8822856,2.9916916,2.4786146,2.1768045,2.335255,2.704972,2.546522,2.2296214,1.9881734,1.4449154,0.7582976,0.62625575,0.663982,0.95447415,1.358145,1.6335466,1.448688,2.2296214,2.052308,1.599593,1.2864652,1.237421,1.4298248,2.3880715,3.399135,3.8254418,3.0822346,2.71629,2.3126192,1.9844007,1.7542707,1.5731846,1.8297231,2.3692086,2.5201135,2.1051247,1.4335974,1.1053791,0.7582976,0.48666862,0.34330887,0.32067314,0.24899325,0.17354076,0.11317875,0.071679875,0.0452715,0.094315626,0.09808825,0.08677038,0.071679875,0.060362,0.071679875,0.094315626,0.11317875,0.1358145,0.18485862,0.2565385,0.4678055,0.754525,0.965792,0.8526133,0.41498876,0.1961765,0.1659955,0.28294688,0.5017591,0.5998474,0.6073926,0.7167987,0.8865669,0.83752275,0.52062225,0.4074435,0.34330887,0.26408374,0.150905,0.12826926,0.120724,0.13958712,0.18485862,0.26031113,0.36971724,0.43385187,0.573439,0.83752275,1.20724,1.2902378,1.1204696,0.9620194,0.90920264,0.8865669,0.9695646,1.1091517,1.2826926,1.50905,1.8599042,2.252257,2.3956168,2.41448,2.493705,2.8822856,3.531177,3.6745367,3.9008942,4.3686996,4.8063245,4.659192,4.640329,5.2288585,6.368191,7.492433,8.311093,8.82417,9.559832,10.714255,12.193124,14.400109,16.539188,17.112627,16.214743,15.516807,13.79649,12.736382,11.121698,9.922004,12.253486,10.872705,11.408418,12.268577,12.034674,9.446653,8.458225,7.624475,6.719045,5.904158,5.723072,4.67051,5.2967653,6.7680893,7.964011,7.4773426,7.1604424,7.6395655,9.084481,11.393328,14.173752,17.640795,19.368656,20.402355,21.202152,21.666185,21.119154,19.764782,18.376457,17.41821,17.029629,16.18456,14.996184,13.257004,11.449917,10.740664,12.012038,13.200415,13.487134,12.528888,10.453944,8.45068,6.7039547,5.409944,4.6214657,4.2404304,4.1574326,3.9159849,3.482133,2.9766011,2.6710186,3.3915899,4.055572,4.4894238,4.6252384,4.515832,3.5160866,1.7354075,0.5772116,0.35462674,0.3055826,0.10940613,0.071679875,0.08677038,0.1358145,0.24522063,0.27917424,0.27917424,0.2867195,0.32821837,0.41121614,0.362172,0.3772625,0.422534,0.4678055,0.5017591,0.5394854,0.62248313,0.76207024,0.9808825,1.297783,1.8221779,2.191895,2.214531,1.9768555,1.8297231,1.7693611,1.8825399,2.0598533,2.123988,1.8297231,1.3807807,1.1657411,1.086516,1.1053791,1.2525115,1.4109617,1.7429527,2.384299,3.4557245,5.0666356,7.3113475,10.355856,13.600313,16.509007,18.58395,19.538425,20.919205,21.820864,21.967995,21.696367,22.22076,21.711456,19.979822,17.444618,15.135772,14.966003,15.335721,15.603577,15.373446,14.494425,14.385019,14.396337,14.200161,13.875714,13.902123,15.158407,15.939341,17.033401,18.87067,21.53037,23.201643,24.197617,26.125427,29.120892,31.844728,33.27455,32.78034,31.184519,29.358568,28.1966,28.136238,27.223263,25.71044,23.907125,22.186808,21.503962,21.047476,20.225042,18.821627,17.014538,16.01102,14.909414,13.585222,12.264804,11.521597,11.140562,10.963248,10.695392,10.0465,8.726082,8.179051,7.6093845,6.8473144,6.0626082,5.7683434,5.80607,5.987156,6.017337,6.043745,6.6662283,6.4738245,5.7570257,5.3646727,5.511805,5.7683434,5.534441,5.7796617,6.3342376,7.0774446,7.91874,8.16396,7.9225125,7.3868,6.771862,6.3342376,6.0626082,5.8136153,5.587258,5.3609,5.081726,2.5993385,2.5616124,2.1881225,1.7731338,1.5467763,1.6637276,1.9278114,2.233394,2.5767028,2.8219235,2.6823363,2.0183544,1.9768555,2.2673476,2.535204,2.3654358,2.305074,2.4182527,2.8709676,3.7763977,5.20245,6.9189944,8.114917,8.692128,9.129752,10.457717,13.671993,16.16947,17.165443,16.343012,13.856852,12.2270775,10.895341,9.891823,9.035437,7.9451485,6.7341356,6.360646,5.8173876,4.957229,4.4516973,4.327201,4.432834,4.606375,4.8629136,5.3986263,5.1458607,4.8553686,4.67051,4.6214657,4.6327834,5.032682,4.7572803,5.1232247,6.7152724,9.4127,11.514051,10.242677,8.541223,8.031919,9.031664,9.49947,10.480352,11.646093,12.400619,11.902632,8.194141,7.2962565,7.8244243,8.631766,8.801534,7.9225125,6.7341356,6.25124,6.549277,6.7869525,6.488915,6.3342376,6.4247804,6.579458,6.3531003,6.7944975,6.560595,6.749226,7.7225633,9.125979,9.914458,10.899114,11.348056,10.846297,9.26934,7.032173,5.300538,3.4594972,2.0447628,2.71629,3.1916409,3.2633207,3.0407357,2.897376,3.4594972,5.80607,5.847569,5.300538,4.859141,4.172523,2.9728284,2.0636258,1.7429527,1.7165444,1.0902886,0.754525,0.6149379,0.5055317,0.36971724,0.25276586,0.26408374,0.30181,0.29803738,0.23767537,0.15467763,0.090543,0.07922512,0.10940613,0.20749438,0.41876137,0.52062225,0.41498876,0.422534,0.66775465,1.0638802,1.0676528,0.9922004,0.8224323,0.59230214,0.38103512,0.23767537,0.09808825,0.05281675,0.12826926,0.27540162,0.181086,0.181086,0.120724,0.011317875,0.0,0.0,0.00754525,0.018863125,0.026408374,0.03772625,0.0452715,0.026408374,0.00754525,0.0,0.0,0.018863125,0.08299775,0.1358145,0.1961765,0.35462674,0.34330887,1.1280149,2.7804246,3.6971724,0.6073926,0.44139713,0.7922512,1.297783,1.6675003,1.6675003,1.2449663,0.80356914,0.452715,0.29803738,0.4376245,0.724344,0.9695646,1.2110126,1.3920987,1.3543724,2.0296721,2.123988,1.7919968,1.3468271,1.2713746,1.1317875,1.0412445,1.0714256,1.2638294,1.6373192,2.0673985,2.2258487,1.991946,1.478869,1.0638802,0.8111144,0.76207024,0.84129536,0.875249,0.58475685,0.5885295,0.97333723,1.2940104,1.3128735,0.9997456,0.6752999,0.80356914,0.95447415,0.8639311,0.44516975,0.15845025,0.08299775,0.06790725,0.033953626,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0150905,0.03772625,0.0452715,0.033953626,0.22258487,0.5017591,0.95447415,1.8372684,2.4899325,2.6974268,2.6785638,2.584248,2.5012503,2.3390274,2.3956168,2.3578906,2.1805773,2.0862615,1.9881734,1.7580433,1.5505489,1.3845534,1.1431054,0.91674787,0.7507524,0.63002837,0.52062225,0.392353,0.271629,0.19240387,0.14713238,0.11317875,0.056589376,0.041498873,0.0452715,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.00754525,0.041498873,0.026408374,0.0150905,0.018863125,0.03772625,0.06790725,0.16222288,0.18485862,0.11317875,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.02263575,0.0150905,0.0150905,0.030181,0.0452715,0.0150905,0.026408374,0.06413463,0.10186087,0.116951376,0.10186087,0.094315626,0.1358145,0.1659955,0.17354076,0.20372175,0.22258487,0.21503963,0.2263575,0.29426476,0.44894236,0.5885295,0.6187105,0.6375736,0.84884065,1.5430037,1.267602,1.8599042,3.1727777,4.6856003,5.511805,4.9421387,5.081726,6.3153744,8.356364,10.242677,9.016574,6.9227667,5.1835866,4.6252384,5.7117543,4.6931453,3.942393,3.3953626,3.0709167,3.048281,2.8181508,2.3390274,1.7014539,1.0902886,0.80734175,0.77716076,0.90543,1.5279131,2.3465726,2.425798,2.4559789,2.1013522,1.7919968,1.7542707,2.0183544,1.1883769,1.6675003,2.6446102,3.440634,3.4972234,2.7125173,2.4371157,2.425798,2.6295197,3.2067313,2.7125173,1.8636768,1.1657411,0.79602385,0.60362,0.77338815,0.77716076,0.7092535,0.6149379,0.49044126,0.25276586,0.15845025,0.116951376,0.08677038,0.08299775,0.10186087,0.1056335,0.094315626,0.08299775,0.10940613,0.10186087,0.09808825,0.10186087,0.120724,0.16976812,0.28294688,0.36594462,0.41121614,0.42630664,0.41498876,0.32821837,0.20372175,0.15845025,0.211267,0.29426476,0.38480774,0.452715,0.5093044,0.52062225,0.41121614,0.33953625,0.32821837,0.32067314,0.29049212,0.24899325,0.24522063,0.18485862,0.13958712,0.15845025,0.26031113,0.4074435,0.513077,0.6073926,0.7205714,0.8526133,1.0638802,1.056335,0.9997456,1.0035182,1.116697,1.0638802,1.1506506,1.2638294,1.4109617,1.7165444,2.252257,2.6597006,2.9615107,3.2482302,3.6783094,3.8254418,3.772625,3.8669407,4.346064,5.330719,5.704209,5.8588867,6.349328,7.1566696,7.673519,7.9451485,8.684583,9.2844305,9.793735,10.899114,12.600568,14.102073,15.0376835,15.618668,16.641048,15.83748,14.075664,11.706455,9.473062,8.492179,8.314865,9.34102,10.140816,9.944639,8.627994,9.239159,10.461489,9.627739,7.224577,6.8925858,6.2625575,5.828706,5.541986,5.4967146,5.926794,5.5985756,7.1906233,9.5183325,11.725319,13.2607765,14.694374,16.550507,18.331184,19.583696,19.908142,19.429018,19.451654,19.885506,19.998686,18.45568,16.746683,15.433809,14.196388,13.053283,12.366665,13.400364,14.339747,14.32843,13.189097,11.415963,9.578695,8.16396,7.462252,7.194396,6.462507,5.624984,4.6931453,3.8593953,3.2444575,2.8898308,2.9841464,3.4142256,3.7688525,3.742444,3.1237335,1.9768555,0.83752275,0.26031113,0.23767537,0.16976812,0.094315626,0.08299775,0.10940613,0.16222288,0.23013012,0.2867195,0.29426476,0.30935526,0.35462674,0.41121614,0.43007925,0.45648763,0.49044126,0.513077,0.49044126,0.44894236,0.44516975,0.5055317,0.633801,0.845068,1.2638294,1.6033657,1.8070874,1.8787673,1.9278114,1.9655377,2.0749438,2.1466236,2.1353056,2.0372176,2.0372176,1.9202662,1.6976813,1.4901869,1.5203679,1.5618668,1.7052265,2.033445,2.5767028,3.31991,3.9348478,5.221313,7.541477,10.61994,13.543724,16.361876,19.579924,22.53389,24.959686,26.996904,27.891016,27.60807,26.09902,23.85808,21.911406,21.175745,19.964731,18.621677,17.286167,15.897841,14.177525,13.762536,13.615403,13.392818,13.43809,13.962485,14.822643,15.939341,17.335213,19.127209,22.311304,24.650331,26.536644,28.347504,30.45263,33.433002,36.156837,36.371876,34.085667,31.531599,29.856554,28.14001,26.495146,24.929506,23.333685,21.967995,20.915434,20.04773,19.372429,19.040438,17.844517,16.803272,15.70921,14.532151,13.43809,12.626976,11.91395,11.427281,11.046246,10.352083,9.4013815,9.020347,9.009028,8.812852,7.5263867,6.9567204,6.5341864,6.258785,6.1418333,6.228604,5.945657,5.983383,6.33801,6.6549106,6.205968,5.8966126,6.0701537,6.307829,6.72659,7.967784,8.171506,8.126234,7.835742,7.3490734,6.771862,6.375736,6.0211096,5.624984,5.168496,4.689373,2.3126192,2.2560298,2.0787163,1.9730829,1.9164935,1.6373192,1.7316349,1.8146327,1.8976303,1.9655377,1.9579924,1.7995421,1.9466745,2.7502437,3.783943,3.8367596,3.451952,3.3350005,3.1124156,3.1765501,4.6554193,5.2779026,6.1305156,7.183078,8.541223,10.435081,11.536687,13.773854,15.328176,15.365902,14.04171,13.083464,13.58145,13.577678,12.566614,11.506506,9.993684,8.654402,7.2358947,6.0211096,5.832478,5.2326307,4.5799665,4.3385186,4.719554,5.674028,5.2665844,4.991183,4.8629136,4.9949555,5.6023483,6.609639,7.039718,7.779153,8.771353,9.012801,7.6886096,6.1078796,5.2892203,5.4476705,5.9720654,6.960493,7.7150183,9.133525,11.431054,14.177525,13.645585,10.103089,7.805561,7.9526935,8.684583,8.213005,6.820906,5.3269467,4.538468,5.2552667,5.1458607,5.1798143,5.4438977,5.753253,5.613666,4.9987283,5.300538,5.5457587,5.59103,6.126743,6.579458,7.2170315,7.183078,6.519096,6.1342883,4.919503,4.5196047,4.4101987,4.221567,3.7613072,3.429316,3.2105038,2.9313297,2.6106565,2.444661,3.0520537,2.9426475,2.6936543,2.6144292,2.7389257,2.3956168,1.8825399,1.6260014,1.478869,0.724344,0.46026024,0.331991,0.271629,0.23013012,0.18863125,0.271629,0.40367088,0.3961256,0.241448,0.124496624,0.094315626,0.090543,0.1056335,0.14713238,0.23013012,0.19994913,0.21881226,0.36971724,0.633801,0.9016574,1.1544232,1.1091517,0.875249,0.58098423,0.3734899,0.21881226,0.10940613,0.09808825,0.16222288,0.20749438,0.120724,0.09808825,0.060362,0.003772625,0.0,0.0,0.003772625,0.00754525,0.0150905,0.018863125,0.02263575,0.13958712,0.19240387,0.13204187,0.0452715,0.018863125,0.041498873,0.06413463,0.16222288,0.52439487,0.513077,0.9922004,1.931584,2.3503454,0.3169005,0.875249,1.1695137,1.3656902,1.50905,1.5241405,1.116697,0.935611,0.7696155,0.59230214,0.56589377,0.62248313,0.73566186,1.0110635,1.4034165,1.720317,2.0372176,2.1579416,2.1202152,2.003264,1.9051756,1.2638294,1.0035182,0.98465514,1.146878,1.5316857,1.9353566,1.931584,1.7014539,1.3694628,1.0148361,0.77338815,0.66775465,0.65643674,0.633801,0.41876137,0.6187105,0.8978847,1.0940613,1.0978339,0.8563859,0.44139713,0.5319401,1.478869,2.4786146,1.569412,0.51684964,0.26031113,0.15845025,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.2263575,0.47157812,0.9695646,1.3505998,1.4939595,1.4864142,1.4147344,1.3317367,1.2940104,1.3355093,1.3204187,1.2298758,1.1619685,1.0751982,0.965792,0.8601585,0.7507524,0.58475685,0.4640329,0.35462674,0.28294688,0.22258487,0.12826926,0.06790725,0.03772625,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.00754525,0.018863125,0.06790725,0.10186087,0.08677038,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.02263575,0.00754525,0.00754525,0.018863125,0.026408374,0.00754525,0.049044125,0.120724,0.18863125,0.1961765,0.09808825,0.060362,0.09808825,0.14713238,0.16222288,0.14335975,0.14713238,0.124496624,0.124496624,0.17354076,0.29426476,0.45648763,0.4376245,0.45648763,0.6488915,1.0487897,1.7467253,2.9916916,3.8707132,4.1197066,4.104616,3.802806,4.0404816,5.1458607,6.9189944,8.650629,8.114917,7.322665,6.677546,6.5945487,7.492433,7.9715567,8.567632,7.496206,5.5759397,6.2323766,5.847569,4.5309224,2.957738,1.9391292,2.4182527,1.991946,1.8184053,1.9504471,2.1805773,2.0485353,1.931584,2.173032,2.1768045,1.8372684,1.5354583,1.0412445,1.6335466,2.8936033,4.044254,3.9499383,3.3651814,3.1425967,3.006782,2.8256962,2.5917933,1.6448646,0.9620194,0.543258,0.33576363,0.27917424,0.46026024,0.70170826,1.0601076,1.2789198,0.77338815,0.3734899,0.18863125,0.116951376,0.1056335,0.120724,0.116951376,0.120724,0.12826926,0.14713238,0.20372175,0.271629,0.2263575,0.18863125,0.21503963,0.2867195,0.36594462,0.3734899,0.33576363,0.29426476,0.31312788,0.32067314,0.271629,0.23013012,0.2263575,0.24522063,0.38103512,0.43007925,0.44894236,0.46026024,0.44139713,0.452715,0.47157812,0.4640329,0.42630664,0.40367088,0.36594462,0.28294688,0.21881226,0.2263575,0.35085413,0.6187105,0.72811663,0.7205714,0.66020936,0.6149379,0.72811663,0.77716076,0.90920264,1.1129243,1.237421,1.2940104,1.3694628,1.3920987,1.4449154,1.7882242,2.3314822,2.8709676,3.289729,3.5500402,3.682082,3.9650288,3.821669,3.8593953,4.406426,5.5080323,6.2889657,6.643593,7.322665,8.280911,8.692128,9.148616,9.65792,9.876732,10.050273,11.050018,11.864905,12.909923,13.932304,14.822643,15.62244,15.098045,14.7170105,13.015556,10.465261,9.484379,9.593785,9.737145,9.914458,9.8239155,8.854351,10.465261,11.121698,10.042727,8.141325,8.039464,6.9869013,5.9418845,5.036454,4.6214657,5.27413,5.7419353,6.3908267,8.239413,10.8576145,12.362892,13.106099,14.505743,16.38451,18.221779,19.15739,18.504726,19.17248,20.209951,20.655123,19.519562,17.889788,16.780636,15.8676605,14.9358225,13.879487,14.117163,14.871688,15.192361,14.66042,13.396591,11.310329,10.008774,9.563604,9.540969,9.016574,7.3679366,5.9607477,4.957229,4.353609,3.9876647,3.62172,3.2218218,2.71629,2.1202152,1.5128226,0.8563859,0.38103512,0.22258487,0.2678564,0.12826926,0.10186087,0.1056335,0.12826926,0.1659955,0.21881226,0.27917424,0.33576363,0.38103512,0.41121614,0.43007925,0.4979865,0.573439,0.59230214,0.543258,0.4979865,0.4376245,0.39989826,0.4074435,0.47157812,0.59607476,0.8601585,1.1883769,1.4071891,1.4977322,1.5958204,1.8259505,2.1541688,2.372981,2.463524,2.6219745,3.0671442,3.2633207,3.0633714,2.6295197,2.4371157,2.0108092,1.8523588,1.901403,2.093807,2.3616633,2.5993385,3.1463692,4.357382,6.25124,8.529905,11.570641,15.264041,19.304522,23.38273,27.211945,28.71345,28.822855,27.811792,26.193335,24.714466,23.665676,22.028357,20.081682,18.082191,16.260014,14.750964,14.520834,14.494425,14.422746,14.86037,15.252723,15.79598,16.497688,17.391802,18.534906,22.699884,25.54067,27.389257,28.807764,30.607307,33.764996,36.50769,37.52253,36.503918,34.149803,31.633461,29.63397,28.109829,26.891272,25.642532,24.054256,22.582933,21.307787,20.326904,19.783646,19.719511,19.266796,18.161417,16.516552,14.841507,13.845533,12.58925,11.846043,11.676274,11.427281,11.415963,11.619685,11.446144,10.450171,8.348819,7.5716586,6.964266,6.609639,6.488915,6.511551,5.994701,6.5228686,6.9491754,6.741681,5.9796104,5.560849,5.594803,5.745708,6.006019,6.688864,6.9152217,7.039718,7.01331,6.8246784,6.515323,6.25124,5.9418845,5.5495315,5.0741806,4.564876,2.1164427,1.8184053,1.8523588,2.0749438,2.1994405,1.8146327,1.6637276,1.7580433,1.7919968,1.780679,2.0636258,2.052308,2.082489,2.9426475,4.2517486,4.459243,4.247976,4.195159,3.8367596,3.5990841,4.7912335,5.7494807,6.2889657,7.032173,8.262049,9.929549,9.359882,9.714509,10.79348,11.747954,11.076427,11.521597,13.792717,15.199906,14.656648,12.668475,11.419736,9.525878,7.665974,6.511551,6.722818,6.470052,5.5382137,4.930821,5.1043615,5.9305663,5.2665844,4.353609,3.9122121,4.6214657,7.111398,8.367682,8.718536,8.820397,8.786444,8.16396,6.952948,6.039973,5.9003854,6.356873,6.5945487,7.3717093,7.201941,7.986647,10.533169,14.539697,15.754482,11.936585,8.620448,8.088508,9.386291,9.307066,7.635793,5.3458095,3.7198083,4.346064,4.504514,4.432834,4.496969,4.745962,4.908185,4.236658,4.666737,4.8402777,4.432834,4.1612053,4.036709,4.1310244,3.953711,3.6254926,3.874486,3.4934506,3.7613072,4.7044635,5.772116,5.836251,5.8702044,4.9345937,3.8405323,2.9124665,2.0372176,1.3166461,1.1393328,1.1317875,1.1544232,1.3241913,1.358145,1.2449663,1.116697,0.9280658,0.4678055,0.33576363,0.23390275,0.16976812,0.15845025,0.18863125,0.33576363,0.5357128,0.6073926,0.4979865,0.27917424,0.1659955,0.120724,0.13958712,0.17731337,0.14713238,0.15467763,0.2678564,0.44516975,0.60362,0.65643674,1.0186088,1.0072908,0.7884786,0.513077,0.3470815,0.19994913,0.124496624,0.124496624,0.1659955,0.18863125,0.124496624,0.056589376,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.124496624,0.1961765,0.150905,0.056589376,0.011317875,0.0,0.0,0.071679875,0.35839936,0.45648763,0.62248313,0.9280658,1.2940104,1.50905,1.8749946,2.0862615,2.0447628,1.7618159,1.3807807,0.9997456,0.94692886,1.0223814,1.0525624,0.8865669,0.7092535,0.66775465,0.84884065,1.2487389,1.7580433,1.8372684,1.9881734,2.2220762,2.3465726,1.9730829,1.2751472,0.9620194,0.88279426,0.97710985,1.2638294,1.5731846,1.5807298,1.4335974,1.2110126,0.9318384,0.7205714,0.5885295,0.513077,0.46026024,0.38103512,0.513077,0.58475685,0.6375736,0.65643674,0.56589377,0.2263575,0.22258487,1.1280149,2.2560298,1.6788181,0.7092535,0.47912338,0.35839936,0.14335975,0.056589376,0.060362,0.0754525,0.0754525,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026408374,0.09808825,0.23767537,0.35462674,0.41121614,0.42630664,0.422534,0.43385187,0.4376245,0.4376245,0.43007925,0.41498876,0.39989826,0.36971724,0.32821837,0.27917424,0.2263575,0.1659955,0.120724,0.0754525,0.05281675,0.041498873,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.003772625,0.003772625,0.018863125,0.026408374,0.030181,0.026408374,0.02263575,0.018863125,0.03772625,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.00754525,0.0,0.0,0.00754525,0.0150905,0.011317875,0.05281675,0.13204187,0.211267,0.241448,0.150905,0.09808825,0.10940613,0.13958712,0.150905,0.10186087,0.07922512,0.05281675,0.0452715,0.0754525,0.14335975,0.23767537,0.21503963,0.32821837,0.6526641,1.0940613,2.3428001,3.1652324,3.380272,3.2444575,3.4444065,3.5953116,3.6783094,4.1612053,5.198677,6.617184,6.6662283,6.5643673,6.417235,6.5228686,7.3868,9.714509,10.989656,9.616421,6.832224,6.72659,6.56814,6.047518,4.6931453,3.2218218,3.5123138,2.8030603,2.3277097,1.9881734,1.7844516,1.81086,1.9164935,2.4899325,2.6295197,2.0749438,1.1732863,1.2298758,2.2748928,3.731126,4.8327327,4.640329,4.221567,3.7763977,3.0218725,2.052308,1.3468271,0.6149379,0.41121614,0.3772625,0.3169005,0.20372175,0.241448,0.46026024,0.9242931,1.327964,0.965792,0.59230214,0.32444575,0.19994913,0.181086,0.1659955,0.1358145,0.116951376,0.11317875,0.1358145,0.181086,0.2678564,0.24522063,0.23013012,0.271629,0.32821837,0.3734899,0.3734899,0.35085413,0.3470815,0.41121614,0.47157812,0.43385187,0.45648763,0.52062225,0.422534,0.46026024,0.482896,0.5394854,0.62248313,0.6752999,0.6752999,0.663982,0.62625575,0.5696664,0.5357128,0.5394854,0.4678055,0.40367088,0.41121614,0.51684964,0.73188925,0.77338815,0.73188925,0.66775465,0.63002837,0.6488915,0.663982,0.8526133,1.1808317,1.3920987,1.6637276,1.7919968,1.8561316,1.9994912,2.3880715,2.897376,3.3576362,3.7386713,4.006528,4.1272516,4.538468,4.459243,4.4705606,4.9534564,6.1116524,6.760544,6.9265394,7.3000293,7.9715567,8.409182,8.892077,8.918486,8.993938,9.57115,11.031156,12.200669,12.879742,13.690856,14.468017,14.230342,13.792717,14.422746,14.124708,12.6345215,11.431054,11.544232,11.129244,10.70671,10.340765,9.654147,10.582213,10.137043,8.797762,7.3905725,7.1000805,6.3945994,6.1342883,5.594803,5.0666356,5.8664317,6.436098,6.0739264,6.9454026,9.359882,11.77059,12.411936,13.35132,14.905642,16.859861,18.45568,18.632996,18.893307,19.33093,19.700647,19.413929,18.719765,18.376457,17.938831,17.074902,15.539442,15.049001,15.607349,16.32792,16.569368,15.961976,13.068373,11.16697,10.235131,9.895596,9.424017,7.7301087,6.4964604,5.7117543,5.2062225,4.666737,3.9612563,3.1425967,2.2711203,1.4335974,0.7394345,0.36594462,0.20372175,0.1961765,0.2263575,0.10940613,0.116951376,0.13958712,0.1659955,0.1961765,0.24522063,0.29426476,0.35839936,0.4074435,0.43007925,0.422534,0.5017591,0.58098423,0.5696664,0.482896,0.44139713,0.41121614,0.38858038,0.392353,0.43007925,0.5093044,0.6488915,0.875249,1.0110635,1.0487897,1.1317875,1.6146835,2.3805263,3.0520537,3.5047686,3.8707132,4.1498876,4.402653,4.29702,3.8103511,3.2482302,2.6408374,2.1843498,1.9278114,1.8825399,2.0070364,2.3918443,2.8106055,3.3312278,4.08198,5.2628117,7.424526,10.567122,14.690601,19.398838,23.903353,27.061039,29.271797,30.188545,29.532108,27.094994,24.137255,22.130219,20.602304,19.349794,18.45568,17.852062,17.286167,16.791954,16.542961,16.867407,16.848543,16.84477,17.169216,18.078419,19.753464,22.737612,25.144547,27.260988,29.222754,31.007204,33.97249,36.45865,38.12992,38.499638,36.88873,33.953625,31.542917,29.784874,28.558771,27.517527,26.276333,25.069094,23.854307,22.590479,21.266287,21.28515,20.95316,19.945868,18.35382,16.690092,15.267814,13.747445,12.83447,12.653384,12.751472,13.000465,12.932558,12.23085,10.823661,8.869441,8.14887,7.575431,7.2170315,7.0812173,7.115171,7.1566696,7.2924843,7.01331,6.247467,5.3986263,5.040227,5.0175915,5.1269975,5.2590394,5.3910813,5.5457587,5.696664,5.794752,5.8211603,5.794752,5.7683434,5.613666,5.3344917,4.949684,4.496969,2.003264,1.6637276,1.8825399,2.2220762,2.3880715,2.2447119,1.8334957,1.9542197,2.0372176,2.0900342,2.674791,2.625747,2.4522061,2.8407867,3.6292653,3.8103511,4.0291634,4.146115,4.195159,4.3913355,5.13077,7.0887623,7.484888,7.2358947,7.17176,8.009283,7.99042,6.8699503,7.0774446,8.390318,7.9451485,9.684328,11.993175,13.6833105,13.547497,10.370946,9.616421,8.307321,7.118943,6.579458,7.0510364,7.6395655,7.001992,6.319147,6.0739264,6.0626082,4.9421387,3.2633207,2.425798,3.5764484,7.598067,9.714509,9.325929,7.91874,6.8058157,7.092535,8.756263,9.220296,9.461743,9.891823,10.378491,10.416218,9.514561,9.7069645,11.668729,14.698147,13.52486,10.955703,8.639311,7.956466,10.020092,10.423763,8.805306,6.719045,5.323174,5.3571277,5.583485,4.983638,4.349837,4.0517993,4.025391,4.085753,3.9386206,3.9310753,4.146115,4.3800178,3.8480775,3.482133,3.5349495,3.874486,3.983892,3.9159849,3.8707132,4.247976,5.3571277,7.413208,9.167479,8.167733,6.205968,4.3724723,3.0331905,1.9768555,1.2826926,0.94692886,0.7997965,0.5357128,0.44516975,0.4074435,0.3734899,0.33953625,0.32821837,0.2678564,0.17354076,0.13958712,0.181086,0.26408374,0.392353,0.5696664,0.7469798,0.7922512,0.47157812,0.32821837,0.28294688,0.32067314,0.34330887,0.18485862,0.2565385,0.38103512,0.47535074,0.5017591,0.46026024,0.62625575,0.6111652,0.5017591,0.3772625,0.3055826,0.14335975,0.13204187,0.13958712,0.14713238,0.26408374,0.23013012,0.20372175,0.181086,0.13204187,0.00754525,0.00754525,0.003772625,0.003772625,0.003772625,0.0150905,0.026408374,0.02263575,0.060362,0.150905,0.26408374,0.211267,0.08677038,0.018863125,0.03772625,0.071679875,0.34330887,0.5470306,0.9393836,1.7391801,3.138824,2.5616124,2.704972,2.6936543,2.2183034,1.5128226,1.0940613,0.9507015,1.146878,1.4071891,1.1242423,0.7922512,0.65643674,0.7507524,1.0299267,1.3807807,1.6448646,1.780679,1.9579924,1.9994912,1.4147344,1.0902886,0.91297525,0.84129536,0.8526133,0.965792,1.1317875,1.2449663,1.2147852,1.0487897,0.8337501,0.6790725,0.58098423,0.5055317,0.43385187,0.34330887,0.31312788,0.33576363,0.4074435,0.49044126,0.5055317,0.2867195,0.124496624,0.13958712,0.33953625,0.633801,0.51684964,0.4640329,0.41121614,0.3169005,0.14335975,0.12826926,0.13958712,0.1358145,0.09808825,0.003772625,0.018863125,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.09808825,0.060362,0.049044125,0.049044125,0.049044125,0.049044125,0.049044125,0.033953626,0.02263575,0.018863125,0.0,0.0,0.0,0.00754525,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.018863125,0.03772625,0.041498873,0.0754525,0.06413463,0.018863125,0.03772625,0.07922512,0.08299775,0.071679875,0.05281675,0.041498873,0.07922512,0.06790725,0.033953626,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.00754525,0.011317875,0.018863125,0.026408374,0.03772625,0.0452715,0.08299775,0.14713238,0.211267,0.20749438,0.124496624,0.116951376,0.13204187,0.1358145,0.090543,0.06790725,0.06413463,0.090543,0.124496624,0.124496624,0.094315626,0.124496624,0.36594462,0.875249,1.6260014,2.3767538,2.123988,1.8674494,2.1768045,3.187868,3.7009451,3.8971217,3.9348478,4.112161,4.8666863,5.3759904,5.1835866,4.9647746,5.198677,6.187105,9.201432,9.835234,8.409182,5.934339,4.0782075,4.274384,5.783434,6.017337,4.715781,3.9574835,3.2218218,2.4710693,1.8485862,1.6033657,2.1013522,2.6068838,3.078462,3.0558262,2.3918443,1.2525115,1.5316857,2.9501927,4.398881,5.2099953,5.1760416,4.376245,3.5387223,2.2673476,0.90920264,0.5583485,0.452715,0.41498876,0.5017591,0.58475685,0.36971724,0.22258487,0.20749438,0.38858038,0.69039035,0.87902164,0.73188925,0.51684964,0.38480774,0.3470815,0.27917424,0.181086,0.10940613,0.0754525,0.071679875,0.071679875,0.10186087,0.15467763,0.23013012,0.29803738,0.2867195,0.30181,0.30935526,0.32821837,0.3772625,0.5017591,0.66020936,0.63002837,0.7394345,0.91674787,0.694163,0.60362,0.62248313,0.73188925,0.8865669,0.9997456,1.0035182,0.91674787,0.80734175,0.724344,0.69793564,0.7997965,0.76584285,0.7130261,0.7092535,0.754525,0.7130261,0.633801,0.6111652,0.6828451,0.8111144,0.9205205,0.9620194,1.1431054,1.4826416,1.8146327,2.2220762,2.4295704,2.516341,2.655928,3.1048703,3.5651307,3.8292143,4.1272516,4.568649,5.160951,5.621211,5.7192993,5.704209,5.9305663,6.862405,6.8359966,6.462507,6.2097406,6.300284,6.72659,7.001992,6.760544,7.1981683,8.805306,11.389555,13.728582,13.86817,13.856852,13.9888935,12.81938,12.483616,12.898605,13.562587,13.551269,11.54046,12.170488,12.698656,12.298758,11.151879,10.453944,9.891823,8.812852,7.333983,5.8588867,5.0741806,5.100589,5.9796104,6.1003346,5.6891184,6.809588,6.8699503,6.277648,6.462507,8.118689,11.204697,11.966766,12.804289,13.928532,15.456445,17.414436,19.063074,18.606586,18.006739,18.101055,18.614132,19.1008,19.493153,19.429018,18.648085,17.006994,16.177015,16.42601,17.195625,17.863379,17.746428,14.32843,11.672502,9.88805,8.778898,7.8508325,6.8133607,6.247467,5.956975,5.6363015,4.8327327,3.7877154,3.0445085,2.4484336,1.7995421,0.875249,0.362172,0.16222288,0.11317875,0.1056335,0.1056335,0.14713238,0.18863125,0.21503963,0.23767537,0.29426476,0.32821837,0.35839936,0.38858038,0.41498876,0.41121614,0.46026024,0.48666862,0.4678055,0.42630664,0.41498876,0.4074435,0.39989826,0.41121614,0.452715,0.52062225,0.5772116,0.6451189,0.68661773,0.7130261,0.7884786,1.4071891,2.6068838,3.8593953,4.7950063,5.198677,4.8742313,4.9421387,4.938366,4.5497856,3.6330378,3.1765501,2.5427492,2.0447628,1.8485862,1.9693103,2.5502944,3.1199608,3.531177,3.783943,4.0593443,4.8742313,6.937857,10.186088,14.222796,18.312323,23.288414,28.588953,32.82561,34.470474,31.856045,26.664913,23.560043,22.213217,22.22076,23.107328,23.16769,21.820864,20.583443,20.160908,20.455173,20.266542,19.685556,19.48561,20.258997,22.401848,23.001694,24.522062,26.86109,29.59247,31.954134,34.587425,37.443302,39.929462,41.129158,39.77101,36.469967,33.383957,30.99966,29.430248,28.430502,27.875927,27.46471,26.898817,25.917934,24.284388,23.05074,22.054766,21.051247,19.97605,18.949896,17.165443,15.569623,14.509516,14.132254,14.407655,14.132254,13.181552,12.091263,11.042474,9.880505,9.325929,8.797762,8.356364,7.997965,7.635793,8.412953,7.7187905,6.6058664,5.6325293,4.8629136,4.666737,4.640329,4.6629643,4.659192,4.6214657,4.644101,4.719554,4.798779,4.878004,4.9760923,5.1458607,5.1798143,5.0553174,4.7874613,4.429062,2.3956168,2.7879698,3.2670932,3.4255435,3.1237335,2.4861598,1.8146327,1.6486372,1.9240388,2.3578906,2.4559789,2.8332415,2.9011486,2.7917426,2.7087448,2.9313297,3.3463185,3.62172,3.7198083,3.8103511,4.2894745,5.1534057,5.6287565,5.6815734,5.594803,5.934339,6.2663302,6.2021956,6.360646,7.141579,8.729855,10.680302,10.767072,9.740918,8.235641,6.7454534,6.156924,6.8737226,7.77538,8.329956,8.575176,7.9526935,6.779407,6.0739264,5.8928404,5.3571277,3.6594462,2.4220252,2.0183544,2.704972,4.610148,10.148361,9.623966,6.802043,4.29702,3.5387223,6.25124,8.375228,9.986138,10.914205,10.7557535,10.220041,10.533169,12.061082,14.245432,15.626213,12.1101265,8.382772,5.515578,4.4894238,6.2097406,8.235641,8.631766,8.322411,7.8319697,7.3075747,7.0774446,6.5530496,5.7079816,4.696918,3.8292143,3.3048196,2.9351022,2.7087448,2.5238862,2.1805773,2.2069857,2.4408884,2.8747404,3.3764994,3.6934,3.4972234,3.5839937,3.5424948,3.5802212,4.5309224,6.670001,8.201687,7.798016,5.915476,4.7912335,3.2670932,1.9504471,1.0902886,0.67152727,0.42630664,0.36594462,0.34330887,0.29803738,0.23013012,0.18485862,0.20749438,0.1659955,0.13204187,0.13204187,0.1659955,0.21503963,0.2565385,0.3169005,0.35085413,0.23013012,0.6187105,0.7884786,0.7582976,0.5885295,0.38103512,0.44139713,0.40367088,0.4074435,0.4979865,0.59607476,0.59607476,0.52062225,0.392353,0.2678564,0.24522063,0.120724,0.27540162,0.27540162,0.1056335,0.150905,0.2867195,0.5583485,0.754525,0.65643674,0.0452715,0.033953626,0.02263575,0.0150905,0.026408374,0.0754525,0.124496624,0.120724,0.23390275,0.58098423,1.20724,1.0336993,0.44139713,0.10186087,0.15845025,0.24522063,0.56212115,1.0072908,1.3845534,1.539231,1.3430545,1.0978339,1.3015556,1.5731846,1.7089992,1.7089992,1.5128226,1.3091009,1.237421,1.1619685,0.68661773,0.44139713,0.47157812,0.7167987,1.0751982,1.4034165,1.8448136,1.9542197,1.9240388,1.8674494,1.8297231,1.3807807,1.1846043,1.086516,1.0148361,0.97710985,0.98842776,1.0110635,1.0601076,1.0525624,0.80734175,0.6752999,0.59607476,0.5394854,0.47535074,0.36594462,0.3772625,0.55457586,0.86770374,1.2034674,1.3732355,0.95824677,0.43385187,0.1358145,0.10940613,0.120724,0.071679875,0.041498873,0.07922512,0.15467763,0.1659955,0.094315626,0.030181,0.0,0.003772625,0.0150905,0.08677038,0.071679875,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.02263575,0.030181,0.049044125,0.09808825,0.18485862,0.15845025,0.3169005,0.27917424,0.049044125,0.0,0.10940613,0.120724,0.0754525,0.030181,0.030181,0.018863125,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.03772625,0.056589376,0.060362,0.060362,0.060362,0.060362,0.05281675,0.08299775,0.15845025,0.24522063,0.16976812,0.181086,0.1659955,0.116951376,0.090543,0.12826926,0.18485862,0.24899325,0.28294688,0.19994913,0.1358145,0.1659955,0.34330887,0.663982,1.0525624,1.3807807,1.237421,1.1996948,1.6222287,2.625747,3.5387223,4.7572803,4.727099,3.561358,3.0369632,3.1840954,3.640583,4.9345937,6.4436436,6.3945994,7.6018395,7.4094353,6.2021956,4.45547,2.746471,2.3201644,4.0517993,5.6513925,6.058836,5.4476705,4.749735,3.682082,2.5616124,1.8674494,2.1956677,3.1727777,3.783943,3.3764994,2.1202152,1.0223814,1.2902378,2.3918443,3.7914882,4.798779,4.5761943,2.4786146,1.4411428,1.0148361,0.8639311,0.77716076,0.8262049,0.6451189,0.83752275,1.2487389,0.9922004,0.55080324,0.32444575,0.23767537,0.24522063,0.3055826,0.452715,0.58098423,0.63002837,0.59607476,0.5357128,0.29049212,0.17354076,0.13204187,0.120724,0.120724,0.120724,0.1961765,0.32821837,0.43385187,0.33576363,0.26408374,0.23390275,0.19994913,0.18485862,0.32067314,0.56589377,0.72811663,0.83752275,0.86770374,0.73188925,0.91674787,0.8978847,0.9393836,1.1431054,1.448688,1.6222287,1.4449154,1.1619685,0.9808825,1.0525624,1.1732863,1.1959221,1.1544232,1.0940613,1.0827434,0.77716076,0.573439,0.49421388,0.58098423,0.8865669,1.3732355,1.7882242,2.2258487,2.6446102,2.8521044,3.0369632,3.3010468,2.886058,2.203213,2.837014,3.169005,3.350091,3.7348988,4.538468,5.8437963,6.7831798,7.001992,6.971811,6.8397694,6.4247804,5.594803,4.8365054,4.719554,5.1873593,5.553304,6.1531515,6.620957,7.9225125,10.608622,14.830189,16.663685,15.675257,13.58145,11.574413,10.329447,10.110635,9.808825,9.2844305,8.601585,8.028146,10.638803,14.275613,15.154634,12.909923,10.589758,10.552032,9.216523,7.6848373,6.5756855,6.0286546,4.7950063,4.1197066,3.9688015,4.478106,5.96452,6.5643673,6.2851934,6.7643166,8.299775,9.827688,10.948157,12.193124,13.170234,14.177525,16.203424,18.010511,18.327412,17.787928,17.463482,18.844261,19.67424,19.368656,18.69713,18.033148,17.350302,16.569368,16.271332,16.478827,16.807045,16.463736,14.607604,12.687338,10.819888,8.99771,7.0812173,6.4436436,6.3153744,6.4436436,6.40969,5.613666,3.9914372,2.9803739,2.3390274,1.7919968,1.0223814,0.362172,0.1358145,0.09808825,0.120724,0.1659955,0.21503963,0.23767537,0.23013012,0.23013012,0.3055826,0.34330887,0.3772625,0.4074435,0.4376245,0.47157812,0.46026024,0.4678055,0.5281675,0.62248313,0.67152727,0.58475685,0.49044126,0.44894236,0.47157812,0.5357128,0.52062225,0.5357128,0.56589377,0.63002837,0.76207024,1.0789708,2.323937,3.8480775,5.0062733,5.1269975,4.7610526,4.878004,4.927048,4.5761943,3.7084904,3.169005,2.6332922,2.1994405,1.931584,1.8448136,2.4559789,3.2029586,3.783943,4.0103,3.8141239,3.5953116,4.7120085,6.2323766,8.145098,11.3669195,15.728074,22.133991,29.867872,37.130177,41.06125,37.703613,32.259716,28.336185,27.355305,28.562544,28.332415,27.01954,26.080156,26.521553,28.913399,30.709167,29.766012,28.038149,26.612097,25.71044,26.27256,27.502436,29.015259,31.233562,35.38345,36.971725,39.714424,42.879654,44.630154,41.993088,37.98656,34.330887,31.512737,29.73583,28.93226,28.845491,28.924715,29.011486,28.909626,28.39655,26.393284,24.31834,22.447119,21.088974,20.598532,19.572378,17.640795,16.195879,15.712983,15.762027,16.007248,15.316857,14.396337,13.483362,12.359119,11.883769,11.197151,10.416218,9.382519,7.6584287,7.2094865,6.7379084,6.0776987,5.3269467,4.851596,4.5950575,4.432834,4.315883,4.2291126,4.1800685,4.2064767,4.293247,4.38379,4.4630156,4.5460134,4.719554,4.870459,4.881777,4.719554,4.4403796,1.1883769,2.093807,2.8596497,3.108643,2.7728794,2.1088974,1.2902378,1.1732863,1.4449154,1.9579924,2.7389257,3.6707642,3.0671442,2.6031113,2.9351022,3.663219,4.244203,4.4894238,4.708236,4.7836885,4.164978,4.5535583,4.8855495,5.093044,5.342037,6.043745,6.3644185,5.66271,5.1571784,5.3873086,6.2021956,7.277394,8.231868,8.299775,7.5490227,6.8774953,7.786698,9.348565,10.144588,9.567377,7.8319697,6.9454026,5.9796104,5.2552667,4.9044123,4.8553686,3.6745367,3.0218725,3.078462,3.942393,5.6325293,7.854605,6.168242,3.9008942,3.1463692,4.772371,7.277394,8.888305,9.446653,9.110889,8.379,7.7150183,8.677037,10.499215,12.121444,12.181807,9.635284,7.3868,5.515578,4.2630663,4.063117,4.957229,5.934339,6.9227667,7.5792036,7.2962565,6.7341356,6.089017,5.455216,4.7421894,3.6594462,2.9011486,2.5389767,2.493705,2.637065,2.8030603,2.957738,3.1124156,3.1652324,3.1954134,3.4859054,3.682082,3.229367,3.0445085,3.4142256,3.99521,4.0404816,4.4441524,5.372218,6.304056,6.013564,4.768598,3.429316,2.203213,1.20724,0.4640329,0.362172,0.482896,0.573439,0.5470306,0.48666862,0.41498876,0.26408374,0.14713238,0.11317875,0.13204187,0.150905,0.17731337,0.21881226,0.27917424,0.362172,0.6752999,0.6526641,0.6111652,0.7130261,0.95447415,0.84884065,0.59230214,0.38858038,0.30935526,0.29049212,0.33953625,0.41498876,0.46026024,0.42630664,0.3055826,0.15467763,0.10186087,0.06413463,0.02263575,0.030181,0.116951376,0.30935526,0.62248313,0.9922004,1.2789198,1.177059,0.91674787,0.86770374,1.0186088,0.9808825,0.7167987,0.58098423,0.5319401,0.5772116,0.77716076,0.68661773,0.663982,0.8639311,1.116697,0.9280658,1.6561824,2.1013522,2.425798,2.6634734,2.7238352,1.8825399,2.04099,2.1654868,1.871222,1.4034165,1.2487389,1.5128226,1.358145,0.724344,0.34330887,0.29426476,0.43385187,0.70170826,1.0450171,1.4034165,1.9127209,2.1692593,2.233394,2.1164427,1.8070874,1.7467253,1.6788181,1.5731846,1.4298248,1.2562841,1.0940613,0.95447415,0.9695646,1.0072908,0.6752999,0.62625575,0.58475685,0.52439487,0.44139713,0.34330887,0.21881226,0.52062225,0.8978847,1.1242423,1.1280149,0.9393836,0.6752999,0.56589377,0.59230214,0.48666862,0.35085413,0.32821837,0.2678564,0.15467763,0.120724,0.06413463,0.02263575,0.0,0.0,0.003772625,0.026408374,0.026408374,0.02263575,0.030181,0.049044125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0150905,0.018863125,0.018863125,0.02263575,0.060362,0.056589376,0.07922512,0.06413463,0.011317875,0.0,0.090543,0.06413463,0.026408374,0.0150905,0.00754525,0.0150905,0.0150905,0.0150905,0.018863125,0.03772625,0.026408374,0.011317875,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.05281675,0.03772625,0.026408374,0.03772625,0.06413463,0.08677038,0.08299775,0.071679875,0.09808825,0.14335975,0.150905,0.120724,0.06790725,0.056589376,0.06413463,0.094315626,0.1659955,0.24899325,0.26031113,0.2263575,0.29426476,0.38480774,0.49044126,0.6752999,0.97333723,1.237421,1.478869,1.7467253,2.11267,2.293756,2.686109,2.7615614,2.4295704,2.0108092,1.8561316,1.9504471,2.5389767,3.440634,4.074435,5.3609,5.723072,5.9494295,5.9796104,4.908185,4.0103,4.2064767,5.0062733,5.824933,5.983383,6.058836,4.889322,3.7537618,3.4330888,4.2102494,3.380272,2.7917426,2.3163917,1.9806281,1.9881734,2.1088974,2.4031622,2.565385,2.3616633,1.6222287,1.0751982,0.8978847,0.8337501,0.7922512,0.814887,0.7092535,0.65643674,0.814887,1.1393328,1.3694628,1.1959221,0.8337501,0.513077,0.32444575,0.21881226,0.18863125,0.23013012,0.35462674,0.47912338,0.4376245,0.32821837,0.23390275,0.150905,0.09808825,0.09808825,0.1056335,0.13958712,0.23767537,0.452715,0.8224323,1.1506506,1.0035182,0.7582976,0.59607476,0.51684964,0.60362,0.8563859,0.9242931,0.784706,0.7582976,1.0374719,1.2261031,1.3166461,1.3619176,1.4600059,1.720317,1.7995421,1.7354075,1.5807298,1.418507,1.5015048,1.4109617,1.2298758,1.0487897,0.9507015,0.7507524,0.784706,1.0789708,1.5203679,1.8749946,2.674791,3.2784111,3.3689542,2.9728284,2.4371157,2.474842,2.3956168,2.214531,2.1315331,2.5314314,3.5462675,4.3385186,5.221313,6.1720147,6.832224,7.1679873,7.432071,7.7112455,7.8734684,7.54525,7.0887623,6.7454534,6.8737226,7.4773426,8.216777,9.107117,9.691874,10.699164,12.238396,13.807808,14.690601,14.6151495,14.034165,13.185325,12.08749,10.831206,9.314611,8.265821,8.52236,11.016065,13.0646,14.93205,16.060064,15.920478,14.019074,12.725064,11.385782,9.967276,8.526133,7.224577,6.1078796,5.624984,5.304311,5.2175403,5.96452,7.1604424,7.877241,8.89585,10.220041,11.072655,10.8576145,10.982111,11.631002,13.041965,15.509261,16.505234,17.048492,17.53139,18.225552,19.28566,19.87796,19.202662,18.16519,17.191853,16.22606,15.524352,15.211224,14.856597,14.019074,12.242168,10.416218,9.514561,9.21275,9.114662,8.75249,7.9225125,7.4697976,7.175533,6.8171334,6.187105,5.2892203,4.2894745,3.2821836,2.2447119,1.0336993,0.38480774,0.1659955,0.14335975,0.17354076,0.20372175,0.21503963,0.211267,0.21881226,0.24522063,0.27917424,0.29803738,0.33576363,0.3961256,0.45648763,0.48666862,0.4640329,0.452715,0.46026024,0.48666862,0.5357128,0.52062225,0.5583485,0.6526641,0.7432071,0.7167987,0.7130261,0.754525,0.80356914,0.875249,1.0186088,1.2185578,2.3163917,3.5123138,4.402653,4.957229,4.9987283,4.429062,3.8707132,3.5236318,3.1840954,2.9086938,2.6068838,2.2069857,1.7618159,1.4298248,1.629774,2.1503963,2.8634224,3.591539,4.1083884,4.055572,4.22534,5.2326307,6.964266,8.586494,10.344538,14.471789,22.224533,33.13119,44.992325,48.266964,45.365814,39.657833,34.515747,33.31228,32.16163,29.954643,28.25319,28.166418,30.343224,34.100758,34.659107,33.712177,32.633205,32.474754,33.72727,34.093212,34.342205,35.115593,36.92268,39.027805,41.114067,42.491074,42.574074,40.906574,37.303715,35.108047,33.810265,33.221737,33.47073,32.848248,32.1654,31.923952,31.908863,31.180746,28.377686,25.435038,23.235598,22.156626,22.08872,21.14179,19.742147,18.33873,17.165443,16.237377,16.0412,15.999702,15.886524,15.55076,14.886778,13.20796,11.921495,10.978339,10.20495,9.2844305,8.14887,7.303802,6.6247296,6.0814714,5.7306175,5.455216,5.1534057,4.8365054,4.52715,4.255521,4.1310244,4.08198,4.06689,4.06689,4.0970707,4.1574326,4.2404304,4.327201,4.402653,4.4516973,0.76584285,1.6335466,2.4182527,2.7351532,2.5238862,2.052308,1.4524606,1.177059,1.0902886,1.2525115,1.9202662,2.6144292,2.5729303,2.674791,3.3425457,4.5422406,4.798779,4.8930945,5.0251365,5.081726,4.666737,4.164978,4.08198,4.1989317,4.466788,5.0213637,5.50426,5.5306683,5.4401255,5.2779026,4.7648253,5.1043615,6.013564,6.828451,7.575431,8.971302,10.612394,11.951676,12.121444,10.801025,8.231868,6.809588,6.0286546,5.7381625,5.881522,6.488915,6.432326,5.832478,5.3910813,5.4288073,5.8626595,6.462507,5.764571,4.930821,4.908185,6.417235,6.6360474,7.0284004,7.3679366,7.5490227,7.598067,7.3075747,7.643338,7.9225125,7.84706,7.515069,6.7077274,5.1458607,3.7084904,2.8747404,2.7087448,4.074435,6.205968,8.484633,9.590013,7.496206,6.2021956,5.5004873,5.1534057,4.8666863,4.266839,3.5802212,3.5236318,3.8480775,4.2819295,4.515832,4.478106,4.715781,4.398881,3.5953116,3.2670932,3.4217708,3.361409,3.361409,3.5689032,3.9989824,3.5274043,3.3161373,3.8141239,4.859141,5.666483,5.028909,3.7009451,2.335255,1.2751472,0.5470306,0.31312788,0.2867195,0.43385187,0.633801,0.7205714,0.6828451,0.5470306,0.3734899,0.211267,0.11317875,0.16976812,0.29426476,0.38480774,0.36971724,0.20372175,0.44516975,0.4376245,0.4678055,0.65643674,0.9507015,0.97333723,0.8186596,0.5696664,0.34330887,0.2867195,0.36971724,0.45648763,0.5017591,0.44894236,0.26408374,0.1961765,0.12826926,0.06413463,0.011317875,0.018863125,0.033953626,0.09808825,0.23767537,0.44516975,0.67152727,0.6752999,0.58098423,0.6073926,0.7507524,0.784706,0.6413463,0.51684964,0.38103512,0.3055826,0.46026024,0.3734899,0.38858038,0.5394854,0.694163,0.58475685,0.9393836,1.5354583,3.3840446,6.228604,8.533678,6.2399216,3.8103511,2.444661,2.142851,1.6675003,1.2411937,1.1280149,0.86770374,0.49044126,0.51684964,0.65643674,0.754525,0.83752275,0.9808825,1.3317367,1.7618159,2.0447628,2.161714,2.1164427,1.9202662,1.9504471,1.81086,1.6033657,1.3996439,1.2713746,1.116697,0.8941121,0.83752275,0.8978847,0.7432071,0.70170826,0.66020936,0.6073926,0.52062225,0.3734899,0.19994913,0.26031113,0.3772625,0.44516975,0.44516975,0.43007925,0.5281675,0.6488915,0.694163,0.55080324,0.241448,0.16222288,0.124496624,0.06413463,0.041498873,0.02263575,0.00754525,0.00754525,0.03772625,0.120724,0.06413463,0.030181,0.030181,0.05281675,0.071679875,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.041498873,0.033953626,0.026408374,0.026408374,0.018863125,0.018863125,0.02263575,0.030181,0.03772625,0.05281675,0.056589376,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.0150905,0.003772625,0.011317875,0.011317875,0.00754525,0.003772625,0.0,0.00754525,0.03772625,0.02263575,0.00754525,0.003772625,0.0,0.003772625,0.011317875,0.011317875,0.00754525,0.018863125,0.0150905,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.018863125,0.02263575,0.0452715,0.14713238,0.16222288,0.12826926,0.07922512,0.041498873,0.0452715,0.0452715,0.03772625,0.033953626,0.060362,0.09808825,0.090543,0.071679875,0.0452715,0.026408374,0.033953626,0.05281675,0.094315626,0.15467763,0.23013012,0.2565385,0.29426476,0.35462674,0.46026024,0.663982,0.97710985,1.177059,1.3770081,1.6750455,2.1654868,2.263575,2.1353056,2.1881225,2.5578396,3.127506,3.2029586,2.9237845,2.463524,1.9994912,1.690136,3.2255943,4.3347464,5.907931,7.9753294,9.740918,10.295494,6.9265394,4.327201,4.074435,4.6252384,5.1647234,4.5497856,3.7198083,3.2670932,3.4255435,2.6898816,2.071171,1.7731338,2.082489,3.380272,4.402653,3.7047176,2.463524,1.3996439,0.77338815,0.6149379,0.5998474,0.70170826,0.8337501,0.8601585,0.69039035,0.6149379,0.58475685,0.6111652,0.724344,0.8186596,0.814887,0.76584285,0.6451189,0.38103512,0.23390275,0.18485862,0.2263575,0.30181,0.30181,0.32444575,0.33953625,0.32444575,0.27917424,0.21881226,0.15845025,0.1358145,0.14713238,0.25276586,0.58098423,0.8111144,0.8299775,0.8563859,0.9695646,1.1053791,0.80356914,0.754525,0.76584285,0.784706,0.9016574,1.0148361,1.2902378,1.5316857,1.6486372,1.6863633,1.780679,1.8636768,1.8259505,1.6863633,1.5845025,1.5316857,1.3732355,1.177059,0.98465514,0.80734175,0.7809334,1.1883769,1.7089992,2.1503963,2.41448,3.5500402,3.832987,3.6481283,3.180323,2.4522061,2.3956168,2.8143783,3.8556228,4.9647746,4.881777,6.0512905,6.8397694,7.01331,6.790725,6.858632,6.458734,6.33801,6.4134626,6.458734,6.115425,5.7192993,6.1795597,6.9454026,7.8017883,8.843033,9.933322,10.499215,11.329193,12.540206,13.558814,13.773854,13.70972,13.649357,13.272095,11.631002,9.993684,8.903395,9.220296,11.3820095,15.418718,15.426264,14.743419,14.958458,15.928022,15.773345,14.18507,12.264804,10.748209,9.756008,8.786444,8.213005,8.050782,7.9828744,7.7225633,7.0548086,7.356619,7.884786,8.854351,10.182315,11.465008,11.517824,11.521597,11.766817,12.457208,13.705947,14.6151495,15.603577,16.70141,17.803017,18.670721,18.863125,18.263277,17.542706,16.965494,16.41092,15.860115,15.328176,14.445381,12.90615,10.461489,8.00551,7.232122,7.673519,8.790216,9.986138,10.001229,8.892077,7.466025,6.2361493,5.406172,4.7836885,4.0103,3.1124156,2.1881225,1.4034165,0.7922512,0.46026024,0.32067314,0.2867195,0.2678564,0.23013012,0.23390275,0.26408374,0.29049212,0.30181,0.31312788,0.3470815,0.41498876,0.48666862,0.48666862,0.47912338,0.49044126,0.47157812,0.452715,0.52062225,0.55080324,0.6149379,0.69793564,0.7696155,0.7809334,0.76584285,0.7809334,0.8111144,0.86770374,0.9922004,1.2525115,1.8825399,2.6898816,3.451952,3.8971217,3.8178966,3.3764994,3.270866,3.5424948,3.5538127,3.3274553,3.048281,2.7011995,2.3126192,1.9504471,1.5505489,1.6071383,2.0447628,2.7125173,3.3953626,3.5802212,3.6368105,4.191386,5.2175403,6.047518,6.779407,8.782671,13.340002,20.515535,29.166164,34.33466,36.654823,36.8095,35.387222,32.863335,30.067822,27.260988,25.118137,24.239115,25.15209,28.596497,30.59599,31.81832,32.833157,34.11962,35.209908,35.2665,36.14552,38.058243,39.57861,41.37438,42.81175,43.51346,43.509686,43.253147,42.649525,41.457375,40.035095,38.714676,37.82811,37.115086,35.598488,34.372387,33.57259,32.361576,29.796192,26.857317,24.34475,22.669704,21.85859,21.383238,21.077656,20.496672,19.270569,17.082445,17.165443,17.591751,17.859608,17.625704,16.72782,14.762281,12.785426,11.34051,10.487898,9.789962,8.835487,8.016829,7.352846,6.8435416,6.4926877,6.1644692,5.7909794,5.372218,4.927048,4.5120597,4.221567,4.006528,3.8556228,3.7575345,3.7160356,3.7386713,3.7990334,3.8707132,3.9574835,4.0970707,0.9242931,1.539231,2.1051247,2.3503454,2.2296214,1.9466745,1.6033657,1.2789198,1.056335,1.0676528,1.5241405,1.7580433,2.3126192,3.0143273,3.821669,4.821415,4.8629136,5.028909,5.138315,5.0515447,4.647874,3.7084904,3.3274553,3.2972744,3.5236318,4.036709,4.610148,5.142088,5.330719,4.927048,3.7198083,4.036709,4.961002,6.3531003,8.194141,10.608622,12.1252165,13.551269,13.43809,11.566868,8.937348,7.2585306,6.5040054,6.017337,5.7683434,6.360646,8.028146,8.567632,8.224322,7.3151197,6.217286,5.6891184,5.8173876,6.126743,6.4549613,6.9793563,5.481624,5.5797124,6.1342883,6.587003,6.9454026,6.900131,6.692637,6.1531515,5.5080323,5.3646727,5.0968165,3.7688525,2.546522,1.9693103,1.9542197,3.270866,5.617439,8.420499,10.321902,9.186342,6.609639,5.198677,4.689373,4.7535076,4.9987283,5.093044,5.3080835,6.089017,6.8661776,6.043745,4.979865,4.7874613,4.67051,4.2630663,3.6594462,3.5160866,3.5575855,3.5990841,3.682082,4.0706625,3.7047176,3.3764994,3.361409,3.8178966,4.798779,4.7233267,3.3840446,1.9579924,0.9997456,0.45648763,0.23013012,0.14335975,0.2565385,0.52439487,0.7809334,0.9016574,0.875249,0.7130261,0.47535074,0.29426476,0.36594462,0.5583485,0.6413463,0.5055317,0.14335975,0.27917424,0.33953625,0.41876137,0.543258,0.694163,0.8337501,0.86770374,0.7394345,0.4979865,0.31312788,0.35839936,0.41498876,0.41876137,0.34330887,0.211267,0.18485862,0.1659955,0.12826926,0.0754525,0.056589376,0.033953626,0.018863125,0.0150905,0.02263575,0.041498873,0.094315626,0.13204187,0.20372175,0.30181,0.38103512,0.35085413,0.2678564,0.15845025,0.10186087,0.24899325,0.6488915,0.8262049,0.84884065,0.77716076,0.6526641,0.56212115,1.1129243,3.138824,6.2323766,8.75249,6.9567204,4.6327834,3.169005,2.6823363,1.9881734,1.3204187,0.8978847,0.633801,0.5357128,0.7054809,0.8186596,0.8186596,0.7809334,0.8526133,1.2261031,1.569412,1.8599042,2.0183544,2.022127,1.9240388,1.8900851,1.6750455,1.4147344,1.2110126,1.1317875,1.0299267,0.845068,0.79602385,0.87147635,0.845068,0.77338815,0.70170826,0.6526641,0.6073926,0.543258,0.32067314,0.15467763,0.0754525,0.0754525,0.12826926,0.1659955,0.35085413,0.59607476,0.76207024,0.66775465,0.24522063,0.056589376,0.003772625,0.003772625,0.0,0.0,0.0,0.011317875,0.06790725,0.22258487,0.10186087,0.033953626,0.018863125,0.03772625,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0452715,0.049044125,0.03772625,0.033953626,0.041498873,0.05281675,0.041498873,0.030181,0.033953626,0.041498873,0.06413463,0.06413463,0.0452715,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.02263575,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.049044125,0.0754525,0.090543,0.11317875,0.1358145,0.150905,0.25276586,0.28294688,0.24899325,0.20372175,0.21503963,0.1659955,0.094315626,0.041498873,0.026408374,0.049044125,0.05281675,0.041498873,0.03772625,0.03772625,0.026408374,0.0452715,0.060362,0.11317875,0.1961765,0.29049212,0.331991,0.33953625,0.38480774,0.5357128,0.83752275,1.2713746,1.7429527,2.1202152,2.354118,2.4710693,2.7615614,3.1954134,3.482133,3.6783094,4.1762958,4.432834,4.112161,3.2218218,2.0145817,0.98842776,1.8221779,3.029418,5.2779026,8.620448,12.468526,13.249459,9.012801,5.251494,4.285702,5.2854476,5.670255,5.587258,5.138315,4.4516973,3.6971724,2.848332,2.1390784,1.7995421,2.11267,3.4179983,4.4894238,3.742444,2.4107075,1.3128735,0.84884065,0.663982,0.63002837,0.784706,1.0412445,1.1657411,0.7884786,0.56212115,0.38858038,0.2565385,0.23013012,0.40367088,0.5998474,0.784706,0.8865669,0.784706,0.59230214,0.33953625,0.181086,0.15845025,0.18485862,0.2565385,0.32821837,0.36971724,0.38480774,0.40367088,0.2678564,0.30181,0.33953625,0.32444575,0.32821837,0.392353,0.543258,0.73188925,0.935611,1.1657411,0.9205205,0.8111144,0.77338815,0.8299775,1.1129243,1.2449663,1.4562333,1.599593,1.6524098,1.7391801,1.7429527,1.7542707,1.7014539,1.5920477,1.5354583,1.2940104,1.1204696,1.026154,1.0487897,1.267602,1.780679,2.1353056,2.384299,2.493705,2.3465726,3.0331905,3.1350515,3.150142,3.0558262,2.3314822,2.1881225,3.1161883,5.119452,7.466025,8.692128,8.062099,7.567886,6.8359966,6.009792,5.7306175,5.1760416,5.081726,5.194905,5.2062225,4.749735,4.293247,4.7535076,5.413717,6.047518,6.8925858,8.560086,9.64283,10.646348,11.808316,13.087236,14.403882,13.837989,12.630749,11.283921,9.574923,9.035437,8.337502,9.046755,11.548005,15.07541,14.830189,14.056801,14.045483,15.0376835,16.22606,15.588487,14.675511,14.234114,14.003984,12.721292,10.902886,10.386037,10.499215,10.397354,9.046755,8.484633,8.175279,8.918486,10.657665,12.472299,12.845788,13.140053,13.45318,13.690856,13.5663595,13.932304,14.84528,16.16947,17.53516,18.297232,17.957695,17.263533,16.663685,16.35433,16.260014,16.244923,15.988385,15.192361,13.641812,11.193378,8.209232,6.470052,6.470052,7.914967,9.718282,10.216269,9.046755,7.2623034,5.704209,5.028909,4.7006907,4.074435,3.1765501,2.2409391,1.690136,1.0751982,0.6790725,0.4640329,0.36594462,0.29803738,0.26408374,0.27917424,0.31312788,0.34330887,0.38103512,0.41876137,0.43007925,0.45648763,0.47912338,0.4376245,0.4376245,0.482896,0.4979865,0.4979865,0.5583485,0.5885295,0.6451189,0.69039035,0.7130261,0.7092535,0.7092535,0.77716076,0.83752275,0.88279426,0.965792,1.2411937,1.5920477,2.1692593,2.8521044,3.2746384,3.199186,2.9916916,3.048281,3.350091,3.500996,3.4368613,3.2444575,2.9954643,2.746471,2.565385,2.2447119,2.0636258,2.3692086,3.1161883,3.874486,3.9008942,3.6556737,3.9310753,4.636556,4.8100967,4.772371,5.2288585,6.760544,9.616421,13.705947,18.150099,23.111101,27.872154,31.199608,31.327879,27.977787,25.291677,22.997923,21.217243,20.485353,22.409393,24.431519,26.827137,29.41893,31.584417,32.384212,32.282352,33.319824,36.036114,39.472977,42.81552,45.448814,46.848457,46.972954,46.24484,46.686234,45.822304,44.35098,42.660843,40.83112,39.642742,37.907337,36.353016,35.08541,33.599,31.527826,29.068075,26.351786,23.741129,21.820864,21.311558,21.560553,21.662413,20.964478,19.051756,19.078165,19.21398,19.236614,18.915941,18.033148,16.127972,13.694629,11.69891,10.435081,9.525878,8.778898,8.096053,7.5075235,7.0246277,6.6360474,6.319147,5.987156,5.617439,5.1835866,4.689373,4.3121104,3.9989824,3.7499893,3.5651307,3.4670424,3.5236318,3.6066296,3.6481283,3.663219,3.7462165,1.2600567,1.6222287,1.8523588,1.931584,1.8787673,1.7467253,1.5165952,1.3845534,1.3166461,1.3732355,1.7089992,1.7127718,2.41448,3.3425457,4.164978,4.689373,4.82896,5.0854983,5.100589,4.7006907,3.904667,3.1652324,2.7691069,2.6634734,2.8785129,3.5047686,3.9612563,4.2291126,4.172523,3.7273536,2.886058,3.8254418,5.1647234,6.911449,8.929804,10.929295,12.140307,14.068119,14.045483,11.857361,9.737145,8.646856,7.798016,6.4210076,4.9723196,5.138315,7.8017883,9.616421,9.933322,8.793989,6.930312,5.2175403,4.949684,5.4250345,5.987156,6.0248823,4.738417,5.4212623,6.006019,5.798525,5.4740787,5.330719,5.13077,5.111907,5.372218,5.8626595,5.3609,4.1536603,2.9313297,2.0636258,1.599593,1.8976303,3.3840446,5.674028,8.13378,9.865415,6.6586833,4.749735,3.9914372,4.164978,4.9647746,6.1531515,6.6549106,7.5301595,8.118689,6.0550632,4.06689,3.3123648,3.783943,4.719554,4.610148,3.9574835,3.4783602,3.3274553,3.5349495,3.983892,3.832987,3.742444,3.663219,3.6707642,3.983892,4.1536603,2.927557,1.5807298,0.724344,0.31312788,0.211267,0.19994913,0.24899325,0.392353,0.73566186,1.0035182,1.1242423,1.0638802,0.86770374,0.66020936,0.73566186,0.86770374,0.845068,0.62625575,0.34330887,0.3961256,0.47157812,0.49044126,0.44516975,0.422534,0.5772116,0.7469798,0.8111144,0.6790725,0.32444575,0.26408374,0.28294688,0.29049212,0.25276586,0.23013012,0.17731337,0.16222288,0.16222288,0.14713238,0.08677038,0.07922512,0.056589376,0.033953626,0.026408374,0.026408374,0.026408374,0.041498873,0.09808825,0.181086,0.21881226,0.15467763,0.094315626,0.07922512,0.13958712,0.30935526,1.2147852,1.8825399,2.173032,2.1164427,1.9202662,1.9881734,1.9768555,2.173032,2.5917933,3.006782,3.2821836,3.712263,3.7009451,3.0709167,2.093807,1.4335974,1.1242423,1.0110635,0.95824677,0.86770374,0.7432071,0.6451189,0.63002837,0.7696155,1.1242423,1.4335974,1.7467253,1.9240388,1.9202662,1.7882242,1.6675003,1.4562333,1.237421,1.0638802,0.965792,0.88279426,0.7997965,0.814887,0.9016574,0.9016574,0.77716076,0.663982,0.6073926,0.63002837,0.72811663,0.46026024,0.25276586,0.1659955,0.19240387,0.2565385,0.23013012,0.25276586,0.482896,0.79602385,0.7997965,0.44139713,0.21503963,0.116951376,0.094315626,0.0452715,0.02263575,0.00754525,0.011317875,0.071679875,0.241448,0.09808825,0.030181,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.018863125,0.030181,0.026408374,0.011317875,0.0,0.018863125,0.018863125,0.011317875,0.0150905,0.02263575,0.06413463,0.0452715,0.018863125,0.011317875,0.011317875,0.02263575,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.011317875,0.07922512,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.018863125,0.049044125,0.116951376,0.15845025,0.17731337,0.21503963,0.2678564,0.27540162,0.3961256,0.5281675,0.51684964,0.41876137,0.52062225,0.41498876,0.27540162,0.150905,0.08299775,0.11317875,0.08299775,0.05281675,0.03772625,0.041498873,0.071679875,0.090543,0.1056335,0.181086,0.29803738,0.3772625,0.39989826,0.40367088,0.44516975,0.59607476,0.94315624,1.5279131,2.5880208,3.5085413,3.8178966,3.1840954,3.429316,4.6290107,5.1760416,4.779916,4.466788,4.8025517,4.715781,4.236658,3.5349495,2.927557,2.282438,2.5729303,4.3347464,7.454707,11.18206,11.204697,9.582467,7.8206515,7.1038527,8.296002,8.145098,8.299775,8.145098,7.3415284,5.836251,4.3121104,3.3689542,2.897376,2.7200627,2.5993385,2.6483827,2.595566,2.233394,1.6373192,1.1581959,0.90543,0.8224323,0.9318384,1.1732863,1.418507,0.8865669,0.5696664,0.38480774,0.27917424,0.24899325,0.29049212,0.3772625,0.58098423,0.875249,1.1355602,0.9620194,0.513077,0.181086,0.09808825,0.124496624,0.1659955,0.20372175,0.24522063,0.31312788,0.4678055,0.32067314,0.45648763,0.59230214,0.5696664,0.3470815,0.35839936,0.5055317,0.66020936,0.754525,0.754525,0.935611,1.0412445,0.97710985,0.9016574,1.2336484,1.5430037,1.6410918,1.5505489,1.4335974,1.5807298,1.5731846,1.50905,1.4335974,1.358145,1.267602,0.9393836,0.84129536,0.91674787,1.2411937,2.0108092,2.9351022,2.8709676,2.5917933,2.3428001,1.8561316,1.6033657,1.7580433,2.1654868,2.4333432,1.9202662,1.8599042,3.059599,5.270357,8.069645,10.872705,8.043237,6.2889657,5.2590394,4.6327834,4.1272516,3.8367596,4.0480266,4.425289,4.5912848,4.142342,3.7952607,3.9008942,4.168751,4.485651,4.8742313,6.5945487,8.273367,9.507015,10.453944,11.830952,14.781145,14.007756,11.400873,8.699674,7.5301595,8.443134,7.745199,7.665974,8.827943,10.231359,11.41219,12.377983,13.04951,13.834216,15.614895,16.131744,17.72002,19.183798,19.270569,16.667458,13.93985,12.683565,12.30253,12.0082655,10.827434,10.008774,9.012801,9.525878,11.555551,13.441863,13.804035,14.456699,15.192361,15.592259,15.026365,14.558559,15.030138,16.271332,17.716248,18.384,17.610613,16.610868,15.773345,15.328176,15.339493,15.999702,16.542961,16.550507,15.633758,13.43809,10.223814,7.1868505,6.009792,6.8058157,8.114917,8.443134,7.828197,6.643593,5.485397,5.168496,5.05909,4.4139714,3.399135,2.3314822,1.6712729,1.0902886,0.72811663,0.513077,0.38858038,0.29803738,0.3055826,0.331991,0.35085413,0.36971724,0.45648763,0.5319401,0.52439487,0.49421388,0.452715,0.3772625,0.36594462,0.41121614,0.47157812,0.5281675,0.5583485,0.56212115,0.6149379,0.65643674,0.6488915,0.5998474,0.65643674,0.845068,0.995973,1.0676528,1.1695137,1.3770081,1.659955,2.0636258,2.584248,3.1576872,3.3274553,3.2029586,2.9237845,2.704972,2.8219235,3.0105548,2.9992368,2.9351022,2.9426475,3.138824,3.338773,3.1312788,3.380272,4.217795,5.0553174,4.957229,4.357382,4.606375,5.458988,5.05909,4.3309736,3.904667,3.9122121,4.6629643,6.6360474,9.371201,13.456953,18.85558,24.880463,30.218727,28.35505,25.891525,23.163918,20.700394,19.198889,19.957186,21.232334,23.201643,25.601034,27.702385,28.54368,28.588953,29.019032,31.195837,36.65105,42.54012,47.59921,50.568264,50.74558,47.984016,46.082615,44.573563,43.40405,42.3364,40.925434,39.46543,38.47323,37.6093,36.624645,35.334404,33.81781,31.810774,28.98885,25.714212,23.020557,21.851044,21.83218,21.994404,21.794455,21.085201,20.62494,20.059048,19.591242,19.221525,18.72731,16.927769,14.449154,12.117672,10.303039,8.956212,8.088508,7.4999785,6.9982195,6.5266414,6.1418333,5.915476,5.726845,5.50426,5.1873593,4.719554,4.3724723,4.044254,3.7537618,3.519859,3.3651814,3.4481792,3.5500402,3.5990841,3.591539,3.5839937,1.1732863,1.3694628,1.3468271,1.3996439,1.5882751,1.7089992,1.4411428,1.6675003,1.6486372,1.3166461,1.2826926,1.599593,2.2447119,3.0709167,4.044254,5.2628117,5.6061206,5.2779026,4.5233774,3.6745367,3.1727777,2.795515,2.5804756,2.5502944,2.7087448,3.0520537,3.187868,2.927557,2.5540671,2.3503454,2.595566,4.1197066,5.9494295,7.5527954,8.937348,10.63503,12.785426,14.456699,14.079436,12.106354,11.031156,11.970539,11.117926,9.114662,7.3717093,8.054554,8.326183,8.073418,7.997965,8.07719,7.5527954,4.696918,2.9954643,2.4861598,3.0105548,4.1800685,5.119452,5.5495315,5.1081343,3.9612563,2.776652,2.3503454,2.3088465,2.8030603,3.8858037,5.5080323,6.862405,5.994701,4.2291126,2.5276587,1.4637785,1.0148361,1.7618159,2.7125173,3.2746384,3.2520027,2.6408374,2.8822856,3.0520537,2.938875,3.0369632,4.4403796,5.66271,5.4665337,4.0782075,3.1727777,2.746471,2.7238352,3.2784111,4.304565,5.4174895,3.953711,2.8822856,2.6068838,3.0709167,3.7537618,3.863168,4.074435,3.7688525,3.1652324,3.3123648,3.2369123,2.625747,1.7693611,0.9808825,0.58098423,0.422534,0.38103512,0.422534,0.55080324,0.80734175,0.9318384,1.1883769,1.3317367,1.2449663,0.97710985,1.1732863,1.0827434,0.8865669,0.73566186,0.7469798,0.90543,0.8639311,0.65643674,0.39989826,0.29049212,0.46026024,0.694163,0.83752275,0.7884786,0.52062225,0.31312788,0.29426476,0.36971724,0.4376245,0.42630664,0.34330887,0.21881226,0.120724,0.0754525,0.0754525,0.0754525,0.08677038,0.07922512,0.06413463,0.0754525,0.0754525,0.1056335,0.1961765,0.3055826,0.3055826,0.21881226,0.16976812,0.21503963,0.44516975,1.0072908,0.935611,2.1805773,3.5274043,4.3347464,4.5309224,5.994701,4.61392,2.5804756,1.1393328,0.56589377,0.9205205,1.4298248,1.9957186,2.323937,1.9240388,1.6524098,1.6675003,1.8297231,1.8674494,1.4034165,1.0374719,0.8903395,0.8978847,0.9808825,1.0525624,1.3694628,1.6788181,1.8297231,1.7995421,1.6788181,1.569412,1.4298248,1.2600567,1.0789708,0.9318384,0.80734175,0.724344,0.724344,0.80734175,0.91674787,0.73188925,0.56589377,0.5017591,0.5357128,0.59607476,0.3734899,0.27540162,0.2565385,0.2565385,0.18485862,0.049044125,0.09808825,0.26408374,0.44516975,0.52062225,0.49421388,0.56212115,0.55457586,0.422534,0.23013012,0.1056335,0.030181,0.00754525,0.0452715,0.1659955,0.08299775,0.05281675,0.026408374,0.0,0.0,0.0,0.018863125,0.018863125,0.0,0.0,0.0,0.0,0.018863125,0.0452715,0.0452715,0.094315626,0.14335975,0.1056335,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.030181,0.030181,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.041498873,0.071679875,0.090543,0.090543,0.1056335,0.116951376,0.13958712,0.19994913,0.33576363,0.70170826,1.2336484,1.237421,0.7884786,0.70170826,0.6149379,0.5017591,0.36971724,0.29426476,0.44139713,0.331991,0.20372175,0.10186087,0.071679875,0.1659955,0.1659955,0.150905,0.13204187,0.13204187,0.1659955,0.241448,0.27917424,0.33953625,0.45648763,0.62625575,1.2110126,2.3390274,3.8895764,5.1760416,4.9421387,4.1989317,3.8556228,3.8405323,4.13857,4.821415,5.613666,5.583485,5.8702044,6.760544,7.673519,6.2097406,4.7346444,4.4139714,5.3948536,6.8359966,8.763808,10.069136,10.510533,10.355856,10.4049,10.148361,10.352083,10.325675,9.537196,7.5829763,6.25124,6.0022464,6.009792,5.492942,3.7235808,3.138824,2.9916916,2.674791,2.0636258,1.5241405,1.1355602,0.7997965,0.6526641,0.68661773,0.7469798,0.77338815,0.7432071,0.6375736,0.47912338,0.32067314,0.19994913,0.22258487,0.35839936,0.573439,0.8563859,0.7205714,0.44894236,0.23390275,0.150905,0.1358145,0.150905,0.14335975,0.14335975,0.150905,0.1358145,0.08677038,0.094315626,0.16976812,0.29803738,0.45648763,0.47157812,0.59230214,0.95824677,1.2902378,0.9016574,1.0223814,1.0638802,1.0299267,0.97710985,0.97710985,1.1581959,1.3053282,1.4222796,1.4939595,1.4939595,1.2638294,1.0789708,0.91674787,0.80356914,0.77716076,0.754525,0.8563859,1.0902886,1.4147344,1.7542707,1.6939086,1.5128226,1.3317367,1.2713746,1.4637785,1.1732863,1.1732863,1.1883769,1.2110126,1.478869,2.0183544,3.6066296,5.541986,6.881268,6.4549613,5.5382137,5.8211603,5.6778007,4.6742826,3.6028569,2.9426475,2.6483827,2.6974268,2.9313297,3.0671442,3.3953626,4.8629136,6.507778,7.752744,8.375228,7.3151197,8.084735,8.786444,8.975075,9.65792,10.831206,11.344283,10.597303,9.031664,8.118689,7.752744,7.6320205,8.043237,8.45068,7.5226145,8.341274,8.345046,9.216523,11.393328,14.053028,13.5663595,16.776863,18.919714,17.814335,13.8870325,17.048492,16.097792,13.766309,11.68382,10.374719,9.544742,9.0543,9.273112,10.231359,11.61214,12.393073,13.377728,14.102073,14.562332,15.196134,15.101818,15.818617,16.788181,17.614386,18.0671,17.369165,16.42601,15.513034,14.815099,14.449154,15.109364,16.35433,17.48989,17.516298,15.135772,11.608367,8.677037,6.820906,6.187105,6.5756855,6.8925858,6.5341864,5.8437963,5.05909,4.304565,3.6556737,2.9615107,2.2862108,1.7089992,1.3430545,1.0638802,0.754525,0.51684964,0.38480774,0.33576363,0.3734899,0.39989826,0.38103512,0.3470815,0.3961256,0.47157812,0.5055317,0.5017591,0.4640329,0.42630664,0.36594462,0.331991,0.32821837,0.35085413,0.41121614,0.422534,0.47157812,0.5281675,0.58475685,0.67152727,0.8186596,1.0299267,1.237421,1.448688,1.7542707,1.9730829,1.9278114,1.8184053,1.8749946,2.3654358,2.5729303,2.5616124,2.463524,2.3956168,2.4559789,2.565385,2.6408374,2.927557,3.4896781,4.2102494,4.0404816,3.5575855,3.1425967,3.1124156,3.7235808,4.908185,5.20245,5.715527,6.4134626,6.1342883,5.7192993,4.8629136,4.1197066,3.7801702,3.8895764,5.0515447,8.160188,13.70972,21.051247,28.411638,30.181,26.378195,21.82841,19.379974,19.881733,21.87368,24.27307,25.408628,25.604805,27.19308,28.607815,29.822601,30.656351,31.852272,35.06655,40.08414,45.769485,49.90428,50.839893,47.47094,41.536602,38.020515,36.307743,35.847485,36.164383,36.688778,37.36785,37.6508,37.371624,36.771774,36.285107,34.093212,31.139246,28.147554,25.634987,23.839218,23.246916,22.816835,21.915178,20.277859,19.779873,19.379974,19.153618,18.97253,18.5085,16.825907,14.7736,12.551523,10.408672,8.650629,7.4811153,6.937857,6.398372,5.7494807,5.43258,5.383536,5.3269467,5.191132,4.9760923,4.7308717,4.4630156,4.183841,3.904667,3.6330378,3.4029078,3.3312278,3.338773,3.4594972,3.6179473,3.6330378,1.2223305,1.1846043,1.2034674,1.177059,1.0902886,1.0374719,1.569412,2.173032,2.1541688,1.5882751,1.3166461,1.6561824,2.4823873,3.451952,4.376245,5.2288585,6.2436943,6.217286,5.6551647,4.9647746,4.45547,3.8820312,3.259548,3.1124156,3.4368613,3.6971724,3.5500402,2.9766011,2.2786655,1.8184053,2.0447628,3.893349,5.594803,6.571913,7.01331,7.888559,10.672756,12.774108,13.766309,13.79649,13.58145,11.955449,10.137043,8.533678,7.5792036,7.7150183,8.062099,7.6282477,7.152897,6.832224,6.356873,5.1232247,4.1310244,3.3350005,2.848332,2.9351022,3.0935526,3.150142,3.0030096,2.9615107,3.7273536,2.8822856,2.6521554,2.6634734,2.6483827,2.4559789,3.0897799,3.863168,4.115934,3.6934,2.9539654,2.6672459,3.4934506,3.821669,3.5123138,3.8971217,3.3727267,3.2142766,3.6896272,4.4705606,4.5988297,4.4101987,4.164978,3.62172,2.8596497,2.2598023,2.3088465,2.1541688,2.3013012,2.837014,3.440634,2.776652,1.81086,1.5769572,2.1881225,2.8143783,3.127506,3.259548,3.1010978,2.7238352,2.384299,2.3503454,2.161714,1.5656394,0.79602385,0.58098423,0.35462674,0.29426476,0.29803738,0.30935526,0.32067314,0.5583485,0.754525,0.9016574,0.9808825,0.91674787,0.8262049,0.875249,0.875249,0.76584285,0.6149379,0.5772116,0.6375736,0.754525,0.7696155,0.422534,0.45648763,0.5281675,0.5696664,0.55457586,0.482896,0.56589377,0.5093044,0.39989826,0.30181,0.21881226,0.1358145,0.120724,0.11317875,0.08677038,0.08677038,0.1358145,0.23767537,0.27540162,0.2263575,0.150905,0.10940613,0.1358145,0.19240387,0.23013012,0.16976812,0.124496624,0.120724,0.15845025,0.24899325,0.4074435,0.6375736,0.8903395,1.1355602,1.3920987,1.7240896,2.546522,2.5012503,2.4295704,2.9124665,4.3121104,5.172269,4.8063245,4.168751,3.9159849,4.398881,3.9763467,3.4972234,3.3312278,3.2633207,2.516341,3.0671442,2.6295197,1.7995421,1.0902886,0.9318384,1.1317875,1.3430545,1.5128226,1.6109109,1.6524098,1.6524098,1.5279131,1.3053282,1.0789708,0.9922004,0.8903395,0.77338815,0.7507524,0.8186596,0.84129536,0.76584285,0.67152727,0.58475685,0.5055317,0.41121614,0.22258487,0.120724,0.08677038,0.094315626,0.10940613,0.120724,0.38480774,0.5583485,0.6111652,0.8111144,1.1393328,1.2147852,1.1204696,0.90920264,0.6073926,0.33953625,0.14713238,0.056589376,0.0754525,0.1659955,0.041498873,0.011317875,0.07922512,0.16976812,0.10940613,0.2565385,0.23013012,0.13958712,0.049044125,0.0,0.0,0.030181,0.033953626,0.00754525,0.00754525,0.018863125,0.030181,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.06790725,0.1961765,0.41121614,0.27917424,0.1056335,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.05281675,0.090543,0.13204187,0.15845025,0.12826926,0.120724,0.181086,0.23013012,0.23013012,0.17731337,0.19994913,0.3470815,0.43007925,0.43385187,0.49421388,0.5055317,0.482896,0.40367088,0.28294688,0.18485862,0.1056335,0.071679875,0.0754525,0.10940613,0.1659955,0.18863125,0.1659955,0.13958712,0.14335975,0.23013012,0.24522063,0.22258487,0.22258487,0.3169005,0.5772116,1.2411937,2.2975287,3.199186,3.5500402,3.1124156,2.9237845,3.229367,3.5085413,3.7084904,4.236658,4.1197066,4.172523,4.8402777,6.013564,7.0284004,6.598321,5.172269,4.266839,4.745962,6.8133607,7.5188417,9.005256,10.751981,12.370438,13.58145,15.022593,13.355092,11.491416,9.955957,6.900131,5.6589375,6.379509,8.09228,9.899368,11.00852,9.114662,7.17176,5.4212623,3.9650288,2.7351532,2.022127,1.4675511,1.0638802,0.814887,0.69793564,0.6073926,0.5319401,0.482896,0.44139713,0.36971724,0.2867195,0.2678564,0.33576363,0.4376245,0.47535074,0.41876137,0.29803738,0.23390275,0.24522063,0.271629,0.24522063,0.3169005,0.38480774,0.36594462,0.19994913,0.18863125,0.16222288,0.15467763,0.18485862,0.2263575,0.2565385,0.331991,0.47157812,0.59607476,0.5470306,0.6111652,0.68661773,0.77338815,0.9318384,1.2826926,1.8561316,1.8863125,1.6448646,1.4373702,1.5920477,1.4298248,1.1883769,0.94692886,0.77338815,0.72811663,0.73566186,0.7884786,0.9507015,1.1808317,1.327964,1.2751472,1.20724,1.1393328,1.1506506,1.4034165,1.5128226,1.3053282,1.448688,1.9655377,2.2258487,2.3428001,3.3350005,4.7421894,6.0211096,6.5530496,6.5756855,6.5002327,6.0022464,5.149633,4.406426,3.6971724,3.3123648,3.0822346,2.9652832,3.029418,3.5160866,4.478106,5.836251,7.3981175,8.83926,10.231359,11.208468,11.6875925,11.68382,11.332966,11.144334,10.989656,10.921749,10.804798,10.291721,8.20546,7.5905213,7.84706,8.371455,8.537451,9.1976595,10.054046,10.895341,11.721546,12.770335,14.64533,15.497944,15.445127,14.181297,10.944386,12.083718,12.702429,12.50248,11.759273,11.302785,12.034674,12.155397,12.117672,12.279895,12.917468,14.264296,14.498198,14.792462,15.4074,15.660167,16.961721,18.451908,18.85558,17.972786,16.675003,15.648849,15.098045,14.5132885,13.7700815,13.12119,14.158662,15.573396,16.644821,16.55428,14.366156,10.974566,8.27714,6.485142,5.696664,5.8928404,6.296511,6.0626082,5.3910813,4.425289,3.229367,2.2711203,1.6146835,1.1431054,0.8186596,0.7092535,0.573439,0.44139713,0.36594462,0.3470815,0.3470815,0.3961256,0.41498876,0.422534,0.41121614,0.3734899,0.3961256,0.41498876,0.47535074,0.5696664,0.62248313,0.58098423,0.5093044,0.4376245,0.3961256,0.38858038,0.38103512,0.41121614,0.4979865,0.6111652,0.66020936,0.7469798,0.875249,1.1129243,1.5882751,2.4974778,2.7879698,2.6332922,2.4333432,2.3390274,2.293756,2.686109,3.240685,3.5387223,3.4444065,3.1161883,3.4029078,3.4217708,3.5387223,3.863168,4.2706113,4.168751,3.8065786,3.3689542,3.1237335,3.440634,3.7198083,3.874486,4.115934,4.3800178,4.3649273,4.45547,3.9574835,3.3953626,3.150142,3.4142256,4.52715,6.752999,10.653893,16.361876,23.578907,27.242125,24.703148,20.028866,16.433554,16.28265,19.07062,21.104065,22.409393,23.8279,27.008223,30.445084,33.938534,36.36056,37.477257,37.933743,38.526047,39.548428,40.446312,40.567036,39.13344,36.960407,35.42495,34.72324,34.859055,35.624897,35.417404,35.236317,35.9003,37.096222,37.348988,36.37942,35.02128,33.229282,31.354286,30.139502,28.14001,26.219744,24.076893,21.835953,20.036411,19.153618,18.738628,18.519815,18.414183,18.546225,17.20317,15.339493,13.185325,11.0613365,9.371201,8.062099,7.145352,6.4436436,5.8664317,5.383536,5.372218,5.3382645,5.2628117,5.1345425,4.949684,4.6818275,4.3686996,4.006528,3.6330378,3.3048196,3.0935526,3.0256453,3.0897799,3.218049,3.289729,1.1996948,0.9922004,0.8186596,0.6752999,0.6526641,0.94315624,1.5279131,1.7278622,1.5769572,1.3241913,1.4298248,1.8448136,2.5540671,3.2821836,3.8895764,4.3686996,5.032682,5.2892203,5.194905,4.9421387,4.8666863,4.4931965,3.9159849,3.6141748,3.7386713,4.0970707,3.8065786,3.1425967,2.463524,2.2183034,2.9501927,6.828451,8.360137,8.45068,8.099826,8.420499,10.834979,12.245941,13.245687,13.754991,13.030646,10.235131,8.322411,6.9982195,6.273875,6.4474163,7.3717093,7.7640624,7.7187905,7.0585814,5.342037,4.6742826,4.5196047,4.429062,4.093298,3.338773,2.9200118,2.7125173,2.9464202,3.6745367,4.7648253,3.6594462,2.9992368,2.9766011,3.2784111,3.0860074,3.0407357,3.5651307,3.682082,3.3350005,3.410453,3.6783094,4.1989317,4.4403796,4.708236,6.1644692,6.470052,6.168242,5.726845,5.1798143,4.1197066,6.0022464,5.7381625,4.7346444,3.802806,3.138824,2.5314314,2.3503454,2.4484336,2.6785638,2.897376,2.6710186,2.1654868,1.6976813,1.569412,2.093807,2.7011995,3.0105548,2.9841464,2.6898816,2.2711203,2.3428001,2.335255,1.9957186,1.3543724,0.7432071,0.7922512,0.663982,0.5055317,0.40367088,0.35462674,0.482896,0.543258,0.60362,0.65643674,0.6149379,0.5394854,0.5998474,0.62248313,0.55080324,0.452715,0.4979865,0.6073926,0.7167987,0.724344,0.513077,0.68661773,0.6790725,0.5583485,0.41498876,0.35462674,0.40367088,0.35839936,0.2867195,0.22258487,0.1659955,0.124496624,0.1358145,0.1358145,0.116951376,0.10940613,0.16222288,0.2867195,0.35085413,0.32821837,0.29426476,0.27540162,0.29049212,0.32067314,0.31312788,0.18485862,0.27917424,0.27540162,0.2565385,0.2867195,0.4074435,0.58475685,0.80734175,1.1921495,1.7165444,2.1843498,2.3088465,2.093807,2.0900342,2.5238862,3.308592,3.5651307,3.2784111,3.429316,3.983892,3.8858037,4.90064,5.0968165,4.504514,3.8556228,4.5950575,3.6066296,2.505023,1.5618668,0.965792,0.8262049,0.9242931,1.0751982,1.2147852,1.3241913,1.4109617,1.4335974,1.3355093,1.1204696,0.875249,0.7507524,0.66020936,0.59607476,0.6111652,0.7054809,0.8526133,1.1091517,1.116697,0.86770374,0.48666862,0.23013012,0.1056335,0.041498873,0.018863125,0.026408374,0.056589376,0.14713238,0.271629,0.31312788,0.32067314,0.5017591,0.8563859,1.0299267,0.935611,0.7507524,0.9016574,0.77338815,0.42630664,0.150905,0.06413463,0.08677038,0.20749438,0.22258487,0.33576363,0.543258,0.63002837,1.3770081,1.1053791,0.5319401,0.1056335,0.0,0.0,0.0150905,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.033953626,0.026408374,0.041498873,0.041498873,0.03772625,0.05281675,0.124496624,0.2678564,0.16976812,0.0754525,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.056589376,0.120724,0.19240387,0.22258487,0.120724,0.08299775,0.1056335,0.150905,0.19994913,0.24899325,0.1358145,0.09808825,0.116951376,0.16222288,0.22258487,0.32444575,0.32067314,0.27917424,0.23013012,0.15845025,0.071679875,0.090543,0.094315626,0.07922512,0.15845025,0.18863125,0.16976812,0.1659955,0.17731337,0.14335975,0.120724,0.1056335,0.10940613,0.15467763,0.27917424,1.3015556,2.0070364,2.2560298,2.0485353,1.539231,1.3128735,1.5316857,1.8184053,2.052308,2.3578906,2.4069347,2.9916916,4.983638,7.281166,6.802043,5.907931,5.6551647,4.8930945,3.8971217,4.3611546,6.3908267,9.246704,12.106354,13.9888935,13.758763,12.762791,11.744182,11.446144,11.34051,9.612649,5.8890676,4.7912335,6.571913,10.227587,13.50977,14.867915,14.524607,12.955194,10.461489,7.145352,4.5497856,2.776652,1.7882242,1.3543724,1.0450171,0.87147635,0.76584285,0.7205714,0.69039035,0.6187105,0.47912338,0.38103512,0.35085413,0.35839936,0.32821837,0.23767537,0.18863125,0.18863125,0.23013012,0.24899325,0.21503963,0.23013012,0.271629,0.28294688,0.17731337,0.23013012,0.29049212,0.30181,0.24899325,0.1961765,0.181086,0.19994913,0.241448,0.30935526,0.41121614,0.80356914,0.8224323,0.88279426,1.1732863,1.6524098,1.8674494,1.8146327,1.6712729,1.5920477,1.7014539,1.5769572,1.3732355,1.177059,1.0374719,0.9808825,1.0110635,1.0902886,1.2185578,1.3091009,1.2034674,1.0299267,0.94692886,0.9507015,1.0638802,1.3355093,1.569412,1.5618668,2.0447628,3.0218725,3.7462165,3.5123138,3.9273026,4.5120597,5.194905,6.300284,6.8359966,6.089017,5.1345425,4.6327834,4.798779,4.606375,4.4894238,4.696918,5.0062733,4.7233267,4.5837393,5.1647234,6.2625575,7.6810646,9.239159,10.751981,11.574413,12.200669,12.721292,12.830698,12.559069,12.510024,13.309821,14.532151,14.68683,12.721292,10.650121,9.529651,9.559832,10.069136,10.435081,11.465008,12.725064,13.788944,14.245432,18.052011,18.980076,17.942604,15.230087,10.518079,9.740918,10.408672,11.174516,11.52537,11.774363,11.864905,12.174261,12.283667,12.23085,12.513797,14.124708,14.947141,15.497944,15.860115,15.660167,16.682549,17.569115,17.437073,16.158154,14.366156,13.747445,13.211733,12.585477,11.921495,11.476325,12.196897,13.340002,14.196388,14.3095665,13.472044,11.608367,9.469289,7.4811153,6.0512905,5.5759397,5.409944,4.8553686,4.0782075,3.1916409,2.2371666,1.5128226,0.9922004,0.59230214,0.331991,0.32067314,0.30181,0.30181,0.331991,0.3772625,0.3961256,0.34330887,0.34330887,0.3961256,0.46026024,0.45648763,0.3961256,0.38103512,0.43007925,0.52062225,0.58098423,0.513077,0.452715,0.4376245,0.44516975,0.39989826,0.36594462,0.3734899,0.43385187,0.52062225,0.573439,0.66775465,0.8111144,1.0525624,1.4675511,2.1541688,2.6446102,2.9200118,3.0331905,3.0181,2.9237845,3.078462,3.350091,3.3727267,3.138824,2.9954643,3.3274553,3.4217708,3.4066803,3.470815,3.893349,4.085753,4.025391,3.7273536,3.2633207,2.757789,3.2821836,3.380272,3.2105038,2.9200118,2.6295197,2.6031113,2.6936543,2.8558772,3.1010978,3.4783602,4.3347464,5.7419353,8.386545,12.58925,18.297232,22.4773,22.299986,19.134754,15.218769,13.679539,14.939595,16.659912,18.580177,20.919205,24.371157,29.04544,33.72727,36.986816,38.239326,37.733795,35.5834,34.025307,32.87088,31.90509,30.88648,30.475266,30.535627,31.60328,33.712177,36.371876,36.126656,35.191048,34.945824,35.779575,37.115086,36.122883,34.73456,33.263233,32.169174,32.071087,30.501673,28.219234,25.763256,23.507227,21.647322,19.749691,18.723537,18.006739,17.384256,16.969267,15.977067,14.781145,13.332457,11.736636,10.284176,8.993938,7.9262853,7.069899,6.405917,5.9003854,5.7570257,5.613666,5.4401255,5.2062225,4.9044123,4.568649,4.22534,3.8820312,3.561358,3.2821836,3.0671442,2.9124665,2.886058,2.9539654,3.0030096,0.80356914,0.62625575,0.47912338,0.47912338,0.69039035,1.1393328,1.4034165,1.2034674,1.1016065,1.3845534,2.093807,2.6106565,2.9501927,3.1199608,3.229367,3.4896781,3.7952607,4.1762958,4.4139714,4.5007415,4.617693,4.52715,4.191386,4.055572,4.3347464,5.0213637,4.4630156,3.663219,3.0709167,3.150142,4.3611546,8.492179,10.235131,9.846551,8.4544525,8.043237,9.167479,9.601331,9.827688,9.812597,9.009028,7.1340337,6.326692,6.0022464,5.66271,4.9157305,6.375736,7.194396,7.2396674,6.379509,4.447925,4.3913355,5.081726,5.59103,5.409944,4.45547,3.9989824,3.874486,3.9989824,4.3422914,4.9534564,4.5988297,4.4630156,4.6554193,5.243949,6.2663302,5.696664,5.191132,4.561104,3.9084394,3.640583,3.7877154,4.221567,4.870459,5.855114,7.496206,8.375228,7.0812173,5.270357,3.8065786,2.7728794,5.281675,5.2854476,4.3913355,3.519859,2.8822856,2.161714,2.1466236,2.3314822,2.4484336,2.4823873,2.5238862,2.3616633,1.780679,1.1129243,1.2638294,1.9806281,2.493705,2.6634734,2.4823873,2.0862615,2.5880208,2.5502944,2.2899833,2.0447628,1.9655377,3.006782,3.0709167,2.3277097,1.237421,0.55457586,0.41498876,0.3961256,0.44139713,0.47157812,0.392353,0.3772625,0.43007925,0.452715,0.41498876,0.3470815,0.44894236,0.58475685,0.6752999,0.6828451,0.5998474,0.7997965,0.7432071,0.5470306,0.33953625,0.24899325,0.27540162,0.29049212,0.30181,0.30181,0.27917424,0.27917424,0.331991,0.3055826,0.20749438,0.1961765,0.24522063,0.36971724,0.5093044,0.5696664,0.4376245,0.41498876,0.482896,0.55457586,0.51684964,0.21881226,0.27917424,0.27917424,0.29049212,0.3961256,0.68661773,1.1242423,1.3166461,1.7580433,2.474842,3.0407357,3.0746894,2.9011486,2.3918443,1.7278622,1.3920987,1.1355602,1.1129243,1.8146327,2.7502437,2.4522061,3.802806,4.538468,4.3724723,3.942393,4.798779,2.7351532,1.539231,0.94315624,0.7432071,0.80734175,0.7809334,1.0450171,1.2336484,1.2185578,1.146878,1.0978339,1.0789708,0.9318384,0.69793564,0.63002837,0.56212115,0.5017591,0.52062225,0.66020936,0.91674787,1.1619685,1.1695137,0.9318384,0.5281675,0.11317875,0.041498873,0.011317875,0.0,0.003772625,0.018863125,0.09808825,0.14335975,0.392353,0.77338815,0.8903395,0.573439,0.5357128,0.52439487,0.5394854,0.8563859,0.875249,0.6375736,0.331991,0.09808825,0.018863125,0.19240387,0.22258487,0.29803738,0.4678055,0.62625575,1.2600567,1.0035182,0.482896,0.10186087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.0452715,0.041498873,0.07922512,0.0754525,0.06790725,0.090543,0.16222288,0.116951376,0.05281675,0.041498873,0.056589376,0.00754525,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.033953626,0.033953626,0.041498873,0.094315626,0.17354076,0.2263575,0.17354076,0.16976812,0.19240387,0.2263575,0.2565385,0.29049212,0.181086,0.1358145,0.13958712,0.14713238,0.094315626,0.15845025,0.150905,0.14713238,0.17354076,0.1961765,0.1056335,0.124496624,0.11317875,0.071679875,0.120724,0.14335975,0.150905,0.16976812,0.181086,0.120724,0.10186087,0.06413463,0.049044125,0.07922512,0.12826926,0.9205205,1.2298758,1.1581959,0.88279426,0.6451189,0.3734899,0.35839936,0.5017591,0.69793564,0.8563859,1.1393328,1.9051756,4.515832,7.9338303,8.726082,5.7494807,5.798525,5.3382645,3.610402,2.6332922,4.678055,8.088508,11.642321,13.758763,12.528888,9.906913,9.559832,11.419736,13.6682205,12.73261,9.016574,6.802043,6.79827,8.643084,10.910432,14.849052,16.908905,17.47857,16.644821,14.18507,8.892077,5.2854476,3.2331395,2.305074,1.7391801,1.3619176,1.2336484,1.2600567,1.2902378,1.1506506,0.8639311,0.6111652,0.4376245,0.33576363,0.271629,0.16976812,0.13958712,0.17731337,0.26408374,0.38480774,0.32821837,0.2565385,0.21503963,0.19240387,0.13958712,0.19994913,0.29426476,0.32821837,0.2867195,0.23013012,0.1961765,0.21503963,0.23767537,0.271629,0.36971724,0.76207024,0.7582976,0.754525,0.935611,1.2600567,1.3166461,1.4109617,1.5807298,1.7995421,1.9881734,1.750498,1.5731846,1.4864142,1.4826416,1.5241405,1.4298248,1.3958713,1.3807807,1.3166461,1.0940613,0.845068,0.8262049,0.9016574,1.0487897,1.358145,1.6788181,1.8938577,2.6106565,3.7613072,4.606375,4.315883,4.2064767,4.0895257,4.45547,6.458734,7.2396674,6.439871,5.4778514,5.198677,5.8928404,5.553304,5.4891696,6.047518,6.907676,7.092535,6.862405,6.930312,7.2623034,7.9413757,9.175024,10.480352,11.510279,13.585222,15.875206,15.388537,14.128481,13.298503,13.45318,14.554788,15.977067,14.913187,13.43809,12.921241,13.547497,14.298248,12.528888,12.687338,13.834216,15.056546,15.471535,18.214233,20.013775,19.791191,17.078674,12.019584,9.2844305,8.91094,9.49947,10.099318,10.197406,9.971047,10.816116,11.932813,12.725064,12.830698,14.298248,15.69412,16.712729,17.078674,16.539188,16.18456,15.63753,14.841507,13.822898,12.702429,12.253486,11.465008,10.665211,10.133271,10.121953,10.785934,11.604594,12.268577,12.725064,13.158916,12.872196,11.544232,9.288202,6.8133607,5.406172,4.534695,3.682082,2.897376,2.1956677,1.5543215,1.1883769,0.875249,0.62248313,0.47157812,0.5281675,0.59230214,0.5696664,0.5017591,0.43385187,0.3772625,0.30181,0.29049212,0.3470815,0.4376245,0.513077,0.49044126,0.49421388,0.5093044,0.51684964,0.48666862,0.44139713,0.4074435,0.3961256,0.3961256,0.34330887,0.32067314,0.30935526,0.32821837,0.38103512,0.45648763,0.59607476,0.7582976,0.965792,1.2449663,1.6109109,2.1692593,2.8747404,3.5500402,3.9688015,3.832987,3.5274043,3.4481792,3.5839937,3.7575345,3.6066296,3.4368613,3.229367,3.0105548,2.9426475,3.2821836,3.5953116,3.5689032,3.289729,2.8181508,2.2107582,2.7351532,2.7502437,2.5201135,2.3013012,2.3201644,2.6446102,2.7691069,3.0331905,3.482133,3.85185,4.4101987,5.1760416,6.485142,8.869441,13.026875,17.297485,19.25925,18.357594,15.335721,12.242168,12.393073,14.083209,16.493916,19.236614,22.36412,28.668177,32.648296,34.73833,35.2665,34.444065,31.848501,30.02255,28.279596,26.438557,24.85028,24.280615,24.58997,26.627188,30.358313,34.832645,36.1757,36.00216,35.289135,34.972233,35.979527,35.70035,34.583652,33.116104,31.93527,31.825865,30.675215,28.939806,27.03463,25.155863,23.29596,21.115381,19.557287,18.13878,16.791954,15.871433,15.24895,14.509516,13.585222,12.47607,11.249968,10.065364,8.986393,8.028146,7.2358947,6.6662283,6.2927384,5.9494295,5.583485,5.168496,4.7044635,4.3309736,3.9876647,3.6896272,3.4330888,3.2067313,3.0445085,2.9086938,2.8407867,2.8294687,2.795515,0.24899325,0.2678564,0.38858038,0.6752999,1.0676528,1.3505998,1.2638294,1.0186088,1.1053791,1.690136,2.6106565,3.2218218,3.3123648,3.1350515,3.0218725,3.3878171,3.7198083,4.0480266,4.3800178,4.640329,4.659192,4.678055,4.5120597,4.61392,5.100589,5.775889,4.9647746,4.146115,3.7386713,4.014073,5.1269975,7.5263867,9.680555,9.574923,7.533932,6.224831,6.0248823,5.836251,5.379763,4.8666863,5.0025005,5.142088,5.511805,5.994701,5.9305663,4.1083884,6.039973,6.571913,6.1795597,5.372218,4.719554,5.4740787,6.4210076,6.8171334,6.3719635,5.2628117,5.062863,5.541986,5.80607,5.847569,6.537959,6.647365,6.851087,6.7643166,6.964266,9.001483,8.4544525,7.3717093,6.398372,5.5268955,4.1197066,3.6179473,4.266839,5.5193505,6.858632,7.7716074,8.201687,5.5495315,2.837014,1.5618668,1.7127718,2.6408374,2.8030603,2.516341,2.0447628,1.5882751,1.4713237,1.6184561,1.7844516,1.8599042,1.9089483,2.1466236,2.0787163,1.6184561,0.9808825,0.663982,1.0978339,1.6750455,2.0636258,2.1051247,1.8448136,2.7804246,2.6974268,2.41448,2.5389767,3.470815,5.4250345,5.9984736,4.8930945,2.7841973,1.3015556,0.754525,0.5470306,0.4979865,0.47157812,0.38858038,0.36594462,0.41498876,0.47157812,0.47535074,0.38103512,0.4074435,0.51684964,0.63002837,0.6790725,0.59607476,0.66020936,0.5885295,0.44894236,0.30935526,0.2263575,0.31312788,0.39989826,0.47535074,0.543258,0.60362,0.7092535,0.845068,0.7205714,0.44139713,0.5017591,0.5281675,0.7432071,1.1091517,1.3091009,0.7394345,0.9695646,1.2223305,1.3128735,1.0714256,0.362172,0.13958712,0.13204187,0.26031113,0.5093044,0.9393836,1.8221779,2.2748928,2.4333432,2.5012503,2.746471,3.1954134,3.731126,3.0822346,1.4713237,0.5998474,0.35839936,0.452715,0.8262049,1.2864652,1.4939595,1.7919968,2.323937,2.8898308,3.1727777,2.7125173,1.1808317,0.58098423,0.44516975,0.52439487,0.77338815,0.6790725,1.0676528,1.297783,1.1883769,0.9808825,0.87902164,0.9393836,0.8639311,0.67152727,0.69039035,0.6413463,0.5394854,0.5394854,0.68661773,0.9016574,0.8262049,0.7507524,0.68661773,0.5281675,0.06413463,0.02263575,0.003772625,0.0,0.00754525,0.033953626,0.15845025,0.26031113,0.77716076,1.4939595,1.5203679,0.4979865,0.150905,0.23013012,0.4979865,0.7130261,0.7997965,0.70170826,0.4376245,0.12826926,0.0,0.0,0.0,0.0,0.018863125,0.09808825,0.018863125,0.02263575,0.041498873,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0150905,0.041498873,0.041498873,0.02263575,0.00754525,0.0150905,0.03772625,0.0452715,0.090543,0.07922512,0.08299775,0.14335975,0.271629,0.1056335,0.08299775,0.07922512,0.0452715,0.026408374,0.0150905,0.02263575,0.0150905,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.003772625,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.049044125,0.049044125,0.018863125,0.026408374,0.07922512,0.15845025,0.23013012,0.2867195,0.35839936,0.4074435,0.41498876,0.38480774,0.43007925,0.43007925,0.42630664,0.3772625,0.17731337,0.090543,0.06790725,0.08299775,0.124496624,0.18485862,0.12826926,0.11317875,0.10940613,0.090543,0.06790725,0.071679875,0.124496624,0.16976812,0.19994913,0.23767537,0.19240387,0.09808825,0.06413463,0.116951376,0.19994913,0.26408374,0.29049212,0.2565385,0.2263575,0.392353,0.25276586,0.1659955,0.1659955,0.23767537,0.32821837,0.573439,1.0676528,3.0030096,6.4738245,10.499215,6.5832305,6.0022464,5.372218,3.7273536,2.5125682,3.0143273,5.7381625,9.193887,11.589504,10.823661,8.7600355,8.511042,11.042474,14.286931,13.132507,12.536433,11.548005,10.001229,8.375228,7.7904706,10.910432,13.551269,16.13929,18.576405,20.270313,13.822898,8.635539,5.198677,3.4255435,2.6597006,2.0598533,1.8787673,1.9391292,1.9957186,1.7467253,1.3241913,0.94692886,0.6451189,0.422534,0.26408374,0.17731337,0.17731337,0.29426476,0.51684964,0.7696155,0.6752999,0.52439487,0.36594462,0.24522063,0.17731337,0.17731337,0.17731337,0.19240387,0.21881226,0.23013012,0.23767537,0.29426476,0.32444575,0.3169005,0.33953625,0.38858038,0.422534,0.40367088,0.3772625,0.46026024,0.6790725,1.0450171,1.4600059,1.8485862,2.1805773,1.8372684,1.6712729,1.6712729,1.8033148,1.9957186,1.7844516,1.569412,1.3807807,1.2034674,0.9620194,0.724344,0.8186596,0.97333723,1.1393328,1.5052774,1.9202662,2.2371666,2.9615107,3.9876647,4.6252384,4.425289,4.187614,4.1498876,4.938366,7.54525,8.160188,8.039464,7.635793,7.4018903,7.816879,6.8473144,6.5341864,6.903904,7.77538,8.75249,9.291975,8.99771,8.329956,8.035691,9.171251,10.502988,11.879996,15.286676,19.032892,17.769064,15.430037,13.355092,11.774363,11.3971,13.396591,12.955194,13.664448,15.23386,17.067356,18.263277,14.913187,14.3095665,14.849052,15.422491,15.422491,14.735873,16.380737,17.618158,17.022083,14.445381,10.401127,8.639311,8.446907,8.858124,8.616675,8.858124,10.250222,12.306303,14.064346,14.117163,15.437581,17.08999,18.451908,18.934805,18.002966,15.961976,13.902123,12.449662,11.781908,11.61214,10.95193,10.050273,9.386291,9.22784,9.635284,10.510533,11.102836,11.638548,12.306303,13.275867,13.6833105,12.947649,10.650121,7.5226145,5.4212623,4.1008434,3.150142,2.4559789,1.9278114,1.478869,1.4298248,1.3430545,1.2562841,1.1959221,1.177059,1.1317875,0.9280658,0.67152727,0.44516975,0.3169005,0.30935526,0.3055826,0.32821837,0.3772625,0.47535074,0.5885295,0.66020936,0.6526641,0.5696664,0.44139713,0.49044126,0.48666862,0.41876137,0.3169005,0.26408374,0.2678564,0.25276586,0.24899325,0.2867195,0.3772625,0.55080324,0.7167987,0.88279426,1.0751982,1.3392819,1.7919968,2.584248,3.7009451,4.678055,4.5912848,4.006528,3.8971217,4.61392,5.541986,5.1081343,4.142342,3.308592,2.795515,2.6332922,2.6634734,2.795515,2.5917933,2.2560298,1.9730829,1.9089483,2.0183544,2.1466236,2.3314822,2.686109,3.3651814,4.236658,3.9876647,3.7990334,4.0480266,4.304565,4.610148,4.881777,4.957229,5.6023483,8.503497,12.30253,15.16218,16.331694,15.335721,11.981857,11.966766,13.604086,15.961976,18.45568,20.847527,27.555252,29.732058,29.826374,29.256706,28.407866,27.027086,26.317833,25.144547,23.280869,21.424738,19.960958,19.606333,21.236107,24.884235,29.747149,33.68577,35.975754,36.537872,35.911617,35.27027,35.477764,34.911873,33.51977,31.79191,30.735577,29.550972,28.622906,27.56657,26.20088,24.525835,23.058285,21.322876,19.247932,17.222033,16.109108,15.784663,15.32063,14.683057,13.819125,12.683565,11.4838705,10.295494,9.171251,8.175279,7.352846,6.7341356,6.2135134,5.723072,5.198677,4.5837393,4.2064767,3.8820312,3.5953116,3.3274553,3.0746894,2.9501927,2.9011486,2.8596497,2.7879698,2.6672459,0.27540162,0.45648763,0.6790725,0.87902164,1.0714256,1.327964,1.1808317,1.1242423,1.1732863,1.2336484,1.0978339,1.7580433,2.4069347,3.0860074,3.863168,4.851596,5.342037,5.59103,5.96452,6.4549613,6.700182,6.4436436,6.085244,5.6325293,5.040227,4.2102494,3.6745367,3.5839937,3.7801702,4.002755,3.904667,5.6513925,7.6282477,8.586494,8.009283,6.1041074,6.224831,6.228604,6.33801,6.8925858,8.345046,8.907167,7.9300575,6.387054,5.2175403,5.342037,8.160188,8.499724,7.91874,7.598067,8.329956,9.2844305,8.809079,8.265821,7.4584794,4.640329,4.1762958,5.8626595,8.60913,11.729091,14.939595,11.763044,8.635539,6.511551,5.8173876,6.439871,7.122716,7.284939,6.851087,5.96452,4.9760923,4.67051,5.4174895,6.9227667,8.552541,9.322156,7.7112455,5.413717,3.338773,2.1164427,2.0900342,2.7879698,3.361409,3.3463185,2.806833,2.3805263,2.233394,2.0673985,1.8599042,1.7278622,1.9240388,2.2748928,2.2748928,2.003264,1.6146835,1.297783,0.9318384,1.3241913,1.8146327,2.1353056,2.4408884,2.9313297,3.1539145,3.048281,2.7992878,2.8219235,3.6669915,4.798779,5.1647234,4.5761943,3.7084904,2.5729303,1.6109109,0.9205205,0.5696664,0.59607476,0.48666862,0.48666862,0.56589377,0.6488915,0.62625575,0.56589377,0.5017591,0.4376245,0.362172,0.29049212,0.362172,0.35462674,0.32444575,0.29803738,0.27540162,0.32444575,0.4376245,0.5998474,0.84884065,1.2525115,1.6788181,1.8485862,1.4750963,0.9393836,1.2826926,1.2336484,1.780679,2.6597006,3.0558262,1.6184561,2.9728284,3.6330378,3.4594972,2.4861598,0.9016574,0.26408374,0.20749438,0.40367088,0.6451189,0.8526133,1.4524606,3.9725742,4.38379,2.3201644,1.0978339,1.5882751,2.6898816,2.8181508,1.8561316,1.1581959,1.1355602,1.3015556,1.4373702,1.5203679,1.7391801,1.7165444,1.388326,0.9318384,0.5281675,0.38103512,0.28294688,0.27917424,0.31312788,0.36971724,0.44139713,0.56589377,0.5583485,0.5998474,0.7507524,0.94692886,1.056335,1.0450171,0.94315624,0.7884786,0.6413463,0.543258,0.5093044,0.5394854,0.58475685,0.5357128,0.4979865,0.44139713,0.362172,0.23390275,0.0150905,0.003772625,0.0,0.0,0.033953626,0.1659955,0.7432071,0.7582976,0.55080324,0.32444575,0.150905,0.116951376,0.16222288,0.22258487,0.45648763,1.2525115,1.3845534,0.6790725,0.10940613,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.07922512,0.19994913,0.19994913,0.11317875,0.0452715,0.033953626,0.071679875,0.1056335,0.08299775,0.041498873,0.0150905,0.0150905,0.0150905,0.0150905,0.2263575,0.2678564,0.11317875,0.0754525,0.06413463,0.033953626,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.00754525,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.03772625,0.060362,0.09808825,0.1358145,0.27917424,0.56589377,0.94692886,1.3619176,1.2713746,0.9808825,0.663982,0.3961256,0.21503963,0.11317875,0.071679875,0.06413463,0.0754525,0.0754525,0.08677038,0.07922512,0.056589376,0.030181,0.056589376,0.124496624,0.23390275,0.35839936,0.45648763,0.18863125,0.1056335,0.12826926,0.19994913,0.27540162,0.13958712,0.1056335,0.14335975,0.20749438,0.24522063,0.24522063,0.271629,0.30935526,0.32821837,0.3055826,0.55080324,0.91297525,1.3468271,2.516341,5.798525,7.7037,7.466025,5.5193505,3.169005,2.6106565,3.3651814,5.342037,7.3905725,8.737399,8.956212,7.432071,7.9753294,8.3525915,7.907422,7.5527954,9.359882,11.69891,13.264549,13.70972,13.626721,12.332711,11.057564,11.019837,13.298503,18.829172,16.716501,11.574413,6.8699503,4.255521,3.5839937,3.1350515,2.7917426,2.5238862,2.2598023,1.8938577,1.539231,1.3128735,1.0487897,0.70170826,0.33576363,0.19994913,0.3055826,0.6828451,1.146878,1.2826926,1.1581959,0.88279426,0.6149379,0.44516975,0.3961256,0.29803738,0.1659955,0.09808825,0.10940613,0.120724,0.1961765,0.241448,0.26408374,0.27917424,0.29049212,0.35085413,0.392353,0.47157812,0.6073926,0.77716076,0.80356914,1.1204696,1.3770081,1.4713237,1.5580941,1.5580941,1.5203679,1.478869,1.4939595,1.6788181,1.7882242,1.7429527,1.6373192,1.448688,1.0223814,0.76584285,0.77338815,1.0072908,1.3694628,1.7240896,2.1390784,2.5087957,3.0935526,3.942393,4.881777,4.357382,5.0515447,6.802043,8.854351,9.842778,9.439108,9.989911,10.427535,10.291721,9.718282,9.220296,8.737399,8.273367,7.9451485,7.9941926,9.473062,9.786189,8.952439,8.341274,10.695392,11.393328,12.068627,12.913695,14.1926155,16.28265,16.58446,15.290449,13.422999,11.747954,10.774617,9.590013,10.133271,11.046246,12.027128,13.8719425,16.007248,17.391802,17.89356,17.240896,15.045229,12.396846,10.872705,11.306557,13.532406,16.388283,13.200415,10.767072,10.26154,11.446144,12.679792,12.570387,13.091009,13.721037,14.177525,14.434063,16.535416,18.889534,20.251451,19.99114,18.112373,15.098045,12.411936,10.740664,10.012547,9.416472,8.854351,8.650629,9.0807085,9.952185,10.574668,10.95193,11.34051,11.714001,12.140307,12.785426,12.483616,11.287694,9.578695,7.6923823,5.934339,4.640329,3.6783094,2.9766011,2.5314314,2.3956168,2.7389257,2.7691069,2.5804756,2.203213,1.6184561,0.94692886,0.52062225,0.33953625,0.32821837,0.36594462,0.36594462,0.3734899,0.39989826,0.41498876,0.36594462,0.48666862,0.59230214,0.58475685,0.49044126,0.44139713,0.6375736,0.6790725,0.5998474,0.45648763,0.33576363,0.31312788,0.331991,0.35085413,0.36594462,0.42630664,0.56212115,0.7582976,0.9318384,1.0940613,1.388326,1.7542707,2.1466236,2.9728284,4.0782075,4.7610526,4.6742826,4.881777,5.726845,6.670001,6.3153744,5.1458607,4.0103,3.1425967,2.6031113,2.2748928,2.1013522,2.04099,1.9504471,1.7731338,1.5430037,1.8938577,2.8898308,3.731126,4.123479,4.255521,4.172523,4.2706113,4.3724723,4.4516973,4.6252384,4.719554,4.4818783,4.2291126,4.436607,5.7079816,7.2698483,9.0807085,11.09529,12.702429,12.725064,11.823407,12.54775,14.037937,15.546988,16.463736,17.931286,19.58747,20.470263,20.474035,20.341993,19.927006,19.655376,19.319613,19.04421,19.28566,18.470772,18.391546,18.62545,19.508244,22.156626,27.528845,32.95388,37.398033,39.529564,37.733795,36.00216,35.028824,34.03285,32.674706,31.052477,29.185026,28.049467,27.559025,27.24967,26.261242,25.650078,23.92976,21.488873,18.980076,17.320122,16.999449,17.40689,17.486116,16.807045,15.562078,13.86817,12.106354,10.453944,8.975075,7.643338,6.802043,6.3342376,6.0550632,5.692891,4.9119577,4.496969,4.1197066,3.7462165,3.3651814,2.9766011,2.8030603,2.7728794,2.757789,2.704972,2.595566,0.6526641,0.7469798,0.9318384,1.1280149,1.2826926,1.3656902,1.20724,1.0336993,1.0978339,1.4034165,1.7089992,2.0862615,2.5691576,3.1840954,3.8971217,4.6214657,5.409944,6.221059,7.1793056,7.937603,7.673519,6.549277,5.624984,5.2175403,5.1571784,4.7836885,4.961002,4.8440504,4.4931965,4.002755,3.5160866,4.293247,5.904158,7.001992,7.1378064,6.72659,7.7376537,7.5829763,7.0284004,6.930312,8.235641,9.424017,9.563604,8.311093,6.488915,6.0739264,6.6850915,6.620957,6.4926877,7.0849895,9.318384,10.310584,9.9257765,8.473316,6.515323,4.847823,3.2482302,5.402399,9.446653,13.641812,16.35433,13.373956,10.238904,7.541477,5.7117543,4.98741,5.7683434,6.1229706,6.258785,6.387054,6.7077274,6.881268,6.277648,5.907931,5.9003854,5.4778514,4.255521,3.2067313,3.2255943,4.5233774,6.6058664,6.571913,5.8513412,4.6742826,3.3727267,2.3805263,1.8221779,1.6146835,1.6373192,1.7769064,1.9353566,2.0447628,2.4069347,2.444661,2.04099,1.5279131,1.2487389,1.1883769,1.3204187,1.6109109,2.0145817,2.5201135,2.9049213,3.0746894,3.0558262,2.9803739,3.6783094,4.123479,3.5764484,2.3277097,1.6939086,3.0105548,3.2255943,2.5691576,1.539231,0.8865669,0.69039035,0.60362,0.663982,0.87147635,1.1883769,1.4977322,1.5052774,1.3656902,1.1732863,0.97333723,0.8224323,0.62625575,0.48666862,0.41498876,0.32444575,0.29426476,0.3734899,0.56589377,0.8224323,1.0299267,2.0145817,3.31991,4.6252384,5.251494,4.187614,3.3161373,2.8445592,2.5729303,2.2975287,1.8259505,2.3578906,2.4974778,2.282438,1.750498,0.9242931,0.29803738,0.14335975,0.17731337,0.29049212,0.5357128,0.9205205,1.4675511,1.539231,1.0902886,0.67152727,0.86770374,1.4637785,1.8825399,2.1466236,2.8558772,4.08198,4.357382,3.519859,2.2220762,1.9240388,1.9844007,1.8636768,1.5920477,1.2562841,1.0035182,0.935611,0.6526641,0.513077,0.63002837,0.87147635,0.9808825,0.8639311,0.90543,1.1883769,1.4826416,1.5543215,1.3807807,1.1355602,0.90543,0.69039035,0.543258,0.49044126,0.543258,0.67152727,0.7922512,0.5772116,0.39989826,0.29049212,0.24899325,0.23390275,0.51684964,0.47535074,0.29426476,0.120724,0.071679875,0.20372175,0.23390275,0.16976812,0.06413463,0.030181,0.02263575,0.1659955,0.25276586,0.26408374,0.33576363,0.29426476,0.1358145,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.02263575,0.02263575,0.0150905,0.026408374,0.026408374,0.049044125,0.08677038,0.08677038,0.060362,0.03772625,0.030181,0.03772625,0.033953626,0.018863125,0.0150905,0.0150905,0.018863125,0.041498873,0.041498873,0.06790725,0.06413463,0.03772625,0.041498873,0.018863125,0.00754525,0.02263575,0.03772625,0.0,0.030181,0.030181,0.018863125,0.011317875,0.003772625,0.011317875,0.041498873,0.0452715,0.011317875,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.011317875,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.08677038,0.21881226,0.422534,0.62625575,0.80734175,0.91297525,0.87147635,0.98465514,0.8224323,0.66020936,0.5885295,0.5055317,0.20749438,0.09808825,0.06413463,0.0452715,0.041498873,0.030181,0.02263575,0.0150905,0.0150905,0.018863125,0.033953626,0.056589376,0.094315626,0.15845025,0.27540162,0.19994913,0.150905,0.13204187,0.13958712,0.150905,0.116951376,0.120724,0.18863125,0.2867195,0.34330887,0.23390275,0.241448,0.29049212,0.32067314,0.3055826,0.422534,0.77716076,1.5316857,2.4861598,3.0633714,3.1539145,3.2142766,2.9237845,2.5616124,3.0256453,3.9650288,5.0062733,5.6891184,5.96452,6.187105,7.2585306,8.507269,8.971302,8.379,7.1868505,5.847569,6.571913,8.0206,9.344792,10.208723,11.227332,12.121444,13.275867,14.603831,15.531898,13.521088,10.95193,9.710737,9.767326,9.163706,6.903904,5.270357,3.9650288,2.916239,2.2598023,2.2748928,2.3163917,1.8636768,0.9997456,0.4074435,0.23390275,0.2263575,0.392353,0.65643674,0.87902164,0.79602385,0.73188925,0.69039035,0.66775465,0.6790725,0.5017591,0.3169005,0.20749438,0.17731337,0.15845025,0.16222288,0.17731337,0.23013012,0.331991,0.46026024,0.5885295,0.6149379,0.6111652,0.6451189,0.76584285,0.87902164,1.1280149,1.2789198,1.3166461,1.4713237,1.3430545,1.2261031,1.1393328,1.1506506,1.3732355,1.5618668,1.599593,1.6146835,1.6146835,1.50905,1.086516,1.026154,1.0978339,1.2525115,1.6260014,2.323937,3.7537618,5.3344917,6.175787,5.0553174,4.715781,6.096562,8.09228,9.944639,11.246195,10.091772,8.805306,8.065872,8.186596,9.0957985,10.578441,11.23865,11.415963,11.495189,11.876224,13.29473,11.932813,9.495697,7.424526,6.900131,7.0585814,7.7716074,8.763808,9.74469,10.386037,11.287694,12.351574,12.691111,12.351574,12.310076,10.442626,9.9257765,10.344538,10.95193,10.646348,13.604086,15.890297,17.425755,18.599041,20.270313,16.633503,14.747191,15.015047,16.859861,18.731083,16.912678,15.509261,15.098045,15.082954,13.679539,13.736128,13.95494,14.139798,14.252977,14.4114275,14.966003,15.377219,15.448899,14.9358225,13.536179,11.955449,10.77839,10.174769,9.865415,9.110889,7.99042,7.809334,8.348819,9.186342,9.684328,9.435335,9.359882,9.525878,9.989911,10.774617,11.133017,10.850069,9.767326,7.99042,5.9117036,4.3422914,3.289729,2.5125682,1.9768555,1.8221779,2.191895,2.41448,2.3277097,1.9429018,1.4449154,0.9205205,0.6526641,0.5281675,0.47912338,0.47535074,0.49421388,0.52439487,0.5281675,0.513077,0.513077,0.56589377,0.6149379,0.6526641,0.66775465,0.6488915,0.66020936,0.66020936,0.55080324,0.3772625,0.32444575,0.3470815,0.38103512,0.43385187,0.4979865,0.55080324,0.633801,0.80734175,0.98842776,1.2110126,1.6335466,1.7655885,1.9542197,2.41448,3.1312788,3.8443048,4.346064,4.7950063,5.4401255,6.115425,6.221059,5.5570765,4.738417,4.085753,3.651901,3.2255943,2.4899325,2.776652,3.1425967,3.1916409,3.0671442,2.8822856,3.772625,4.395108,4.3385186,4.112161,4.014073,4.014073,4.006528,4.036709,4.293247,4.3913355,4.2592936,4.0593443,4.1272516,4.98741,5.855114,6.8246784,8.171506,9.695646,10.736891,10.612394,11.570641,12.925014,13.917213,13.717264,13.317367,14.1926155,14.943368,15.192361,15.614895,16.373192,16.199652,15.897841,16.052519,17.029629,17.569115,18.504726,18.961214,18.859352,18.919714,21.371922,26.332922,31.99186,36.439785,37.662117,36.258698,35.077866,33.87063,32.542664,31.124157,29.501928,28.038149,26.872408,26.061293,25.601034,25.733074,24.699375,22.4358,19.749691,18.293459,17.625704,17.108854,16.769318,16.505234,16.101564,15.135772,13.86817,12.095036,10.050273,8.375228,7.2698483,6.6058664,6.1531515,5.7381625,5.2288585,4.8440504,4.5196047,4.217795,3.92353,3.610402,3.410453,3.3161373,3.2331395,3.0860074,2.837014,0.77338815,0.8865669,1.0148361,1.2034674,1.3920987,1.3920987,1.2261031,1.237421,1.4034165,1.6939086,2.082489,2.5238862,2.9652832,3.4444065,3.8556228,3.9122121,4.82896,6.0022464,7.356619,8.465771,8.560086,7.2698483,5.8966126,5.2288585,5.481624,6.273875,7.1906233,6.643593,5.8136153,5.221313,4.7346444,5.149633,7.8432875,9.25425,8.707218,8.439363,9.027891,8.7751255,7.4018903,6.3719635,8.888305,9.205205,8.386545,6.971811,5.7117543,5.5797124,5.4212623,5.492942,6.1078796,7.54525,10.061591,8.98262,7.7150183,6.2663302,4.8930945,4.08198,3.6896272,6.405917,10.065364,12.913695,13.59654,10.284176,8.213005,6.9227667,6.205968,6.1342883,6.4474163,5.80607,5.304311,5.4363527,6.096562,7.277394,7.484888,6.722818,5.2628117,3.6179473,2.5917933,2.837014,4.1989317,6.115425,7.643338,6.1644692,4.8553686,3.9273026,3.4444065,3.3425457,2.3013012,1.8599042,1.7995421,2.003264,2.4408884,2.9313297,2.9049213,2.493705,1.9278114,1.5430037,1.5430037,1.5958204,1.4109617,1.116697,1.2562841,1.8523588,2.3692086,2.5993385,2.7728794,3.561358,4.044254,3.8405323,3.0445085,2.2409391,2.516341,2.4597516,2.6785638,2.6597006,2.2183034,1.4750963,0.98465514,0.90920264,1.116697,1.5203679,2.1164427,2.7804246,3.0445085,2.8709676,2.4069347,1.9693103,1.6712729,1.4600059,1.3807807,1.3392819,1.1053791,1.026154,0.9695646,0.84129536,0.76207024,1.0601076,1.6750455,2.625747,3.6556737,4.22534,3.4670424,2.927557,2.372981,1.8221779,1.3317367,0.9997456,1.1016065,1.086516,0.9695646,0.76207024,0.4640329,0.19994913,0.17731337,0.18863125,0.18863125,0.27540162,0.41498876,0.452715,0.49421388,0.5394854,0.52062225,0.5885295,0.7432071,0.9242931,1.2902378,2.2183034,2.584248,2.5389767,2.1692593,1.8938577,2.463524,2.0485353,2.123988,2.191895,2.0447628,1.7731338,2.6785638,1.7354075,0.76207024,0.5017591,0.6375736,0.724344,0.7507524,0.9393836,1.3053282,1.6448646,1.690136,1.4411428,1.1619685,1.0374719,1.177059,0.9242931,0.6488915,0.65643674,0.935611,1.1846043,0.73566186,0.45648763,0.40367088,0.48666862,0.4640329,0.5696664,0.4640329,0.27917424,0.11317875,0.0452715,0.120724,0.10186087,0.0452715,0.0,0.0,0.23390275,0.41876137,0.663982,0.8299775,0.5357128,0.11317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.026408374,0.033953626,0.03772625,0.033953626,0.02263575,0.033953626,0.02263575,0.0150905,0.018863125,0.02263575,0.02263575,0.018863125,0.018863125,0.018863125,0.011317875,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.018863125,0.018863125,0.0150905,0.026408374,0.041498873,0.030181,0.0150905,0.00754525,0.018863125,0.026408374,0.0,0.0150905,0.0150905,0.0150905,0.0150905,0.00754525,0.00754525,0.030181,0.03772625,0.018863125,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.06790725,0.17354076,0.36594462,0.56212115,0.56212115,0.70170826,0.83752275,0.7582976,0.52062225,0.46026024,0.4376245,0.3470815,0.28294688,0.271629,0.241448,0.10940613,0.060362,0.0452715,0.03772625,0.041498873,0.056589376,0.056589376,0.05281675,0.0452715,0.05281675,0.041498873,0.033953626,0.033953626,0.05281675,0.10940613,0.10186087,0.07922512,0.06790725,0.0754525,0.0754525,0.08677038,0.116951376,0.19240387,0.27917424,0.31312788,0.32444575,0.38103512,0.44894236,0.5281675,0.62625575,0.59230214,0.65643674,0.9280658,1.2751472,1.3091009,1.6109109,2.1315331,2.916239,4.0216184,5.5268955,6.1418333,6.3116016,5.7570257,4.825187,4.459243,6.017337,7.594294,8.963757,10.186088,11.581959,10.736891,9.522105,7.865923,6.3644185,6.270103,7.0246277,8.194141,9.850324,11.695138,13.072145,13.132507,12.706201,12.808062,13.505998,13.947394,12.064855,10.401127,8.60913,6.696409,5.0062733,4.402653,4.0216184,3.0709167,1.6373192,0.6828451,0.35462674,0.23767537,0.23767537,0.33576363,0.59607476,0.5885295,0.5772116,0.67152727,0.8186596,0.8224323,0.6752999,0.5281675,0.44139713,0.4376245,0.48666862,0.4376245,0.3772625,0.35462674,0.43007925,0.63002837,0.8865669,0.87902164,0.7809334,0.7130261,0.73566186,0.87147635,1.056335,1.177059,1.20724,1.2110126,1.0902886,1.0676528,1.1129243,1.2034674,1.3317367,1.4600059,1.5580941,1.6561824,1.7014539,1.5241405,1.2789198,1.3204187,1.388326,1.4600059,1.7655885,2.8596497,4.3309736,5.907931,7.0284004,6.828451,6.115425,6.217286,7.17176,8.518587,9.288202,7.696155,7.250985,7.816879,9.0957985,10.63503,11.917723,12.004493,11.872451,12.019584,12.491161,13.947394,13.196642,10.868933,8.122461,6.6549106,6.006019,5.8400235,5.8173876,5.956975,6.6322746,7.7904706,9.208978,10.18986,10.63503,11.065109,11.465008,11.691365,11.434827,10.589758,9.265567,11.649866,13.79649,15.607349,17.372938,19.779873,18.71222,18.19537,18.519815,19.628967,21.122927,21.209698,21.047476,20.477808,19.28566,17.199398,15.452672,14.524607,14.11339,13.898351,13.536179,13.736128,13.898351,13.902123,13.600313,12.800517,11.77059,10.838752,10.1294985,9.5032425,8.5563135,7.4773426,7.232122,7.5716586,8.084735,8.197914,7.7225633,7.4207535,7.6395655,8.333729,9.06939,9.691874,9.891823,9.469289,8.311093,6.3908267,5.66271,5.032682,4.2706113,3.3764994,2.565385,2.191895,1.8636768,1.4826416,1.0751982,0.7922512,0.63002837,0.6073926,0.59607476,0.56589377,0.56589377,0.58475685,0.5772116,0.543258,0.5017591,0.47535074,0.44516975,0.49044126,0.5470306,0.59607476,0.6187105,0.6187105,0.59607476,0.52439487,0.4376245,0.4376245,0.41121614,0.42630664,0.5055317,0.6111652,0.6526641,0.66775465,0.7394345,0.8563859,1.0525624,1.4109617,1.7693611,1.9844007,2.4182527,3.2746384,4.5950575,5.7192993,5.7117543,5.7607985,6.066381,5.836251,5.0968165,4.587512,4.13857,3.6934,3.308592,3.1161883,3.4444065,3.8292143,3.9876647,3.832987,3.4783602,3.6066296,3.7386713,3.772625,3.9725742,3.9197574,3.8971217,3.8971217,3.953711,4.1008434,4.2064767,4.0895257,3.9876647,4.115934,4.659192,5.3269467,6.2097406,7.2094865,8.130007,8.699674,8.627994,9.224068,10.370946,11.532914,11.732863,11.52537,12.14408,12.808062,13.128735,13.124963,12.804289,12.325166,12.479843,13.521088,15.165953,16.29774,16.878725,16.984358,16.825907,16.739138,17.7502,21.104065,25.431265,29.494383,32.169174,32.78411,32.618114,31.871136,30.829891,29.87919,28.939806,27.672205,26.468737,25.476536,24.612606,24.454155,23.77131,22.379211,20.53817,18.987621,18.119919,17.4333,16.991903,16.648594,16.044973,16.007248,15.422491,14.068119,12.121444,10.144588,8.590267,7.5075235,6.760544,6.205968,5.6853456,5.372218,5.1571784,4.919503,4.610148,4.244203,3.9876647,3.893349,3.7462165,3.4594972,3.0897799,1.3920987,1.3468271,1.2336484,1.2562841,1.4600059,1.7316349,1.2902378,1.3807807,1.750498,2.2409391,2.776652,3.3236825,3.9159849,4.7308717,5.5080323,5.572167,4.870459,5.3344917,6.187105,6.937857,7.413208,6.94163,5.613666,4.749735,4.983638,6.2625575,7.360391,7.069899,6.9491754,7.111398,6.2436943,6.1908774,8.488406,9.933322,9.616421,8.914713,8.805306,8.578949,7.61693,7.0170827,9.593785,8.59404,7.281166,6.1229706,5.3873086,5.1081343,5.2137675,5.5797124,6.349328,7.462252,8.646856,6.5455046,5.0854983,4.617693,4.82896,4.749735,5.3646727,8.069645,10.646348,11.966766,11.989402,9.740918,8.914713,9.4127,10.487898,10.748209,9.842778,8.0206,6.488915,5.7909794,5.798525,8.028146,9.5183325,9.522105,8.065872,5.975838,4.0782075,4.168751,4.9760923,5.594803,5.50426,4.06689,3.0822346,2.7615614,3.0369632,3.572676,2.8747404,2.3956168,2.1654868,2.2899833,2.9313297,3.3727267,2.848332,2.082489,1.569412,1.5882751,2.3654358,3.169005,3.3689542,2.655928,1.0186088,1.2261031,1.6109109,1.9127209,2.3277097,3.5236318,4.0178456,3.4745877,2.5691576,1.9655377,2.3163917,1.8146327,1.7052265,1.8033148,1.8523588,1.5165952,1.1619685,1.0714256,1.2562841,1.6976813,2.3390274,3.0897799,3.531177,3.4481792,2.9313297,2.4031622,2.082489,1.9768555,2.1164427,2.3503454,2.372981,2.5125682,2.1881225,1.4335974,0.7432071,1.0940613,1.1317875,1.3543724,1.6448646,1.8221779,1.6373192,1.5845025,1.2826926,0.90543,0.56212115,0.30181,0.23390275,0.20749438,0.181086,0.14335975,0.09808825,0.08677038,0.16222288,0.21881226,0.24522063,0.32444575,0.5055317,0.66020936,0.6111652,0.44894236,0.52439487,0.98465514,1.4222796,1.7165444,1.7995421,1.6448646,1.0035182,0.66020936,0.6790725,1.086516,1.8787673,2.0258996,2.3503454,2.41448,2.123988,1.7354075,3.2029586,2.3767538,1.3166461,0.8865669,0.754525,0.5885295,0.58098423,0.79602385,1.1996948,1.6524098,1.720317,1.3694628,0.9997456,0.8978847,1.1846043,1.1506506,1.0827434,1.2298758,1.50905,1.4713237,1.2261031,0.995973,0.9620194,1.2902378,2.142851,1.2110126,0.6451189,0.33576363,0.18485862,0.11317875,0.124496624,0.15845025,0.30935526,0.5093044,0.5357128,0.35085413,0.35839936,0.56212115,0.7469798,0.49421388,0.1056335,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.0452715,0.041498873,0.026408374,0.02263575,0.0452715,0.049044125,0.033953626,0.018863125,0.011317875,0.00754525,0.00754525,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.033953626,0.02263575,0.02263575,0.026408374,0.02263575,0.011317875,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0452715,0.08677038,0.10186087,0.060362,0.02263575,0.003772625,0.003772625,0.00754525,0.02263575,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.041498873,0.090543,0.19994913,0.38858038,0.56212115,0.49421388,0.5319401,0.5696664,0.41498876,0.15845025,0.16222288,0.124496624,0.094315626,0.071679875,0.060362,0.041498873,0.041498873,0.03772625,0.049044125,0.0754525,0.11317875,0.10940613,0.11317875,0.1358145,0.15467763,0.124496624,0.08299775,0.0452715,0.026408374,0.030181,0.03772625,0.030181,0.02263575,0.026408374,0.041498873,0.0452715,0.08299775,0.124496624,0.23767537,0.3961256,0.4640329,0.49421388,0.5055317,0.59607476,0.7582976,0.88279426,0.7884786,0.6752999,0.6187105,0.6149379,0.6187105,1.2487389,1.8636768,2.6898816,3.92353,5.726845,7.3453007,7.914967,7.405663,6.296511,5.613666,5.8626595,7.5112963,9.235386,10.56335,11.876224,12.310076,11.77059,9.533423,6.749226,6.4210076,7.911195,7.484888,7.696155,9.0957985,10.26154,10.816116,11.197151,11.846043,13.075918,15.082954,14.916959,14.758509,14.683057,13.422999,8.397863,6.63982,5.4476705,4.006528,2.3163917,1.1883769,0.67152727,0.39989826,0.2678564,0.25276586,0.43007925,0.44139713,0.482896,0.60362,0.7507524,0.7469798,0.7394345,0.6413463,0.73188925,1.0110635,1.177059,1.0525624,0.87902164,0.6752999,0.5281675,0.6149379,0.8224323,0.8262049,0.754525,0.7092535,0.76584285,0.9016574,1.0827434,1.2751472,1.3958713,1.3091009,1.146878,1.086516,1.1016065,1.1581959,1.2298758,1.1959221,1.2902378,1.4373702,1.5316857,1.4260522,1.5015048,2.0787163,2.5578396,2.7879698,3.0558262,3.6971724,4.172523,5.2967653,6.9152217,7.9262853,7.54525,7.115171,7.3113475,7.911195,7.786698,6.5530496,6.673774,7.375482,8.213005,9.035437,9.763554,9.710737,9.57115,9.57115,9.480607,10.86516,11.5857315,10.895341,9.0957985,7.533932,6.436098,5.59103,4.8063245,4.2894745,4.678055,5.5985756,7.5603404,9.325929,10.529396,11.680047,13.558814,14.445381,14.022847,12.577931,11.004747,11.593277,12.604341,14.313339,17.206944,21.96045,22.141537,22.250942,22.662159,22.7942,21.1267,22.04722,22.711203,22.356575,20.877707,18.848034,16.414692,14.981093,14.226569,13.819125,13.407909,13.841762,14.1926155,14.317112,14.086982,13.407909,12.291212,11.18206,10.069136,9.001483,8.062099,7.273621,6.907676,6.881268,6.9152217,6.519096,6.058836,5.8664317,6.228604,7.0585814,7.9036493,8.431817,8.692128,8.601585,8.028146,6.7869525,6.590776,6.2436943,5.587258,4.617693,3.4632697,2.4522061,1.7127718,1.1619685,0.784706,0.5998474,0.5583485,0.58475685,0.6073926,0.6111652,0.62248313,0.59607476,0.51684964,0.45648763,0.43385187,0.41498876,0.3470815,0.3470815,0.3961256,0.47912338,0.5696664,0.58098423,0.55080324,0.51684964,0.5017591,0.513077,0.44894236,0.4376245,0.49044126,0.58098423,0.62248313,0.6187105,0.65643674,0.7582976,0.935611,1.2034674,1.6260014,1.9202662,2.444661,3.3953626,4.8100967,6.043745,6.0701537,6.0512905,6.156924,5.594803,4.851596,4.5724216,4.357382,3.9725742,3.3576362,3.229367,3.240685,3.3764994,3.5764484,3.7160356,3.6066296,3.410453,3.2670932,3.3161373,3.6745367,4.142342,4.327201,4.323428,4.2102494,4.0404816,4.0517993,3.9612563,4.0216184,4.2706113,4.5497856,4.8365054,5.406172,6.2436943,7.152897,7.7376537,7.5905213,7.2962565,7.6018395,8.480861,9.107117,9.484379,10.084227,10.751981,11.151879,10.733118,9.831461,9.537196,10.291721,12.0724,14.369928,14.769827,14.547242,14.234114,14.151116,14.426518,15.124454,16.72782,19.074392,21.881226,24.752193,26.70264,27.604298,27.69484,27.366621,27.1629,27.136492,26.642279,26.166927,25.623669,24.337204,23.544952,22.813063,21.911406,20.775846,19.519562,18.75372,18.172735,17.723793,17.316349,16.848543,17.067356,16.912678,16.06761,14.48688,12.408164,10.416218,9.050528,8.062099,7.2887115,6.6360474,6.368191,6.1003346,5.726845,5.2326307,4.696918,4.304565,4.1536603,4.002755,3.742444,3.4029078,2.2598023,2.2107582,1.9579924,1.7693611,1.841041,2.305074,1.5580941,1.6184561,2.1390784,2.8219235,3.4217708,3.9197574,4.7648253,6.1078796,7.5490227,8.126234,5.4778514,4.727099,4.5724216,4.5724216,5.1647234,5.704209,4.817642,3.9650288,3.9725742,5.0515447,6.1041074,6.6662283,7.665974,8.507269,7.092535,6.458734,7.1868505,8.443134,9.137298,7.9300575,7.2660756,6.983129,7.281166,8.186596,9.525878,7.8961043,7.175533,6.673774,6.013564,5.1232247,5.4476705,5.6476197,5.938112,6.1003346,5.4891696,4.1574326,3.4783602,4.274384,5.8626595,6.0814714,6.677546,8.899622,10.823661,11.744182,12.193124,11.529142,11.283921,12.536433,14.468017,14.373701,12.721292,10.759526,8.846806,7.2660756,6.205968,8.477088,10.367173,11.498961,11.548005,10.220041,7.277394,5.7909794,4.659192,3.4142256,2.203213,2.1466236,2.033445,2.1805773,2.595566,2.987919,3.199186,2.9766011,2.6521554,2.5389767,2.9464202,2.8898308,2.2183034,1.5467763,1.3053282,1.7618159,3.3840446,4.8553686,5.6023483,4.772371,1.2223305,0.8262049,0.91297525,1.2713746,1.8297231,2.637065,3.338773,2.8521044,1.931584,1.1317875,0.79602385,1.4713237,1.177059,0.86770374,0.8941121,1.0299267,1.1129243,1.0110635,1.0148361,1.2600567,1.7316349,2.3314822,2.806833,2.8898308,2.5917933,2.1994405,2.0749438,2.1315331,2.4559789,3.0105548,3.6707642,3.7047176,3.4594972,2.71629,1.8070874,1.6071383,0.8941121,0.63002837,0.55080324,0.4979865,0.452715,0.48666862,0.35839936,0.22258487,0.150905,0.116951376,0.041498873,0.033953626,0.041498873,0.041498873,0.041498873,0.060362,0.120724,0.19994913,0.31312788,0.51684964,0.91297525,1.2261031,1.0525624,0.573439,0.56589377,1.539231,2.474842,3.0143273,2.7992878,1.478869,0.80734175,0.48666862,0.422534,0.5357128,0.7696155,2.252257,2.8332415,2.6182017,1.9391292,1.358145,2.5427492,2.7125173,2.3767538,1.8448136,1.2525115,0.72811663,0.513077,0.5998474,0.9507015,1.4600059,1.5656394,1.1657411,0.77338815,0.62625575,0.69039035,1.1355602,1.750498,2.3993895,2.7502437,2.282438,2.0108092,1.690136,1.5580941,2.0183544,3.6292653,1.8863125,1.026154,0.66020936,0.47912338,0.2678564,0.16976812,0.29803738,0.663982,1.0676528,1.0978339,0.23767537,0.011317875,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.02263575,0.018863125,0.011317875,0.018863125,0.041498873,0.08299775,0.0754525,0.05281675,0.033953626,0.0150905,0.011317875,0.011317875,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.033953626,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.0,0.003772625,0.07922512,0.15467763,0.18485862,0.1358145,0.05281675,0.011317875,0.003772625,0.0150905,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.03772625,0.071679875,0.08299775,0.06790725,0.08677038,0.10186087,0.1056335,0.120724,0.090543,0.07922512,0.0754525,0.08677038,0.09808825,0.10186087,0.07922512,0.056589376,0.0452715,0.033953626,0.030181,0.03772625,0.071679875,0.12826926,0.18485862,0.12826926,0.124496624,0.18485862,0.25276586,0.1961765,0.120724,0.06790725,0.049044125,0.056589376,0.071679875,0.05281675,0.033953626,0.02263575,0.033953626,0.05281675,0.10940613,0.14335975,0.29049212,0.52439487,0.6526641,0.5998474,0.573439,0.69793564,0.8903395,0.88279426,0.8563859,0.7884786,0.80356914,0.8865669,0.87147635,1.3694628,1.6524098,2.0070364,2.6823363,3.9084394,6.598321,8.09228,8.635539,8.431817,7.6131573,6.255012,7.8206515,9.623966,10.140816,8.99771,9.910686,11.438599,11.1782875,9.601331,10.035183,12.838243,11.012292,9.6051035,9.955957,9.676784,7.9338303,8.054554,9.042982,10.469034,12.449662,13.249459,14.64533,16.795727,16.991903,9.673011,7.4811153,5.9532022,4.3686996,2.6936543,1.599593,0.97710985,0.58475685,0.3772625,0.31312788,0.32067314,0.29426476,0.38103512,0.44516975,0.46026024,0.48666862,0.59607476,0.5281675,0.784706,1.3241913,1.5618668,1.4298248,1.3430545,1.1242423,0.77338815,0.452715,0.452715,0.49421388,0.5394854,0.63002837,0.84884065,1.0714256,1.3128735,1.6146835,1.8787673,1.8485862,1.5430037,1.20724,0.9808825,0.9280658,1.026154,0.8639311,0.875249,0.965792,1.0902886,1.2185578,1.6448646,2.9539654,4.2517486,5.089271,5.455216,5.3269467,4.5535583,4.715781,6.047518,7.4282985,8.054554,8.488406,8.835487,8.907167,8.231868,8.114917,8.243186,7.673519,6.360646,5.1232247,5.3910813,6.089017,6.6020937,6.571913,5.8928404,7.092535,8.907167,10.103089,10.054046,8.7600355,7.624475,6.488915,5.379763,4.5950575,4.6856003,5.221313,7.696155,10.1294985,11.872451,13.63804,15.633758,16.957949,17.135263,16.03743,13.86817,12.879742,12.657157,14.071891,18.052011,25.593489,25.186045,24.774828,24.771055,23.767538,18.549997,19.534653,20.496672,20.492899,19.338476,17.591751,16.233604,15.109364,14.268067,13.807808,13.845533,14.64533,15.203679,15.335721,14.909414,13.875714,12.400619,11.0613365,9.718282,8.511042,7.8696957,7.3490734,6.820906,6.379509,5.938112,5.198677,4.8930945,4.9345937,5.2854476,5.9192486,6.79827,7.1793056,7.360391,7.322665,7.0510364,6.541732,6.0739264,5.613666,5.089271,4.425289,3.5689032,2.5502944,1.8485862,1.3958713,1.1091517,0.9016574,0.724344,0.6187105,0.58475685,0.6073926,0.63002837,0.55080324,0.422534,0.3772625,0.41876137,0.422534,0.35839936,0.29426476,0.32067314,0.44516975,0.59230214,0.56589377,0.5357128,0.513077,0.5017591,0.47912338,0.43385187,0.41121614,0.41121614,0.43385187,0.47535074,0.51684964,0.6187105,0.76584285,0.9507015,1.1732863,1.4222796,1.8033148,2.384299,3.169005,4.085753,4.991183,5.564622,5.9796104,6.119198,5.5268955,4.9760923,4.772371,4.745962,4.587512,3.8593953,3.0369632,2.535204,2.3503454,2.493705,2.9803739,3.308592,3.4066803,3.3463185,3.259548,3.3425457,4.3800178,4.957229,5.0477724,4.7346444,4.217795,3.9650288,3.8971217,4.0970707,4.4101987,4.4705606,4.2781568,4.4705606,5.3269467,6.628502,7.673519,7.4282985,6.3153744,5.5985756,5.6778007,6.058836,6.530414,7.0849895,7.7716074,8.280911,7.9338303,7.6093845,7.854605,8.914713,10.853842,13.562587,13.060828,12.457208,11.993175,11.857361,12.178034,12.789199,13.143826,13.9888935,15.629986,17.927513,20.108091,21.907633,22.941332,23.371412,23.918442,24.827644,25.212452,25.661396,25.933023,24.971004,23.809036,22.620659,21.466236,20.496672,19.945868,19.557287,19.123436,18.599041,18.131235,18.09351,17.961468,18.014284,17.644567,16.52787,14.6151495,12.434572,11.031156,9.940866,8.963757,8.167733,7.665974,7.039718,6.3229194,5.5759397,4.8855495,4.398881,4.191386,4.112161,4.0216184,3.8103511,2.1353056,3.1614597,3.610402,3.572676,3.1840954,2.6106565,2.2899833,2.6446102,2.9237845,2.8709676,2.7011995,2.957738,3.863168,4.870459,5.587258,5.783434,5.281675,4.7912335,4.6214657,4.9119577,5.6287565,5.485397,4.851596,4.1762958,4.134797,5.66271,7.699928,8.439363,8.273367,7.5792036,6.7152724,6.0286546,7.5905213,8.986393,8.956212,7.3717093,6.1003346,5.1873593,5.4703064,6.7341356,7.7225633,7.3792543,7.073672,6.670001,6.089017,5.292993,4.025391,2.7728794,2.7125173,3.5123138,3.3425457,2.8785129,2.8709676,3.7613072,4.825187,4.164978,4.557331,6.7039547,9.676784,11.706455,10.193633,7.9828744,6.862405,6.5568223,6.7831798,7.232122,7.9526935,8.333729,7.937603,6.802043,5.4476705,5.142088,5.515578,6.907676,8.729855,9.476834,7.937603,5.0062733,2.7313805,1.7882242,1.4939595,1.6524098,2.003264,2.516341,2.9992368,3.097325,3.3651814,3.5236318,3.2670932,2.6521554,2.0900342,2.052308,1.8787673,1.6109109,1.4939595,1.9693103,3.3463185,3.9310753,3.6368105,2.5389767,0.8563859,0.694163,0.77338815,0.935611,1.1355602,1.4637785,2.2447119,2.1315331,1.7014539,1.3468271,1.237421,1.3468271,1.1091517,0.98465514,1.0299267,0.87147635,0.79602385,0.90543,0.9016574,0.8299775,1.0978339,1.6486372,2.123988,2.293756,2.1881225,2.0900342,2.5314314,2.7313805,2.8219235,3.1576872,4.3196554,2.5238862,3.6783094,5.4363527,5.9305663,3.7688525,1.50905,1.0827434,1.2110126,1.1959221,0.91674787,0.5017591,0.22258487,0.071679875,0.018863125,0.030181,0.041498873,0.10940613,0.14713238,0.1358145,0.1358145,0.19994913,0.26031113,0.23390275,0.17354076,0.26031113,0.49044126,0.694163,0.7507524,0.6526641,0.52062225,0.9808825,0.9695646,0.543258,0.026408374,0.0150905,0.55080324,0.73188925,0.84884065,1.146878,1.8297231,3.2821836,3.9763467,3.8556228,3.1765501,2.516341,3.0671442,4.191386,4.0895257,2.595566,1.1883769,0.6790725,0.48666862,0.49044126,0.6073926,0.77716076,0.80356914,0.7092535,0.72811663,0.7997965,0.58098423,1.2525115,2.4974778,4.055572,5.27413,5.1269975,2.795515,1.4901869,1.0978339,1.0299267,0.19994913,0.41876137,0.91297525,1.2298758,1.1091517,0.48666862,0.5357128,0.5017591,0.4074435,0.2678564,0.120724,0.02263575,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.06413463,0.0754525,0.06413463,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.018863125,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.02263575,0.056589376,0.0754525,0.071679875,0.060362,0.03772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.05281675,0.1056335,0.15467763,0.1659955,0.14335975,0.1358145,0.14335975,0.1659955,0.23013012,0.14335975,0.08677038,0.056589376,0.049044125,0.060362,0.08677038,0.08299775,0.071679875,0.056589376,0.0452715,0.033953626,0.030181,0.049044125,0.071679875,0.060362,0.03772625,0.030181,0.08677038,0.16976812,0.18485862,0.10940613,0.06413463,0.056589376,0.094315626,0.1659955,0.13204187,0.0754525,0.033953626,0.026408374,0.0754525,0.124496624,0.15467763,0.181086,0.21503963,0.27540162,0.3470815,0.6790725,0.8978847,0.8563859,0.62625575,0.784706,0.77716076,0.83752275,1.1280149,1.7391801,2.4220252,2.354118,3.218049,4.798779,5.0213637,4.508287,4.7006907,5.670255,6.3531003,4.5460134,3.9725742,5.3571277,8.929804,12.940104,13.671993,13.951167,13.547497,12.370438,11.106608,11.231105,11.536687,12.593022,14.203933,16.03743,17.621931,11.936585,12.189351,13.158916,12.079946,8.650629,6.307829,6.0626082,5.938112,5.3382645,5.0213637,5.20245,5.2590394,4.2328854,2.3918443,1.2223305,0.7582976,0.4678055,0.32067314,0.24899325,0.1358145,0.10186087,0.08299775,0.071679875,0.08299775,0.1659955,0.14335975,0.090543,0.071679875,0.120724,0.24522063,0.40367088,1.0186088,1.5505489,1.5015048,0.42630664,0.34330887,0.32821837,0.3961256,0.56589377,0.8865669,1.4600059,1.7580433,2.082489,2.4220252,2.4710693,1.9730829,1.2336484,0.8111144,0.8299775,0.97710985,0.9507015,0.754525,0.5885295,0.5357128,0.5357128,1.3015556,2.8219235,5.062863,7.273621,7.9941926,8.763808,8.07719,6.1305156,4.425289,5.7683434,6.7454534,8.024373,9.122208,9.748463,9.797507,11.016065,12.97783,12.875969,10.020092,5.8437963,4.8327327,5.9418845,7.194396,7.798016,8.16396,9.273112,10.797253,11.717773,11.725319,11.200924,9.918231,8.122461,6.1041074,5.1043615,7.322665,8.179051,8.503497,9.235386,10.427535,11.246195,14.626467,17.769064,19.108345,17.565342,12.574159,12.951422,13.185325,14.049255,16.143063,19.866644,20.85507,20.43631,18.659403,16.414692,15.411173,17.95015,19.078165,18.45568,16.77309,15.746937,15.418718,14.283158,13.238141,12.759018,12.894833,13.856852,15.060319,15.535669,14.988639,13.777626,12.106354,10.38981,9.046755,8.296002,8.16396,7.6622014,6.960493,6.1606965,5.4174895,4.927048,4.8666863,4.779916,4.640329,4.515832,4.5761943,5.2967653,5.8437963,6.0512905,5.8211603,5.111907,4.002755,3.1840954,2.6710186,2.384299,2.1503963,1.8938577,1.4750963,1.1393328,0.9507015,0.7922512,0.6828451,0.5998474,0.5394854,0.52062225,0.59607476,0.5357128,0.49044126,0.5357128,0.60362,0.52062225,0.44516975,0.4074435,0.44516975,0.543258,0.6413463,0.56589377,0.52062225,0.48666862,0.44139713,0.38103512,0.34330887,0.35462674,0.35839936,0.35462674,0.36594462,0.47535074,0.66775465,0.83752275,0.97710985,1.1581959,1.478869,2.0145817,2.5389767,3.059599,3.8292143,4.647874,5.1081343,5.5193505,5.7570257,5.292993,4.6856003,4.3121104,4.2517486,4.496969,4.957229,3.7273536,2.8785129,2.493705,2.4182527,2.2748928,2.7389257,3.0445085,3.2029586,3.2821836,3.4029078,3.7575345,4.678055,5.349582,5.3910813,4.851596,4.1197066,3.9273026,4.085753,4.3121104,4.22534,4.2894745,5.3646727,6.511551,7.145352,7.0510364,6.270103,5.534441,5.111907,4.8968673,4.4101987,4.38379,4.644101,5.1534057,5.6891184,5.8588867,5.836251,5.828706,6.273875,7.5301595,9.88805,11.242422,11.461235,11.291467,11.234878,11.566868,10.868933,10.751981,10.970794,11.642321,13.230596,16.060064,19.353567,21.153109,21.454918,22.186808,23.846762,24.205162,24.491882,25.155863,25.865116,25.129456,23.114874,21.281378,20.33822,20.26277,20.311813,20.085455,19.334703,18.251959,17.471025,17.399347,17.91997,18.19537,17.689838,16.188334,14.369928,13.026875,11.940358,10.978339,10.084227,8.631766,7.3188925,6.224831,5.3986263,4.8365054,4.5422406,4.52715,4.587512,4.564876,4.3347464,4.1989317,4.1310244,4.1310244,3.9574835,3.5160866,2.8521044,2.7917426,3.0633714,3.4745877,3.8367596,4.0178456,4.557331,6.047518,7.6131573,8.480861,7.9941926,8.575176,8.620448,8.27714,7.779153,7.424526,7.5226145,7.567886,7.201941,6.7454534,7.1868505,8.677037,9.016574,8.299775,7.1076255,6.507778,6.673774,7.111398,7.01331,6.145606,4.8440504,4.4139714,5.198677,6.56814,7.7678347,7.914967,7.3000293,6.8850408,6.911449,7.2283497,7.284939,7.911195,8.224322,8.424272,8.182823,6.6247296,5.251494,4.074435,3.6594462,4.0178456,4.617693,6.609639,7.7376537,8.75249,9.552286,9.178797,6.677546,5.9532022,5.8173876,5.772116,5.9984736,6.7680893,8.416726,9.103344,8.29223,6.752999,5.413717,4.817642,4.6026025,4.4705606,4.191386,3.4029078,2.4484336,1.7580433,1.5015048,1.569412,2.3314822,3.31991,4.2328854,4.708236,4.3196554,4.478106,4.429062,3.9801195,3.1312788,2.052308,1.901403,1.6675003,1.418507,1.2487389,1.2864652,2.0862615,2.4974778,2.493705,2.1541688,1.6712729,1.358145,1.1129243,1.1732863,1.5316857,1.9391292,2.233394,2.0485353,1.6675003,1.3732355,1.418507,1.3807807,1.1732863,1.1695137,1.3619176,1.358145,1.6184561,1.8334957,1.9391292,1.9278114,1.8448136,2.4220252,2.9049213,3.2029586,3.4368613,3.9461658,4.406426,4.6856003,4.9534564,5.4665337,6.5756855,7.0170827,6.4247804,5.8173876,5.3759904,4.4177437,1.4260522,0.9997456,1.3468271,1.6033657,1.8297231,1.9542197,1.3053282,0.6451189,0.3169005,0.24899325,0.26408374,0.24899325,0.21881226,0.18863125,0.19994913,0.21881226,0.20749438,0.14335975,0.071679875,0.08677038,0.17354076,0.24522063,0.27540162,0.28294688,0.33576363,0.331991,0.27540162,0.181086,0.094315626,0.11317875,0.43385187,0.5394854,0.7809334,1.3166461,2.0862615,2.2220762,3.059599,3.5236318,3.2633207,2.6634734,2.1881225,1.8938577,1.8523588,1.7693611,0.9695646,0.7809334,0.47912338,0.3470815,0.5093044,0.9242931,1.0676528,0.9507015,0.9393836,1.0487897,0.94692886,1.901403,2.867195,3.380272,3.399135,3.3312278,2.0258996,1.6071383,1.7919968,1.9353566,1.0299267,0.663982,0.5998474,0.6111652,0.5319401,0.27917424,0.27917424,0.2867195,0.2565385,0.18863125,0.120724,0.150905,0.08677038,0.026408374,0.018863125,0.041498873,0.0452715,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0,0.003772625,0.018863125,0.05281675,0.0754525,0.07922512,0.060362,0.033953626,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.011317875,0.011317875,0.003772625,0.0,0.0,0.003772625,0.0,0.003772625,0.018863125,0.0452715,0.08677038,0.120724,0.12826926,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.08299775,0.20372175,0.35085413,0.47535074,0.4979865,0.41498876,0.31312788,0.1961765,0.10940613,0.13204187,0.1056335,0.090543,0.094315626,0.10186087,0.08677038,0.071679875,0.049044125,0.041498873,0.0452715,0.033953626,0.09808825,0.08677038,0.056589376,0.03772625,0.03772625,0.011317875,0.0150905,0.02263575,0.03772625,0.049044125,0.0452715,0.03772625,0.03772625,0.049044125,0.08299775,0.08299775,0.0452715,0.0150905,0.00754525,0.026408374,0.03772625,0.041498873,0.049044125,0.06413463,0.1056335,0.1659955,0.28294688,0.36594462,0.41876137,0.5281675,0.6752999,0.72811663,0.80356914,1.1129243,1.9466745,3.059599,4.036709,5.406172,7.141579,8.669493,8.333729,6.79827,5.342037,4.485651,3.9989824,3.0822346,4.0103,5.583485,6.688864,6.2851934,5.560849,6.296511,6.9152217,7.009537,7.3377557,8.707218,9.948412,9.87296,8.880759,8.944894,9.710737,10.978339,12.00072,11.631002,8.296002,5.828706,4.647874,4.0480266,3.5387223,2.8596497,2.757789,2.384299,1.7655885,1.0676528,0.6111652,0.4678055,0.3470815,0.27917424,0.26031113,0.24899325,0.16222288,0.10940613,0.09808825,0.11317875,0.13204187,0.08677038,0.14713238,0.19240387,0.17731337,0.1358145,0.17731337,0.331991,0.5017591,0.56212115,0.36594462,0.38858038,0.42630664,0.51684964,0.65643674,0.7884786,1.0186088,1.4147344,1.991946,2.5880208,2.8521044,2.173032,1.6335466,1.418507,1.5279131,1.780679,1.8259505,1.4826416,1.0789708,0.814887,0.76584285,1.6712729,3.4594972,5.704209,7.5527954,7.7150183,7.956466,7.9526935,7.6018395,7.2698483,7.7829256,8.428044,9.088254,9.178797,8.631766,7.8810134,7.8319697,8.326183,8.495952,8.345046,8.748717,8.918486,8.726082,7.4697976,5.904158,6.270103,7.020855,8.820397,11.2650585,13.58145,14.618922,12.340257,9.522105,6.903904,5.66271,7.3981175,8.416726,10.114408,11.068882,10.714255,9.367428,12.355347,15.482853,16.516552,14.954685,12.012038,12.283667,14.275613,16.769318,18.934805,20.357084,20.866388,18.851807,17.554024,17.448391,16.24115,16.124199,15.878979,15.516807,15.109364,14.807553,13.766309,12.487389,11.7894535,12.091263,13.419228,15.954432,18.202915,18.923487,17.625704,14.57365,12.136535,10.250222,8.907167,8.103599,7.8206515,7.4773426,7.2170315,6.8473144,6.4964604,6.6134114,6.1229706,5.5985756,5.2326307,5.1156793,5.2250857,5.515578,5.6551647,5.621211,5.3646727,4.7836885,3.8367596,2.848332,2.071171,1.5769572,1.237421,0.9808825,0.76207024,0.663982,0.66020936,0.66020936,0.6752999,0.6488915,0.5998474,0.5470306,0.47157812,0.41121614,0.49421388,0.56589377,0.58475685,0.6149379,0.6111652,0.5394854,0.513077,0.5357128,0.5055317,0.5885295,0.62625575,0.5696664,0.45648763,0.4074435,0.39989826,0.36971724,0.362172,0.40367088,0.52439487,0.73188925,0.88279426,0.9620194,0.98465514,0.9997456,1.5807298,2.0372176,2.493705,3.1199608,4.123479,4.5497856,4.8855495,5.0213637,4.961002,4.817642,4.776143,4.8440504,4.8968673,4.847823,4.666737,4.2064767,4.0480266,3.8782585,3.482133,2.7502437,3.006782,3.199186,3.1539145,2.969056,3.0105548,3.3350005,3.9084394,4.557331,5.2779026,6.19465,7.1604424,7.84706,7.8961043,7.2057137,5.9607477,5.485397,6.096562,6.5228686,6.156924,5.0854983,4.115934,3.4444065,3.2972744,3.6669915,4.3121104,4.659192,5.1798143,5.926794,6.7039547,7.0812173,6.6850915,5.8664317,5.4363527,5.7607985,6.79827,7.61693,7.907422,7.8621507,7.756517,7.9300575,8.60913,9.25425,9.74469,10.269085,11.299012,12.96274,15.554533,18.063328,19.794964,20.37972,21.160654,21.967995,22.526344,22.737612,22.665932,21.737865,21.013521,20.55326,20.447628,20.813572,20.655123,19.99114,19.123436,18.23687,17.384256,17.538933,18.51227,18.915941,18.048239,15.882751,14.943368,14.268067,13.528633,12.585477,11.491416,9.5183325,7.805561,6.485142,5.594803,5.0439997,4.870459,4.9459114,5.036454,4.961002,4.6026025,5.1647234,5.1081343,4.9459114,4.7233267,4.45547,4.1310244,4.3083377,4.878004,5.583485,6.1003346,6.0248823,5.7683434,6.7341356,7.9828744,8.782671,8.590267,8.382772,8.246958,8.096053,8.050782,8.431817,8.801534,8.246958,7.17176,6.296511,6.643593,7.7942433,8.3525915,8.084735,7.356619,7.141579,7.2924843,7.394345,7.164215,6.643593,6.205968,6.828451,7.7942433,8.280911,7.835742,6.3531003,6.330465,7.1378064,8.544995,10.054046,10.884023,10.616167,10.774617,10.480352,9.273112,7.1000805,5.4778514,4.7421894,4.98741,5.7607985,6.0776987,6.2361493,7.5490227,8.348819,8.262049,8.213005,7.122716,6.802043,6.809588,6.8850408,6.9454026,8.028146,10.035183,11.3820095,11.208468,9.386291,7.6848373,6.3908267,5.172269,3.942393,2.886058,2.6182017,2.4559789,2.2748928,2.052308,1.8448136,2.5691576,3.3953626,4.055572,4.3007927,3.9273026,4.0895257,4.247976,3.9574835,3.1425967,2.071171,1.961765,1.9844007,1.7618159,1.3091009,1.0601076,1.4750963,1.7391801,1.8184053,1.7354075,1.5279131,1.2110126,0.965792,1.056335,1.4600059,1.8599042,2.0070364,1.8787673,1.7127718,1.6071383,1.5467763,1.4901869,1.358145,1.2826926,1.3204187,1.4524606,2.2484846,2.9124665,3.3878171,3.6066296,3.4557245,3.802806,3.7650797,3.5462675,3.4029078,3.6594462,3.9197574,4.3309736,4.878004,5.553304,6.3342376,6.48137,4.930821,4.564876,5.7607985,6.436098,4.432834,3.1463692,2.4672968,2.1994405,2.033445,1.8561316,1.3241913,0.7884786,0.43385187,0.3055826,0.26031113,0.211267,0.1659955,0.13204187,0.120724,0.11317875,0.090543,0.056589376,0.026408374,0.026408374,0.060362,0.08677038,0.11317875,0.1659955,0.26408374,0.5281675,0.5319401,0.42630664,0.3169005,0.23767537,0.36594462,0.68661773,1.3355093,2.214531,2.9954643,2.5201135,3.3161373,3.8103511,3.500996,2.957738,2.625747,2.173032,2.1013522,2.2598023,1.8297231,1.6486372,1.6146835,1.3241913,0.875249,0.8526133,0.91297525,0.8903395,0.8224323,0.7884786,0.88279426,1.5430037,2.1881225,2.595566,2.8521044,3.361409,2.2371666,1.7127718,1.7127718,1.8900851,1.6222287,2.4107075,2.5616124,2.1315331,1.2562841,0.18485862,0.392353,0.39989826,0.33953625,0.28294688,0.24899325,0.23767537,0.15467763,0.0754525,0.033953626,0.026408374,0.033953626,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.026408374,0.02263575,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.00754525,0.011317875,0.02263575,0.033953626,0.033953626,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.056589376,0.094315626,0.10940613,0.08677038,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.090543,0.10940613,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.049044125,0.14335975,0.2678564,0.362172,0.35085413,0.2678564,0.241448,0.2263575,0.20749438,0.18863125,0.15467763,0.1358145,0.124496624,0.116951376,0.090543,0.0754525,0.056589376,0.03772625,0.018863125,0.011317875,0.090543,0.11317875,0.10186087,0.071679875,0.02263575,0.003772625,0.003772625,0.00754525,0.0150905,0.033953626,0.030181,0.041498873,0.05281675,0.056589376,0.041498873,0.056589376,0.041498873,0.030181,0.030181,0.041498873,0.041498873,0.06413463,0.094315626,0.116951376,0.124496624,0.1056335,0.10940613,0.124496624,0.15845025,0.23767537,0.35462674,0.44894236,0.482896,0.6828451,1.5505489,2.214531,2.8181508,3.6481283,4.768598,6.039973,6.6850915,6.2625575,5.4476705,4.938366,5.455216,5.9682927,6.7869525,7.828197,8.922258,9.805053,9.5032425,8.612903,7.9828744,8.156415,9.393836,10.729345,10.374719,9.280658,8.4544525,8.963757,7.7904706,9.125979,10.902886,11.41219,9.288202,6.9265394,5.8890676,5.221313,4.395108,3.3161373,2.3616633,1.6184561,1.086516,0.73566186,0.513077,0.422534,0.362172,0.32067314,0.29426476,0.28294688,0.19240387,0.124496624,0.094315626,0.10186087,0.120724,0.08677038,0.1358145,0.18863125,0.20749438,0.181086,0.17731337,0.20749438,0.26031113,0.31312788,0.32444575,0.4376245,0.5093044,0.5696664,0.633801,0.69039035,0.754525,0.9922004,1.4373702,1.9579924,2.2296214,1.8825399,1.6825907,1.6976813,1.8372684,1.8561316,1.7919968,1.6071383,1.4449154,1.4298248,1.6863633,3.0558262,4.5309224,5.2892203,5.4740787,6.1720147,7.7829256,8.831716,9.34102,9.789962,11.140562,12.400619,12.053536,10.684074,9.027891,7.9489207,10.103089,10.212496,9.009028,7.6207023,7.5792036,10.133271,10.748209,9.525878,7.432071,6.319147,6.270103,8.431817,11.151879,13.396591,14.766054,13.894578,11.491416,8.571404,6.8473144,8.714764,10.955703,11.861133,11.725319,11.321648,11.887542,14.188843,16.33924,16.207197,14.162435,13.087236,14.154889,15.184815,16.686321,17.976559,17.210714,16.346785,15.46399,15.015047,14.7736,13.841762,14.019074,14.136025,14.566105,15.147089,15.196134,14.656648,14.456699,15.101818,16.675003,18.840488,20.956932,21.934042,20.839981,17.746428,13.728582,10.676529,8.7751255,7.779153,7.466025,7.61693,7.4509344,7.3792543,7.111398,6.7341356,6.730363,6.0626082,5.458988,5.1269975,5.0515447,4.9760923,4.8930945,4.957229,5.0062733,4.881777,4.432834,3.8820312,2.9011486,1.871222,1.0751982,0.694163,0.52062225,0.4640329,0.4678055,0.4979865,0.543258,0.63002837,0.65643674,0.66775465,0.65643674,0.56212115,0.5583485,0.62625575,0.6375736,0.59607476,0.6413463,0.56589377,0.44139713,0.38858038,0.41498876,0.42630664,0.513077,0.56589377,0.55080324,0.482896,0.45648763,0.4640329,0.42630664,0.38858038,0.3961256,0.5017591,0.62248313,0.68661773,0.724344,0.754525,0.7884786,1.0450171,1.7316349,2.5238862,3.3312278,4.304565,5.330719,5.715527,5.6287565,5.2628117,4.82896,4.772371,4.9459114,4.90064,4.5422406,4.134797,4.014073,4.063117,4.3649273,4.610148,4.112161,3.4632697,3.2972744,3.1652324,2.9501927,2.8521044,2.9766011,3.3312278,3.9801195,5.0062733,6.4926877,7.6093845,8.394091,8.695901,8.356364,7.2283497,6.579458,6.6058664,6.7114997,6.417235,5.3609,4.1800685,3.4972234,3.2784111,3.4896781,4.0970707,4.90064,5.753253,6.6850915,7.4207535,7.3868,6.590776,6.0248823,5.7004366,5.643847,5.926794,6.5228686,6.356873,5.8513412,5.379763,5.2892203,6.217286,7.33021,8.43559,9.397609,10.148361,11.517824,13.675766,15.950659,17.836971,18.983849,19.621422,20.52308,21.119154,21.11161,20.492899,20.277859,20.228815,20.413673,20.790936,21.205925,20.632486,19.534653,18.23687,17.180534,16.94286,17.591751,18.534906,18.402864,16.965494,15.1395445,14.867915,15.128226,14.641558,13.177779,11.54046,9.827688,8.348819,7.1340337,6.198423,5.553304,5.3344917,5.300538,5.27413,5.1043615,4.67051,5.6287565,5.956975,6.058836,6.006019,5.8626595,5.7004366,5.938112,6.530414,7.0812173,7.375482,7.3717093,7.149124,7.752744,8.571404,9.21275,9.49947,8.831716,8.337502,8.175279,8.405409,9.001483,8.907167,8.001738,6.9567204,6.387054,6.8699503,7.2924843,7.54525,7.496206,7.3151197,7.4999785,7.5565677,8.103599,8.420499,8.246958,7.7829256,8.160188,8.6732645,8.541223,7.443389,5.541986,5.2326307,6.647365,9.103344,11.532914,12.50248,10.899114,9.869187,8.899622,7.6320205,5.847569,4.7006907,4.8025517,6.0362,7.394345,6.960493,6.1003346,7.443389,8.541223,8.560086,8.29223,7.6923823,7.277394,7.2057137,7.2396674,6.7756343,7.8131065,9.703192,11.374464,11.796998,9.978593,9.669238,8.582722,6.990674,5.240176,3.772625,3.410453,3.5538127,3.5575855,3.138824,2.372981,2.5276587,2.7879698,2.9992368,3.0671442,2.9501927,3.2331395,3.85185,4.22534,4.0706625,3.4142256,3.1199608,3.31991,2.795515,1.5920477,1.0223814,1.2411937,1.5543215,1.7467253,1.7467253,1.6071383,1.2826926,1.0336993,1.1506506,1.5807298,1.9240388,1.9542197,1.841041,1.7882242,1.7957695,1.6825907,1.5731846,1.5769572,1.5882751,1.569412,1.5430037,2.8709676,3.8254418,4.485651,4.8742313,4.9647746,5.032682,4.346064,3.5424948,3.0445085,3.0746894,3.3463185,3.6707642,4.104616,4.647874,5.2250857,5.281675,4.3121104,4.1762958,5.160951,5.9720654,5.2590394,4.093298,3.0935526,2.444661,1.8938577,1.539231,1.3053282,0.91297525,0.42630664,0.2565385,0.18485862,0.13958712,0.094315626,0.05281675,0.03772625,0.03772625,0.030181,0.02263575,0.018863125,0.041498873,0.049044125,0.056589376,0.07922512,0.13958712,0.26408374,1.0186088,1.0035182,0.95824677,1.1883769,1.569412,0.9695646,0.98465514,1.8863125,3.31991,4.3007927,3.1312788,3.6179473,4.2819295,4.398881,4.014073,3.591539,3.561358,3.9273026,4.1536603,3.1840954,2.11267,1.8221779,1.4449154,0.8563859,0.6375736,0.6413463,0.66775465,0.59607476,0.7507524,1.8938577,2.3918443,2.7238352,3.0181,3.2935016,3.4444065,2.3013012,1.599593,1.3355093,1.3430545,1.2525115,2.203213,2.4031622,1.9806281,1.1280149,0.120724,0.45648763,0.4376245,0.33576363,0.29426476,0.29803738,0.18863125,0.120724,0.0754525,0.041498873,0.02263575,0.011317875,0.00754525,0.00754525,0.00754525,0.00754525,0.0,0.0,0.003772625,0.011317875,0.011317875,0.011317875,0.003772625,0.0,0.00754525,0.030181,0.041498873,0.056589376,0.060362,0.06790725,0.116951376,0.10186087,0.06413463,0.033953626,0.0150905,0.00754525,0.0,0.0,0.00754525,0.0150905,0.00754525,0.02263575,0.026408374,0.02263575,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.13204187,0.2263575,0.241448,0.1358145,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.05281675,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.049044125,0.10186087,0.13958712,0.120724,0.0754525,0.11317875,0.18485862,0.25276586,0.2678564,0.26408374,0.2263575,0.181086,0.14713238,0.116951376,0.094315626,0.08677038,0.06790725,0.0452715,0.049044125,0.09808825,0.11317875,0.1056335,0.07922512,0.02263575,0.00754525,0.003772625,0.003772625,0.0150905,0.041498873,0.041498873,0.060362,0.071679875,0.06790725,0.06790725,0.060362,0.056589376,0.06413463,0.071679875,0.08677038,0.0754525,0.1358145,0.2565385,0.41876137,0.6073926,0.4376245,0.2867195,0.17354076,0.1056335,0.090543,0.1358145,0.19994913,0.23013012,0.35085413,0.87902164,1.0110635,1.2298758,1.6071383,2.1541688,2.8407867,3.7575345,4.2706113,4.4139714,4.4743333,4.983638,5.9494295,6.79827,7.99042,9.567377,11.159425,11.283921,9.918231,9.329701,10.201178,11.634775,12.106354,10.902886,9.574923,9.224068,10.495442,8.805306,9.488152,10.208723,9.967276,9.06939,6.8435416,6.398372,6.379509,6.0022464,5.0439997,3.470815,2.444661,1.7354075,1.2147852,0.8601585,0.84884065,0.8186596,0.7130261,0.5357128,0.3734899,0.241448,0.16222288,0.124496624,0.10940613,0.12826926,0.11317875,0.12826926,0.18485862,0.24899325,0.27917424,0.27917424,0.31312788,0.35839936,0.38480774,0.33576363,0.39989826,0.47157812,0.5470306,0.6111652,0.633801,0.7394345,1.1393328,1.7165444,2.1466236,1.901403,1.6222287,1.5580941,1.6825907,1.8297231,1.690136,1.6033657,1.5203679,1.6335466,2.0636258,2.8747404,4.6856003,5.5382137,5.1760416,4.3875628,4.991183,7.039718,8.880759,10.148361,11.046246,12.344029,12.966512,12.370438,11.544232,10.891568,10.220041,12.325166,12.147853,10.110635,7.77538,7.854605,11.329193,12.498707,12.00072,10.521852,8.76758,8.035691,9.424017,11.234878,12.687338,13.8719425,15.773345,14.709465,11.661184,8.929804,10.148361,13.041965,13.336229,12.51757,12.091263,13.592768,16.301512,17.425755,16.244923,13.79649,12.887287,14.509516,15.245177,16.448645,17.603067,16.316603,13.721037,12.755245,12.1252165,11.3669195,10.819888,11.661184,12.774108,14.234114,15.520579,15.501716,15.403628,16.13929,17.644567,19.595015,21.398329,22.186808,21.651094,19.383747,15.690348,11.589504,8.790216,7.333983,6.8925858,7.062354,7.3792543,7.4396167,7.194396,6.700182,6.1908774,6.0776987,5.455216,4.957229,4.67051,4.5233774,4.2894745,4.195159,4.1762958,4.221567,4.236658,4.025391,3.6556737,2.6710186,1.6146835,0.84129536,0.5017591,0.38480774,0.40367088,0.47157812,0.543258,0.6149379,0.6790725,0.66020936,0.6488915,0.6488915,0.59230214,0.56589377,0.5696664,0.5696664,0.56589377,0.5998474,0.482896,0.36971724,0.32067314,0.34330887,0.35839936,0.392353,0.4376245,0.47157812,0.482896,0.45648763,0.44894236,0.422534,0.38858038,0.3772625,0.42630664,0.422534,0.43385187,0.4678055,0.5357128,0.633801,0.70170826,1.3166461,2.1881225,3.1614597,4.214022,5.2062225,5.696664,5.6778007,5.2779026,4.7535076,4.610148,4.678055,4.610148,4.3083377,3.9461658,3.863168,3.942393,4.4403796,5.0175915,4.7308717,3.9084394,3.5990841,3.3123648,2.9086938,2.6182017,2.595566,2.8143783,3.3425457,4.2517486,5.5985756,6.5040054,7.164215,7.699928,8.0206,7.8244243,7.2358947,6.9869013,6.9982195,6.971811,6.398372,5.198677,4.436607,4.002755,3.8895764,4.168751,4.817642,5.621211,6.4436436,6.94163,6.56814,5.6589375,5.20245,4.9647746,4.90064,5.1647234,5.7117543,5.481624,4.9723196,4.6026025,4.715781,5.3458095,6.2323766,7.3981175,8.567632,9.178797,10.272858,12.0082655,14.019074,16.03743,17.863379,19.093256,20.26277,20.904116,20.715485,19.564833,19.662922,19.40261,19.1423,19.029121,18.97253,18.58395,17.969013,16.980585,15.939341,15.626213,16.35433,17.380484,17.493662,16.542961,15.452672,15.222542,15.339493,14.675511,13.075918,11.3669195,10.084227,9.050528,8.00551,6.9567204,6.1644692,5.772116,5.5193505,5.3080835,5.0251365,4.5460134,5.9720654,6.7379084,7.4811153,7.91874,7.9715567,7.7602897,8.07719,8.416726,8.492179,8.503497,9.107117,9.635284,10.272858,10.789707,11.114153,11.336739,11.348056,10.61994,9.914458,9.484379,9.107117,8.495952,7.914967,7.575431,7.567886,7.8998766,7.6018395,6.862405,6.2851934,6.149379,6.4021444,6.470052,7.594294,8.480861,8.458225,7.4999785,6.809588,6.7756343,6.752999,6.368191,5.50426,4.3422914,5.191132,7.6131573,10.186088,10.49167,8.571404,6.72659,5.6551647,5.191132,4.293247,3.8254418,4.538468,6.5040054,8.624221,8.6581745,8.084735,8.439363,9.0957985,9.367428,8.503497,7.5905213,6.94163,6.609639,6.2399216,5.0854983,5.828706,7.4697976,9.148616,9.918231,8.741172,10.3634,10.170997,8.741172,6.7869525,5.1571784,4.357382,4.534695,4.568649,3.9876647,2.938875,2.5087957,2.2598023,2.2107582,2.2711203,2.252257,2.5238862,3.4444065,4.5799665,5.451443,5.5495315,5.142088,5.251494,4.2328854,2.2258487,1.177059,1.1732863,1.5656394,1.9353566,2.1315331,2.2899833,1.8636768,1.5467763,1.6335466,2.0145817,2.1654868,2.003264,1.9164935,1.9844007,2.1654868,2.323937,2.003264,1.9542197,2.0372176,2.0636258,1.8033148,3.218049,4.063117,4.6290107,5.1232247,5.6778007,5.8626595,4.930821,3.7877154,3.0143273,2.9011486,3.399135,3.7084904,3.7462165,3.7914882,4.466788,5.594803,6.3908267,5.6287565,3.863168,3.4481792,3.31991,2.9615107,2.463524,1.9240388,1.4373702,1.2751472,1.2562841,0.9016574,0.31312788,0.1659955,0.124496624,0.10186087,0.060362,0.011317875,0.003772625,0.030181,0.041498873,0.03772625,0.033953626,0.0754525,0.0754525,0.124496624,0.1659955,0.22258487,0.39989826,1.8976303,1.6637276,1.750498,2.8294687,4.195159,2.5087957,1.8146327,2.425798,3.904667,5.062863,3.8858037,3.863168,4.4139714,4.938366,4.825187,4.274384,4.768598,5.66271,5.945657,4.266839,2.2711203,1.3128735,0.7809334,0.44516975,0.43007925,0.56589377,0.6451189,0.56589377,0.97710985,3.2821836,3.7650797,3.9159849,4.0782075,4.085753,3.2482302,2.1994405,1.50905,1.086516,0.76207024,0.26408374,0.19994913,0.13204187,0.07922512,0.056589376,0.0754525,0.35839936,0.30181,0.18863125,0.16222288,0.19994913,0.049044125,0.026408374,0.03772625,0.03772625,0.02263575,0.003772625,0.011317875,0.018863125,0.0150905,0.0150905,0.011317875,0.02263575,0.049044125,0.0754525,0.060362,0.0452715,0.030181,0.060362,0.124496624,0.1659955,0.150905,0.1659955,0.1961765,0.23767537,0.27540162,0.21503963,0.13204187,0.06413463,0.030181,0.011317875,0.003772625,0.0,0.0150905,0.030181,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.02263575,0.0452715,0.17731337,0.29049212,0.29426476,0.1358145,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.030181,0.090543,0.16976812,0.2565385,0.31312788,0.27917424,0.23390275,0.21503963,0.21503963,0.1961765,0.19240387,0.18485862,0.17354076,0.18485862,0.20749438,0.17731337,0.1358145,0.094315626,0.06413463,0.03772625,0.0150905,0.003772625,0.00754525,0.02263575,0.0452715,0.06790725,0.071679875,0.06790725,0.1056335,0.07922512,0.071679875,0.08299775,0.10186087,0.1056335,0.07922512,0.15845025,0.34330887,0.6451189,1.0676528,0.8526133,0.6488915,0.49421388,0.38480774,0.26408374,0.17354076,0.17731337,0.29426476,0.41498876,0.3055826,0.1961765,0.44139713,0.7922512,1.1431054,1.5430037,1.8825399,2.3277097,2.8030603,3.1539145,3.138824,3.078462,3.9876647,5.3571277,6.6549106,7.2924843,6.79827,6.587003,7.8017883,10.001229,11.1782875,10.997202,9.9257765,8.903395,8.763808,10.231359,10.993429,10.616167,8.892077,6.7831798,6.432326,4.7421894,4.8629136,5.7004366,6.3417826,6.085244,4.6856003,3.6141748,2.6785638,1.8561316,1.3015556,1.4034165,1.4034165,1.2298758,0.9016574,0.5357128,0.32821837,0.24522063,0.20749438,0.18485862,0.15845025,0.14335975,0.15467763,0.21503963,0.3055826,0.35462674,0.3772625,0.43007925,0.5055317,0.55080324,0.47157812,0.38858038,0.44139713,0.55080324,0.6375736,0.6073926,0.8262049,1.5618668,2.4710693,2.9728284,2.2862108,1.8523588,1.7957695,1.9202662,2.0070364,1.8259505,1.720317,1.5505489,1.6788181,2.282438,3.3463185,5.372218,6.217286,6.198423,5.723072,5.304311,6.1305156,7.8696957,9.608876,10.823661,11.348056,10.367173,10.057818,10.880251,12.264804,12.600568,12.253486,11.962994,11.012292,10.578441,13.762536,14.505743,14.351066,13.751218,12.826925,11.393328,11.212241,11.0613365,11.16697,11.619685,12.404391,16.535416,17.255987,14.916959,11.6875925,11.570641,13.992666,14.332202,13.385274,12.287439,12.525115,16.007248,16.927769,15.645076,13.223051,11.419736,12.67602,14.003984,15.75071,17.414436,17.629477,14.981093,13.000465,11.193378,9.839006,9.993684,10.616167,11.7894535,13.166461,14.222796,14.302021,14.403882,15.418718,16.833452,18.09351,18.62545,18.221779,17.135263,15.294222,12.691111,9.386291,7.5716586,6.7341356,6.617184,6.8246784,6.8359966,6.9265394,6.466279,5.915476,5.587258,5.6476197,5.0138187,4.610148,4.2819295,3.942393,3.5953116,3.591539,3.4255435,3.3463185,3.3840446,3.3538637,2.9200118,2.0183544,1.1996948,0.69793564,0.47157812,0.3961256,0.43007925,0.5394854,0.6790725,0.77338815,0.7809334,0.68661773,0.5885295,0.5357128,0.5357128,0.43385187,0.41121614,0.47535074,0.55080324,0.5055317,0.4640329,0.41876137,0.3961256,0.392353,0.40367088,0.3169005,0.30935526,0.362172,0.43007925,0.41876137,0.35085413,0.32821837,0.32444575,0.32821837,0.34330887,0.29426476,0.30181,0.35462674,0.44894236,0.5998474,0.80356914,1.0676528,1.6109109,2.5238862,3.7688525,4.2291126,4.6856003,4.8025517,4.5837393,4.3686996,4.2781568,4.1989317,4.2706113,4.3913355,4.221567,3.9914372,3.9461658,4.1800685,4.4403796,4.112161,3.9310753,3.8065786,3.470815,2.9237845,2.463524,2.3616633,2.444661,2.7087448,3.187868,3.9688015,4.696918,5.2137675,5.7419353,6.3531003,6.9491754,6.5643673,6.507778,6.6247296,6.7341356,6.6360474,5.7117543,5.028909,4.508287,4.183841,4.1762958,4.221567,4.715781,5.1798143,5.27413,4.7874613,4.0970707,3.500996,3.2105038,3.3538637,3.9725742,4.45547,4.5309224,4.504514,4.666737,5.2967653,5.643847,5.987156,6.7077274,7.665974,8.20546,8.744945,9.857869,11.634775,13.849306,15.98084,18.097282,19.83269,20.847527,20.919205,19.934551,19.153618,17.931286,16.62973,15.535669,14.841507,15.120681,15.426264,15.245177,14.5283785,13.660675,14.147344,15.241405,16.13929,16.459963,16.229834,15.99593,15.158407,14.003984,12.73261,11.457462,10.480352,9.748463,8.797762,7.624475,6.6813188,6.039973,5.515578,5.1269975,4.776143,4.2706113,6.3644185,7.6923823,9.216523,10.559577,11.3971,11.457462,12.411936,12.879742,13.072145,13.43809,14.649103,14.562332,14.796235,14.86037,14.437836,13.411682,14.634012,13.856852,12.00072,9.910686,8.360137,9.314611,9.031664,8.194141,7.364164,6.971811,7.3377557,5.7570257,4.112161,3.180323,2.595566,2.3993895,2.9086938,3.7160356,4.4705606,4.8968673,4.776143,4.2592936,3.8141239,3.6594462,3.7688525,3.5387223,3.4896781,4.617693,6.0739264,5.1571784,4.496969,4.3422914,4.67051,4.9647746,4.195159,3.5123138,4.606375,7.492433,11.551778,15.516807,13.283413,11.268831,9.476834,7.7942433,6.013564,6.8774953,7.0774446,6.5756855,5.5495315,4.3649273,5.402399,6.960493,8.280911,9.058073,9.461743,10.057818,10.3634,9.4127,7.352846,5.462761,4.7912335,4.4403796,3.9650288,3.3538637,3.0369632,2.938875,2.795515,2.9615107,3.169005,2.5314314,2.1805773,2.5578396,3.5877664,4.9647746,6.149379,6.6850915,6.462507,5.323174,3.5349495,1.7995421,1.1431054,1.1129243,1.5656394,2.3163917,3.1576872,2.535204,2.2711203,2.2899833,2.323937,1.9240388,1.6410918,1.8636768,2.505023,3.4217708,4.4101987,3.591539,2.8181508,2.2748928,2.0598533,2.1805773,2.5616124,2.9313297,3.410453,4.1272516,5.1873593,6.5568223,6.4474163,5.2326307,3.6330378,2.7313805,3.218049,4.4403796,4.538468,3.8443048,4.881777,7.3981175,9.718282,8.341274,4.376245,3.5689032,2.727608,1.4373702,0.5696664,0.35085413,0.35085413,0.26408374,0.16976812,0.10940613,0.090543,0.090543,0.090543,0.10186087,0.08677038,0.05281675,0.0150905,0.003772625,0.026408374,0.05281675,0.06413463,0.0754525,0.11317875,0.36971724,0.5357128,0.59607476,0.83752275,3.9386206,3.2029586,3.1010978,4.991183,7.1264887,4.8930945,4.142342,3.5538127,3.0256453,3.6481283,5.4778514,4.957229,3.5764484,2.5427492,2.7615614,3.874486,4.67051,4.8553686,4.5120597,4.1197066,3.4745877,2.5804756,1.4449154,0.4678055,0.44139713,1.0148361,1.388326,1.1129243,0.80734175,2.1353056,2.052308,2.3578906,3.3048196,4.285702,3.8443048,3.0030096,2.142851,1.3355093,0.63002837,0.0452715,0.20372175,0.16976812,0.07922512,0.026408374,0.0754525,0.271629,0.21881226,0.1056335,0.030181,0.030181,0.00754525,0.026408374,0.041498873,0.02263575,0.0,0.0,0.018863125,0.02263575,0.0150905,0.0150905,0.05281675,0.116951376,0.19994913,0.2565385,0.18485862,0.09808825,0.1056335,0.3055826,0.56589377,0.52062225,0.3470815,0.24899325,0.36594462,0.52062225,0.21503963,0.06790725,0.011317875,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.033953626,0.02263575,0.060362,0.071679875,0.0754525,0.08299775,0.10186087,0.1358145,0.06413463,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.041498873,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.003772625,0.0,0.00754525,0.02263575,0.060362,0.09808825,0.1358145,0.19994913,0.31312788,0.45648763,0.52062225,0.5055317,0.4640329,0.43007925,0.44139713,0.49044126,0.48666862,0.41876137,0.30935526,0.19994913,0.11317875,0.056589376,0.02263575,0.011317875,0.0,0.0,0.026408374,0.0452715,0.0452715,0.0452715,0.056589376,0.060362,0.06790725,0.071679875,0.0452715,0.00754525,0.018863125,0.041498873,0.1056335,0.27540162,0.47157812,0.7092535,1.0412445,1.2261031,0.76207024,0.47157812,0.52439487,0.8111144,0.9393836,0.24522063,0.1358145,0.271629,0.58475685,0.9808825,1.3732355,1.4939595,2.2748928,3.338773,4.3347464,4.957229,4.164978,5.138315,6.187105,6.300284,5.142088,2.335255,1.9730829,3.31991,5.613666,8.043237,9.224068,7.213259,6.40969,7.752744,8.744945,8.20546,6.771862,4.5460134,2.3088465,1.5279131,1.7089992,2.0673985,2.6031113,3.2520027,3.874486,3.7650797,3.1237335,2.2748928,1.5354583,1.20724,1.1695137,1.177059,1.1657411,1.0336993,0.65643674,0.46026024,0.35839936,0.32821837,0.3169005,0.24522063,0.16976812,0.18863125,0.24899325,0.3169005,0.36594462,0.392353,0.47912338,0.6073926,0.7394345,0.8224323,0.7130261,0.7884786,0.7997965,0.6790725,0.5357128,0.6451189,1.0186088,1.690136,2.4672968,2.9464202,2.9803739,3.31991,3.4896781,3.3010468,2.837014,2.3126192,1.9353566,1.6788181,1.5430037,1.5430037,3.5085413,6.5341864,8.6581745,8.990166,7.7225633,7.073672,7.2057137,8.096053,9.627739,11.581959,10.774617,9.695646,9.024119,9.258021,10.695392,10.902886,11.815862,14.43029,19.621422,28.166418,20.794708,16.561823,13.822898,11.54046,9.291975,12.540206,12.098808,10.370946,9.046755,9.0957985,12.121444,14.618922,15.275358,14.392565,13.853079,15.222542,14.815099,12.879742,10.582213,10.008774,11.7555,14.11339,14.369928,12.593022,11.627231,11.359374,11.23865,11.34051,12.272349,15.150862,17.67852,18.28214,15.735619,12.434572,14.388792,13.973803,12.276122,10.012547,8.601585,10.163452,11.114153,12.132762,13.041965,13.570132,13.35132,12.898605,12.540206,11.955449,10.899114,9.216523,8.152642,7.2094865,6.4738245,5.956975,5.613666,5.040227,5.0439997,5.587258,6.330465,6.6360474,5.3684454,4.847823,4.4705606,3.9386206,3.2670932,2.6672459,2.535204,2.505023,2.3654358,2.0598533,1.6939086,1.3468271,0.8526133,0.3470815,0.27540162,0.33576363,0.3961256,0.48666862,0.59230214,0.6413463,0.7130261,0.73188925,0.66020936,0.5583485,0.59607476,0.58475685,0.633801,0.7205714,0.7130261,0.3961256,0.52062225,0.5319401,0.5055317,0.55080324,0.7922512,0.41498876,0.23767537,0.21881226,0.30935526,0.44139713,0.26031113,0.17731337,0.150905,0.16222288,0.19994913,0.28294688,0.3055826,0.3470815,0.4678055,0.68661773,1.0148361,1.327964,1.478869,1.780679,2.9766011,4.293247,4.285702,3.9197574,3.7198083,3.7688525,3.8178966,3.7650797,4.0480266,4.5497856,4.6252384,4.1612053,3.5839937,3.2520027,3.150142,2.9313297,2.8936033,3.048281,3.3350005,3.4745877,2.9766011,2.7087448,2.5314314,2.4522061,2.4899325,2.686109,2.8181508,3.0558262,3.2859564,3.3840446,3.187868,3.1161883,3.6028569,4.1574326,4.4743333,4.425289,4.0593443,4.085753,3.9348478,3.4670424,2.9916916,3.0256453,3.6594462,3.8367596,3.2972744,2.5804756,2.1994405,2.2258487,2.505023,2.9237845,3.3878171,3.5462675,3.3312278,3.2746384,3.5877664,4.1498876,4.7610526,5.3910813,6.126743,6.900131,7.462252,7.413208,7.5490227,8.29223,9.691874,11.41219,13.807808,16.143063,18.244415,20.02132,21.4851,18.372684,15.954432,14.332202,13.377728,12.740154,13.12119,12.921241,12.487389,12.1101265,12.0233555,12.792972,13.087236,13.385274,13.947394,14.800008,16.071383,15.354584,14.000212,12.725064,11.627231,10.846297,10.0465,9.0807085,7.9753294,6.911449,5.9984736,5.198677,4.719554,4.432834,3.904667,7.3377557,9.031664,10.212496,11.027383,11.532914,11.691365,11.529142,11.981857,12.725064,13.705947,15.147089,16.146835,16.346785,15.648849,14.139798,12.068627,10.917976,10.589758,10.408672,9.993684,9.265567,8.654402,7.454707,6.1531515,5.243949,5.2137675,5.3382645,4.768598,3.7386713,2.637065,2.033445,1.7391801,1.7127718,1.8863125,2.2069857,2.6031113,2.6068838,2.5578396,2.5729303,2.7125173,2.938875,2.746471,2.686109,2.987919,3.4859054,3.6066296,3.5538127,3.682082,3.8971217,4.0178456,3.7575345,3.4632697,4.425289,7.4471617,12.027128,16.38451,14.120935,10.827434,8.937348,8.967529,9.491924,9.733373,8.624221,6.9265394,5.2326307,3.9612563,4.5007415,6.719045,8.443134,8.9788475,9.107117,9.216523,9.239159,9.129752,8.677037,7.488661,6.417235,5.458988,4.568649,3.874486,3.6971724,3.802806,3.6971724,3.229367,2.8785129,3.7273536,3.7462165,3.5349495,3.3425457,3.4481792,4.183841,4.6327834,5.20245,5.462761,5.0553174,3.6934,3.2784111,2.8294687,2.4974778,2.4069347,2.6332922,2.8709676,2.746471,2.6710186,2.7615614,2.837014,2.1466236,2.1881225,2.5993385,3.1539145,3.7499893,3.832987,3.4896781,3.1199608,2.938875,2.9615107,3.048281,2.7728794,2.897376,3.5651307,4.285702,4.5007415,3.5274043,2.6295197,2.6634734,4.074435,5.198677,5.4778514,4.930821,4.085753,3.9914372,4.006528,3.7499893,2.7238352,1.358145,0.9695646,0.68661773,0.362172,0.1659955,0.13204187,0.13204187,0.14335975,0.1961765,0.2678564,0.29426476,0.17731337,0.98842776,1.1204696,0.8337501,0.4074435,0.124496624,0.6413463,0.724344,0.56212115,0.362172,0.34330887,1.2298758,1.2751472,1.5618668,2.3314822,2.987919,2.2220762,1.4713237,1.780679,3.0860074,4.2102494,3.2255943,3.4745877,3.3878171,2.6898816,2.41448,3.0445085,3.6556737,4.2291126,4.644101,4.678055,4.617693,4.568649,5.062863,5.6589375,4.938366,4.191386,3.6707642,2.9728284,2.41448,2.9954643,2.6672459,2.41448,2.7841973,3.399135,2.9539654,3.0633714,3.0331905,3.0256453,3.6745367,6.066381,4.8063245,4.696918,4.9119577,4.112161,0.46026024,0.3169005,0.24522063,0.19240387,0.12826926,0.05281675,0.19994913,0.18485862,0.12826926,0.0754525,0.00754525,0.0,0.150905,0.22258487,0.17731337,0.18485862,0.0452715,0.00754525,0.05281675,0.12826926,0.1358145,0.094315626,0.241448,0.44516975,0.633801,0.80734175,0.8865669,0.7884786,0.58475685,0.46026024,0.7130261,0.67152727,0.29049212,0.071679875,0.1056335,0.041498873,0.0150905,0.003772625,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.026408374,0.02263575,0.018863125,0.0150905,0.02263575,0.08677038,0.30935526,0.2263575,0.08299775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.049044125,0.094315626,0.06413463,0.041498873,0.03772625,0.041498873,0.060362,0.09808825,0.22258487,0.32444575,0.3772625,0.4074435,0.5055317,0.56589377,0.6149379,0.68661773,0.7582976,0.7092535,0.70170826,0.7394345,0.7884786,0.7582976,0.49044126,0.26031113,0.11317875,0.03772625,0.011317875,0.0,0.0,0.011317875,0.02263575,0.030181,0.056589376,0.090543,0.08299775,0.06413463,0.0452715,0.02263575,0.003772625,0.003772625,0.0150905,0.033953626,0.06790725,0.116951376,0.15845025,0.241448,0.32821837,0.32444575,0.31312788,0.32067314,0.35839936,0.3734899,0.24522063,0.23013012,0.25276586,0.2867195,0.35839936,0.55457586,0.9620194,1.5580941,1.9391292,2.2220762,3.029418,4.112161,5.59103,7.062354,8.126234,8.401636,8.337502,8.126234,7.937603,7.997965,8.601585,7.707473,6.9265394,7.5112963,9.390063,11.159425,9.869187,8.748717,7.0284004,4.768598,2.8445592,2.354118,1.9353566,1.6788181,1.6109109,1.6788181,1.7542707,1.6712729,1.4335974,1.1317875,0.9507015,1.1355602,1.1431054,0.97710985,0.6790725,0.35085413,0.271629,0.38103512,0.5055317,0.543258,0.4376245,0.30935526,0.24522063,0.23390275,0.24522063,0.2565385,0.26031113,0.29426476,0.35839936,0.44139713,0.52062225,0.6526641,0.814887,0.91297525,0.90543,0.8262049,0.84884065,1.2600567,2.0485353,2.8294687,2.8332415,3.006782,3.240685,3.4066803,3.3915899,3.0822346,2.8030603,2.8936033,3.0520537,2.9652832,2.3088465,3.9159849,6.1342883,8.126234,9.537196,10.502988,10.7557535,11.272603,11.676274,11.680047,11.106608,8.82417,9.046755,10.472807,12.0233555,12.808062,11.3669195,12.027128,15.064092,19.353567,22.382984,20.066593,19.376202,16.610868,12.581704,12.600568,15.116908,15.339493,13.283413,10.789707,11.510279,13.358865,14.600059,15.147089,15.652621,17.516298,18.874443,18.45568,16.388283,14.056801,14.086982,16.252468,17.293713,16.071383,13.404137,12.079946,11.653639,11.815862,12.672247,14.479335,17.655886,18.832945,18.293459,16.244923,13.86817,13.340002,13.645585,13.777626,12.909923,11.219787,9.880505,9.759781,10.842525,12.291212,13.422999,13.743673,13.106099,12.253486,11.374464,10.631257,10.167224,10.121953,9.337247,8.382772,7.4773426,6.470052,5.4967146,5.089271,5.2175403,5.6589375,6.0022464,5.7796617,5.2628117,4.508287,3.6556737,2.9351022,2.2975287,1.8146327,1.50905,1.3053282,1.0110635,0.7507524,0.6149379,0.5093044,0.44139713,0.49421388,0.4678055,0.47157812,0.5470306,0.6413463,0.59230214,0.5394854,0.5319401,0.543258,0.5470306,0.5470306,0.56212115,0.5696664,0.59230214,0.6073926,0.55457586,0.56212115,0.55080324,0.5055317,0.43385187,0.35462674,0.27917424,0.22258487,0.19240387,0.20749438,0.28294688,0.2867195,0.2565385,0.19994913,0.14713238,0.17354076,0.26031113,0.30181,0.35085413,0.4376245,0.5885295,0.8224323,0.90920264,0.94692886,1.1581959,1.9240388,3.2444575,4.1574326,4.6252384,4.5120597,3.572676,3.2029586,3.229367,3.5839937,4.0970707,4.5007415,3.8820312,3.259548,2.848332,2.7502437,2.9803739,3.1652324,3.1576872,3.0105548,2.8558772,2.9011486,3.0331905,3.361409,3.5802212,3.5047686,3.0633714,3.3538637,4.044254,4.659192,4.9534564,4.9232755,4.3422914,3.7273536,3.4066803,3.380272,3.3010468,2.8106055,2.6295197,2.3880715,2.1013522,2.161714,2.674791,3.3463185,3.3538637,2.5804756,1.6146835,1.569412,2.4597516,3.1614597,3.218049,2.8634224,2.8634224,2.806833,3.0935526,3.893349,5.1269975,6.0701537,6.2814207,6.156924,6.0512905,6.2889657,6.387054,6.647365,7.2962565,8.420499,9.937095,11.781908,14.102073,16.58446,18.8254,20.300495,19.500698,18.214233,16.735365,15.222542,13.6682205,13.189097,12.951422,12.857106,12.804289,12.672247,13.370183,12.657157,11.6875925,11.193378,11.491416,12.54775,13.211733,13.35132,13.000465,12.370438,11.45369,11.117926,10.310584,8.7600355,6.9869013,5.6098933,4.6629643,4.06689,3.6934,3.3463185,8.179051,9.374973,10.559577,10.982111,10.593531,10.072908,9.325929,8.869441,9.21275,10.54826,12.728837,14.758509,16.007248,16.146835,14.837734,11.706455,10.035183,9.34102,9.186342,9.14107,8.786444,7.6622014,6.1720147,4.8855495,4.2404304,4.52715,4.429062,3.7763977,2.8407867,2.0145817,1.8372684,1.5128226,1.2713746,1.1506506,1.177059,1.3619176,1.4260522,1.5052774,1.6976813,1.9881734,2.2371666,2.1994405,2.1881225,2.1881225,2.2409391,2.4522061,2.8106055,3.0331905,2.987919,2.7389257,2.5389767,2.7841973,3.9122121,7.0057645,11.159425,13.505998,12.136535,10.484125,10.144588,11.129244,11.853588,11.593277,10.544487,9.367428,8.420499,7.7678347,7.3717093,7.756517,8.22055,8.75249,10.005001,10.110635,9.87296,9.276885,8.612903,8.461998,8.60913,8.5563135,8.280911,7.8696957,7.496206,6.7077274,5.5797124,4.3347464,3.5877664,4.3385186,4.5007415,4.1574326,3.904667,4.146115,5.0854983,4.7648253,4.979865,5.3571277,5.5759397,5.383536,5.481624,4.606375,3.6330378,3.0633714,3.0407357,3.5877664,3.5462675,3.3840446,3.2444575,2.957738,2.1503963,2.305074,2.8936033,3.6066296,4.3649273,4.5950575,4.036709,3.4255435,3.1425967,3.1954134,3.3161373,2.9803739,2.6483827,2.6219745,3.006782,2.8822856,2.161714,1.5731846,1.629774,2.625747,3.6858547,3.983892,3.308592,2.233394,2.1013522,1.7278622,1.1846043,0.6375736,0.241448,0.12826926,0.18863125,0.23767537,0.26408374,0.26408374,0.24899325,0.47912338,0.543258,0.48666862,0.36594462,0.271629,1.8863125,1.9127209,1.297783,0.7469798,0.7205714,1.3732355,2.3654358,2.6898816,2.1503963,1.3355093,2.546522,2.0749438,2.0183544,2.8256962,3.3048196,1.4977322,0.97333723,1.5920477,3.0709167,4.9723196,6.3342376,6.741681,6.3116016,5.3458095,4.3121104,3.7763977,4.0178456,4.798779,5.832478,6.7869525,6.9982195,6.5530496,6.4511886,6.828451,6.9454026,5.2175403,3.3274553,2.938875,3.5651307,2.5691576,1.8900851,1.9693103,2.9841464,4.0517993,3.240685,3.0709167,3.029418,3.0746894,3.2821836,3.8480775,4.063117,4.2894745,4.1800685,3.2670932,0.995973,0.49044126,0.91297525,0.9318384,0.3470815,0.08299775,0.29803738,0.17731337,0.05281675,0.06413463,0.14713238,0.16222288,0.21503963,0.22258487,0.181086,0.19240387,0.211267,0.08677038,0.13204187,0.35839936,0.47912338,0.52062225,0.62625575,0.76207024,0.90920264,1.0638802,1.1053791,0.6488915,0.331991,0.36971724,0.5885295,0.55457586,0.21881226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.00754525,0.0,0.0,0.0150905,0.090543,0.31312788,0.2867195,0.11317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.124496624,0.2263575,0.26408374,0.20372175,0.17354076,0.35085413,0.5055317,0.5319401,0.47157812,0.43007925,0.392353,0.3772625,0.39989826,0.4640329,0.5470306,0.63002837,0.7997965,0.95824677,0.814887,0.66775465,0.67152727,0.754525,0.80734175,0.694163,0.47535074,0.271629,0.120724,0.03772625,0.018863125,0.011317875,0.00754525,0.00754525,0.026408374,0.116951376,0.094315626,0.08299775,0.060362,0.033953626,0.0150905,0.003772625,0.003772625,0.011317875,0.0150905,0.00754525,0.018863125,0.011317875,0.0150905,0.041498873,0.094315626,0.120724,0.12826926,0.13204187,0.14713238,0.181086,0.26408374,0.29049212,0.29049212,0.33576363,0.48666862,0.965792,1.3807807,1.4901869,1.4675511,1.9240388,2.969056,4.9119577,7.1906233,9.016574,9.382519,9.374973,9.439108,9.484379,9.325929,8.688355,7.039718,6.149379,7.020855,9.544742,12.506252,12.012038,9.559832,6.820906,4.749735,3.5839937,3.1237335,2.5201135,1.7655885,1.0638802,0.845068,0.8639311,0.8639311,0.7997965,0.7130261,0.72811663,0.94315624,0.94315624,0.784706,0.51684964,0.19240387,0.15845025,0.2678564,0.3772625,0.41121614,0.35839936,0.3470815,0.362172,0.3961256,0.43385187,0.44894236,0.44139713,0.4074435,0.3961256,0.41121614,0.422534,0.46026024,0.543258,0.7507524,1.0638802,1.3845534,1.1657411,1.6788181,2.5729303,3.3312278,3.2935016,3.127506,3.1652324,3.2142766,3.2142766,3.2255943,3.4368613,4.0480266,4.478106,4.798779,5.723072,7.1302614,8.416726,8.518587,8.141325,9.752235,11.827179,13.985121,14.966003,14.203933,11.838497,9.7069645,10.416218,13.079691,15.32063,13.298503,11.434827,11.6008215,13.060828,15.524352,19.112118,18.648085,18.12369,16.124199,13.434318,13.023102,14.18507,14.377474,13.472044,12.261031,12.427027,13.502225,14.5132885,14.894323,14.871688,15.475307,17.659658,19.232841,19.221525,17.757746,16.094019,17.354074,18.255732,17.482344,15.264041,13.3626375,11.962994,12.057309,12.777881,13.65313,14.64533,13.928532,13.517315,13.324911,13.302276,13.407909,13.822898,13.660675,12.728837,11.1631975,9.435335,9.676784,10.902886,12.393073,13.419228,13.226823,11.649866,10.005001,9.110889,9.280658,10.325675,11.080199,10.925522,10.182315,9.058073,7.635793,6.247467,5.3571277,5.1571784,5.4891696,5.881522,5.8513412,5.2552667,4.3309736,3.3538637,2.6521554,2.1277604,1.6675003,1.2826926,0.9695646,0.72811663,0.5696664,0.4376245,0.36971724,0.38858038,0.5017591,0.52062225,0.5583485,0.6187105,0.67152727,0.6451189,0.5281675,0.51684964,0.5357128,0.56589377,0.62625575,0.67152727,0.7130261,0.7167987,0.69039035,0.694163,0.7167987,0.7092535,0.6375736,0.52439487,0.49044126,0.62248313,0.44139713,0.23390275,0.14335975,0.150905,0.19994913,0.241448,0.241448,0.20749438,0.18485862,0.241448,0.29049212,0.33576363,0.38103512,0.42630664,0.51684964,0.55080324,0.58098423,0.7092535,1.0789708,2.0673985,3.0860074,3.7763977,4.195159,4.798779,4.1310244,3.3915899,3.1840954,3.5689032,4.085753,3.712263,3.2935016,3.0860074,3.0633714,2.9351022,3.229367,3.3727267,3.218049,2.8936033,2.7841973,2.7879698,3.5689032,4.4215164,4.8365054,4.485651,4.8138695,5.2137675,5.6551647,6.017337,6.0776987,5.413717,4.459243,3.7914882,3.4330888,2.8294687,2.9615107,2.9992368,2.6785638,2.2183034,2.3201644,2.776652,3.3651814,3.2784111,2.3993895,1.3091009,1.146878,1.6146835,2.0975795,2.3428001,2.4484336,2.4899325,2.5691576,2.927557,3.7235808,5.0213637,6.013564,6.6662283,6.832224,6.5945487,6.307829,6.304056,6.749226,7.5112963,8.43559,9.374973,10.902886,12.97783,15.045229,16.724047,17.80679,17.799244,17.274849,16.365646,15.211224,13.966258,13.158916,12.759018,12.679792,12.740154,12.657157,12.604341,11.646093,10.521852,9.673011,9.246704,9.623966,10.567122,11.419736,11.8045435,11.604594,11.23865,11.02361,10.487898,9.435335,7.937603,6.205968,4.957229,4.0517993,3.429316,3.1048703,7.4169807,7.779153,8.3525915,8.552541,8.518587,9.103344,8.526133,8.028146,8.182823,9.099571,10.408672,12.377983,13.943622,14.588741,13.875714,11.438599,10.167224,9.639057,9.488152,9.288202,8.560086,6.5266414,5.160951,4.3611546,4.1197066,4.52715,4.38379,3.2218218,2.0447628,1.418507,1.4411428,1.2525115,1.0450171,0.8903395,0.814887,0.8111144,0.8224323,0.9016574,1.086516,1.327964,1.4939595,1.5580941,1.6146835,1.6033657,1.5618668,1.5882751,1.9806281,2.2258487,2.123988,1.7731338,1.5618668,2.704972,4.3875628,6.8737226,9.288202,9.612649,9.1825695,9.076936,9.673011,10.502988,10.265312,10.521852,10.419991,10.140816,9.952185,10.212496,9.031664,8.107371,7.9715567,9.084481,11.838497,11.570641,10.665211,9.4127,8.499724,9.012801,9.64283,10.091772,10.140816,9.733373,8.967529,7.8810134,7.01331,6.149379,5.413717,5.2665844,5.028909,4.851596,4.9459114,5.4174895,6.270103,5.9984736,5.7607985,5.6891184,5.8211603,6.092789,6.304056,5.455216,4.538468,3.983892,3.6669915,3.6745367,3.380272,3.1916409,3.1350515,2.867195,2.41448,2.595566,3.006782,3.5990841,4.67051,5.0779533,4.5422406,3.5990841,2.8332415,2.8822856,2.9766011,2.7313805,2.2107582,1.7278622,1.8448136,1.750498,1.5354583,1.3619176,1.3619176,1.6486372,1.9353566,2.04099,1.599593,0.86770374,0.7469798,0.5772116,0.38103512,0.20749438,0.090543,0.06790725,0.38858038,0.4979865,0.49421388,0.4678055,0.5017591,0.724344,1.2487389,1.9881734,2.837014,3.682082,3.3727267,2.8030603,2.5087957,2.6974268,3.218049,2.6936543,4.7006907,6.0324273,5.534441,4.1083884,4.432834,3.1010978,2.3314822,2.6446102,2.8521044,1.7165444,1.4109617,2.7351532,5.3571277,7.809334,9.0807085,8.054554,7.01331,6.858632,7.0774446,7.3868,7.854605,8.137552,8.345046,9.058073,8.726082,7.435844,6.2436943,6.0022464,7.360391,5.6476197,3.1840954,2.4823873,3.2067313,2.161714,1.5241405,1.8297231,3.0445085,4.1612053,3.180323,3.0369632,3.078462,3.1312788,2.927557,2.0975795,2.7087448,2.727608,2.3088465,1.7580433,1.5203679,1.2147852,1.4864142,1.2298758,0.422534,0.124496624,0.392353,0.18485862,0.0,0.030181,0.14713238,0.16222288,0.14335975,0.11317875,0.094315626,0.10186087,0.19240387,0.13958712,0.211267,0.41876137,0.5017591,0.4979865,0.51684964,0.56212115,0.6187105,0.6790725,0.67152727,0.2678564,0.06790725,0.1961765,0.28294688,0.25276586,0.09808825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.0,0.0150905,0.06413463,0.181086,0.181086,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.041498873,0.041498873,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.13204187,0.21881226,0.24522063,0.23013012,0.24522063,0.47157812,0.6375736,0.6451189,0.55080324,0.47912338,0.38480774,0.3470815,0.36971724,0.40367088,0.422534,0.47535074,0.633801,0.80734175,0.7582976,0.7167987,0.8299775,0.9242931,0.90920264,0.76584285,0.6187105,0.44139713,0.2678564,0.12826926,0.060362,0.030181,0.0150905,0.011317875,0.030181,0.09808825,0.060362,0.056589376,0.049044125,0.033953626,0.02263575,0.02263575,0.041498873,0.0452715,0.041498873,0.06790725,0.20749438,0.3169005,0.29426476,0.1659955,0.10186087,0.056589376,0.05281675,0.071679875,0.1056335,0.150905,0.23390275,0.27917424,0.3734899,0.6187105,1.1242423,1.7316349,2.0183544,1.9768555,1.7919968,1.8636768,2.4295704,3.6971724,5.281675,6.628502,7.0359454,7.699928,8.627994,9.0807085,8.578949,6.888813,5.300538,4.6856003,5.904158,8.809079,12.242168,12.0233555,8.661947,5.515578,4.025391,3.7386713,3.519859,2.9803739,2.1692593,1.3468271,0.965792,0.72811663,0.5281675,0.42630664,0.44516975,0.55080324,0.69793564,0.6790725,0.573439,0.40367088,0.14335975,0.09808825,0.14713238,0.20749438,0.241448,0.24522063,0.32067314,0.42630664,0.5319401,0.62625575,0.724344,0.76584285,0.724344,0.6828451,0.68661773,0.7582976,0.663982,0.5998474,0.8224323,1.388326,2.1654868,1.81086,2.123988,2.7992878,3.5085413,3.8782585,3.3425457,3.138824,3.0897799,3.150142,3.440634,3.5500402,3.9801195,4.3649273,5.0175915,6.9152217,9.465516,11.276376,10.978339,9.329701,9.205205,11.393328,14.196388,15.871433,15.467763,12.81938,10.653893,11.77059,14.634012,16.74291,14.622695,13.615403,12.759018,12.445889,13.392818,16.641048,16.923996,16.4826,15.411173,14.060574,13.023102,13.407909,13.875714,14.581196,15.116908,14.524607,13.52486,12.664702,12.08749,12.200669,13.645585,15.999702,16.576914,16.77309,16.795727,15.679029,16.87118,17.80679,17.757746,16.735365,15.467763,13.807808,12.936331,12.306303,11.627231,10.850069,10.4049,10.967021,12.061082,13.124963,13.50977,12.913695,11.729091,10.77839,10.544487,11.18206,11.578186,12.947649,14.622695,15.705438,15.082954,12.321393,9.797507,8.60913,9.046755,10.56335,11.646093,11.729091,11.083972,9.944639,8.507269,7.1679873,6.5756855,6.228604,5.9117036,5.66271,5.515578,4.9345937,4.134797,3.31991,2.6634734,2.1353056,1.6033657,1.146878,0.83752275,0.724344,0.69039035,0.543258,0.42630664,0.41498876,0.5093044,0.543258,0.5772116,0.63002837,0.6828451,0.68661773,0.5772116,0.5319401,0.5319401,0.5696664,0.6488915,0.69039035,0.7696155,0.80356914,0.784706,0.7809334,0.79602385,0.8299775,0.83752275,0.8111144,0.79602385,1.0450171,0.8941121,0.5696664,0.26408374,0.120724,0.1358145,0.17731337,0.19994913,0.181086,0.1358145,0.17731337,0.2263575,0.26408374,0.27540162,0.24899325,0.2678564,0.3055826,0.35839936,0.43385187,0.5772116,1.1317875,1.9768555,2.8332415,3.7801702,5.2665844,4.878004,3.8669407,3.229367,3.2633207,3.5689032,3.5462675,3.270866,3.048281,2.9351022,2.7389257,3.0709167,3.169005,3.0520537,2.8106055,2.6446102,2.5804756,3.1576872,3.9688015,4.5799665,4.534695,4.779916,5.0779533,5.455216,5.8626595,6.175787,5.80607,5.221313,4.45547,3.5877664,2.7615614,2.8332415,2.897376,2.8634224,2.7841973,2.8445592,3.2821836,3.5424948,3.2633207,2.4107075,1.2902378,0.91674787,0.9280658,1.2411937,1.7240896,2.214531,2.505023,2.6672459,2.938875,3.4745877,4.3196554,5.247721,6.349328,7.2170315,7.6207023,7.492433,7.3792543,7.6207023,8.141325,8.865668,9.710737,10.850069,12.253486,13.607859,14.694374,15.414946,15.573396,15.362129,14.7736,13.947394,13.185325,12.449662,12.038446,12.034674,12.204442,12.019584,11.34051,10.657665,9.899368,9.046755,8.111144,7.937603,8.469543,9.224068,9.835234,10.038955,10.140816,9.982366,9.631512,9.073163,8.216777,6.9454026,5.613666,4.3913355,3.4594972,2.9992368,5.27413,5.3080835,5.138315,5.4363527,6.7341356,9.416472,9.725827,10.133271,10.480352,10.54826,10.061591,11.068882,11.959221,12.057309,11.336739,10.401127,9.537196,9.601331,9.673011,9.201432,7.9753294,5.3269467,4.398881,4.1989317,4.236658,4.52715,4.504514,3.1539145,1.7354075,0.9318384,0.8563859,0.86770374,0.784706,0.70170826,0.6451189,0.55457586,0.482896,0.5470306,0.6375736,0.7130261,0.77716076,0.8601585,0.97333723,1.0601076,1.0789708,0.9695646,1.1431054,1.3996439,1.478869,1.3505998,1.2147852,3.0407357,5.1269975,6.530414,6.8397694,6.1908774,6.1833324,6.488915,6.9944468,7.2170315,6.307829,7.5603404,8.194141,8.179051,8.009283,8.699674,7.7716074,7.250985,7.7716074,9.676784,13.026875,12.238396,10.555805,9.099571,8.544995,9.122208,9.186342,9.012801,8.692128,8.156415,7.2057137,6.647365,7.326438,7.8508325,7.5905213,6.700182,5.772116,5.583485,5.9682927,6.620957,7.0887623,7.5188417,7.194396,6.722818,6.3644185,6.043745,5.824933,5.3759904,5.0666356,4.859141,4.2894745,3.4557245,2.6974268,2.3088465,2.3880715,2.867195,2.9992368,2.9954643,2.8332415,2.8785129,3.8782585,4.4894238,4.3385186,3.3576362,2.1881225,2.1805773,2.082489,1.8674494,1.4750963,1.0638802,1.0223814,1.0525624,1.146878,1.3468271,1.599593,1.750498,1.2411937,0.8865669,0.7582976,0.724344,0.43007925,0.35085413,0.3470815,0.3734899,0.38858038,0.35085413,0.7432071,0.8224323,0.7507524,0.6752999,0.7205714,0.7394345,2.093807,4.032936,6.043745,7.8621507,5.304311,3.9612563,3.9688015,4.881777,5.670255,3.8782585,6.258785,8.397863,8.786444,8.816625,9.303293,6.7114997,4.1762958,2.9728284,2.5012503,2.3465726,2.2069857,4.0970707,7.635793,10.023865,9.6201935,7.020855,5.8664317,6.9944468,8.469543,9.854096,10.767072,10.570895,9.699419,9.635284,8.07719,5.7909794,3.8895764,3.6481283,6.5002327,5.7494807,3.8971217,2.7426984,2.8030603,3.3048196,2.6332922,2.4899325,3.229367,4.123479,3.3915899,3.6745367,3.7537618,3.519859,3.059599,2.6446102,2.546522,2.2258487,1.8561316,1.6260014,1.7542707,2.2975287,1.9466745,1.1996948,0.482896,0.14713238,0.39989826,0.29426476,0.17731337,0.150905,0.05281675,0.02263575,0.056589376,0.0754525,0.05281675,0.0150905,0.02263575,0.211267,0.362172,0.3734899,0.23767537,0.056589376,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.056589376,0.02263575,0.00754525,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.003772625,0.003772625,0.00754525,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.049044125,0.17354076,0.29803738,0.16222288,0.033953626,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.041498873,0.056589376,0.08677038,0.17354076,0.26408374,0.35462674,0.392353,0.35462674,0.27917424,0.32821837,0.3169005,0.3055826,0.31312788,0.30181,0.21503963,0.20372175,0.2678564,0.38480774,0.52439487,0.7167987,1.0110635,1.1695137,1.0940613,0.8299775,0.8299775,0.7469798,0.58475685,0.38103512,0.19994913,0.07922512,0.041498873,0.033953626,0.026408374,0.018863125,0.0150905,0.02263575,0.030181,0.03772625,0.030181,0.05281675,0.0754525,0.071679875,0.06790725,0.13958712,0.41498876,0.66020936,0.66775465,0.47157812,0.32821837,0.1659955,0.10940613,0.116951376,0.1659955,0.241448,0.271629,0.27540162,0.5281675,1.1355602,2.022127,2.5804756,2.6446102,2.4974778,2.4220252,2.704972,3.0030096,2.6785638,2.4069347,2.6031113,3.4142256,5.2590394,6.771862,7.17176,6.175787,3.9876647,3.048281,3.4179983,5.093044,7.5792036,9.88805,9.050528,6.2399216,4.0593443,3.4368613,3.6028569,3.5689032,3.108643,2.4899325,1.9240388,1.5430037,1.0601076,0.6187105,0.3772625,0.3470815,0.3734899,0.43385187,0.42630664,0.38480774,0.30181,0.124496624,0.0754525,0.08299775,0.124496624,0.16976812,0.19240387,0.271629,0.41498876,0.5583485,0.69793564,0.8865669,0.9922004,0.995973,0.9922004,1.0638802,1.2902378,1.2449663,1.0902886,1.2487389,1.871222,2.8445592,2.5691576,2.4559789,2.6898816,3.2821836,4.0480266,3.4179983,3.0331905,2.927557,3.0860074,3.4444065,3.0633714,2.8521044,2.9501927,3.5877664,5.0439997,9.367428,13.502225,15.181043,13.928532,11.057564,11.2801485,13.124963,15.0376835,15.513034,13.117417,10.269085,11.400873,13.800262,15.746937,16.516552,16.463736,14.562332,13.445636,13.88326,14.769827,15.347038,15.735619,15.656394,14.984866,13.728582,14.136025,15.328176,17.316349,19.010258,18.229324,15.245177,11.510279,8.990166,9.148616,12.96274,14.452927,12.155397,10.887795,11.970539,13.215506,15.256495,16.418465,17.003222,17.21826,17.165443,16.16947,14.286931,12.185578,10.416218,9.382519,11.246195,12.66093,13.588995,13.898351,13.332457,11.548005,9.495697,8.975075,10.676529,14.154889,14.060574,15.603577,17.780382,19.281887,18.500954,14.713238,11.721546,10.197406,10.159679,10.9594755,11.721546,11.491416,10.702937,9.673011,8.624221,7.673519,7.496206,6.937857,5.80607,4.878004,4.7120085,4.293247,3.863168,3.4179983,2.71629,2.0862615,1.4713237,1.0525624,0.8601585,0.80734175,0.84884065,0.724344,0.59607476,0.5394854,0.55080324,0.5357128,0.5281675,0.58475685,0.694163,0.77338815,0.724344,0.62625575,0.58098423,0.62248313,0.7054809,0.7054809,0.73566186,0.7696155,0.7997965,0.83752275,0.79602385,0.84884065,0.965792,1.0638802,1.0223814,1.3015556,1.3166461,0.995973,0.482896,0.150905,0.124496624,0.120724,0.10940613,0.08299775,0.041498873,0.08299775,0.120724,0.14335975,0.14335975,0.1056335,0.12826926,0.181086,0.23767537,0.30181,0.392353,0.5998474,1.2034674,2.1692593,3.3274553,4.38379,4.7950063,4.398881,3.7650797,3.2821836,3.169005,3.3878171,3.1916409,2.8143783,2.4974778,2.4974778,2.6672459,2.5578396,2.4710693,2.5427492,2.746471,2.916239,2.9049213,2.9351022,3.0558262,3.138824,3.2218218,3.651901,4.074435,4.429062,4.9119577,5.040227,5.2137675,4.659192,3.5236318,2.867195,2.282438,2.0862615,2.3465726,2.8030603,2.867195,3.6971724,3.7688525,3.3274553,2.5389767,1.4901869,0.875249,0.754525,1.0374719,1.5165952,1.8900851,2.565385,2.8898308,3.180323,3.5538127,3.9348478,4.7006907,5.794752,7.1264887,8.412953,9.167479,9.137298,8.835487,8.744945,9.175024,10.257768,10.861387,11.400873,12.102581,12.925014,13.562587,14.015302,13.913441,13.336229,12.513797,11.84227,11.185833,10.819888,10.921749,11.193378,10.876478,10.144588,9.861642,9.567377,9.031664,8.239413,7.9489207,7.816879,7.8696957,8.073418,8.341274,8.431817,8.303548,7.99042,7.5905213,7.277394,6.94163,5.8890676,4.640329,3.5764484,2.9351022,3.663219,5.0553174,5.934339,6.8661776,8.145098,9.782416,11.393328,12.042219,12.140307,12.113899,12.404391,13.004238,13.517315,12.498707,10.035183,7.752744,6.4210076,5.934339,5.3269467,4.496969,4.164978,4.0178456,3.8556228,3.682082,3.5538127,3.5387223,3.6141748,3.2482302,2.0372176,0.62248313,0.67152727,0.6451189,0.5319401,0.38480774,0.24899325,0.150905,0.18863125,0.2263575,0.24522063,0.27917424,0.41121614,0.5357128,0.6828451,0.8111144,0.8224323,0.58098423,0.76207024,0.9922004,1.1883769,1.2864652,1.2525115,2.1805773,3.3463185,4.2064767,4.346064,3.4783602,3.150142,3.6179473,4.4403796,5.2967653,5.96452,6.760544,6.1908774,5.0854983,4.085753,3.6481283,5.149633,6.1003346,7.432071,9.22784,10.740664,10.570895,9.027891,7.8998766,7.7904706,8.13378,8.303548,6.862405,5.983383,6.092789,5.873977,5.4212623,6.590776,7.884786,8.458225,8.118689,7.043491,5.8400235,6.304056,8.114917,8.835487,8.786444,8.627994,8.29223,7.643338,6.470052,5.6778007,5.3684454,5.342037,5.372218,5.20245,4.617693,3.6934,2.3918443,1.5731846,2.9766011,3.2557755,2.987919,2.516341,2.1202152,1.9994912,2.071171,1.9994912,1.7316349,1.4109617,1.3732355,1.1280149,0.8865669,0.6790725,0.5357128,0.47157812,0.6187105,0.80356914,0.95447415,1.0035182,0.87147635,0.965792,0.90920264,0.7922512,0.68661773,0.62625575,0.62625575,0.73566186,0.8865669,1.0223814,1.0827434,0.98465514,1.1242423,1.1921495,1.0601076,0.7922512,0.7922512,2.595566,3.9084394,4.13857,4.395108,6.7869525,5.406172,3.6443558,2.9351022,2.776652,2.9954643,4.3347464,5.828706,8.379,14.724555,21.594505,17.301258,10.487898,5.613666,2.9313297,2.3918443,2.5238862,3.2670932,4.859141,7.8131065,9.4127,8.7600355,8.933576,9.457971,6.270103,3.440634,2.1466236,1.901403,2.6634734,4.8365054,3.8858037,1.961765,1.0789708,2.704972,7.7829256,6.964266,5.1760416,4.870459,6.013564,6.089017,4.4894238,3.1916409,2.7238352,3.31991,4.9421387,5.4212623,5.4740787,5.2137675,4.7535076,4.2404304,5.2665844,5.451443,4.7648253,3.3048196,1.267602,2.867195,2.9464202,2.1390784,1.026154,0.120724,0.3169005,0.68661773,0.8941121,0.7582976,0.26031113,0.11317875,0.27917424,0.36971724,0.26031113,0.0754525,0.06413463,0.52062225,0.7696155,0.60362,0.27540162,0.1056335,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056589376,0.27540162,0.116951376,0.030181,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.18485862,0.56589377,1.0902886,0.5998474,0.12826926,0.041498873,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.041498873,0.090543,0.17354076,0.32067314,0.38103512,0.41498876,0.41498876,0.35085413,0.1659955,0.13204187,0.13958712,0.1659955,0.15467763,0.0452715,0.00754525,0.00754525,0.026408374,0.049044125,0.060362,0.049044125,0.28294688,0.63002837,0.965792,1.1581959,1.5505489,1.5203679,1.2751472,0.94692886,0.58098423,0.21503963,0.0754525,0.041498873,0.030181,0.030181,0.018863125,0.00754525,0.00754525,0.018863125,0.030181,0.041498873,0.026408374,0.00754525,0.00754525,0.030181,0.090543,0.16976812,0.4074435,0.7054809,0.7167987,0.362172,0.21881226,0.21503963,0.31312788,0.5357128,0.6451189,0.46026024,0.97333723,2.033445,2.3503454,1.9353566,1.3355093,1.2562841,2.093807,3.9348478,4.0216184,2.7087448,2.003264,2.5616124,3.6481283,3.682082,3.308592,3.5085413,3.953711,2.9766011,3.3048196,4.3309736,5.5004873,6.0550632,5.0062733,3.9914372,3.218049,2.7728794,2.8596497,3.7990334,3.8254418,3.3538637,2.6144292,1.9844007,1.9844007,1.6675003,1.2223305,0.73188925,0.31312788,0.090543,0.1056335,0.21503963,0.30181,0.26031113,0.0150905,0.05281675,0.08677038,0.124496624,0.15467763,0.1659955,0.23013012,0.3734899,0.5319401,0.663982,0.76207024,0.8111144,0.8224323,0.8978847,1.0714256,1.327964,1.6335466,1.5882751,1.7655885,2.282438,2.806833,2.806833,2.5691576,2.5993385,2.9351022,3.1425967,2.886058,2.5201135,2.354118,2.4333432,2.516341,2.516341,2.3993895,2.293756,2.4672968,3.3123648,7.4018903,14.747191,19.31584,19.066847,15.992157,14.011529,14.388792,15.860115,16.120426,11.812089,8.552541,7.9451485,10.084227,13.660675,15.992157,14.611377,12.913695,12.50248,13.562587,14.830189,14.441608,14.754736,16.177015,17.30503,14.924504,15.399856,17.029629,19.444109,21.583187,21.681276,21.31533,17.670975,12.540206,8.59404,9.4013815,9.703192,9.880505,9.876732,9.771099,9.797507,11.615912,14.211478,16.263786,16.957949,16.007248,15.467763,14.815099,13.622949,12.242168,11.763044,14.973549,15.603577,15.128226,14.332202,13.321139,12.551523,10.182315,9.857869,12.053536,14.068119,13.604086,15.456445,18.202915,20.002459,18.58395,14.203933,11.962994,11.091517,10.899114,10.789707,10.506761,9.944639,9.039209,8.073418,7.6584287,6.719045,4.919503,3.4444065,2.8785129,3.218049,3.4029078,3.218049,3.187868,3.1048703,2.0447628,1.5316857,1.5052774,1.5731846,1.478869,1.0978339,0.965792,0.8563859,0.72811663,0.5885295,0.5017591,0.4678055,0.48666862,0.5772116,0.77338815,1.1280149,1.1657411,1.0450171,0.9016574,0.875249,1.1431054,1.0940613,0.90920264,0.7394345,0.7167987,0.9620194,0.8865669,0.8224323,0.7922512,0.8526133,1.0827434,1.3166461,1.20724,0.8865669,0.47157812,0.090543,0.1056335,0.116951376,0.10940613,0.07922512,0.030181,0.030181,0.02263575,0.02263575,0.033953626,0.0452715,0.056589376,0.1056335,0.17354076,0.24899325,0.32067314,0.41876137,0.5696664,1.0450171,1.931584,3.127506,4.2894745,4.878004,4.4894238,3.5123138,3.1576872,3.3651814,3.4896781,3.4557245,3.1539145,2.4710693,2.0070364,2.0485353,2.293756,2.7238352,3.6028569,4.2102494,4.346064,3.742444,2.795515,2.565385,2.5012503,2.4333432,2.3578906,2.2786655,2.1654868,2.704972,3.3953626,3.8065786,3.6707642,2.916239,2.7313805,2.3918443,1.8674494,1.3505998,1.267602,3.0860074,3.9989824,3.863168,2.9916916,2.1353056,1.0751982,0.5696664,0.46026024,0.59607476,0.83752275,1.9240388,2.7917426,3.5802212,4.376245,5.2175403,5.572167,6.138061,7.115171,8.484633,10.008774,10.401127,9.793735,9.220296,9.1825695,9.65792,9.7069645,9.865415,10.220041,10.827434,11.717773,13.196642,13.555041,13.230596,12.487389,11.41219,10.193633,9.457971,9.250477,9.386291,9.461743,9.265567,8.9788475,9.001483,9.397609,9.88805,9.948412,9.367428,8.5563135,7.779153,7.1566696,6.741681,6.3908267,6.0626082,5.764571,5.5683947,5.251494,4.7610526,4.1800685,3.5575855,2.897376,5.0175915,6.5341864,7.960239,9.2995205,10.26154,10.257768,9.525878,9.235386,9.691874,10.631257,11.257513,12.762791,12.751472,11.099063,8.575176,6.858632,4.8365054,3.8971217,3.4142256,2.8709676,1.8599042,1.9164935,2.2296214,2.505023,2.5578396,2.2711203,2.9992368,2.584248,1.5845025,0.6451189,0.48666862,0.5319401,0.45648763,0.33953625,0.23390275,0.17731337,0.14713238,0.1659955,0.18485862,0.181086,0.181086,0.22258487,0.29426476,0.331991,0.30935526,0.24899325,0.33576363,0.43007925,0.56212115,0.724344,0.87147635,1.1959221,1.4034165,1.5467763,1.6222287,1.5882751,1.8146327,2.4182527,4.0970707,6.4021444,7.748972,8.013056,8.001738,7.798016,7.3490734,6.4436436,6.888813,9.1976595,11.487643,12.702429,12.585477,10.616167,7.956466,6.862405,7.699928,8.952439,9.22784,8.511042,8.043237,8.224322,8.60913,8.5563135,8.850578,10.020092,10.9594755,8.948667,7.9715567,7.9225125,9.076936,11.114153,13.094781,12.449662,10.868933,8.869441,6.8246784,4.979865,4.0216184,3.5990841,3.6028569,3.874486,4.2027044,4.3083377,4.274384,3.904667,3.1237335,1.9994912,2.2107582,2.474842,2.7502437,3.029418,3.3161373,2.1994405,1.6146835,1.3656902,1.3128735,1.3732355,1.5015048,1.3770081,1.1506506,0.9280658,0.7922512,0.94692886,1.146878,1.3241913,1.4637785,1.6146835,2.2786655,1.9957186,1.9127209,2.3616633,2.848332,1.4524606,1.2110126,1.4524606,1.780679,2.0975795,2.252257,2.7426984,2.6031113,2.082489,2.625747,5.1232247,4.3800178,3.4934506,3.5424948,3.6141748,4.4818783,7.2396674,8.231868,7.069899,6.6586833,7.798016,9.993684,12.162943,13.004238,11.000975,8.20546,5.3609,3.5274043,3.0030096,3.2972744,4.3121104,5.8400235,9.0807085,12.713746,12.913695,10.891568,8.080963,6.0701537,5.111907,4.123479,3.9574835,4.112161,3.7499893,3.0218725,3.0671442,2.282438,2.1881225,4.006528,7.7037,11.981857,12.2270775,10.091772,6.488915,3.5953116,4.8327327,4.587512,4.0480266,3.5462675,3.4255435,4.0517993,3.983892,3.4179983,2.8747404,3.187868,5.485397,7.432071,9.291975,9.997457,8.326183,2.938875,3.0633714,3.2557755,3.187868,2.6106565,1.3656902,0.91674787,0.88279426,1.056335,1.267602,1.3807807,0.814887,0.6111652,0.5017591,0.35462674,0.16222288,0.041498873,0.1056335,0.15467763,0.15845025,0.24899325,0.09808825,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.0452715,0.011317875,0.056589376,0.02263575,0.00754525,0.0,0.003772625,0.011317875,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.00754525,0.018863125,0.018863125,0.0,0.011317875,0.030181,0.033953626,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.049044125,0.15845025,0.36971724,0.6111652,1.2487389,1.3015556,0.6413463,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.05281675,0.120724,0.150905,0.13958712,0.150905,0.16222288,0.14713238,0.120724,0.090543,0.033953626,0.026408374,0.026408374,0.033953626,0.030181,0.00754525,0.0,0.0,0.003772625,0.011317875,0.011317875,0.011317875,0.094315626,0.21503963,0.31312788,0.3055826,0.5093044,0.6526641,0.6790725,0.55457586,0.27540162,0.16222288,0.10940613,0.0754525,0.03772625,0.018863125,0.00754525,0.0,0.0,0.003772625,0.00754525,0.026408374,0.030181,0.02263575,0.011317875,0.00754525,0.018863125,0.120724,0.30181,0.47912338,0.52062225,0.3055826,0.17354076,0.116951376,0.124496624,0.181086,0.211267,0.3470815,0.68661773,1.1129243,1.2751472,0.9695646,0.66020936,0.56589377,0.784706,1.3015556,1.3770081,1.1431054,1.0638802,1.327964,1.8297231,2.0975795,2.6408374,3.2255943,3.5651307,3.2935016,3.2331395,5.330719,6.9567204,6.930312,5.5306683,3.6858547,3.1124156,3.0746894,3.1312788,3.1539145,2.757789,2.505023,2.0598533,1.5203679,1.4335974,1.5769572,1.6410918,1.3543724,0.80356914,0.45648763,0.3055826,0.23767537,0.22258487,0.20749438,0.08677038,0.056589376,0.06790725,0.0754525,0.071679875,0.08299775,0.16222288,0.29049212,0.4074435,0.49421388,0.543258,0.91297525,1.2638294,1.2487389,0.94315624,0.83752275,0.9393836,1.116697,1.4939595,2.2748928,3.7462165,3.3878171,2.9916916,3.0897799,3.482133,3.240685,2.897376,2.8445592,3.0897799,3.4896781,3.7499893,4.093298,4.6214657,5.0062733,4.7572803,3.2369123,4.61392,7.224577,9.457971,11.019837,12.96274,12.4307995,13.70972,15.218769,15.475307,13.079691,9.088254,8.533678,10.495442,13.717264,16.625957,12.551523,11.261286,11.717773,13.038192,14.5132885,15.792209,15.505488,15.192361,15.207452,14.739646,14.8339615,13.660675,14.147344,16.735365,19.349794,20.587215,18.176508,14.4152,11.249968,10.27663,10.193633,11.657412,13.057055,13.781399,14.226569,14.7170105,16.610868,16.984358,15.580941,14.7736,15.290449,15.588487,15.343266,14.920732,15.354584,16.11288,15.716756,14.437836,12.506252,10.148361,9.318384,9.220296,9.442881,9.839006,10.518079,11.751727,14.015302,15.569623,15.264041,12.51757,9.669238,8.107371,7.462252,7.3792543,7.492433,7.699928,7.6584287,7.201941,6.4549613,5.8664317,4.689373,3.440634,2.444661,1.8334957,1.5241405,1.4147344,1.3996439,1.5430037,1.6750455,1.3732355,1.4562333,1.5920477,1.6260014,1.5316857,1.4298248,1.3619176,1.3015556,1.2110126,1.0789708,0.90543,0.73188925,0.67152727,0.7054809,0.79602385,0.8978847,0.8639311,0.9997456,1.2147852,1.4260522,1.5467763,1.2826926,1.1393328,1.0186088,0.8978847,0.83752275,0.94315624,0.9507015,0.9016574,0.8526133,0.9016574,1.0525624,1.1242423,0.97710985,0.633801,0.27540162,0.19994913,0.1659955,0.14335975,0.1056335,0.06790725,0.03772625,0.02263575,0.0150905,0.033953626,0.094315626,0.1659955,0.13204187,0.13204187,0.19240387,0.24899325,0.32444575,0.46026024,0.7582976,1.418507,2.7125173,3.7650797,3.9197574,3.6481283,3.4330888,3.7801702,3.9499383,3.7047176,3.5424948,3.4745877,3.0331905,2.6974268,2.5540671,2.5201135,2.6144292,2.9652832,3.3727267,3.651901,3.4745877,3.0143273,2.9803739,2.546522,2.052308,1.7693611,1.7127718,1.6410918,2.052308,2.5012503,2.6219745,2.4484336,2.41448,2.203213,1.81086,1.3656902,0.97710985,0.76584285,1.267602,1.8636768,2.5012503,3.1954134,4.0404816,3.2029586,2.123988,1.0827434,0.43007925,0.59607476,1.1544232,2.123988,3.180323,4.032936,4.425289,5.451443,6.009792,6.7756343,8.062099,9.80128,10.691619,10.427535,9.710737,9.06939,8.83926,9.767326,10.148361,10.197406,10.1294985,10.133271,11.140562,11.838497,12.3289385,12.581704,12.415709,11.487643,10.472807,9.74469,9.420244,9.374973,9.5032425,9.367428,9.291975,9.333474,9.314611,8.937348,8.254503,7.5188417,6.851087,6.228604,5.73439,5.3269467,5.2175403,5.2364035,4.825187,4.2328854,3.8141239,3.4632697,3.127506,2.7879698,7.7904706,9.348565,9.80128,10.099318,10.570895,10.914205,11.559323,12.483616,12.611885,11.7894535,10.797253,12.385528,12.623203,11.261286,8.850578,6.719045,5.1081343,4.2064767,3.9084394,3.8593953,3.4594972,3.5764484,4.002755,4.06689,3.482133,2.3654358,1.9655377,1.5128226,0.9620194,0.46026024,0.331991,0.41498876,0.35839936,0.26408374,0.1961765,0.18485862,0.22258487,0.29049212,0.271629,0.16222288,0.094315626,0.09808825,0.13204187,0.14335975,0.12826926,0.120724,0.14713238,0.17731337,0.23390275,0.33953625,0.52062225,0.633801,0.633801,0.66020936,0.7582976,0.8865669,1.0374719,1.3505998,2.4333432,4.0216184,4.9723196,5.6551647,6.379509,6.8359966,6.8133607,6.198423,6.432326,8.246958,10.604849,12.415709,12.506252,9.74469,6.9944468,5.7683434,6.175787,6.9227667,7.9300575,8.578949,8.98262,9.26934,9.593785,9.337247,9.446653,10.201178,10.751981,9.137298,9.114662,9.808825,11.148107,12.936331,14.864142,11.993175,9.469289,7.466025,6.013564,5.0025005,4.353609,3.8141239,3.4632697,3.3727267,3.6141748,4.195159,4.4630156,4.6214657,4.61392,4.142342,3.3727267,2.9728284,2.8106055,2.7653341,2.7238352,2.1202152,1.5052774,1.1129243,1.0035182,1.0902886,1.2638294,1.1846043,1.026154,0.8903395,0.80734175,0.8337501,0.965792,1.1581959,1.3958713,1.690136,2.2258487,2.493705,2.6785638,2.8634224,3.0445085,2.5238862,2.8634224,3.821669,5.05909,6.149379,6.851087,7.333983,5.7796617,3.1425967,3.1463692,5.5683947,4.221567,3.470815,4.22534,3.9574835,3.4066803,4.7421894,5.481624,5.413717,6.6134114,8.469543,10.231359,11.106608,10.367173,7.322665,3.9725742,2.3088465,2.4710693,3.531177,3.5047686,3.6368105,4.22534,5.7494807,7.360391,6.8850408,5.5004873,4.315883,4.0216184,4.4403796,4.5196047,3.6934,2.746471,2.0145817,1.6486372,1.6071383,1.750498,2.2786655,3.8593953,6.1003346,7.5490227,8.088508,7.6282477,6.2361493,4.9157305,5.613666,7.5075235,7.779153,6.4247804,4.244203,2.8407867,3.731126,4.032936,3.9310753,3.9989824,5.1835866,6.458734,7.805561,8.265821,6.752999,2.0560806,2.8106055,3.8405323,4.534695,4.376245,2.9426475,1.539231,1.0374719,0.9695646,0.98842776,0.8865669,0.784706,0.7130261,0.6413463,0.5394854,0.40367088,0.16222288,0.094315626,0.07922512,0.071679875,0.09808825,0.03772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.018863125,0.05281675,0.071679875,0.0452715,0.0754525,0.090543,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.0,0.003772625,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.030181,0.030181,0.049044125,0.090543,0.1659955,0.21881226,0.573439,0.6375736,0.32067314,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.094315626,0.1358145,0.12826926,0.08299775,0.018863125,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.011317875,0.02263575,0.030181,0.033953626,0.1056335,0.16976812,0.181086,0.1358145,0.08677038,0.06790725,0.03772625,0.018863125,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.0452715,0.060362,0.03772625,0.10186087,0.17354076,0.211267,0.181086,0.07922512,0.060362,0.06790725,0.13204187,0.23013012,0.3169005,0.32067314,0.15467763,0.03772625,0.02263575,0.00754525,0.011317875,0.011317875,0.0150905,0.011317875,0.0,0.00754525,0.06413463,0.14713238,0.23013012,0.27917424,0.19994913,0.124496624,0.07922512,0.071679875,0.08299775,0.10186087,0.23390275,0.44894236,0.6375736,0.6149379,0.41876137,0.28294688,0.24522063,0.29049212,0.3470815,0.38480774,0.3961256,0.422534,0.5093044,0.68661773,1.0827434,1.8674494,2.6634734,3.0181,2.4031622,2.916239,5.2552667,7.4018903,8.190369,7.3075747,5.534441,4.666737,4.1498876,3.5953116,2.7804246,1.9730829,1.6033657,1.3468271,1.1091517,1.0148361,1.086516,1.2223305,1.1280149,0.77338815,0.40367088,0.33953625,0.33576363,0.33576363,0.2867195,0.14335975,0.13958712,0.14335975,0.13204187,0.1056335,0.08677038,0.1659955,0.27540162,0.3734899,0.47157812,0.62625575,0.965792,1.3091009,1.297783,0.9393836,0.5885295,0.62248313,0.8299775,1.4600059,2.637065,4.3385186,4.9647746,4.689373,4.247976,3.8443048,3.138824,2.6408374,2.5616124,2.9464202,3.62172,4.195159,4.749735,5.43258,5.938112,6.1795597,6.296511,7.884786,7.745199,8.756263,10.899114,11.2650585,8.171506,8.692128,11.080199,13.313594,13.094781,10.216269,8.9788475,9.737145,12.098808,14.909414,13.109872,11.69891,10.653893,10.401127,11.815862,14.471789,16.199652,16.708956,16.22606,15.490398,15.226315,14.339747,14.766054,16.622187,18.191597,18.368912,16.539188,14.030393,11.92904,11.057564,12.359119,14.698147,16.286423,16.912678,17.942604,16.946632,16.01102,14.452927,12.81938,12.853333,14.456699,15.671484,16.576914,16.678776,14.913187,14.366156,13.6682205,12.491161,10.853842,9.107117,8.616675,8.397863,8.171506,7.9451485,8.016829,10.49167,12.483616,12.974057,11.838497,9.839006,7.745199,6.609639,6.017337,5.6551647,5.311856,5.6589375,5.6363015,5.240176,4.689373,4.429062,3.8895764,3.0897799,2.3201644,1.7354075,1.3091009,1.0299267,1.2449663,1.6825907,2.1503963,2.5238862,3.0030096,2.7841973,2.2899833,1.8599042,1.7127718,1.7655885,1.7429527,1.6561824,1.5165952,1.327964,1.1846043,1.0525624,0.935611,0.84884065,0.8224323,0.9242931,1.267602,1.6486372,1.901403,1.8749946,1.5882751,1.5430037,1.6637276,1.7429527,1.4298248,1.0789708,0.8903395,0.784706,0.7205714,0.69793564,0.79602385,1.0186088,0.98842776,0.66020936,0.32821837,0.32067314,0.2867195,0.26408374,0.241448,0.1659955,0.10940613,0.06413463,0.049044125,0.071679875,0.1056335,0.19994913,0.30935526,0.32067314,0.2565385,0.28294688,0.32067314,0.41876137,0.62248313,1.1883769,2.5729303,3.9725742,4.3686996,4.1536603,3.7348988,3.5349495,3.531177,3.4859054,3.6556737,3.9197574,3.7688525,3.229367,2.8709676,2.6521554,2.6031113,2.8181508,3.1350515,3.2520027,3.0822346,2.8521044,3.0822346,2.6446102,2.123988,1.8259505,1.7844516,1.7655885,1.9240388,2.0787163,2.0070364,1.7542707,1.6033657,1.3770081,1.2713746,1.388326,1.720317,2.1805773,1.9542197,1.7655885,1.7354075,1.9353566,2.384299,2.123988,1.4713237,0.7432071,0.27917424,0.43385187,0.814887,1.5316857,2.4786146,3.4896781,4.327201,5.2967653,5.9230213,6.651138,7.6320205,8.726082,10.133271,10.144588,9.5183325,8.963757,9.129752,9.752235,9.865415,9.710737,9.49947,9.431562,9.869187,10.435081,11.242422,12.23085,13.151371,12.815607,11.593277,10.291721,9.424017,9.1976595,9.325929,9.061845,8.6732645,8.333729,8.126234,7.6093845,6.9869013,6.3945994,5.87775,5.3910813,4.9987283,4.659192,4.485651,4.3686996,4.006528,3.5236318,3.1576872,2.8898308,2.6823363,2.516341,11.921495,13.200415,13.000465,12.593022,12.657157,13.29473,14.456699,15.373446,14.66042,12.47607,10.502988,10.785934,10.33322,8.952439,7.073672,5.7494807,5.2665844,4.82896,4.5497856,4.38379,4.1498876,4.274384,4.644101,4.8138695,4.285702,2.5238862,1.448688,1.0525624,0.7432071,0.38480774,0.30181,0.3734899,0.35839936,0.29426476,0.23390275,0.2263575,0.24522063,0.30181,0.331991,0.29049212,0.17354076,0.11317875,0.090543,0.090543,0.090543,0.090543,0.0754525,0.07922512,0.090543,0.14335975,0.28294688,0.32821837,0.35085413,0.422534,0.55080324,0.6790725,0.67152727,0.7092535,1.0412445,1.629774,2.1692593,3.9273026,5.292993,6.085244,6.304056,6.149379,6.217286,6.937857,8.333729,9.891823,10.552032,8.661947,6.881268,6.0701537,6.368191,7.220804,7.8508325,8.846806,9.522105,9.673011,9.574923,9.435335,9.910686,10.461489,10.567122,9.7296,9.778644,10.31813,11.000975,11.676274,12.37421,9.661693,7.809334,6.6247296,5.956975,5.6778007,5.560849,5.6589375,5.3571277,4.6214657,3.9725742,4.221567,4.315883,4.429062,4.6252384,4.889322,4.353609,3.802806,3.2331395,2.6483827,2.082489,1.9278114,1.8825399,1.5920477,1.1091517,0.875249,0.87902164,0.8262049,0.8337501,0.91297525,0.9695646,0.9205205,0.90920264,0.97710985,1.1506506,1.4637785,1.9504471,2.637065,2.9351022,2.8030603,2.746471,3.0558262,3.8405323,5.4438977,7.2698483,7.798016,7.752744,7.8206515,5.836251,2.7087448,2.41448,3.6896272,2.8445592,3.2633207,4.8440504,4.014073,3.8895764,5.379763,6.6322746,7.3981175,9.035437,9.937095,9.808825,8.492179,6.432326,4.689373,3.1124156,2.2107582,2.5880208,3.5953116,3.3236825,2.637065,2.214531,2.2107582,2.3918443,2.123988,2.282438,2.7841973,3.5877664,4.244203,3.8782585,2.5201135,1.3468271,1.0751982,1.4939595,1.4750963,1.9240388,2.263575,3.108643,4.0970707,3.8895764,4.3686996,5.0062733,5.6589375,6.273875,6.8925858,9.510788,10.061591,8.507269,5.8211603,3.9650288,4.561104,5.270357,5.7796617,5.885295,5.485397,6.368191,7.3188925,7.7112455,6.888813,4.142342,4.715781,5.7004366,6.5266414,6.677546,5.692891,3.1199608,1.9655377,1.4977322,1.1695137,0.63002837,0.6790725,1.086516,1.4373702,1.4713237,1.056335,0.58475685,0.32067314,0.17354076,0.0754525,0.0,0.0,0.02263575,0.06413463,0.12826926,0.20749438,0.23013012,0.15845025,0.10186087,0.1056335,0.1358145,0.08677038,0.094315626,0.094315626,0.06413463,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0,0.00754525,0.03772625,0.094315626,0.15845025,0.120724,0.08299775,0.049044125,0.030181,0.03772625,0.02263575,0.00754525,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.094315626,0.1358145,0.12826926,0.08299775,0.018863125,0.011317875,0.003772625,0.011317875,0.049044125,0.120724,0.11317875,0.0754525,0.041498873,0.02263575,0.026408374,0.07922512,0.124496624,0.150905,0.15845025,0.14335975,0.20749438,0.21881226,0.181086,0.11317875,0.05281675,0.026408374,0.00754525,0.003772625,0.00754525,0.02263575,0.056589376,0.06413463,0.060362,0.06413463,0.07922512,0.030181,0.00754525,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.1056335,0.25276586,0.41498876,0.58475685,0.38103512,0.17731337,0.10940613,0.0754525,0.060362,0.03772625,0.018863125,0.00754525,0.00754525,0.0150905,0.026408374,0.0452715,0.06790725,0.09808825,0.090543,0.071679875,0.06413463,0.07922512,0.094315626,0.1056335,0.15845025,0.271629,0.38103512,0.331991,0.2678564,0.241448,0.24522063,0.23767537,0.16976812,0.124496624,0.1056335,0.1056335,0.12826926,0.19994913,0.58475685,1.3543724,2.0560806,2.2711203,1.6448646,2.444661,4.2328854,6.247467,7.677292,7.6697464,6.888813,6.277648,5.4703064,4.293247,2.7540162,1.6976813,1.1959221,1.0148361,0.97710985,0.9393836,0.94315624,1.0336993,0.95447415,0.6526641,0.2867195,0.25276586,0.2867195,0.32821837,0.31312788,0.17354076,0.18485862,0.19240387,0.19240387,0.17354076,0.14335975,0.2263575,0.33576363,0.43385187,0.5281675,0.6790725,0.845068,0.995973,0.97333723,0.7507524,0.44139713,0.44894236,0.58098423,1.1695137,2.3126192,3.85185,4.9157305,4.8742313,4.168751,3.240685,2.516341,2.4408884,2.776652,3.451952,4.104616,4.074435,4.436607,4.908185,5.3759904,6.1003346,7.7301087,10.861387,10.785934,10.842525,11.193378,8.827943,5.7494807,5.915476,7.9451485,10.280403,11.185833,9.582467,8.047009,8.001738,9.797507,12.728837,13.404137,12.027128,10.035183,8.91094,10.212496,13.170234,15.546988,16.980585,17.53139,17.682293,17.886015,17.587978,17.584206,18.025602,18.406637,18.089737,16.094019,14.102073,12.974057,12.736382,14.5283785,15.946886,16.618414,17.13149,19.047983,19.149845,16.558052,13.788944,12.3893,12.928786,14.728328,15.380992,15.62244,15.226315,12.996693,12.1101265,12.117672,12.128989,11.695138,10.785934,9.857869,8.741172,8.031919,7.960239,8.382772,10.797253,12.00072,12.245941,12.064855,12.298758,11.4838705,10.552032,9.001483,6.907676,4.9044123,4.4931965,4.3422914,4.187614,4.055572,4.2328854,4.315883,4.025391,3.482133,2.8596497,2.3880715,2.0145817,2.0787163,2.5993385,3.3953626,4.055572,4.4931965,4.002755,3.1237335,2.3428001,2.0787163,2.123988,2.1202152,2.0598533,1.9429018,1.7542707,1.6335466,1.4750963,1.2902378,1.116697,1.0035182,1.1883769,1.5430037,1.841041,1.9164935,1.6939086,1.4071891,1.418507,1.659955,1.8636768,1.5769572,1.1619685,0.935611,0.7922512,0.694163,0.65643674,0.65643674,0.8337501,0.86770374,0.67152727,0.422534,0.38858038,0.3055826,0.24899325,0.21881226,0.16222288,0.1659955,0.15845025,0.13958712,0.116951376,0.11317875,0.1961765,0.34330887,0.3772625,0.31312788,0.33953625,0.331991,0.3961256,0.5281675,0.91297525,1.901403,3.338773,4.06689,4.1762958,3.9008942,3.6066296,3.308592,3.2067313,3.4179983,3.7952607,3.9461658,3.4896781,2.9992368,2.6106565,2.4522061,2.6597006,3.108643,3.361409,3.2482302,2.9615107,3.0822346,2.886058,2.4823873,2.1202152,1.8938577,1.7354075,1.5882751,1.4562333,1.3241913,1.1732863,0.9808825,0.76207024,0.8563859,1.3656902,2.1390784,2.757789,2.2673476,1.6939086,1.2562841,1.0789708,1.20724,1.1846043,0.9393836,0.6752999,0.52062225,0.5357128,0.8224323,1.3505998,2.1805773,3.2142766,4.187614,4.9949555,5.7117543,6.3342376,6.900131,7.492433,9.016574,9.559832,9.382519,9.110889,9.710737,9.695646,9.522105,9.344792,9.2844305,9.450426,9.57115,9.782416,10.355856,11.393328,12.864652,12.860879,11.680047,10.272858,9.307066,9.1976595,9.246704,8.82417,8.2507305,7.7225633,7.333983,6.790725,6.228604,5.696664,5.2288585,4.8365054,4.5233774,4.2404304,3.9612563,3.6745367,3.3764994,3.0369632,2.727608,2.493705,2.3428001,2.2447119,15.788436,16.576914,16.675003,16.693865,16.950403,17.463482,17.025856,15.882751,13.864397,11.506506,10.016319,8.8618965,7.0887623,5.1534057,3.783943,3.9801195,5.1647234,5.4665337,4.9987283,4.044254,3.0709167,3.078462,3.5538127,4.327201,4.557331,2.7087448,1.5807298,1.146878,0.8111144,0.4376245,0.3470815,0.3734899,0.392353,0.36594462,0.30935526,0.2867195,0.20372175,0.18485862,0.29049212,0.4074435,0.271629,0.15845025,0.08299775,0.06413463,0.08299775,0.08677038,0.060362,0.049044125,0.049044125,0.0754525,0.150905,0.150905,0.17731337,0.24522063,0.362172,0.52062225,0.52439487,0.5017591,0.633801,1.0450171,1.7919968,4.4215164,6.126743,7.020855,7.3377557,7.413208,7.009537,6.749226,6.647365,6.7944975,7.322665,7.164215,6.8774953,7.1566696,8.216777,9.808825,9.035437,9.627739,10.178542,10.114408,9.684328,9.997457,10.902886,11.521597,11.570641,11.363147,10.989656,10.970794,10.518079,9.457971,8.190369,7.3981175,7.3188925,7.141579,6.722818,6.5832305,6.964266,7.8734684,7.8206515,6.5266414,4.9421387,4.3686996,3.953711,3.6934,3.6292653,3.8405323,4.568649,4.5799665,4.08198,3.2935016,2.4522061,2.1843498,2.848332,2.886058,1.9957186,1.1431054,0.76207024,0.6451189,0.80734175,1.1091517,1.2789198,1.2261031,1.0751982,0.98465514,1.0223814,1.1732863,1.7127718,2.3465726,2.6295197,2.5616124,2.584248,2.837014,3.4670424,4.961002,6.4436436,5.696664,4.3347464,3.8292143,2.6823363,1.3807807,2.425798,2.505023,1.8863125,3.1539145,5.2892203,3.6669915,5.040227,8.741172,11.257513,11.800771,12.306303,11.231105,9.092027,6.4021444,3.9876647,2.987919,2.2711203,1.8674494,2.0372176,2.5540671,2.7011995,2.1390784,1.6675003,1.8485862,2.535204,2.8332415,3.6066296,4.3121104,4.485651,3.85185,2.323937,1.4222796,1.2034674,1.6825907,2.3013012,1.931584,1.9881734,1.9164935,2.444661,3.3236825,3.3048196,4.214022,5.0515447,5.7419353,6.304056,6.8699503,8.722309,9.35611,8.809079,7.567886,6.5568223,5.4967146,5.847569,6.9152217,7.6848373,6.828451,7.8961043,9.133525,9.899368,9.5183325,7.303802,7.152897,7.201941,7.360391,7.5112963,7.533932,4.7120085,3.361409,2.806833,2.493705,1.9957186,1.1544232,1.5769572,2.2107582,2.3578906,1.7014539,1.1129243,0.62625575,0.29049212,0.11317875,0.056589376,0.026408374,0.06790725,0.1659955,0.30935526,0.4640329,0.47912338,0.3169005,0.16976812,0.11317875,0.120724,0.08299775,0.03772625,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.003772625,0.0150905,0.09808825,0.23013012,0.33953625,0.27917424,0.16222288,0.056589376,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.09808825,0.24899325,0.2263575,0.15467763,0.0754525,0.026408374,0.03772625,0.15467763,0.2263575,0.26031113,0.26031113,0.23013012,0.26031113,0.211267,0.13204187,0.06413463,0.011317875,0.003772625,0.0,0.003772625,0.0150905,0.026408374,0.116951376,0.12826926,0.124496624,0.12826926,0.15845025,0.060362,0.018863125,0.011317875,0.033953626,0.090543,0.10186087,0.094315626,0.05281675,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.071679875,0.20749438,0.5281675,0.452715,0.28294688,0.17731337,0.13958712,0.26408374,0.25276586,0.16976812,0.071679875,0.033953626,0.03772625,0.03772625,0.026408374,0.018863125,0.0150905,0.0150905,0.02263575,0.0452715,0.08299775,0.10940613,0.09808825,0.10940613,0.14713238,0.20372175,0.2565385,0.2867195,0.33953625,0.362172,0.32067314,0.20749438,0.08299775,0.0452715,0.0452715,0.0754525,0.1659955,0.4376245,1.0978339,1.5165952,1.5279131,1.4449154,2.0975795,2.9728284,4.2064767,5.541986,6.33801,6.6134114,6.6134114,5.945657,4.5761943,2.8332415,1.9391292,1.4222796,1.1921495,1.146878,1.1846043,1.2487389,1.3166461,1.116697,0.6526641,0.23390275,0.12826926,0.10940613,0.16222288,0.21881226,0.16222288,0.15845025,0.181086,0.20372175,0.211267,0.1961765,0.27917424,0.392353,0.49044126,0.56212115,0.6073926,0.62248313,0.58475685,0.51684964,0.43007925,0.33953625,0.31312788,0.33953625,0.6149379,1.2789198,2.4220252,3.097325,3.3236825,2.8822856,2.0900342,1.7957695,2.444661,3.350091,4.2328854,4.5837393,3.6443558,3.6066296,3.6858547,3.9725742,4.708236,6.273875,10.284176,11.868678,11.400873,9.593785,7.4811153,7.9791017,7.9941926,8.043237,8.431817,9.239159,8.443134,7.1000805,6.8850408,8.409182,11.242422,12.355347,11.2801485,9.661693,8.884532,10.057818,12.249713,13.124963,14.494425,16.818363,19.191343,20.643805,20.583443,19.862871,19.357338,19.930779,20.57967,18.65563,16.659912,15.739391,15.667711,16.003475,14.996184,14.0983,14.437836,16.795727,19.364883,17.508753,14.962231,13.9888935,15.384765,16.708956,15.811071,13.9888935,12.525115,12.694883,12.381755,13.287186,14.4114275,14.890551,13.973803,12.045992,10.344538,9.450426,9.646602,10.884023,12.687338,13.932304,15.531898,17.542706,19.191343,19.772327,18.72731,15.430037,10.593531,6.247467,4.7006907,4.515832,4.938366,5.587258,6.4549613,6.470052,6.33801,5.7872066,4.930821,4.285702,3.7348988,3.2935016,3.5651307,4.447925,5.1269975,5.168496,4.659192,3.772625,2.8898308,2.595566,2.565385,2.5389767,2.4861598,2.3880715,2.252257,2.0636258,1.8976303,1.7354075,1.5769572,1.418507,1.5279131,1.7052265,1.7542707,1.5807298,1.1883769,0.8978847,0.9280658,1.1280149,1.3166461,1.2864652,1.2638294,1.1581959,0.97333723,0.77716076,0.7092535,0.6111652,0.6149379,0.6526641,0.6413463,0.48666862,0.35085413,0.211267,0.120724,0.08299775,0.07922512,0.18863125,0.2565385,0.23767537,0.15845025,0.124496624,0.17731337,0.211267,0.24522063,0.27540162,0.31312788,0.29426476,0.34330887,0.42630664,0.56589377,0.87147635,1.8599042,2.7200627,3.361409,3.8065786,4.191386,3.8065786,3.3312278,3.1312788,3.3010468,3.6481283,3.5839937,3.0181,2.4371157,2.1881225,2.4861598,3.2633207,3.8367596,3.7990334,3.2784111,2.9615107,3.0709167,2.9426475,2.5238862,1.9240388,1.4147344,1.0374719,0.76584285,0.72811663,0.8563859,0.87147635,0.59230214,0.6451189,1.1204696,1.7693611,1.9881734,1.6071383,1.1619685,0.94692886,1.1053791,1.6146835,1.5354583,1.2826926,1.20724,1.2864652,1.1242423,1.0978339,1.4977322,2.203213,3.0181,3.6669915,4.485651,5.27413,5.7494807,6.0211096,6.587003,7.8206515,8.944894,9.491924,9.64283,10.208723,9.774872,9.484379,9.469289,9.7220545,10.069136,10.174769,10.125726,10.197406,10.702937,11.989402,11.846043,10.812344,9.676784,9.0543,9.390063,9.442881,8.933576,8.269594,7.6282477,6.9491754,6.40969,5.8966126,5.3986263,4.927048,4.5460134,4.2291126,3.9461658,3.640583,3.308592,2.9916916,2.6898816,2.4484336,2.263575,2.1466236,2.082489,16.188334,16.712729,17.497435,18.912169,20.70794,22.00195,19.927006,16.388283,12.506252,9.590013,9.125979,9.465516,8.096053,5.885295,3.832987,3.0520537,6.4926877,7.564113,6.851087,5.119452,3.3274553,2.886058,4.06689,5.300538,5.5193505,4.1498876,1.720317,0.70170826,0.392353,0.32444575,0.27540162,0.24899325,0.23390275,0.23013012,0.23767537,0.27540162,0.24899325,0.21503963,0.17354076,0.124496624,0.0754525,0.041498873,0.030181,0.03772625,0.05281675,0.0754525,0.0754525,0.056589376,0.041498873,0.026408374,0.0150905,0.026408374,0.049044125,0.071679875,0.116951376,0.21503963,0.3961256,0.46026024,1.0714256,2.41448,4.195159,6.0626082,7.665974,8.703445,9.0957985,8.986393,7.8998766,6.934085,5.9494295,4.930821,3.9688015,4.13857,4.749735,6.360646,8.4544525,9.431562,8.099826,9.752235,11.272603,11.54046,11.442371,11.627231,12.193124,12.774108,13.355092,14.283158,15.490398,16.003475,14.977322,12.427027,9.216523,6.8246784,7.462252,8.039464,7.6810646,7.707473,8.29223,8.311093,7.4811153,6.1531515,5.311856,4.640329,3.5387223,3.2633207,3.9725742,4.7308717,5.2552667,5.221313,4.9534564,4.587512,4.074435,3.9159849,4.425289,4.534695,3.7914882,2.3654358,1.2789198,0.79602385,0.87147635,1.20724,1.267602,1.1431054,1.0223814,1.1016065,1.237421,0.9318384,0.8941121,1.2525115,1.8070874,2.2786655,2.305074,2.2447119,2.2560298,2.2183034,2.2296214,2.6106565,2.3767538,1.7354075,1.0450171,1.901403,7.1264887,6.5040054,3.8858037,4.2894745,6.7039547,4.104616,4.727099,6.511551,7.2283497,6.688864,6.7756343,5.50426,4.044254,3.1954134,2.6597006,1.0223814,0.52062225,0.83752275,1.8561316,2.7125173,1.7844516,1.5165952,1.7618159,2.4861598,3.6141748,5.0062733,5.1760416,5.247721,5.3571277,5.1345425,3.6934,2.4974778,1.5731846,0.9393836,0.5885295,0.5055317,0.68661773,0.77716076,0.7922512,0.80356914,0.9620194,4.085753,6.2021956,6.8925858,5.9796104,3.5236318,5.1232247,6.9227667,8.216777,8.254503,6.2399216,4.689373,5.2628117,6.937857,8.379,7.964011,8.4544525,9.5183325,9.805053,7.877241,2.214531,4.2517486,4.093298,3.0935526,2.493705,3.4330888,3.482133,3.7763977,4.346064,5.1081343,5.8890676,2.8521044,1.3770081,0.9016574,0.965792,1.237421,1.1732863,0.8563859,0.5281675,0.32821837,0.29049212,0.13204187,0.120724,0.181086,0.24522063,0.24522063,0.071679875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.10186087,0.27917424,0.47157812,0.47157812,0.24522063,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.018863125,0.060362,0.1659955,0.3961256,0.44516975,0.4376245,0.2678564,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.018863125,0.030181,0.7394345,0.8978847,0.694163,0.35085413,0.1056335,0.13204187,0.120724,0.0754525,0.026408374,0.0150905,0.0150905,0.00754525,0.00754525,0.02263575,0.060362,0.049044125,0.0452715,0.0452715,0.049044125,0.060362,0.060362,0.14335975,0.23390275,0.27917424,0.24522063,0.15845025,0.10186087,0.08299775,0.116951376,0.21503963,0.35839936,0.7167987,1.0450171,1.237421,1.3128735,2.372981,2.757789,3.2821836,4.2517486,5.4476705,5.119452,4.61392,3.904667,3.1048703,2.4559789,2.4672968,2.04099,1.6222287,1.4298248,1.4637785,1.4411428,1.4901869,1.2826926,0.7582976,0.1358145,0.08677038,0.0754525,0.071679875,0.06413463,0.0754525,0.10186087,0.150905,0.17731337,0.16976812,0.18485862,0.20749438,0.2678564,0.35462674,0.44894236,0.5357128,0.5583485,0.5357128,0.4640329,0.362172,0.29049212,0.25276586,0.19994913,0.27917424,0.56589377,1.0676528,1.8485862,2.4031622,2.372981,2.003264,2.1353056,2.5993385,2.8822856,3.0105548,3.0709167,3.2029586,3.218049,2.9539654,2.7540162,3.0030096,4.1498876,5.983383,7.5565677,8.179051,8.98262,12.940104,15.965749,13.5663595,11.32542,11.23865,11.7026825,11.691365,10.103089,9.408927,10.133271,10.86516,10.718028,9.7296,8.428044,7.665974,8.605357,9.752235,9.363655,9.95973,12.279895,15.260268,17.84829,19.1423,19.828917,20.65135,22.447119,24.069347,24.484337,23.043194,20.60985,19.56106,17.097536,14.0907545,11.759273,10.838752,11.581959,12.815607,13.223051,12.796744,13.309821,18.327412,19.828917,18.85558,16.407146,14.796235,17.637022,18.859352,18.953669,18.62545,17.80679,15.671484,13.754991,12.359119,11.291467,10.933067,12.253486,15.207452,19.855326,25.302996,29.128437,27.359077,27.332668,25.65385,21.092747,14.475562,8.650629,7.175533,7.1906233,8.2507305,10.080454,12.559069,11.374464,10.023865,8.529905,7.115171,6.224831,5.1873593,4.3611546,4.112161,4.5422406,5.492942,5.2137675,4.6290107,3.9574835,3.4255435,3.2821836,3.4142256,3.2935016,3.0407357,2.8521044,2.9615107,2.655928,2.3880715,2.1654868,2.003264,1.9089483,1.8599042,1.7995421,1.6863633,1.4826416,1.1883769,0.995973,1.0940613,1.3355093,1.5920477,1.7391801,1.6675003,1.4109617,1.0676528,0.7469798,0.56589377,0.5017591,0.48666862,0.482896,0.422534,0.23013012,0.19240387,0.17354076,0.1659955,0.1659955,0.150905,0.19994913,0.241448,0.241448,0.19994913,0.1358145,0.150905,0.16222288,0.14335975,0.1056335,0.1056335,0.15467763,0.22258487,0.30935526,0.43385187,0.6413463,1.0940613,1.9202662,2.848332,3.7160356,4.485651,4.90064,4.38379,3.7763977,3.5500402,3.7688525,3.8405323,3.0445085,2.2899833,2.1315331,2.7917426,3.9386206,4.1536603,3.7084904,2.987919,2.4861598,2.7313805,3.3048196,3.1652324,2.2183034,1.327964,1.0110635,0.9205205,1.177059,1.539231,1.418507,0.8224323,0.72811663,0.8601585,1.1204696,1.5731846,1.6675003,1.1883769,0.8865669,1.1016065,1.7844516,2.1277604,1.6712729,1.7769064,2.4672968,2.4559789,1.5769572,1.448688,1.6561824,2.0673985,2.837014,3.7537618,4.561104,5.149633,5.624984,6.270103,7.213259,8.216777,9.442881,10.54826,10.695392,10.291721,9.963503,10.238904,10.948157,11.216014,11.363147,11.498961,11.46878,11.491416,12.162943,11.54046,10.284176,9.144843,8.729855,9.537196,9.74469,9.163706,8.122461,6.9491754,5.9984736,5.4967146,5.168496,4.9119577,4.644101,4.304565,3.9386206,3.663219,3.380272,3.0520537,2.686109,2.4031622,2.2258487,2.1202152,2.0673985,2.0447628,13.773854,15.69412,15.931795,14.792462,13.068373,12.019584,12.336484,13.837989,14.230342,12.974057,11.310329,9.231613,6.6624556,4.285702,2.848332,3.150142,5.7306175,6.6549106,6.326692,5.292993,4.2404304,3.9386206,4.870459,5.3948536,4.776143,3.1727777,1.2147852,0.51684964,0.32821837,0.241448,0.19994913,0.18863125,0.1659955,0.13958712,0.116951376,0.116951376,0.10186087,0.08299775,0.0754525,0.071679875,0.05281675,0.033953626,0.02263575,0.030181,0.0452715,0.05281675,0.041498873,0.030181,0.026408374,0.030181,0.026408374,0.018863125,0.02263575,0.030181,0.056589376,0.1056335,0.19994913,0.3055826,0.5055317,0.8186596,1.1921495,2.0560806,3.500996,5.1835866,6.228604,5.240176,4.006528,3.7499893,3.6179473,3.2520027,2.795515,2.848332,3.429316,4.8025517,6.5530496,7.598067,7.567886,7.877241,8.639311,9.6051035,10.163452,10.725573,11.272603,11.197151,10.623712,10.401127,12.272349,15.199906,17.135263,17.014538,14.781145,12.487389,11.0613365,9.797507,8.631766,8.156415,8.050782,7.937603,7.7037,7.515069,7.8244243,7.786698,7.1981683,6.1908774,5.311856,5.523123,5.3344917,4.749735,3.953711,3.289729,3.2444575,3.62172,4.29702,4.9345937,5.1571784,4.538468,3.2746384,2.142851,1.5958204,1.5430037,1.3505998,1.3958713,1.5580941,1.8221779,1.9353566,1.3958713,1.0827434,1.0789708,1.3770081,1.8599042,2.305074,2.6446102,2.8596497,2.8785129,2.7841973,2.7917426,2.5616124,2.142851,1.6448646,1.6637276,3.2935016,3.6481283,3.3538637,3.399135,3.7613072,3.410453,3.4255435,3.2784111,2.6031113,1.8787673,2.4408884,2.2069857,1.7429527,1.2826926,0.8639311,0.35085413,0.4074435,0.9620194,1.8787673,2.6219745,2.2484846,1.8448136,1.9881734,2.7426984,4.0593443,5.772116,6.228604,6.0626082,5.4967146,4.82896,4.425289,3.863168,2.7426984,1.3543724,0.26031113,0.28294688,0.84884065,1.0789708,1.0940613,1.146878,1.6071383,3.169005,4.3347464,4.8138695,4.3422914,2.6710186,2.3767538,2.9841464,3.942393,4.5460134,3.9461658,2.2409391,4.115934,6.617184,7.6395655,5.926794,5.20245,5.2628117,5.5759397,5.5759397,4.678055,5.4363527,5.873977,5.9117036,5.4740787,4.4705606,3.7952607,3.4066803,3.1576872,2.916239,2.546522,1.6335466,1.599593,1.7316349,1.4713237,0.43007925,0.331991,0.35462674,0.38480774,0.33953625,0.15467763,0.094315626,0.1056335,0.13204187,0.14713238,0.15845025,0.15467763,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08677038,0.071679875,0.033953626,0.011317875,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.06413463,0.0452715,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.018863125,0.056589376,0.1056335,0.09808825,0.049044125,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.003772625,0.0,0.003772625,0.0,0.011317875,0.011317875,0.00754525,0.0,0.003772625,0.003772625,0.003772625,0.0,0.003772625,0.02263575,0.033953626,0.033953626,0.03772625,0.060362,0.116951376,0.124496624,0.124496624,0.16976812,0.19994913,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.14713238,0.19994913,0.18485862,0.19240387,0.38858038,0.43007925,0.271629,0.116951376,0.0452715,0.0150905,0.0150905,0.02263575,0.02263575,0.018863125,0.02263575,0.02263575,0.0150905,0.00754525,0.011317875,0.02263575,0.02263575,0.049044125,0.094315626,0.1358145,0.09808825,0.060362,0.03772625,0.030181,0.06413463,0.18863125,0.29803738,0.5772116,1.1921495,1.8334957,1.750498,1.9240388,2.4522061,3.9763467,5.7192993,5.5193505,4.8100967,3.9763467,2.916239,2.0673985,2.3956168,2.4371157,2.2296214,2.1051247,2.0296721,1.599593,1.5958204,1.5958204,1.2902378,0.7092535,0.23390275,0.116951376,0.08677038,0.08299775,0.11317875,0.271629,0.44139713,0.5470306,0.5470306,0.47535074,0.4376245,0.3772625,0.32067314,0.271629,0.24522063,0.241448,0.21503963,0.20372175,0.2263575,0.2867195,0.38858038,0.38858038,0.36594462,0.3470815,0.38103512,0.5319401,0.9808825,1.5430037,2.1013522,2.5125682,2.637065,3.470815,4.979865,6.72659,7.356619,4.6214657,4.2027044,3.8480775,3.5538127,3.802806,5.564622,6.507778,6.696409,6.2323766,5.828706,6.8246784,8.171506,9.042982,10.427535,12.457208,14.377474,12.849561,11.310329,10.876478,12.291212,15.894069,13.098554,9.793735,7.1264887,6.439871,9.25425,10.401127,9.97482,9.231613,9.21275,10.718028,15.316857,17.467255,17.889788,17.452164,17.184307,18.429274,20.153362,21.130472,20.428764,17.425755,16.094019,14.607604,13.343775,12.608112,12.630749,15.8676605,16.67123,16.248695,15.99593,17.508753,18.715992,19.685556,20.398582,21.130472,22.46221,22.862108,21.892544,20.14959,17.96524,15.437581,13.58145,13.505998,14.452927,15.965749,17.87847,19.455427,22.515026,25.623669,27.5213,27.128946,27.423212,26.578144,24.012758,19.915688,15.256495,13.52486,13.717264,14.354838,14.494425,13.743673,10.759526,9.337247,8.518587,7.779153,7.0057645,5.8136153,5.100589,4.8402777,4.938366,5.2250857,5.0515447,4.927048,4.696918,4.3309736,3.953711,3.9008942,3.8405323,3.8065786,3.7763977,3.6934,3.006782,2.686109,2.505023,2.335255,2.1390784,1.8561316,1.6222287,1.448688,1.3204187,1.2034674,1.0072908,0.8941121,0.87147635,0.935611,1.0450171,1.2336484,1.2336484,1.0827434,0.84884065,0.6375736,0.5093044,0.42630664,0.43007925,0.47912338,0.46026024,0.33576363,0.32444575,0.331991,0.31312788,0.24899325,0.17354076,0.181086,0.1961765,0.18485862,0.17354076,0.15845025,0.14713238,0.13204187,0.124496624,0.14335975,0.19240387,0.25276586,0.32444575,0.42630664,0.60362,0.995973,1.8448136,2.7917426,3.572676,4.0103,3.9461658,3.731126,3.2369123,2.7653341,3.0746894,4.074435,4.1083884,4.1008434,4.323428,4.4139714,4.244203,4.1272516,3.5500402,2.6031113,1.9730829,1.9051756,1.9127209,1.6524098,1.146878,0.754525,0.63002837,0.56212115,0.6828451,0.91674787,0.9922004,0.95824677,1.146878,1.2411937,1.1431054,0.9620194,0.6790725,0.44139713,0.754525,1.5882751,2.372981,2.7426984,2.625747,3.1199608,4.1989317,4.715781,4.255521,3.2859564,2.5087957,2.3390274,2.9124665,3.6896272,4.1762958,4.7044635,5.3759904,6.0512905,6.8850408,7.854605,8.68081,9.405154,10.38981,11.170743,11.604594,12.019584,12.219532,11.472552,10.718028,10.412445,10.567122,10.880251,10.733118,10.314357,9.808825,8.431817,6.8397694,7.1076255,7.6848373,7.8734684,7.488661,6.617184,5.6061206,5.0779533,4.881777,4.5950575,4.1498876,3.8254418,3.5500402,3.3236825,3.059599,2.7200627,2.3428001,2.1315331,1.9693103,1.8825399,1.8561316,1.7995421,14.68683,15.399856,14.577423,12.5326605,10.121953,8.744945,9.307066,11.155652,12.245941,11.653639,9.548513,7.062354,4.644101,2.6672459,1.6033657,1.991946,3.1463692,3.7084904,3.92353,3.8292143,3.270866,4.0593443,5.0025005,4.738417,3.2746384,1.9957186,0.8941121,0.42630664,0.28294688,0.241448,0.17354076,0.15467763,0.14335975,0.116951376,0.07922512,0.06790725,0.06413463,0.06413463,0.060362,0.049044125,0.03772625,0.03772625,0.03772625,0.033953626,0.03772625,0.03772625,0.03772625,0.030181,0.02263575,0.02263575,0.02263575,0.0150905,0.0150905,0.02263575,0.03772625,0.06790725,0.1056335,0.181086,0.25276586,0.29803738,0.32444575,0.60362,1.5052774,2.957738,4.2819295,4.191386,3.9574835,3.9989824,3.8103511,3.3764994,3.180323,3.3350005,3.893349,4.8666863,6.0324273,6.9491754,6.349328,6.145606,6.990674,8.416726,8.835487,9.948412,10.789707,10.812344,10.050273,9.125979,9.590013,11.351829,13.328684,14.664193,14.7170105,14.317112,12.917468,10.657665,8.484633,8.179051,7.4584794,6.9982195,6.820906,6.8171334,6.741681,7.6018395,8.186596,8.371455,8.3525915,8.650629,6.9152217,6.356873,6.7680893,7.201941,5.96452,5.4476705,5.353355,5.4212623,5.243949,4.266839,3.4594972,2.8256962,2.5201135,2.4672968,2.335255,2.0447628,1.9164935,1.9542197,2.0183544,1.8221779,1.3996439,1.2298758,1.3468271,1.6939086,2.11267,2.9086938,3.187868,3.0331905,2.897376,3.5802212,2.746471,1.9353566,1.3656902,1.3694628,2.3805263,3.2331395,4.0517993,4.61392,4.7006907,4.0970707,3.783943,3.1954134,2.3616633,1.5430037,1.2298758,1.2525115,1.0676528,0.73566186,0.41121614,0.33953625,0.6073926,1.2525115,2.0673985,2.6446102,2.372981,2.0145817,2.1088974,2.7540162,3.9989824,5.873977,6.4738245,6.149379,5.3609,4.7421894,5.1043615,5.1835866,4.3121104,2.8219235,1.2298758,0.24899325,0.452715,0.56589377,0.62625575,0.7582976,1.1581959,1.6976813,2.5427492,3.2369123,3.2557755,1.9881734,1.8221779,1.8221779,2.1315331,2.4861598,2.2183034,1.6071383,3.1237335,4.8968673,5.594803,4.429062,5.1232247,5.0968165,4.8365054,4.8440504,5.6325293,6.138061,6.790725,6.911449,5.847569,2.9803739,2.806833,2.8294687,2.7917426,2.4597516,1.6260014,1.086516,1.1657411,1.3505998,1.2298758,0.49421388,1.1883769,1.2751472,0.995973,0.58098423,0.24899325,0.23390275,0.13204187,0.060362,0.049044125,0.056589376,0.09808825,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.060362,0.056589376,0.041498873,0.0,0.0,0.003772625,0.00754525,0.011317875,0.011317875,0.030181,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.011317875,0.0150905,0.011317875,0.00754525,0.0,0.0,0.003772625,0.003772625,0.003772625,0.02263575,0.041498873,0.049044125,0.071679875,0.120724,0.18485862,0.1961765,0.14713238,0.15845025,0.24899325,0.30181,0.44894236,0.21503963,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.00754525,0.0,0.0,0.02263575,0.056589376,0.12826926,0.30181,0.29803738,0.18863125,0.09808825,0.07922512,0.07922512,0.06413463,0.05281675,0.03772625,0.02263575,0.0150905,0.02263575,0.041498873,0.056589376,0.05281675,0.041498873,0.041498873,0.033953626,0.041498873,0.060362,0.060362,0.05281675,0.033953626,0.02263575,0.03772625,0.090543,0.1659955,0.41876137,0.9393836,1.5052774,1.5958204,1.4373702,1.7769064,3.0860074,4.7836885,5.247721,4.617693,3.640583,2.7125173,2.191895,2.3993895,2.2786655,1.9127209,1.720317,1.7316349,1.6222287,1.6976813,1.7919968,1.5241405,0.8941121,0.31312788,0.1659955,0.124496624,0.11317875,0.14335975,0.29426476,0.5357128,0.83752275,0.995973,0.97710985,0.91674787,0.7997965,0.6752999,0.5583485,0.45648763,0.35839936,0.23390275,0.18863125,0.19994913,0.26031113,0.3470815,0.35462674,0.3734899,0.3772625,0.3772625,0.41498876,0.56212115,0.8224323,1.3015556,1.9579924,2.6144292,3.9989824,4.6290107,5.13077,5.2364035,3.802806,3.7386713,3.4859054,3.2142766,3.2821836,4.244203,4.7912335,5.564622,5.6325293,5.036454,4.8100967,5.281675,6.4738245,7.907422,9.235386,10.220041,9.424017,8.526133,9.122208,11.653639,15.403628,14.260523,12.208215,9.103344,6.4549613,7.4094353,10.336992,10.906659,10.54826,9.955957,9.06939,10.042727,13.830443,16.524097,16.867407,16.263786,16.090246,17.271078,18.342503,18.146326,15.848798,14.418973,13.309821,13.389046,14.4114275,15.045229,16.218515,15.396083,14.535924,14.279386,13.970031,13.355092,15.588487,17.772837,18.908396,19.866644,19.24416,18.991394,18.614132,17.742655,16.11288,14.679284,14.290704,14.136025,14.43029,16.38451,18.402864,19.138527,19.65915,20.474035,21.541689,22.877197,23.390276,23.292187,22.669704,21.4851,21.130472,21.994404,21.575642,19.029121,15.135772,11.978085,10.442626,9.684328,9.178797,8.710991,8.197914,7.5603404,7.1076255,6.858632,6.549277,6.066381,5.6853456,5.3194013,4.991183,4.851596,5.0779533,5.1534057,5.2288585,5.2250857,4.817642,3.832987,3.2067313,2.8294687,2.5691576,2.2598023,1.8976303,1.6184561,1.4260522,1.2940104,1.177059,1.0638802,0.94692886,0.84884065,0.784706,0.77716076,0.9016574,1.0827434,1.2638294,1.3770081,1.3317367,1.2298758,0.9280658,0.9393836,1.2638294,1.3694628,0.94692886,0.60362,0.41876137,0.35839936,0.29426476,0.211267,0.19240387,0.181086,0.16976812,0.18485862,0.17354076,0.15467763,0.18863125,0.26408374,0.32821837,0.33953625,0.3055826,0.3055826,0.3734899,0.48666862,0.8563859,1.659955,2.6672459,3.6330378,4.304565,4.3913355,4.2894745,3.5990841,2.625747,2.3692086,3.1539145,3.6707642,4.0480266,4.2102494,3.8707132,3.229367,3.0860074,3.0218725,2.837014,2.5502944,2.1051247,1.599593,1.1506506,0.8337501,0.7205714,0.7507524,0.8111144,0.94692886,1.116697,1.1883769,1.1959221,1.4260522,1.6561824,1.6637276,1.2110126,0.8903395,1.0186088,1.7467253,2.686109,2.9313297,2.625747,2.757789,3.5274043,4.636556,5.2967653,5.1043615,4.3309736,3.482133,2.9954643,3.2029586,3.6179473,3.832987,4.2592936,5.0175915,5.9494295,6.881268,7.884786,8.8618965,9.80128,10.763299,11.638548,12.58925,13.773854,14.694374,14.200161,12.679792,10.770844,9.484379,8.956212,8.424272,8.213005,7.7602897,6.647365,5.349582,5.2552667,5.723072,5.987156,5.8890676,5.458988,4.9232755,4.5007415,4.266839,3.9461658,3.5085413,3.138824,2.8709676,2.6597006,2.4484336,2.2183034,1.991946,1.8334957,1.7278622,1.6863633,1.6788181,1.6486372,17.780382,15.90916,14.335975,12.777881,11.193378,9.774872,8.914713,8.899622,8.850578,8.156415,6.462507,4.6742826,3.1161883,1.841041,1.0487897,1.0601076,1.2110126,1.5015048,1.8900851,2.1692593,1.9655377,2.938875,3.4745877,2.9954643,1.8259505,1.1959221,0.70170826,0.3961256,0.2565385,0.2263575,0.181086,0.1358145,0.10940613,0.08299775,0.056589376,0.056589376,0.06413463,0.071679875,0.06790725,0.05281675,0.030181,0.049044125,0.049044125,0.03772625,0.026408374,0.030181,0.033953626,0.02263575,0.018863125,0.0150905,0.0150905,0.0150905,0.0150905,0.018863125,0.026408374,0.041498873,0.056589376,0.090543,0.14335975,0.20749438,0.27540162,0.31312788,0.88279426,1.9164935,3.0369632,3.5839937,3.7273536,3.8141239,3.6254926,3.2482302,3.0520537,3.150142,3.7235808,4.6214657,5.6363015,6.5341864,5.541986,5.1835866,5.726845,6.647365,6.643593,7.798016,8.726082,9.231613,9.265567,8.937348,8.356364,8.080963,8.582722,9.884277,11.563096,12.223305,11.631002,9.952185,8.058327,7.5075235,6.8473144,6.387054,6.387054,6.779407,7.1793056,8.741172,10.453944,11.917723,12.698656,12.332711,10.137043,8.695901,8.371455,8.416726,7.0057645,5.764571,5.1534057,4.8968673,4.6931453,4.22534,4.036709,3.7348988,3.429316,3.1539145,2.897376,2.5993385,2.3088465,2.1088974,2.033445,2.0485353,1.6146835,1.4147344,1.3996439,1.478869,1.5316857,2.1202152,2.323937,2.2220762,2.214531,3.0369632,2.2862108,1.4637785,0.9242931,0.97710985,1.8749946,2.6785638,3.5538127,4.2291126,4.3121104,3.289729,3.5085413,3.3915899,3.0105548,2.41448,1.6373192,1.5543215,1.4411428,1.2411937,0.97710985,0.7582976,1.0638802,1.7014539,2.3956168,2.8030603,2.5201135,2.1768045,2.3428001,2.957738,4.014073,5.5268955,5.847569,5.3684454,4.6290107,4.2328854,4.8629136,5.462761,5.100589,3.9574835,2.2899833,0.41121614,0.2263575,0.2678564,0.40367088,0.5319401,0.5885295,0.94692886,1.5203679,2.0673985,2.252257,1.6373192,1.8184053,1.6863633,1.6750455,1.8372684,1.841041,1.8938577,2.4107075,3.048281,3.5500402,3.7575345,5.0741806,5.0062733,4.402653,4.123479,5.05909,5.5495315,6.1116524,6.1606965,5.1081343,2.3654358,2.4069347,2.5616124,2.5427492,2.1805773,1.4260522,1.2525115,1.1883769,1.1053791,0.98842776,0.94692886,1.5882751,1.4939595,1.0336993,0.55080324,0.35462674,0.2867195,0.150905,0.08299775,0.08677038,0.049044125,0.094315626,0.071679875,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.0754525,0.03772625,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.00754525,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0150905,0.0452715,0.056589376,0.08677038,0.15467763,0.2678564,0.33576363,0.271629,0.18863125,0.18863125,0.33953625,0.5470306,0.331991,0.090543,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.011317875,0.011317875,0.0,0.030181,0.094315626,0.16976812,0.23390275,0.26408374,0.1961765,0.14713238,0.116951376,0.1056335,0.10940613,0.1056335,0.1056335,0.10940613,0.1056335,0.056589376,0.041498873,0.0754525,0.10940613,0.11317875,0.09808825,0.094315626,0.090543,0.10940613,0.15845025,0.23013012,0.15467763,0.08677038,0.06413463,0.071679875,0.049044125,0.07922512,0.271629,0.62248313,1.0148361,1.2411937,1.0676528,1.20724,1.931584,3.127506,4.2819295,4.236658,3.6254926,2.927557,2.4974778,2.5691576,2.1390784,1.6524098,1.4298248,1.5165952,1.7165444,1.7542707,1.8334957,1.690136,1.2110126,0.4376245,0.25276586,0.21881226,0.24899325,0.29426476,0.3772625,0.5357128,0.80356914,0.995973,1.056335,1.0638802,0.97333723,0.87147635,0.784706,0.7167987,0.6451189,0.49421388,0.3961256,0.35085413,0.33576363,0.33576363,0.28294688,0.29049212,0.32444575,0.36971724,0.4376245,0.47535074,0.5357128,0.7809334,1.3128735,2.1994405,3.1463692,3.0822346,2.9464202,3.0218725,2.9464202,3.0256453,2.8785129,2.71629,2.7992878,3.4444065,3.3878171,3.92353,4.1612053,3.9273026,3.7537618,4.1574326,4.7610526,5.05909,4.983638,4.8855495,5.824933,6.156924,6.911449,8.616675,11.276376,12.185578,11.785681,9.450426,6.217286,4.7836885,10.997202,13.890805,14.053028,12.30253,9.669238,7.4396167,10.106862,13.309821,14.8339615,14.6151495,13.675766,13.902123,14.479335,14.68683,13.88326,13.830443,13.909668,14.603831,15.214996,13.856852,14.064346,13.302276,12.079946,10.929295,10.423763,9.009028,10.816116,13.140053,14.84528,16.380737,15.841252,16.38451,17.225805,17.693611,17.237123,17.003222,16.724047,15.920478,14.886778,14.652876,15.275358,15.030138,14.916959,15.46399,16.724047,18.565088,20.145817,21.779364,23.352549,24.314568,25.038912,25.865116,24.910643,21.790682,17.614386,14.796235,13.068373,12.132762,11.69891,11.495189,11.257513,10.570895,9.869187,9.231613,8.386545,7.454707,6.677546,6.1229706,5.8626595,5.9796104,6.515323,6.983129,7.183078,6.907676,5.9305663,4.617693,3.712263,3.1350515,2.7426984,2.3277097,1.9353566,1.6448646,1.4373702,1.2751472,1.1053791,1.0789708,1.0148361,0.91297525,0.7997965,0.73566186,0.7432071,0.91674787,1.20724,1.5052774,1.6373192,1.569412,1.4562333,1.6712729,2.093807,2.0975795,1.5241405,1.0035182,0.65643674,0.49044126,0.392353,0.32444575,0.2867195,0.2565385,0.241448,0.24899325,0.20749438,0.17731337,0.23013012,0.35085413,0.43007925,0.392353,0.30181,0.26408374,0.31312788,0.41121614,0.7507524,1.5015048,2.5578396,3.7613072,4.919503,4.930821,4.5309224,3.6669915,2.6332922,2.0862615,2.3805263,2.8445592,3.2821836,3.5462675,3.5274043,2.9803739,2.686109,2.7728794,3.0369632,2.9351022,2.354118,1.7693611,1.297783,1.026154,1.0487897,1.3128735,1.5015048,1.5203679,1.3807807,1.2223305,1.3053282,1.569412,1.7957695,1.8070874,1.4675511,1.2940104,1.5920477,2.263575,2.9200118,2.8936033,2.2711203,2.252257,2.8106055,3.7348988,4.6026025,4.7572803,4.5422406,3.9197574,3.2218218,3.1727777,3.4330888,3.6745367,4.1310244,4.90064,5.934339,6.8058157,7.858378,9.001483,10.152134,11.246195,12.064855,12.717519,13.736128,14.898096,15.245177,13.585222,11.197151,9.235386,8.084735,7.4018903,7.0849895,6.3153744,5.3458095,4.4931965,4.1310244,4.2404304,4.2781568,4.187614,3.99521,3.7801702,3.4934506,3.2444575,2.9615107,2.625747,2.2786655,2.0485353,1.871222,1.7316349,1.6260014,1.5543215,1.4637785,1.4071891,1.3845534,1.3807807,1.3807807,21.737865,17.165443,14.818871,14.11339,13.8719425,12.344029,9.740918,7.7376537,6.300284,5.2288585,4.1762958,3.229367,2.5729303,2.1013522,1.7316349,1.3996439,1.0751982,1.116697,1.2449663,1.3241913,1.3694628,1.539231,1.3543724,1.1393328,1.0299267,0.965792,0.66775465,0.41498876,0.2565385,0.18863125,0.1961765,0.1358145,0.08299775,0.049044125,0.03772625,0.0452715,0.071679875,0.08299775,0.08299775,0.06790725,0.026408374,0.0452715,0.0452715,0.033953626,0.02263575,0.030181,0.02263575,0.011317875,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.018863125,0.018863125,0.026408374,0.041498873,0.08299775,0.1659955,0.2867195,0.31312788,0.8639311,1.5656394,2.1654868,2.4974778,2.2560298,2.3277097,2.384299,2.2673476,1.9844007,1.9957186,2.6672459,3.8141239,5.172269,6.3832817,6.3153744,5.847569,5.43258,5.1345425,4.61392,4.82896,5.27413,6.1418333,7.3453007,8.544995,8.443134,7.1566696,6.2851934,6.692637,8.503497,8.899622,8.820397,8.4544525,7.8395147,6.858632,6.8359966,6.6850915,7.009537,8.050782,9.699419,11.200924,12.917468,14.441608,15.116908,14.045483,13.091009,10.54826,7.8734684,5.994701,5.2967653,4.4101987,3.904667,3.783943,4.044254,4.6931453,5.0779533,4.8025517,4.2291126,3.5990841,3.0181,3.0143273,2.8558772,2.5578396,2.214531,1.9844007,1.599593,1.418507,1.3128735,1.1581959,0.8526133,0.7130261,0.80734175,0.98465514,1.1695137,1.3656902,1.3430545,0.9922004,0.6451189,0.56212115,0.91674787,1.3204187,1.6675003,1.8749946,1.7844516,1.177059,2.033445,2.5012503,2.6710186,2.6106565,2.3428001,2.1277604,2.04099,1.9429018,1.6863633,1.1506506,1.4939595,2.1881225,2.8407867,3.1425967,2.8596497,2.3578906,2.565385,3.169005,3.9348478,4.6818275,4.4403796,3.9273026,3.470815,3.3915899,3.9612563,4.7044635,4.7346444,4.044254,2.6672459,0.6488915,0.3961256,0.422534,0.5394854,0.56212115,0.32821837,0.9808825,1.2034674,1.267602,1.3505998,1.5241405,1.6222287,1.6410918,1.750498,2.0145817,2.4107075,2.2107582,1.8749946,1.7580433,2.1654868,3.350091,3.802806,3.6368105,3.2859564,3.187868,3.7914882,4.093298,4.2592936,4.2064767,3.7952607,2.8445592,2.5880208,2.4182527,2.1202152,1.7693611,1.750498,2.1541688,1.9730829,1.4411428,1.0487897,1.5656394,1.1959221,0.80734175,0.48666862,0.30935526,0.34330887,0.18863125,0.13204187,0.150905,0.17731337,0.09808825,0.12826926,0.11317875,0.071679875,0.030181,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.00754525,0.0,0.003772625,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0452715,0.060362,0.0754525,0.124496624,0.23767537,0.3470815,0.31312788,0.19994913,0.10186087,0.14713238,0.26408374,0.3055826,0.20372175,0.033953626,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.06413463,0.18863125,0.31312788,0.38858038,0.3772625,0.30181,0.22258487,0.15845025,0.11317875,0.1056335,0.13958712,0.18863125,0.2565385,0.30181,0.21881226,0.13204187,0.12826926,0.13958712,0.14335975,0.14713238,0.1358145,0.14713238,0.19994913,0.30181,0.44139713,0.29049212,0.150905,0.116951376,0.15845025,0.116951376,0.10186087,0.20749438,0.46026024,0.76584285,0.94315624,0.84884065,0.87902164,1.1393328,1.7655885,2.9124665,3.6594462,3.7084904,3.1916409,2.5917933,2.7389257,2.1654868,1.7127718,1.5618668,1.6976813,1.8900851,1.7995421,1.7089992,1.6260014,1.3732355,0.5583485,0.33953625,0.31312788,0.3961256,0.4979865,0.543258,0.5319401,0.543258,0.5998474,0.69793564,0.784706,0.7469798,0.7092535,0.69793564,0.7167987,0.7507524,0.65643674,0.55457586,0.5017591,0.47912338,0.4074435,0.2678564,0.2263575,0.26031113,0.35085413,0.47535074,0.58098423,0.65643674,0.7507524,1.0148361,1.6637276,1.6448646,1.7165444,2.173032,2.7653341,2.7125173,2.5993385,2.5540671,2.493705,2.6710186,3.6330378,3.229367,2.4899325,2.0975795,2.214531,2.5012503,3.0935526,3.2935016,2.8407867,2.0447628,1.7995421,3.983892,5.3194013,5.342037,4.9232755,6.2436943,7.9489207,8.314865,7.383027,5.4438977,3.0407357,10.469034,15.562078,16.493916,13.973803,11.276376,8.661947,7.6848373,8.75249,10.850069,11.521597,10.910432,10.552032,10.714255,11.302785,11.830952,14.400109,15.577168,15.7657995,14.464244,10.253995,10.842525,12.442118,12.215759,10.295494,9.763554,8.431817,8.854351,10.555805,12.894833,15.052773,15.762027,16.550507,17.248442,17.682293,17.663431,18.51227,18.908396,18.71222,17.497435,14.543469,12.404391,12.608112,13.622949,14.64533,15.596032,17.693611,19.968504,22.303759,24.310795,25.333178,26.32915,26.740366,26.215971,24.729557,22.571615,19.987368,17.969013,16.573141,15.682802,15.01882,14.222796,13.419228,12.536433,11.465008,10.065364,8.7600355,7.779153,7.2283497,7.1302614,7.435844,8.13378,8.831716,8.888305,8.062099,6.507778,5.0138187,4.055572,3.4142256,2.9086938,2.3993895,1.9768555,1.6788181,1.4600059,1.267602,1.0299267,1.0223814,0.95824677,0.87147635,0.7884786,0.754525,0.7130261,0.7469798,0.8865669,1.1091517,1.3355093,1.388326,1.750498,2.2069857,2.5125682,2.3956168,1.9504471,1.5882751,1.2751472,0.98842776,0.72811663,0.543258,0.46026024,0.41876137,0.38858038,0.35839936,0.2565385,0.2263575,0.27540162,0.38480774,0.47157812,0.38103512,0.27540162,0.241448,0.29803738,0.43007925,0.7054809,1.3694628,2.3654358,3.6481283,5.198677,4.8742313,4.134797,3.3463185,2.7238352,2.293756,2.3126192,2.4069347,2.7087448,3.2520027,3.9310753,3.9688015,3.429316,3.0256453,2.9237845,2.7125173,2.3578906,2.082489,1.7278622,1.3694628,1.3015556,1.690136,1.8825399,1.7165444,1.2902378,0.9620194,1.3015556,1.6561824,1.7429527,1.5731846,1.4675511,1.4071891,1.6260014,1.9391292,2.203213,2.3277097,1.9768555,1.6825907,1.7769064,2.3805263,3.4029078,4.112161,4.3913355,4.0103,3.2935016,3.1463692,3.3840446,3.772625,4.3083377,4.991183,5.828706,6.4474163,7.4773426,8.59404,9.759781,11.204697,11.978085,11.800771,11.664956,12.030901,12.811834,11.8045435,10.612394,9.495697,8.597813,7.91874,7.2660756,6.119198,4.9685473,4.085753,3.519859,3.2859564,3.0746894,2.8747404,2.6634734,2.4371157,2.2296214,2.0447628,1.8485862,1.6335466,1.4147344,1.267602,1.1506506,1.0789708,1.0487897,1.0487897,1.0299267,0.995973,0.9620194,0.935611,0.935611,25.069094,18.964987,14.347293,13.053283,14.030393,13.321139,10.891568,8.43559,6.809588,5.847569,4.3347464,3.308592,2.9313297,3.2369123,3.7801702,3.6481283,2.546522,1.9542197,1.7882242,1.8938577,2.0296721,2.1013522,1.780679,1.4600059,1.2713746,1.1129243,0.88279426,0.5319401,0.2867195,0.20749438,0.18485862,0.16976812,0.13204187,0.08677038,0.056589376,0.0452715,0.071679875,0.11317875,0.11317875,0.06413463,0.0150905,0.0150905,0.02263575,0.03772625,0.041498873,0.030181,0.030181,0.030181,0.02263575,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.030181,0.030181,0.041498873,0.05281675,0.07922512,0.150905,0.2867195,0.68661773,1.0336993,1.2261031,1.3732355,1.4449154,1.6863633,1.6222287,1.2864652,1.1883769,1.7391801,2.6182017,3.863168,5.492942,7.5075235,9.899368,9.235386,7.8961043,6.8473144,5.613666,3.663219,2.8256962,3.270866,4.8100967,6.8963585,8.68081,8.465771,8.182823,8.616675,9.382519,9.797507,9.114662,8.360137,7.9941926,7.91874,8.345046,8.13378,8.333729,9.224068,10.284176,10.321902,9.461743,9.027891,9.5032425,10.529396,11.812089,10.79348,8.537451,5.9796104,3.9688015,4.6629643,4.478106,4.0593443,3.742444,3.5689032,4.5233774,4.979865,4.9760923,4.5912848,3.983892,3.712263,3.591539,3.2067313,2.4710693,1.6184561,1.3015556,1.0638802,0.9507015,0.91297525,0.83752275,0.4979865,0.6413463,0.86770374,0.9620194,0.9016574,0.9016574,0.7092535,0.48666862,0.34330887,0.3055826,0.42630664,0.44894236,0.5281675,0.72811663,1.0072908,0.55457586,0.6451189,1.0601076,1.6222287,2.1956677,2.0862615,1.8033148,1.4449154,1.0902886,0.80734175,1.4071891,2.463524,3.361409,3.712263,3.3727267,2.4672968,2.335255,2.5616124,2.8521044,3.0218725,2.5087957,2.372981,2.565385,3.0445085,3.7537618,3.9008942,3.6707642,3.0445085,2.0296721,0.68661773,0.68661773,0.48666862,0.26031113,0.14713238,0.24522063,0.67152727,0.77716076,0.8639311,1.0601076,1.327964,1.388326,1.5580941,1.8033148,2.082489,2.3503454,1.690136,1.2336484,1.1657411,1.4449154,1.7995421,1.9579924,2.293756,2.7125173,3.1425967,3.5085413,3.410453,2.8106055,2.052308,1.4901869,1.4637785,1.4524606,1.5128226,1.6222287,2.1654868,3.9348478,3.802806,2.9803739,1.8749946,1.2864652,2.3956168,1.5165952,0.95824677,0.6451189,0.452715,0.18485862,0.09808825,0.06790725,0.03772625,0.0,0.0,0.0,0.0,0.071679875,0.150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030181,0.150905,0.030181,0.0,0.0,0.003772625,0.0150905,0.003772625,0.0,0.0,0.003772625,0.0150905,0.026408374,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.026408374,0.049044125,0.07922512,0.116951376,0.150905,0.1659955,0.15845025,0.150905,0.15845025,0.18485862,0.27917424,0.35839936,0.3169005,0.17354076,0.0754525,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.10186087,0.181086,0.27917424,0.42630664,0.52439487,0.30181,0.120724,0.1056335,0.1659955,0.23013012,0.33576363,0.49421388,0.633801,0.6111652,0.41498876,0.27540162,0.1659955,0.09808825,0.120724,0.120724,0.0754525,0.071679875,0.1358145,0.26031113,0.271629,0.14713238,0.12826926,0.23767537,0.27540162,0.24899325,0.32821837,0.5470306,0.79602385,0.80734175,0.68661773,0.58475685,0.6451189,1.056335,2.0447628,3.1425967,3.4368613,3.150142,2.655928,2.4710693,2.5201135,2.0560806,1.7995421,1.9127209,1.9994912,1.901403,1.6373192,1.2789198,0.8865669,0.5357128,0.31312788,0.22258487,0.29049212,0.45648763,0.58098423,0.56589377,0.49044126,0.4678055,0.49044126,0.44139713,0.34330887,0.26408374,0.23390275,0.23767537,0.21503963,0.17731337,0.18485862,0.35839936,0.58098423,0.52062225,0.3470815,0.35085413,0.39989826,0.452715,0.55080324,0.73188925,0.79602385,0.8224323,0.95447415,1.418507,1.9579924,2.0372176,2.0975795,2.2371666,2.2107582,2.335255,2.5578396,2.4408884,2.1579416,2.4861598,3.5839937,2.9464202,2.2183034,2.0108092,1.8749946,1.8146327,1.9579924,1.8599042,1.6788181,2.1654868,3.3161373,3.8480775,3.8556228,3.6669915,3.874486,5.7079816,6.56814,6.255012,5.070408,3.7990334,3.470815,7.462252,11.208468,12.619431,12.068627,10.578441,7.443389,6.2889657,7.9791017,10.604849,10.627484,10.186088,9.593785,9.574923,11.246195,14.517061,12.955194,11.7026825,12.083718,11.59705,9.216523,12.989148,17.191853,18.323639,15.07541,11.876224,12.396846,13.536179,14.237886,15.456445,17.384256,18.289686,18.02183,16.87118,15.565851,15.173498,15.030138,14.735873,14.053028,12.894833,11.185833,11.378237,12.721292,14.864142,17.867151,21.798227,25.069094,27.687294,29.603788,30.716713,32.131447,33.591454,34.22148,33.632954,31.93527,29.309525,26.925224,24.337204,21.439827,18.463226,16.618414,15.856343,14.984866,13.445636,11.321648,9.869187,8.993938,8.60913,8.714764,9.397609,10.20495,9.948412,8.918486,7.4509344,5.934339,4.8629136,4.191386,3.6669915,3.1312788,2.5314314,2.082489,1.8485862,1.659955,1.4109617,1.0676528,0.935611,0.77338815,0.68661773,0.694163,0.7167987,0.65643674,0.6488915,0.66775465,0.7469798,0.9922004,1.5052774,1.8334957,2.0673985,2.2975287,2.6408374,2.4672968,2.4823873,2.474842,2.2409391,1.5580941,0.935611,0.694163,0.59230214,0.49044126,0.38103512,0.32067314,0.34330887,0.43385187,0.56589377,0.70170826,0.543258,0.392353,0.331991,0.38103512,0.5017591,0.69793564,1.1053791,1.780679,2.8030603,4.255521,4.1612053,3.942393,3.6481283,3.259548,2.686109,2.7841973,2.7992878,3.006782,3.4179983,3.783943,5.0553174,4.6290107,3.5500402,2.6031113,2.335255,2.505023,2.4559789,2.0598533,1.3996439,0.77716076,0.66775465,0.60362,0.62248313,0.72811663,0.9016574,1.4373702,1.8561316,1.9844007,1.8221779,1.5430037,1.2864652,1.4034165,1.6486372,1.8523588,1.9391292,1.841041,2.0258996,2.2107582,2.3880715,2.8521044,4.3422914,4.8327327,4.8025517,4.5761943,4.3196554,4.085753,4.13857,4.425289,4.8629136,5.342037,5.80607,6.590776,7.6395655,8.82417,9.933322,10.091772,9.673011,8.858124,7.964011,7.4773426,7.7716074,8.216777,8.627994,8.7600355,8.345046,7.564113,6.307829,4.8327327,3.5047686,2.8219235,2.5314314,2.293756,2.0598533,1.8146327,1.5731846,1.3656902,1.1921495,1.0450171,0.9242931,0.83752275,0.754525,0.68661773,0.6375736,0.6111652,0.6111652,0.6111652,0.573439,0.52062225,0.45648763,0.3961256,26.657368,20.368402,15.211224,12.113899,11.159425,11.563096,10.080454,8.322411,6.752999,5.723072,5.4703064,4.561104,4.0517993,4.123479,4.617693,5.0515447,4.98741,4.3649273,3.2105038,1.8938577,1.1506506,1.3392819,1.7542707,2.2296214,2.3088465,1.2110126,0.65643674,0.31312788,0.14713238,0.11317875,0.14713238,0.18485862,0.18485862,0.14335975,0.07922512,0.0452715,0.060362,0.094315626,0.10940613,0.090543,0.05281675,0.033953626,0.02263575,0.02263575,0.033953626,0.030181,0.02263575,0.011317875,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.00754525,0.018863125,0.018863125,0.026408374,0.0452715,0.06790725,0.1056335,0.15845025,0.27540162,0.35085413,0.3734899,0.422534,0.7884786,1.3920987,1.6675003,1.5354583,1.3958713,1.6146835,2.214531,3.4444065,4.908185,5.5683947,6.9227667,8.650629,9.344792,8.318638,5.59103,3.6292653,3.8443048,4.768598,5.4476705,5.455216,5.764571,6.8963585,6.903904,5.764571,5.379763,5.696664,6.255012,7.3000293,8.262049,7.748972,6.368191,5.221313,5.247721,6.5455046,8.379,10.427535,12.581704,12.743927,10.93684,9.307066,8.60913,8.729855,9.224068,9.4127,8.375228,6.541732,5.036454,3.8556228,3.138824,3.1916409,4.123479,4.3649273,4.1310244,3.7160356,3.5047686,3.6594462,3.3350005,2.8181508,2.3692086,2.2296214,2.5238862,1.6825907,0.91297525,0.6790725,0.7054809,0.80356914,0.72811663,0.63002837,0.58475685,0.5696664,0.66020936,0.5093044,0.33576363,0.23013012,0.1961765,0.23013012,0.30181,0.45648763,0.6828451,0.935611,0.9997456,1.116697,1.3392819,1.6939086,2.161714,2.6936543,2.0975795,1.3996439,1.1393328,1.3468271,2.2371666,3.006782,3.5538127,3.7801702,3.6028569,2.7087448,2.6144292,2.625747,2.4333432,2.1051247,2.3654358,3.410453,4.22534,4.304565,3.6556737,3.1954134,2.384299,1.5128226,0.7582976,0.19994913,0.21881226,0.18863125,0.150905,0.124496624,0.1358145,0.24899325,0.29803738,0.38103512,0.5394854,0.77716076,1.0751982,1.4713237,1.8863125,2.1164427,1.8485862,1.8523588,1.5543215,1.267602,1.1581959,1.237421,1.3091009,1.2902378,1.3053282,1.4524606,1.7882242,1.5543215,1.3656902,1.2449663,1.1657411,1.0751982,1.6561824,1.7429527,1.5128226,1.3694628,1.9579924,1.9504471,1.5656394,0.98842776,0.51684964,0.56589377,0.32067314,0.19240387,0.12826926,0.090543,0.03772625,0.018863125,0.0150905,0.16222288,0.31312788,0.0,0.0,0.0,0.0150905,0.033953626,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.060362,0.07922512,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.030181,0.00754525,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.00754525,0.041498873,0.060362,0.10186087,0.08299775,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.018863125,0.02263575,0.033953626,0.049044125,0.06790725,0.060362,0.071679875,0.09808825,0.1358145,0.16976812,0.18863125,0.19240387,0.16976812,0.15845025,0.23390275,0.44894236,0.23013012,0.033953626,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.060362,0.124496624,0.18485862,0.20372175,0.120724,0.049044125,0.041498873,0.094315626,0.14713238,0.29426476,0.67152727,1.2826926,1.9881734,2.282438,1.6863633,0.9205205,0.392353,0.16976812,0.14335975,0.10940613,0.094315626,0.10186087,0.1358145,0.13958712,0.1358145,0.2263575,0.422534,0.663982,0.44516975,0.5772116,0.7432071,0.7394345,0.4678055,0.43385187,0.3961256,0.41121614,0.5583485,0.9205205,2.022127,2.3956168,2.3277097,2.0900342,1.9466745,1.9844007,1.931584,2.0900342,2.595566,3.4029078,2.757789,2.1088974,1.5052774,1.0110635,0.7167987,0.36971724,0.1961765,0.1961765,0.33953625,0.56589377,0.52439487,0.47912338,0.45648763,0.452715,0.44139713,0.38480774,0.34330887,0.31312788,0.27917424,0.2263575,0.15845025,0.124496624,0.14335975,0.19240387,0.18863125,0.31312788,0.3961256,0.41498876,0.3961256,0.42630664,0.47535074,0.5696664,0.724344,0.91674787,1.0902886,1.2638294,1.4222796,1.6222287,1.7618159,1.5882751,1.9164935,2.0975795,1.9466745,1.6712729,1.8636768,2.2107582,2.2484846,2.2862108,2.263575,1.7316349,1.4750963,1.4335974,1.5279131,1.6976813,1.9240388,2.474842,2.9992368,3.4896781,3.85185,3.9122121,4.8063245,5.7683434,6.7567716,6.809588,4.055572,2.9464202,4.214022,7.145352,9.797507,8.993938,7.5829763,6.221059,6.2097406,8.035691,11.374464,11.52537,9.876732,7.854605,6.48137,6.387054,9.465516,12.781653,15.011275,15.203679,12.781653,9.861642,9.246704,10.552032,12.528888,13.060828,12.344029,12.098808,13.060828,14.743419,15.456445,16.293968,16.893814,16.51278,15.39231,14.758509,14.388792,14.071891,14.252977,14.928277,15.652621,15.916705,16.018566,15.999702,16.21097,17.320122,19.598787,22.515026,25.585943,28.490864,31.093975,33.693314,36.194565,37.258446,36.786865,35.9418,34.847736,33.77631,32.086174,29.64906,26.838455,24.1448,21.915178,19.21398,15.999702,13.151371,11.310329,10.336992,10.167224,10.469034,10.646348,10.238904,9.0957985,7.907422,6.9227667,5.9494295,5.1571784,4.870459,4.689373,4.346064,3.7160356,2.886058,2.2711203,1.8636768,1.5845025,1.3015556,1.0374719,0.88279426,0.8337501,0.8639311,0.8865669,0.8262049,0.7997965,0.8865669,1.1091517,1.4298248,1.8372684,2.0447628,2.4220252,2.9615107,3.2746384,2.6332922,2.6106565,2.6446102,2.4295704,1.9089483,1.1808317,0.784706,0.5885295,0.4979865,0.4678055,0.45648763,0.5017591,0.5998474,0.7167987,0.8111144,0.73188925,0.62248313,0.5772116,0.633801,0.784706,1.0487897,1.3694628,1.9089483,2.7351532,3.8065786,4.402653,4.2781568,3.9122121,3.5387223,3.150142,3.0633714,3.4783602,4.032936,4.432834,4.45547,4.3686996,4.1762958,3.772625,3.1727777,2.505023,3.0369632,3.138824,2.8634224,2.2862108,1.4864142,1.3958713,1.5618668,1.7429527,1.780679,1.6222287,1.8938577,1.9466745,1.8561316,1.7127718,1.6260014,1.3317367,1.2223305,1.2223305,1.2940104,1.448688,1.6335466,2.0900342,2.6295197,3.1652324,3.7084904,4.5422406,5.0477724,5.323174,5.323174,4.8327327,4.5196047,4.4931965,4.6856003,4.9685473,5.168496,5.300538,5.5570765,5.956975,6.5228686,7.273621,7.61693,7.5829763,7.183078,6.4926877,5.6325293,5.1345425,5.0553174,5.3646727,5.938112,6.587003,5.8966126,4.8365054,3.6556737,2.637065,2.0900342,1.7693611,1.4713237,1.177059,0.9016574,0.7054809,0.58475685,0.5017591,0.44516975,0.40367088,0.38858038,0.38103512,0.44894236,0.6073926,0.7130261,0.48666862,0.34330887,0.25276586,0.19994913,0.15845025,0.116951376,20.168453,16.682549,13.162688,10.246449,8.495952,8.394091,8.865668,8.461998,7.3981175,6.1305156,5.349582,4.821415,4.478106,4.247976,4.0895257,4.0103,4.191386,3.9273026,3.097325,1.9806281,1.2525115,1.8221779,2.4182527,2.9011486,2.9539654,2.0673985,0.8978847,0.41498876,0.24522063,0.17354076,0.120724,0.1659955,0.17354076,0.14335975,0.094315626,0.071679875,0.07922512,0.08299775,0.08299775,0.071679875,0.033953626,0.02263575,0.011317875,0.00754525,0.0150905,0.02263575,0.0150905,0.011317875,0.00754525,0.00754525,0.00754525,0.00754525,0.003772625,0.003772625,0.00754525,0.00754525,0.0150905,0.018863125,0.033953626,0.060362,0.090543,0.09808825,0.120724,0.14713238,0.17354076,0.21881226,0.41121614,0.724344,0.94692886,1.0110635,1.0110635,1.9655377,3.097325,4.395108,5.4363527,5.402399,5.8702044,7.092535,8.111144,7.937603,5.5495315,5.0175915,5.745708,6.56814,6.9755836,7.1302614,6.043745,5.4288073,4.8063245,4.38379,5.0741806,6.7831798,8.763808,10.665211,11.317875,8.741172,6.820906,5.379763,4.821415,5.6815734,8.601585,10.687846,11.932813,11.3971,9.424017,7.647111,6.145606,5.4665337,6.3719635,8.084735,8.284684,6.983129,5.5495315,4.5950575,4.0895257,3.361409,3.500996,4.0706625,4.036709,3.308592,2.7389257,2.584248,2.4786146,2.6182017,2.8407867,2.637065,2.2899833,1.4600059,0.79602385,0.5319401,0.47157812,0.5319401,0.482896,0.41876137,0.38480774,0.3772625,0.422534,0.3734899,0.29426476,0.23390275,0.20372175,0.1961765,0.20372175,0.33576363,0.58098423,0.79602385,0.8903395,0.8262049,0.965792,1.4034165,1.9693103,2.6332922,2.5993385,2.2975287,2.003264,1.8297231,1.9051756,2.565385,3.2557755,3.651901,3.6330378,2.8106055,2.6144292,2.584248,2.5389767,2.5917933,3.4029078,4.187614,4.5233774,4.214022,3.31991,2.4522061,1.4977322,0.77716076,0.41876137,0.36971724,0.18863125,0.20372175,0.2565385,0.271629,0.25276586,0.49421388,0.5055317,0.47912338,0.51684964,0.62248313,0.814887,1.1355602,1.5052774,1.7919968,1.8146327,1.5769572,1.2411937,0.98465514,0.9393836,1.20724,0.9205205,0.77716076,0.814887,1.086516,1.6788181,1.2940104,1.2336484,1.3166461,1.327964,1.0035182,1.6335466,1.8033148,1.6222287,1.2600567,0.9507015,0.83752275,0.70170826,0.5470306,0.36971724,0.14335975,0.07922512,0.07922512,0.10940613,0.124496624,0.06413463,0.21881226,0.3055826,0.36594462,0.33576363,0.056589376,0.09808825,0.14335975,0.09808825,0.003772625,0.0150905,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.049044125,0.060362,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.026408374,0.049044125,0.041498873,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.026408374,0.0452715,0.071679875,0.03772625,0.03772625,0.060362,0.10186087,0.15845025,0.1358145,0.12826926,0.124496624,0.12826926,0.14713238,0.3169005,0.24522063,0.14713238,0.094315626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.049044125,0.049044125,0.03772625,0.02263575,0.018863125,0.041498873,0.10940613,0.20749438,0.43385187,0.88279426,1.6486372,2.3578906,2.3126192,1.6637276,0.8299775,0.513077,0.38103512,0.2867195,0.20749438,0.15467763,0.150905,0.17354076,0.20749438,0.27540162,0.38858038,0.543258,0.43007925,0.44516975,0.4640329,0.41876137,0.32821837,0.4376245,0.5583485,0.6111652,0.663982,0.91674787,1.6410918,2.0560806,2.2183034,2.2371666,2.263575,2.1390784,1.9655377,2.3013012,3.1237335,3.8254418,3.3538637,2.505023,1.7731338,1.3128735,0.9280658,0.5357128,0.331991,0.29803738,0.392353,0.5470306,0.56212115,0.5583485,0.5394854,0.5281675,0.543258,0.56212115,0.5885295,0.6111652,0.59607476,0.52062225,0.38103512,0.23767537,0.13958712,0.10186087,0.1056335,0.20749438,0.271629,0.29049212,0.28294688,0.2867195,0.3055826,0.35085413,0.5281675,0.7809334,0.87147635,0.72811663,0.76584285,0.90543,1.0186088,0.9205205,0.94692886,1.1091517,1.2713746,1.4411428,1.7919968,2.0447628,2.082489,2.1013522,2.0862615,1.7957695,1.4071891,1.3807807,1.6184561,2.0070364,2.3918443,2.7087448,3.169005,3.6707642,4.06689,4.187614,4.606375,4.8855495,5.4665337,5.938112,5.0175915,2.9916916,2.727608,4.244203,6.549277,7.6282477,5.9230213,5.515578,5.8702044,6.537959,7.152897,7.492433,7.1868505,6.730363,6.198423,5.2628117,6.175787,8.729855,11.302785,12.823153,12.766563,10.740664,9.224068,9.129752,10.831206,14.158662,12.449662,11.23865,11.355601,12.815607,14.815099,14.713238,14.735873,14.720782,14.656648,14.68683,14.581196,14.999957,16.244923,18.116146,19.911915,20.406128,19.934551,18.749947,17.206944,15.754482,15.878979,16.991903,18.685812,20.719257,23.02433,25.204908,26.962952,27.642023,27.46471,27.540163,28.275824,29.071848,29.317068,28.645542,26.936543,24.623924,22.149082,19.323385,16.4411,14.27184,12.913695,12.166716,11.902632,11.736636,11.046246,9.835234,8.416726,7.333983,6.6624556,6.0248823,5.5457587,5.270357,4.90064,4.3083377,3.519859,2.7313805,2.1541688,1.7580433,1.478869,1.2487389,1.0487897,0.9507015,0.9318384,0.97333723,1.0412445,1.0751982,1.1317875,1.2751472,1.5203679,1.8259505,2.1466236,2.3277097,2.5767028,2.9237845,3.259548,3.0822346,2.8143783,2.5804756,2.323937,1.7882242,1.0450171,0.7167987,0.6073926,0.5885295,0.6073926,0.63002837,0.6828451,0.77716076,0.8865669,0.9507015,0.90920264,0.87902164,0.8978847,0.9808825,1.1016065,1.2298758,1.3732355,1.7655885,2.4672968,3.3727267,4.112161,4.0593443,3.7613072,3.440634,2.9803739,2.5238862,2.7841973,3.5236318,4.4101987,5.0062733,4.696918,4.2592936,3.6971724,3.029418,2.282438,2.4371157,2.516341,2.5087957,2.3767538,2.082489,2.1164427,2.0636258,1.9127209,1.6825907,1.4147344,1.5128226,1.5618668,1.5618668,1.5165952,1.4298248,1.2411937,1.086516,1.0072908,1.0638802,1.3468271,1.8599042,2.5691576,3.3274553,4.0291634,4.636556,4.6554193,4.568649,4.5535583,4.61392,4.5912848,4.8402777,4.7912335,4.5912848,4.406426,4.432834,4.3121104,4.2328854,4.2328854,4.3800178,4.776143,5.0854983,5.304311,5.402399,5.383536,5.27413,4.5837393,4.1083884,3.9763467,4.217795,4.7308717,4.1536603,3.3161373,2.41448,1.6410918,1.1921495,0.90920264,0.6790725,0.48666862,0.33576363,0.23013012,0.17731337,0.15467763,0.14335975,0.1358145,0.12826926,0.13204187,0.17354076,0.2565385,0.31312788,0.19994913,0.120724,0.07922512,0.05281675,0.033953626,0.018863125,13.140053,11.800771,9.884277,8.013056,6.7869525,6.7831798,7.877241,7.888559,7.4169807,6.647365,5.349582,4.715781,4.304565,3.92353,3.5236318,3.218049,3.4368613,3.6707642,3.9461658,4.172523,4.168751,4.2328854,3.7537618,3.3048196,2.9615107,2.3314822,1.0978339,0.4979865,0.2565385,0.16976812,0.08299775,0.1056335,0.1056335,0.10186087,0.094315626,0.08677038,0.07922512,0.06790725,0.05281675,0.041498873,0.0150905,0.011317875,0.003772625,0.011317875,0.026408374,0.041498873,0.041498873,0.026408374,0.0150905,0.0150905,0.02263575,0.0150905,0.011317875,0.011317875,0.011317875,0.0,0.00754525,0.011317875,0.033953626,0.071679875,0.120724,0.094315626,0.08299775,0.09808825,0.13958712,0.1961765,0.26031113,0.38858038,0.58098423,0.8299775,1.1317875,2.8709676,4.214022,5.119452,5.4438977,4.949684,4.647874,5.149633,6.0022464,6.2625575,4.515832,5.3986263,6.2399216,6.749226,6.9944468,7.4282985,6.1229706,4.825187,4.2781568,4.9119577,6.862405,10.242677,12.396846,13.275867,13.124963,12.449662,9.812597,7.6584287,6.0550632,5.994701,9.386291,10.216269,10.099318,9.469289,8.744945,8.345046,6.888813,5.5570765,5.541986,6.779407,7.9753294,7.575431,6.4549613,5.5004873,4.6856003,3.0256453,2.4710693,2.9351022,3.127506,2.6936543,2.2258487,1.991946,2.0560806,2.3767538,2.655928,2.323937,1.720317,1.2298758,0.80356914,0.4640329,0.29803738,0.241448,0.241448,0.24899325,0.24899325,0.2565385,0.271629,0.29426476,0.30935526,0.3055826,0.29426476,0.271629,0.241448,0.29426476,0.44894236,0.6375736,0.7696155,0.7432071,0.9393836,1.4298248,1.9693103,2.463524,2.7200627,2.6672459,2.354118,1.9730829,1.690136,2.3126192,3.0407357,3.429316,3.3727267,2.674791,2.535204,2.6219745,2.8106055,3.2067313,4.085753,4.376245,4.244203,3.7914882,3.0709167,2.1503963,1.20724,0.58098423,0.362172,0.41121614,0.18863125,0.17731337,0.2678564,0.38103512,0.47912338,0.67152727,0.633801,0.56212115,0.55080324,0.5998474,0.694163,0.8903395,1.1129243,1.3128735,1.4562333,1.2638294,0.9997456,0.8262049,0.86770374,1.2449663,0.724344,0.633801,0.80356914,1.1431054,1.6184561,1.1393328,1.0186088,1.1091517,1.2449663,1.2600567,1.3468271,1.4034165,1.3807807,1.1581959,0.573439,0.5281675,0.47912338,0.38480774,0.24522063,0.120724,0.29426476,0.392353,0.3470815,0.20372175,0.10186087,0.29049212,0.38480774,0.33576363,0.1961765,0.1358145,0.11317875,0.14335975,0.09808825,0.0,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.0,0.003772625,0.011317875,0.018863125,0.02263575,0.018863125,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.018863125,0.02263575,0.02263575,0.02263575,0.026408374,0.02263575,0.026408374,0.03772625,0.060362,0.056589376,0.071679875,0.0754525,0.06790725,0.1056335,0.090543,0.1056335,0.116951376,0.10186087,0.049044125,0.1056335,0.1659955,0.27917424,0.362172,0.19994913,0.060362,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.02263575,0.0452715,0.120724,0.13958712,0.17354076,0.40367088,1.116697,2.1881225,2.5729303,2.3654358,1.7882242,1.1959221,0.814887,0.6149379,0.47535074,0.36971724,0.3470815,0.3734899,0.482896,0.59230214,0.663982,0.70170826,0.6413463,0.48666862,0.35839936,0.31312788,0.35839936,0.42630664,0.56212115,0.67152727,0.80356914,1.1657411,1.7542707,2.082489,2.2447119,2.3503454,2.5314314,2.4786146,2.1390784,2.3088465,3.0369632,3.6368105,3.7047176,2.9728284,2.173032,1.6184561,1.1959221,0.6752999,0.4640329,0.4640329,0.59230214,0.7884786,0.8186596,0.7582976,0.67152727,0.6073926,0.6149379,0.663982,0.7167987,0.7696155,0.7884786,0.73566186,0.5583485,0.3772625,0.25276586,0.19994913,0.20372175,0.241448,0.2867195,0.32821837,0.362172,0.3734899,0.3772625,0.36594462,0.452715,0.59607476,0.6149379,0.4074435,0.35839936,0.4074435,0.482896,0.48666862,0.3734899,0.5055317,0.814887,1.2298758,1.6863633,2.0108092,2.0258996,1.8825399,1.720317,1.6712729,1.4637785,1.5618668,1.8334957,2.1956677,2.625747,2.9237845,3.361409,3.7688525,4.074435,4.2894745,4.4215164,4.2328854,4.2894745,4.61392,4.7006907,3.1312788,2.5578396,2.9501927,4.1612053,5.934339,4.979865,4.821415,5.062863,5.111907,4.191386,4.402653,4.983638,5.6551647,5.926794,5.119452,4.647874,5.3156285,7.073672,9.359882,11.106608,9.661693,8.303548,7.7225633,8.635539,11.781908,10.299266,9.288202,9.1976595,10.1294985,11.830952,11.6008215,11.861133,12.570387,13.411682,13.819125,14.283158,15.596032,17.440845,19.38752,20.89657,20.972023,20.232588,18.85558,17.067356,15.124454,14.388792,14.498198,15.184815,16.305285,17.803017,18.976303,19.68933,19.817598,19.557287,19.447882,20.323132,21.4851,22.454664,22.790428,22.096264,20.492899,18.580177,16.603323,14.852824,13.6833105,12.955194,12.479843,12.049765,11.431054,10.38981,9.058073,7.8810134,7.0585814,6.507778,5.885295,5.481624,4.9987283,4.349837,3.572676,2.8294687,2.293756,1.8863125,1.5807298,1.3543724,1.1732863,1.0902886,1.0902886,1.1657411,1.2713746,1.3468271,1.4675511,1.6146835,1.780679,1.961765,2.173032,2.5201135,2.7992878,2.9803739,3.1048703,3.259548,3.270866,2.897376,2.5201135,2.191895,1.629774,1.0676528,0.90543,0.875249,0.845068,0.8262049,0.8337501,0.8941121,0.995973,1.0940613,1.1091517,1.0525624,1.0450171,1.0714256,1.1242423,1.1808317,1.20724,1.237421,1.5203679,2.142851,3.029418,3.8820312,4.1989317,4.1536603,3.8405323,3.2670932,2.5804756,2.2862108,2.6031113,3.4368613,4.3724723,4.7535076,4.5497856,3.8971217,3.0105548,2.1843498,1.9466745,1.9164935,2.0636258,2.2862108,2.3880715,2.2748928,2.0447628,1.7769064,1.5203679,1.2864652,1.2487389,1.2789198,1.297783,1.2826926,1.237421,1.1619685,1.0601076,1.0223814,1.1242423,1.4373702,2.305074,3.1463692,3.8178966,4.274384,4.587512,4.5460134,4.561104,4.768598,5.0779533,5.1835866,5.2137675,4.7572803,4.115934,3.5651307,3.3764994,3.3425457,3.2029586,2.9954643,2.8332415,2.897376,3.2935016,3.8707132,4.402653,4.8327327,5.2552667,4.821415,4.1800685,3.6066296,3.2520027,3.1539145,2.6219745,1.9579924,1.3015556,0.77338815,0.47157812,0.29426476,0.17731337,0.10940613,0.071679875,0.041498873,0.02263575,0.02263575,0.026408374,0.026408374,0.018863125,0.018863125,0.018863125,0.018863125,0.018863125,0.018863125,0.011317875,0.00754525,0.003772625,0.0,0.0,9.87296,9.118435,7.805561,6.643593,6.1833324,6.8435416,7.2094865,6.8850408,6.934085,7.1604424,6.119198,4.8968673,4.0404816,3.482133,3.1916409,3.169005,3.5500402,4.3724723,5.9494295,7.960239,9.495697,8.424272,6.1116524,4.0216184,2.71629,1.8863125,1.0827434,0.452715,0.1358145,0.0754525,0.041498873,0.030181,0.026408374,0.041498873,0.06413463,0.06413463,0.05281675,0.03772625,0.030181,0.026408374,0.018863125,0.00754525,0.003772625,0.02263575,0.056589376,0.0754525,0.07922512,0.041498873,0.018863125,0.02263575,0.030181,0.018863125,0.0150905,0.0150905,0.011317875,0.003772625,0.003772625,0.011317875,0.041498873,0.094315626,0.1659955,0.13204187,0.090543,0.071679875,0.08299775,0.124496624,0.23390275,0.43007925,0.7884786,1.3807807,2.252257,4.2328854,4.9723196,4.949684,4.508287,3.8405323,3.2520027,3.7575345,4.5196047,4.745962,3.7198083,4.8930945,5.8664317,6.2323766,6.017337,5.6778007,4.9949555,4.7912335,5.0175915,5.873977,7.805561,11.446144,12.740154,12.249713,11.921495,15.082954,11.54046,9.439108,7.798016,7.1906233,9.733373,9.408927,8.884532,8.771353,9.337247,10.502988,9.627739,8.548768,7.5226145,7.1679873,8.465771,8.382772,7.4584794,6.1305156,4.5233774,2.4710693,1.7127718,1.5882751,1.7769064,2.04099,2.2183034,2.293756,2.3314822,2.2409391,1.9768555,1.5430037,1.3128735,1.1695137,0.8639311,0.44894236,0.26408374,0.17354076,0.14335975,0.13958712,0.15467763,0.181086,0.20749438,0.24899325,0.3055826,0.36594462,0.38858038,0.36971724,0.35462674,0.32821837,0.33953625,0.5017591,0.7884786,1.0450171,1.3430545,1.6976813,2.071171,2.3126192,2.263575,2.123988,1.9994912,1.931584,2.0070364,2.4069347,2.8181508,3.0218725,2.8596497,2.41448,2.5578396,2.886058,3.2255943,3.6481283,4.2064767,4.3121104,4.115934,3.7160356,3.1161883,2.3088465,1.3694628,0.65643674,0.29426476,0.16976812,0.120724,0.10940613,0.21881226,0.4376245,0.67152727,0.5357128,0.452715,0.44516975,0.513077,0.6149379,0.69793564,0.8224323,0.9205205,0.9507015,0.8978847,1.1204696,1.056335,0.95824677,0.9695646,1.1581959,0.6413463,0.66020936,0.87147635,1.0450171,1.086516,0.754525,0.60362,0.6451189,0.90543,1.4071891,0.8186596,0.6413463,0.76584285,0.875249,0.44516975,0.5885295,0.58475685,0.4074435,0.17354076,0.13958712,0.5093044,0.66020936,0.5055317,0.18485862,0.07922512,0.14713238,0.16222288,0.09808825,0.030181,0.15845025,0.030181,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.011317875,0.011317875,0.003772625,0.00754525,0.02263575,0.030181,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.03772625,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.018863125,0.026408374,0.026408374,0.026408374,0.041498873,0.041498873,0.030181,0.0150905,0.011317875,0.06413463,0.120724,0.11317875,0.049044125,0.026408374,0.049044125,0.0754525,0.090543,0.07922512,0.033953626,0.03772625,0.07922512,0.30935526,0.58475685,0.49044126,0.29426476,0.12826926,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.02263575,0.033953626,0.07922512,0.124496624,0.094315626,0.060362,0.20749438,0.8262049,1.9542197,2.3013012,2.474842,2.4522061,1.5882751,1.0336993,0.77716076,0.633801,0.5319401,0.5319401,0.59607476,0.8111144,0.9922004,1.0714256,1.0827434,0.98842776,0.7469798,0.5394854,0.452715,0.47157812,0.34330887,0.35085413,0.482896,0.7696155,1.2826926,1.9278114,2.0900342,2.1353056,2.3314822,2.8521044,2.9615107,2.4823873,2.2296214,2.5201135,3.187868,3.772625,3.4217708,2.6144292,1.81086,1.478869,0.8563859,0.58098423,0.56589377,0.7507524,1.0789708,1.0978339,0.995973,0.8262049,0.66775465,0.633801,0.6413463,0.6526641,0.66775465,0.6828451,0.6752999,0.5319401,0.42630664,0.36971724,0.35839936,0.38103512,0.41876137,0.46026024,0.51684964,0.5696664,0.5885295,0.573439,0.5470306,0.52062225,0.48666862,0.41876137,0.33953625,0.29049212,0.29803738,0.35462674,0.42630664,0.4979865,0.56212115,0.7092535,0.9620194,1.3053282,1.6184561,1.7354075,1.5845025,1.3317367,1.358145,1.5505489,1.8485862,2.1164427,2.3126192,2.4974778,2.7502437,3.127506,3.4670424,3.7386713,4.0178456,4.002755,3.8707132,3.8669407,3.8669407,3.3953626,3.3048196,3.1124156,2.969056,3.0897799,3.7386713,4.1310244,4.0291634,4.1612053,4.52715,4.3800178,4.187614,4.327201,4.6629643,4.930821,4.749735,4.395108,4.2328854,5.0779533,6.809588,8.371455,6.9793563,5.836251,5.3344917,5.624984,6.598321,7.0359454,7.115171,7.413208,7.8696957,7.779153,8.050782,9.020347,10.178542,11.136789,11.619685,12.596795,14.264296,15.875206,16.984358,17.421982,17.240896,16.784409,16.165699,15.558306,15.214996,15.147089,15.592259,16.305285,17.123945,17.96524,18.331184,18.636768,18.693357,18.35382,17.512526,17.154125,17.184307,17.335213,17.346529,16.969267,15.777118,14.532151,13.449409,12.630749,12.076173,11.69891,11.336739,10.79348,10.054046,9.242931,8.29223,7.54525,6.9567204,6.379509,5.564622,4.9459114,4.214022,3.451952,2.7804246,2.3578906,2.0183544,1.7127718,1.4939595,1.358145,1.2600567,1.2449663,1.3317367,1.5128226,1.7089992,1.780679,1.9466745,2.1390784,2.3088465,2.4333432,2.5389767,2.9426475,3.361409,3.610402,3.610402,3.3953626,3.0935526,2.7841973,2.4522061,2.0598533,1.5656394,1.3053282,1.2713746,1.237421,1.146878,1.0789708,1.056335,1.1204696,1.2185578,1.2751472,1.2110126,1.1280149,1.0978339,1.086516,1.0827434,1.1016065,1.1393328,1.1657411,1.388326,1.9202662,2.795515,3.7952607,4.5309224,4.708236,4.3385186,3.7386713,3.1048703,2.3578906,2.0183544,2.2975287,3.1199608,4.3649273,4.7836885,4.3724723,3.4330888,2.546522,2.11267,2.003264,2.1768045,2.444661,2.5012503,2.0636258,1.8070874,1.6712729,1.5618668,1.3505998,1.2525115,1.2110126,1.1657411,1.1280149,1.1732863,1.1317875,1.0751982,1.086516,1.2147852,1.4939595,2.5502944,3.399135,3.821669,3.8971217,4.0103,4.6327834,5.3194013,6.092789,6.620957,6.2323766,5.372218,4.3686996,3.4934506,2.8634224,2.4371157,2.5540671,2.4522061,2.1843498,1.8863125,1.7693611,2.3465726,3.3425457,4.112161,4.4705606,4.6856003,4.5837393,3.9801195,3.218049,2.5087957,1.9504471,1.418507,0.9016574,0.482896,0.20372175,0.08677038,0.03772625,0.011317875,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,11.457462,11.544232,10.1294985,8.039464,6.247467,5.8437963,6.3945994,6.9869013,7.54525,7.8508325,7.5829763,6.0701537,4.610148,3.2633207,2.293756,2.1805773,2.9011486,4.538468,7.009537,10.325675,14.588741,13.415455,10.201178,6.379509,3.229367,1.8599042,1.0186088,0.38858038,0.08677038,0.056589376,0.030181,0.018863125,0.00754525,0.00754525,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.030181,0.030181,0.030181,0.011317875,0.00754525,0.026408374,0.0754525,0.08677038,0.056589376,0.03772625,0.041498873,0.030181,0.018863125,0.0150905,0.00754525,0.003772625,0.0150905,0.0150905,0.0150905,0.041498873,0.090543,0.150905,0.17731337,0.1358145,0.1056335,0.11317875,0.1358145,0.19994913,0.241448,0.8941121,2.323937,4.2404304,5.7570257,5.2552667,4.168751,3.410453,3.3878171,3.7650797,4.2064767,4.8855495,5.7570257,6.5756855,6.187105,7.9941926,8.778898,7.4509344,5.0213637,4.044254,4.002755,4.063117,3.8895764,3.6330378,3.9008942,5.20245,6.9793563,8.22055,7.4773426,4.2781568,6.428553,8.771353,9.307066,9.186342,9.955957,9.322156,8.439363,8.254503,9.537196,9.461743,8.986393,8.3525915,7.7942433,7.537705,7.9526935,7.5716586,6.368191,4.7044635,3.3274553,2.7540162,2.463524,2.335255,2.3654358,2.6710186,2.8030603,2.8294687,2.7389257,2.3503454,1.3128735,0.94692886,0.77338815,0.6187105,0.44516975,0.33576363,0.23767537,0.1659955,0.15467763,0.181086,0.1659955,0.1659955,0.17731337,0.21881226,0.29049212,0.35085413,0.35085413,0.34330887,0.33576363,0.35462674,0.42630664,0.694163,1.1393328,1.3505998,1.388326,1.7542707,1.8749946,1.4147344,1.3656902,1.8825399,2.2748928,2.4069347,1.991946,1.8636768,2.1503963,2.2748928,2.335255,2.8332415,3.470815,4.063117,4.561104,4.878004,4.98741,4.8025517,4.3121104,3.5538127,2.505023,1.4826416,0.7205714,0.29426476,0.120724,0.20749438,0.31312788,0.4640329,0.62248313,0.67152727,0.32821837,0.25276586,0.36971724,0.58098423,0.76207024,0.7394345,0.7696155,0.8903395,1.0676528,1.1883769,1.1280149,1.1506506,1.20724,1.20724,1.0374719,0.5998474,0.6073926,0.62625575,0.55080324,0.6111652,0.9507015,1.1393328,1.1581959,0.9808825,0.56589377,0.11317875,0.0,0.32821837,0.69039035,0.150905,0.090543,0.27917424,0.6073926,0.8224323,0.52062225,0.31312788,0.1961765,0.14713238,0.116951376,0.030181,0.018863125,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.041498873,0.06413463,0.05281675,0.011317875,0.0,0.011317875,0.05281675,0.056589376,0.026408374,0.0150905,0.026408374,0.030181,0.02263575,0.02263575,0.0452715,0.071679875,0.056589376,0.0754525,0.18485862,0.44139713,0.88279426,0.543258,0.14713238,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.041498873,0.056589376,0.041498873,0.030181,0.018863125,0.0150905,0.0150905,0.033953626,0.1056335,0.46026024,0.73188925,0.8903395,0.8299775,0.36594462,0.23013012,0.124496624,0.08677038,0.13958712,0.27540162,0.55457586,0.77338815,0.80356914,0.7167987,0.77716076,0.83752275,0.754525,0.5696664,0.422534,0.5357128,0.3734899,0.3169005,0.422534,0.7432071,1.3430545,1.5505489,1.6373192,1.9391292,2.7426984,4.3196554,4.025391,3.0746894,2.41448,2.4031622,2.806833,3.440634,3.500996,2.7992878,1.81086,1.6637276,1.3317367,0.7922512,0.482896,0.51684964,0.68661773,0.88279426,1.0676528,1.026154,0.7922512,0.67152727,0.6111652,0.52062225,0.4376245,0.36971724,0.32067314,0.29426476,0.30935526,0.362172,0.44139713,0.5017591,0.5394854,0.5394854,0.52062225,0.5017591,0.5017591,0.51684964,0.52062225,0.56212115,0.62625575,0.62625575,0.5281675,0.4678055,0.47157812,0.56212115,0.73188925,0.98842776,0.9620194,0.8262049,0.7205714,0.73188925,0.97710985,0.935611,0.9016574,1.0035182,1.237421,1.6637276,2.2183034,2.6710186,2.8634224,2.71629,2.5201135,2.5729303,2.7691069,3.0445085,3.3727267,3.531177,3.5990841,3.5990841,3.5877664,3.663219,3.904667,3.6556737,3.259548,2.9313297,2.7615614,2.7728794,3.4179983,4.1310244,4.696918,5.2326307,4.8063245,4.478106,4.398881,4.504514,4.515832,4.45547,4.3309736,4.3121104,4.745962,6.149379,5.587258,5.172269,5.2099953,5.7419353,6.560595,6.85486,6.983129,6.8850408,6.730363,6.911449,7.303802,7.647111,7.865923,8.069645,8.544995,9.22784,10.023865,10.887795,11.638548,11.917723,12.1252165,12.261031,12.528888,13.004238,13.626721,14.418973,15.396083,16.275105,16.905132,17.255987,17.610613,18.523588,19.647831,20.549488,20.723028,20.353312,19.83269,19.217752,18.48209,17.516298,16.11288,14.64533,13.392818,12.464753,11.793225,11.427281,10.861387,10.287949,9.718282,8.986393,8.231868,7.5565677,6.934085,6.270103,5.4174895,4.429062,3.6028569,2.9954643,2.6521554,2.6408374,2.1013522,1.750498,1.5769572,1.5543215,1.6033657,1.5769572,1.6260014,1.750498,1.9240388,2.1202152,2.3163917,2.5125682,2.7389257,2.9539654,3.0520537,3.259548,3.742444,3.9612563,3.7348988,3.2331395,2.8558772,2.516341,2.11267,1.6863633,1.418507,1.3468271,1.2449663,1.1883769,1.1996948,1.237421,1.2713746,1.3468271,1.3656902,1.2864652,1.1129243,1.0902886,1.1091517,1.1544232,1.2110126,1.297783,1.3807807,1.4600059,1.6373192,2.003264,2.625747,3.429316,3.8254418,3.731126,3.2746384,2.7615614,2.4333432,2.1843498,2.1353056,2.4710693,3.4481792,4.5120597,4.7572803,4.538468,4.08198,3.5085413,2.7653341,2.7992878,3.0407357,3.1124156,2.806833,2.4295704,2.033445,1.6410918,1.2525115,0.8224323,0.8865669,1.0299267,1.1695137,1.2336484,1.1581959,1.0487897,0.91297525,0.814887,0.87147635,1.237421,1.931584,2.8030603,3.270866,3.5953116,4.851596,5.8664317,6.2927384,6.511551,6.4134626,5.402399,4.6214657,3.8480775,3.2331395,2.7540162,2.2447119,1.7429527,1.3694628,1.1581959,1.1091517,1.2223305,1.659955,2.8143783,3.4896781,3.3538637,2.916239,2.6446102,2.1202152,1.6260014,1.2525115,0.9016574,0.4979865,0.23013012,0.07922512,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,13.619176,14.358611,13.705947,11.747954,9.159933,7.224577,6.5228686,6.5341864,6.670001,6.7869525,7.194396,7.748972,5.9003854,3.731126,2.3390274,1.841041,2.2371666,2.3201644,3.361409,5.6023483,8.239413,7.9753294,5.5457587,2.927557,1.2110126,0.6149379,0.33953625,0.15845025,0.06790725,0.041498873,0.00754525,0.003772625,0.00754525,0.00754525,0.003772625,0.003772625,0.02263575,0.03772625,0.041498873,0.033953626,0.00754525,0.00754525,0.011317875,0.018863125,0.033953626,0.05281675,0.05281675,0.056589376,0.056589376,0.049044125,0.018863125,0.026408374,0.018863125,0.0150905,0.011317875,0.0150905,0.0150905,0.02263575,0.03772625,0.06790725,0.13958712,0.18485862,0.19240387,0.181086,0.18863125,0.271629,0.32444575,0.36971724,0.62625575,1.3015556,2.5804756,3.802806,4.4215164,4.0895257,3.2369123,3.1048703,3.8367596,5.1081343,5.836251,5.994701,6.5756855,7.6508837,10.042727,10.684074,8.990166,6.862405,5.624984,5.696664,6.0814714,6.3455553,6.647365,7.1604424,8.194141,8.314865,7.0472636,4.878004,3.572676,4.7610526,6.375736,7.726336,9.480607,11.310329,11.548005,11.004747,10.306811,9.891823,10.295494,9.522105,8.778898,8.729855,9.476834,10.510533,10.038955,8.461998,6.187105,3.6556737,2.6898816,2.1881225,1.9693103,1.8636768,1.6675003,1.8523588,1.8599042,1.7052265,1.3732355,0.8224323,0.70170826,0.7205714,0.77716076,0.754525,0.52062225,0.35462674,0.2565385,0.23013012,0.241448,0.23013012,0.23767537,0.24899325,0.271629,0.30181,0.31312788,0.31312788,0.35462674,0.4678055,0.56212115,0.4376245,0.6488915,1.0186088,1.1732863,1.0827434,1.0601076,1.0525624,0.9997456,1.1921495,1.6109109,1.8825399,1.8900851,1.6184561,1.5015048,1.569412,1.4675511,1.6675003,2.6332922,3.5877664,4.236658,4.7572803,5.1156793,5.251494,4.9685473,4.266839,3.3840446,2.3654358,1.3355093,0.5998474,0.24899325,0.14713238,0.211267,0.24522063,0.35085413,0.5093044,0.58475685,0.331991,0.31312788,0.3772625,0.45648763,0.58098423,0.69039035,0.91674787,1.116697,1.1544232,0.8978847,0.8865669,0.7432071,0.573439,0.44139713,0.3772625,0.5357128,0.5696664,0.59230214,0.7809334,1.3807807,0.44139713,0.2263575,0.23013012,0.1961765,0.11317875,0.02263575,0.0,0.1358145,0.27540162,0.030181,0.018863125,0.056589376,0.120724,0.1659955,0.1056335,0.06413463,0.03772625,0.030181,0.02263575,0.00754525,0.003772625,0.1056335,0.1056335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.030181,0.041498873,0.033953626,0.030181,0.018863125,0.003772625,0.0,0.003772625,0.018863125,0.05281675,0.116951376,0.211267,0.15467763,0.090543,0.03772625,0.0150905,0.00754525,0.06413463,0.071679875,0.06790725,0.06790725,0.10186087,0.2678564,0.2565385,0.14335975,0.02263575,0.02263575,0.003772625,0.00754525,0.030181,0.05281675,0.026408374,0.026408374,0.033953626,0.0452715,0.056589376,0.056589376,0.041498873,0.026408374,0.011317875,0.00754525,0.033953626,0.1056335,0.17354076,0.21503963,0.20372175,0.120724,0.0754525,0.033953626,0.02263575,0.0452715,0.090543,0.362172,0.7092535,0.8111144,0.7205714,0.8526133,0.9507015,0.91297525,0.7130261,0.4678055,0.41121614,0.41876137,0.4979865,0.62248313,0.875249,1.4637785,2.1013522,2.233394,2.4333432,2.9426475,3.6594462,3.6896272,2.7351532,1.9994912,2.0296721,2.7351532,4.217795,3.953711,3.0181,2.1277604,1.6524098,1.5052774,1.0412445,0.6790725,0.573439,0.6375736,0.77338815,0.9242931,1.026154,1.0638802,1.0374719,1.0336993,0.77716076,0.482896,0.29426476,0.28294688,0.3169005,0.38103512,0.4376245,0.46026024,0.44139713,0.392353,0.362172,0.34330887,0.331991,0.32067314,0.34330887,0.3772625,0.41876137,0.46026024,0.47912338,0.392353,0.331991,0.35839936,0.5281675,0.91674787,1.0638802,1.1431054,1.1996948,1.2638294,1.3543724,1.4524606,1.418507,1.4600059,1.6184561,1.7731338,1.8976303,2.0108092,2.173032,2.354118,2.4220252,2.4333432,2.3880715,2.3201644,2.3163917,2.5314314,2.9049213,3.3764994,3.8707132,4.244203,4.3083377,4.093298,3.7650797,3.6066296,3.6141748,3.482133,3.338773,3.4444065,3.682082,4.0404816,4.636556,5.05909,4.8138695,4.564876,4.5761943,4.6742826,4.8666863,4.821415,4.8025517,4.991183,5.4665337,5.753253,5.9230213,6.224831,6.696409,7.17176,6.8774953,7.073672,7.356619,7.5603404,7.7414265,7.91874,7.914967,7.7829256,7.6131573,7.54525,8.111144,8.677037,9.152389,9.405154,9.25425,9.416472,9.733373,10.148361,10.555805,10.804798,11.151879,11.61214,12.045992,12.310076,12.264804,12.464753,13.117417,14.177525,15.486626,16.780636,17.644567,18.331184,18.806536,19.021576,18.908396,18.206688,17.127718,15.833707,14.479335,13.223051,11.959221,10.801025,9.903141,9.280658,8.793989,8.209232,7.537705,6.6850915,5.7004366,4.7572803,4.236658,4.0216184,3.640583,3.0218725,2.493705,2.142851,1.9089483,1.7693611,1.7391801,1.8448136,1.9579924,2.0108092,2.1013522,2.2560298,2.463524,2.71629,2.9049213,3.1237335,3.4066803,3.6971724,3.8858037,4.025391,4.025391,3.8178966,3.3576362,2.6446102,2.082489,1.6788181,1.4222796,1.2713746,1.2185578,1.2411937,1.3204187,1.4524606,1.6260014,1.7618159,1.659955,1.4939595,1.358145,1.2864652,1.3770081,1.448688,1.5015048,1.5430037,1.5882751,1.7052265,1.9579924,2.3880715,2.987919,3.6971724,4.006528,4.29702,4.406426,4.1272516,3.2142766,2.9916916,2.8596497,3.1312788,3.85185,4.7912335,4.9760923,4.6516466,4.357382,4.2630663,4.168751,4.0895257,4.044254,3.8405323,3.4972234,3.270866,2.727608,2.1353056,1.6863633,1.4335974,1.3015556,1.2940104,1.2562841,1.0902886,0.86770374,0.8563859,0.8526133,0.8526133,0.9922004,1.3128735,1.750498,2.1013522,2.4786146,3.0445085,4.036709,5.7419353,6.647365,6.228604,5.6815734,5.3156285,4.534695,3.85185,3.1765501,2.516341,1.8825399,1.2902378,0.87902164,0.6828451,0.6451189,0.7432071,0.9997456,1.3996439,1.6750455,1.7127718,1.539231,1.3015556,1.1317875,0.8941121,0.66020936,0.45648763,0.27917424,0.13958712,0.056589376,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,13.264549,14.298248,14.003984,12.393073,10.220041,8.9788475,7.567886,6.511551,5.696664,5.27413,5.6476197,5.7192993,4.402653,2.9351022,2.022127,1.8297231,1.7278622,1.2487389,1.3845534,2.2409391,3.0105548,2.8558772,1.8485862,0.8903395,0.38480774,0.2678564,0.21503963,0.1056335,0.030181,0.0150905,0.0,0.0,0.003772625,0.003772625,0.0,0.00754525,0.026408374,0.030181,0.02263575,0.0150905,0.00754525,0.00754525,0.018863125,0.030181,0.041498873,0.0452715,0.05281675,0.060362,0.06790725,0.08299775,0.09808825,0.060362,0.033953626,0.02263575,0.0150905,0.0150905,0.030181,0.041498873,0.071679875,0.1358145,0.24899325,0.33953625,0.35085413,0.30935526,0.2565385,0.26031113,0.3169005,0.6073926,1.0978339,1.7014539,2.305074,3.1652324,3.9725742,4.266839,3.7348988,2.2107582,2.5389767,3.3463185,3.712263,3.5274043,3.482133,4.0216184,5.3344917,6.4247804,6.6020937,5.50426,5.383536,6.3229194,7.352846,8.00551,8.296002,9.031664,10.193633,9.061845,5.9909286,4.4101987,4.715781,6.0286546,6.56814,6.466279,7.756517,9.797507,10.646348,11.106608,11.41219,11.242422,10.846297,9.25425,7.9300575,7.5905213,8.224322,9.612649,8.963757,7.273621,5.240176,3.2633207,2.9049213,2.2862108,1.750498,1.4260522,1.2261031,1.50905,1.4977322,1.3355093,1.1204696,0.875249,0.66020936,0.6413463,0.694163,0.7054809,0.5470306,0.47157812,0.39989826,0.34330887,0.31312788,0.30935526,0.2678564,0.241448,0.23013012,0.23390275,0.24899325,0.24899325,0.29049212,0.36971724,0.44139713,0.3961256,0.46026024,0.6187105,0.7432071,0.7582976,0.6375736,0.63002837,0.69039035,0.83752275,1.056335,1.2638294,1.267602,1.1355602,1.0714256,1.1242423,1.146878,1.5769572,2.5578396,3.3953626,3.9650288,4.696918,5.281675,5.4401255,4.8930945,3.7914882,2.6898816,1.7429527,0.9808825,0.47535074,0.2263575,0.16222288,0.23013012,0.20749438,0.27540162,0.44139713,0.55457586,0.43385187,0.5772116,0.6526641,0.56589377,0.47912338,0.47157812,0.5583485,0.6488915,0.66775465,0.5772116,0.663982,0.6073926,0.5055317,0.4376245,0.452715,0.97710985,0.8526133,0.5696664,0.5394854,1.0940613,0.6451189,0.6187105,0.7054809,0.70170826,0.513077,0.10186087,0.0,0.05281675,0.116951376,0.06413463,0.011317875,0.0,0.03772625,0.09808825,0.12826926,0.026408374,0.0,0.033953626,0.08299775,0.090543,0.0754525,0.10186087,0.071679875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.026408374,0.02263575,0.011317875,0.003772625,0.0,0.0,0.00754525,0.018863125,0.030181,0.056589376,0.11317875,0.08299775,0.049044125,0.026408374,0.018863125,0.026408374,0.08299775,0.1056335,0.090543,0.0452715,0.0150905,0.0452715,0.08299775,0.124496624,0.14335975,0.08677038,0.018863125,0.003772625,0.0150905,0.030181,0.02263575,0.02263575,0.02263575,0.033953626,0.056589376,0.071679875,0.056589376,0.03772625,0.018863125,0.011317875,0.0150905,0.0150905,0.02263575,0.02263575,0.02263575,0.033953626,0.0150905,0.0150905,0.02263575,0.033953626,0.06413463,0.23013012,0.41121614,0.5394854,0.6526641,0.91674787,0.90920264,0.8563859,0.73188925,0.5696664,0.47157812,0.513077,0.5772116,0.6790725,0.8978847,1.358145,2.1088974,2.516341,2.8445592,3.199186,3.5387223,3.350091,2.565385,1.7957695,1.6071383,2.516341,5.323174,6.1606965,4.8063245,2.4786146,1.81086,1.4600059,1.0601076,0.7922512,0.70170826,0.7167987,0.7809334,0.8526133,0.87147635,0.86770374,0.965792,0.9997456,0.814887,0.543258,0.32067314,0.29426476,0.362172,0.4678055,0.573439,0.6451189,0.6451189,0.543258,0.43385187,0.35085413,0.30935526,0.32067314,0.38858038,0.41876137,0.42630664,0.41876137,0.4074435,0.3734899,0.34330887,0.35839936,0.44894236,0.6413463,0.69039035,0.8865669,1.1544232,1.4675511,1.841041,2.354118,2.384299,2.2899833,2.2598023,2.282438,2.4333432,2.282438,2.1088974,2.0862615,2.2598023,2.4597516,2.6785638,2.8106055,2.7653341,2.4559789,2.655928,3.0256453,3.470815,3.8405323,3.9310753,3.682082,3.4481792,3.3651814,3.4029078,3.361409,3.4330888,3.561358,3.6971724,3.9008942,4.357382,4.7572803,4.847823,5.0515447,5.4174895,5.613666,5.847569,5.9720654,6.115425,6.3153744,6.5228686,6.722818,6.771862,6.8774953,7.1076255,7.3981175,7.2358947,7.164215,7.277394,7.5301595,7.756517,7.9753294,8.09228,7.9791017,7.7112455,7.5792036,7.937603,8.465771,8.967529,9.250477,9.103344,8.699674,9.061845,9.457971,9.552286,9.386291,9.193887,9.224068,9.337247,9.4127,9.322156,9.144843,9.386291,9.97482,10.819888,11.793225,12.642066,13.396591,14.060574,14.626467,15.0905,15.24895,14.928277,14.252977,13.340002,12.31762,11.272603,10.272858,9.382519,8.631766,7.9828744,7.2924843,6.5455046,5.7381625,4.98741,4.5196047,4.3083377,4.146115,3.742444,3.108643,2.565385,2.3201644,2.161714,2.033445,1.9429018,1.961765,2.1013522,2.2409391,2.3578906,2.5087957,2.8407867,3.1539145,3.3463185,3.4972234,3.682082,3.9801195,4.1197066,4.014073,3.8367596,3.6179473,3.240685,2.7200627,2.3163917,2.003264,1.7618159,1.5731846,1.4750963,1.5505489,1.6863633,1.8070874,1.8900851,1.8787673,1.7542707,1.6410918,1.5958204,1.6222287,1.7278622,1.8033148,1.8863125,1.9806281,2.0749438,2.1466236,2.5012503,2.938875,3.3463185,3.6745367,4.1574326,4.3724723,4.3309736,3.983892,3.2331395,2.8709676,2.8785129,3.308592,4.036709,4.7610526,4.315883,3.893349,3.7650797,3.9159849,4.0480266,4.2517486,4.2328854,3.9310753,3.5085413,3.3123648,2.757789,2.1353056,1.6184561,1.358145,1.4637785,1.3166461,1.0412445,0.76207024,0.58098423,0.56589377,0.62248313,0.7167987,0.9016574,1.1280149,1.2713746,1.4449154,1.7919968,2.584248,3.7575345,4.930821,5.4288073,5.13077,4.6554193,4.164978,3.3463185,2.4974778,2.022127,1.569412,1.0487897,0.6149379,0.41498876,0.45648763,0.543258,0.633801,0.845068,1.2940104,1.1506506,0.84884065,0.60362,0.43385187,0.33953625,0.26408374,0.19240387,0.116951376,0.049044125,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,12.419481,13.70972,13.6682205,12.626976,11.32542,10.917976,9.175024,7.2170315,5.59103,4.6554193,4.587512,3.953711,3.108643,2.354118,1.9164935,1.9391292,1.4826416,0.9507015,0.69039035,0.6526641,0.41498876,0.25276586,0.124496624,0.09808825,0.15845025,0.23013012,0.1961765,0.08677038,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.02263575,0.018863125,0.018863125,0.041498873,0.041498873,0.033953626,0.03772625,0.0452715,0.0452715,0.05281675,0.06413463,0.0754525,0.09808825,0.116951376,0.06413463,0.033953626,0.02263575,0.02263575,0.026408374,0.03772625,0.049044125,0.08677038,0.16222288,0.27917424,0.39989826,0.41121614,0.35462674,0.27917424,0.23013012,0.29426476,0.60362,1.1053791,1.6825907,2.1654868,2.9954643,3.7386713,4.395108,4.5950575,3.572676,3.270866,3.1916409,2.987919,2.6182017,2.3767538,1.7014539,1.8184053,2.8181508,3.953711,3.6179473,4.025391,5.0477724,6.2663302,7.515069,8.8769865,9.87296,10.846297,9.857869,7.1868505,5.3269467,5.6853456,6.730363,6.8246784,6.066381,6.2927384,7.7716074,8.926031,9.688101,10.291721,11.291467,11.185833,9.654147,7.835742,6.6662283,6.888813,8.07719,7.3188925,5.666483,3.9159849,2.595566,2.4522061,2.1051247,1.690136,1.3656902,1.2940104,1.6260014,1.4864142,1.2110126,0.98465514,0.8337501,0.6073926,0.56212115,0.59230214,0.6111652,0.5696664,0.55457586,0.482896,0.3961256,0.331991,0.32067314,0.34330887,0.29049212,0.21881226,0.18485862,0.20749438,0.23013012,0.2678564,0.3055826,0.331991,0.35462674,0.35462674,0.38103512,0.4678055,0.58475685,0.6187105,0.55457586,0.5394854,0.59607476,0.8186596,1.3656902,1.2487389,0.94315624,0.7696155,0.90920264,1.3656902,1.9693103,2.6823363,3.2369123,3.6745367,4.353609,5.0515447,5.451443,4.8327327,3.3764994,2.1541688,1.2789198,0.66775465,0.3169005,0.16976812,0.13204187,0.18863125,0.19994913,0.28294688,0.4376245,0.52062225,0.38103512,0.5470306,0.6526641,0.5885295,0.47157812,0.36971724,0.44139713,0.4979865,0.4640329,0.392353,0.41498876,0.5055317,0.5772116,0.60362,0.6111652,1.2185578,1.1431054,0.7997965,0.55457586,0.73566186,0.6790725,0.754525,0.8563859,0.8601585,0.62248313,0.124496624,0.0,0.049044125,0.116951376,0.1056335,0.02263575,0.0,0.07922512,0.1961765,0.18485862,0.056589376,0.011317875,0.08677038,0.22258487,0.24899325,0.19240387,0.094315626,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.011317875,0.026408374,0.03772625,0.03772625,0.0452715,0.030181,0.02263575,0.018863125,0.018863125,0.033953626,0.07922512,0.1358145,0.17731337,0.19994913,0.211267,0.16976812,0.10940613,0.120724,0.17731337,0.15845025,0.22258487,0.20749438,0.15467763,0.08677038,0.02263575,0.02263575,0.026408374,0.041498873,0.06413463,0.08299775,0.090543,0.090543,0.094315626,0.094315626,0.06413463,0.0754525,0.071679875,0.06413463,0.0452715,0.0150905,0.00754525,0.02263575,0.033953626,0.041498873,0.071679875,0.12826926,0.17731337,0.3055826,0.52062225,0.7809334,0.80356914,0.814887,0.7809334,0.7130261,0.66775465,0.69039035,0.6790725,0.7205714,0.9280658,1.4147344,2.203213,2.8181508,3.3764994,3.8971217,4.285702,3.9763467,3.0897799,2.071171,1.5052774,2.11267,4.8063245,6.8246784,6.1003346,3.3350005,2.003264,1.3656902,0.98842776,0.7884786,0.69039035,0.663982,0.7394345,0.7394345,0.65643674,0.573439,0.6526641,0.69793564,0.59607476,0.42630664,0.27540162,0.24899325,0.32067314,0.4376245,0.5772116,0.7092535,0.7809334,0.70170826,0.573439,0.44894236,0.36594462,0.35839936,0.43007925,0.44894236,0.44139713,0.44139713,0.47157812,0.4678055,0.44894236,0.43385187,0.42630664,0.41498876,0.41121614,0.5885295,0.88279426,1.2713746,1.7731338,2.6106565,3.108643,3.0143273,2.5276587,2.2899833,2.463524,2.5012503,2.4069347,2.2862108,2.3314822,2.3503454,2.6634734,2.9237845,2.9313297,2.6144292,2.6823363,2.746471,2.938875,3.2255943,3.3689542,3.2218218,3.3161373,3.4896781,3.6443558,3.7613072,4.0706625,4.29702,4.4177437,4.508287,4.7233267,4.957229,5.27413,5.753253,6.2851934,6.5643673,6.930312,7.273621,7.5905213,7.854605,7.997965,7.809334,7.5565677,7.3905725,7.3792543,7.4999785,7.4396167,7.145352,6.9567204,7.0246277,7.3377557,7.677292,7.964011,8.043237,7.907422,7.6923823,7.8244243,8.243186,8.771353,9.1825695,9.201432,8.684583,8.831716,8.944894,8.748717,8.379,7.9338303,7.7112455,7.6320205,7.6018395,7.5226145,7.250985,7.2698483,7.4584794,7.745199,8.099826,8.488406,8.892077,9.322156,9.808825,10.378491,10.917976,11.234878,11.18206,10.733118,9.989911,9.325929,8.537451,7.7338815,6.971811,6.273875,5.617439,4.979865,4.432834,4.074435,4.044254,3.9386206,3.8103511,3.5274043,3.0897799,2.625747,2.4899325,2.3880715,2.2484846,2.1051247,2.082489,2.2862108,2.5238862,2.7125173,2.8747404,3.1652324,3.3651814,3.4557245,3.5462675,3.7198083,4.0291634,4.093298,3.9159849,3.6934,3.4481792,3.0520537,2.7238352,2.535204,2.3805263,2.2183034,2.0372176,1.9730829,2.052308,2.142851,2.173032,2.1088974,1.9730829,1.8863125,1.871222,1.9164935,1.9730829,2.0183544,2.0598533,2.123988,2.2183034,2.3390274,2.4295704,2.969056,3.451952,3.6443558,3.6179473,4.1310244,4.2706113,4.06689,3.6066296,3.0407357,2.6672459,3.0709167,3.7499893,4.2291126,4.0480266,3.8405323,3.610402,3.5349495,3.6254926,3.7273536,3.8858037,3.9386206,3.8254418,3.5651307,3.240685,2.6446102,2.0673985,1.5769572,1.2789198,1.3128735,1.146878,0.8601585,0.573439,0.38103512,0.3470815,0.4376245,0.5394854,0.6413463,0.7130261,0.72811663,0.8865669,1.3241913,2.2409391,3.399135,4.0895257,4.1197066,3.772625,3.2972744,2.8256962,2.372981,1.8297231,1.478869,1.1204696,0.73566186,0.4979865,0.48666862,0.56212115,0.55080324,0.45648763,0.4678055,0.76584285,0.6073926,0.35839936,0.1961765,0.08677038,0.03772625,0.026408374,0.02263575,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,12.196897,13.505998,13.985121,13.739901,13.0646,12.427027,10.529396,8.190369,6.228604,5.0062733,4.432834,3.7688525,3.0407357,2.4559789,2.1277604,2.082489,1.6750455,1.2298758,0.8186596,0.47157812,0.15845025,0.1056335,0.0754525,0.08677038,0.13958712,0.19994913,0.124496624,0.060362,0.02263575,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.011317875,0.02263575,0.026408374,0.033953626,0.06413463,0.06790725,0.0452715,0.041498873,0.049044125,0.056589376,0.056589376,0.06790725,0.07922512,0.07922512,0.056589376,0.03772625,0.02263575,0.02263575,0.030181,0.0452715,0.03772625,0.0452715,0.071679875,0.12826926,0.23013012,0.36594462,0.41498876,0.3734899,0.2867195,0.23767537,0.29803738,0.3961256,0.56212115,0.8903395,1.5656394,2.505023,3.338773,4.172523,5.0666356,6.043745,5.4740787,4.606375,3.8141239,3.3840446,3.482133,2.2484846,2.0749438,2.5616124,3.108643,2.927557,2.9124665,3.2105038,3.9763467,5.413717,7.786698,8.99771,9.623966,9.884277,9.235386,6.379509,5.764571,5.9682927,6.224831,6.156924,5.7683434,6.360646,7.394345,7.6886096,7.594294,9.012801,10.072908,9.6051035,7.865923,6.013564,6.0626082,6.643593,5.9682927,4.5120597,2.8898308,1.8561316,1.4298248,1.5543215,1.629774,1.50905,1.50905,1.7693611,1.4977322,1.1129243,0.8224323,0.6488915,0.5583485,0.543258,0.5583485,0.573439,0.58098423,0.5583485,0.482896,0.392353,0.32067314,0.29049212,0.422534,0.36594462,0.24899325,0.17354076,0.19240387,0.2678564,0.32067314,0.34330887,0.33953625,0.32821837,0.3772625,0.3961256,0.4376245,0.56212115,0.83752275,0.6451189,0.5093044,0.5470306,0.95447415,2.0296721,1.7316349,1.1091517,0.7092535,0.8526133,1.6448646,2.3163917,2.8445592,3.3161373,3.7763977,4.195159,4.8063245,5.4740787,4.961002,3.3651814,2.1088974,1.2223305,0.5394854,0.21881226,0.19994913,0.1659955,0.16222288,0.241448,0.36971724,0.47912338,0.44516975,0.19994913,0.241448,0.36971724,0.4640329,0.482896,0.392353,0.56589377,0.66020936,0.543258,0.29426476,0.15467763,0.32067314,0.55457586,0.73188925,0.8337501,1.1242423,1.2223305,1.1204696,0.8865669,0.66775465,0.5470306,0.5093044,0.49421388,0.44516975,0.29049212,0.056589376,0.0,0.060362,0.1358145,0.08677038,0.018863125,0.026408374,0.15467763,0.29049212,0.150905,0.1056335,0.0754525,0.16222288,0.30935526,0.3169005,0.23013012,0.08299775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.02263575,0.03772625,0.026408374,0.018863125,0.02263575,0.026408374,0.018863125,0.0150905,0.0150905,0.011317875,0.00754525,0.003772625,0.0,0.011317875,0.030181,0.056589376,0.07922512,0.08299775,0.049044125,0.033953626,0.026408374,0.02263575,0.02263575,0.056589376,0.14713238,0.2678564,0.38480774,0.45648763,0.46026024,0.32444575,0.181086,0.116951376,0.1961765,0.45648763,0.5017591,0.44894236,0.32067314,0.041498873,0.03772625,0.049044125,0.06413463,0.08299775,0.090543,0.124496624,0.16222288,0.1961765,0.19994913,0.1358145,0.15467763,0.16222288,0.15845025,0.12826926,0.03772625,0.02263575,0.02263575,0.033953626,0.049044125,0.056589376,0.056589376,0.090543,0.19994913,0.35839936,0.5055317,0.7054809,0.88279426,0.94315624,0.8941121,0.8639311,0.8337501,0.754525,0.73188925,0.91674787,1.4864142,2.2711203,2.8785129,3.5953116,4.436607,5.1345425,5.1647234,4.036709,2.6446102,1.6939086,1.7240896,3.006782,5.492942,6.375736,4.889322,2.3088465,1.3920987,0.9318384,0.68661773,0.5319401,0.45648763,0.58475685,0.56589377,0.47535074,0.3772625,0.33953625,0.35839936,0.27540162,0.18863125,0.14713238,0.150905,0.19240387,0.28294688,0.40367088,0.5394854,0.6752999,0.6752999,0.6073926,0.5055317,0.40367088,0.35462674,0.38480774,0.38858038,0.39989826,0.44894236,0.56589377,0.56212115,0.56589377,0.5583485,0.51684964,0.4678055,0.452715,0.5055317,0.6488915,0.8903395,1.2261031,1.9240388,2.8521044,2.9313297,2.1956677,1.8033148,1.8863125,2.323937,2.6634734,2.7540162,2.7426984,2.252257,2.3277097,2.535204,2.7087448,2.9615107,3.1425967,3.0407357,3.0331905,3.187868,3.2670932,3.169005,3.5462675,4.032936,4.429062,4.689373,5.010046,5.172269,5.2364035,5.2552667,5.2892203,5.492942,5.8136153,6.2097406,6.6247296,6.9869013,7.5603404,8.058327,8.492179,8.82417,8.959985,8.616675,8.265821,7.997965,7.8432875,7.786698,7.5565677,7.1868505,6.828451,6.7039547,7.0774446,7.496206,7.8508325,8.099826,8.13378,7.7602897,7.6697464,7.8734684,8.273367,8.695901,8.873214,8.703445,8.477088,8.179051,7.8244243,7.454707,7.069899,6.79827,6.6360474,6.5341864,6.40969,6.3832817,6.398372,6.405917,6.405917,6.4511886,6.458734,6.4964604,6.5568223,6.673774,6.9227667,7.281166,7.8206515,8.084735,7.8734684,7.2585306,6.688864,5.9909286,5.3156285,4.7308717,4.2517486,3.8443048,3.5047686,3.3350005,3.3463185,3.4444065,3.289729,3.2255943,3.1425967,2.957738,2.6031113,2.6408374,2.5691576,2.4182527,2.293756,2.372981,2.625747,2.8822856,3.1199608,3.308592,3.4029078,3.3425457,3.3312278,3.4859054,3.7914882,4.085753,4.074435,3.9499383,3.7386713,3.429316,2.9652832,2.7200627,2.6710186,2.6823363,2.6634734,2.5804756,2.6182017,2.655928,2.6446102,2.565385,2.4182527,2.2484846,2.1956677,2.2258487,2.2748928,2.2598023,2.214531,2.191895,2.1843498,2.214531,2.3201644,2.5917933,3.3651814,3.983892,4.2027044,4.1762958,4.3800178,4.357382,4.032936,3.5047686,3.0407357,2.9200118,3.7235808,4.6214657,4.870459,3.8103511,4.183841,4.1800685,4.036709,3.85185,3.5764484,3.5764484,3.6028569,3.6292653,3.5160866,3.0105548,2.372981,1.8976303,1.539231,1.2562841,1.0299267,0.94692886,0.8111144,0.55457586,0.26408374,0.19994913,0.29049212,0.3470815,0.35839936,0.3734899,0.49421388,0.73566186,1.2110126,2.0636258,3.0558262,3.591539,3.270866,2.5767028,1.8976303,1.5430037,1.750498,2.0296721,1.9881734,1.6863633,1.2261031,0.7507524,0.7469798,0.6752999,0.46026024,0.1659955,0.0,0.011317875,0.018863125,0.03772625,0.05281675,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.00754525,0.0,0.0,12.770335,13.162688,14.852824,15.660167,14.709465,12.449662,10.38981,8.231868,6.40969,5.13077,4.4101987,3.8103511,3.240685,2.686109,2.2748928,2.2899833,2.546522,2.033445,1.2562841,0.56212115,0.120724,0.10940613,0.07922512,0.08677038,0.12826926,0.150905,0.1056335,0.056589376,0.02263575,0.0150905,0.0150905,0.003772625,0.0,0.00754525,0.0150905,0.0150905,0.0150905,0.00754525,0.00754525,0.0150905,0.0150905,0.026408374,0.041498873,0.05281675,0.071679875,0.1056335,0.1056335,0.08677038,0.071679875,0.056589376,0.0452715,0.0452715,0.03772625,0.02263575,0.02263575,0.0452715,0.056589376,0.071679875,0.08299775,0.1358145,0.3055826,0.48666862,0.6451189,0.5885295,0.3734899,0.27540162,0.2867195,0.4074435,0.47157812,0.4678055,0.56589377,0.965792,2.1956677,3.2859564,3.9310753,4.45547,4.640329,3.2105038,2.0258996,1.81086,2.1503963,2.372981,3.3312278,4.2064767,4.52715,4.195159,4.074435,4.3083377,4.398881,4.123479,3.5236318,4.696918,5.8513412,6.888813,7.232122,5.828706,5.5495315,5.4212623,5.4401255,5.4740787,5.2779026,5.462761,5.7570257,6.0248823,5.873977,4.6554193,4.9345937,5.3910813,4.719554,3.4255435,3.8141239,3.9989824,3.6783094,2.6936543,1.4637785,0.97710985,0.9393836,1.1053791,1.20724,1.1883769,1.1883769,1.2261031,1.1355602,1.0299267,0.95447415,0.87147635,0.7582976,0.66020936,0.55457586,0.45648763,0.3961256,0.43385187,0.46026024,0.44894236,0.39989826,0.35085413,0.33953625,0.27917424,0.21503963,0.1659955,0.1659955,0.30181,0.362172,0.3734899,0.35462674,0.3055826,0.392353,0.41121614,0.43007925,0.5319401,0.8224323,0.59230214,0.47912338,0.5583485,0.9808825,1.9693103,1.7957695,1.3619176,0.91674787,0.7054809,0.9620194,1.6825907,2.6295197,3.712263,4.6856003,5.172269,5.6363015,5.9909286,5.406172,3.9386206,2.546522,1.4373702,0.6375736,0.41876137,0.59607476,0.5357128,0.362172,0.38480774,0.47535074,0.5055317,0.33576363,0.17731337,0.211267,0.32067314,0.3961256,0.33576363,0.27540162,0.17731337,0.08677038,0.02263575,0.0,0.0,0.08299775,0.392353,0.965792,1.7240896,1.1242423,0.965792,0.965792,0.91297525,0.65643674,1.1317875,1.20724,0.98465514,0.63002837,0.35085413,0.071679875,0.0,0.0,0.0,0.0,0.0,0.12826926,0.33576363,0.45648763,0.21503963,0.21503963,0.27917424,0.271629,0.15845025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.08299775,0.1358145,0.1358145,0.08677038,0.0754525,0.06413463,0.041498873,0.0150905,0.0150905,0.033953626,0.041498873,0.02263575,0.0,0.0,0.00754525,0.02263575,0.033953626,0.0452715,0.033953626,0.030181,0.03772625,0.049044125,0.060362,0.071679875,0.120724,0.18863125,0.24899325,0.27540162,0.63002837,0.62625575,0.38858038,0.120724,0.120724,0.20749438,0.41121614,0.68661773,0.7507524,0.090543,0.06790725,0.07922512,0.090543,0.090543,0.090543,0.116951376,0.150905,0.1659955,0.15845025,0.120724,0.1358145,0.17354076,0.20372175,0.1961765,0.120724,0.049044125,0.02263575,0.026408374,0.0452715,0.0452715,0.033953626,0.030181,0.07922512,0.19994913,0.3961256,0.6526641,1.0374719,1.237421,1.1431054,0.83752275,0.694163,0.59230214,0.55457586,0.63002837,0.9016574,1.448688,1.8523588,2.41448,3.240685,4.2404304,5.1345425,4.3309736,2.9011486,1.7844516,1.7844516,2.5804756,4.52715,6.620957,7.0170827,3.0520537,1.6976813,0.9280658,0.55457586,0.4074435,0.32067314,0.34330887,0.41498876,0.41498876,0.33953625,0.29049212,0.241448,0.19994913,0.150905,0.1056335,0.090543,0.1056335,0.124496624,0.1659955,0.23390275,0.32067314,0.36971724,0.3734899,0.3470815,0.3169005,0.3055826,0.3055826,0.2867195,0.29803738,0.3470815,0.3961256,0.4074435,0.56589377,0.7092535,0.7582976,0.7469798,0.724344,0.7432071,0.77338815,0.7884786,0.76207024,0.77338815,0.8526133,1.0035182,1.1921495,1.327964,1.3015556,1.5807298,2.1353056,2.867195,3.5839937,2.6936543,2.4371157,2.7087448,3.3161373,3.953711,4.4516973,4.7233267,4.7120085,4.4516973,4.074435,3.8782585,3.8480775,4.134797,4.5912848,4.776143,4.7648253,4.7346444,4.7044635,4.715781,4.8365054,4.983638,5.221313,5.587258,6.058836,6.5455046,7.0849895,7.5188417,8.001738,8.507269,8.850578,9.031664,9.042982,8.944894,8.786444,8.590267,8.224322,7.7376537,7.4509344,7.492433,7.798016,8.175279,8.571404,8.778898,8.726082,8.469543,8.16396,8.224322,8.473316,8.7751255,9.016574,8.710991,8.269594,7.805561,7.3717093,6.94163,6.6247296,6.436098,6.2851934,6.126743,5.9796104,6.1531515,6.1229706,5.987156,5.8890676,6.013564,5.9494295,5.715527,5.330719,4.919503,4.7006907,4.7836885,5.0553174,5.3646727,5.511805,5.2175403,4.5724216,4.1612053,3.85185,3.5802212,3.3727267,3.138824,3.0633714,3.2784111,3.6179473,3.6179473,3.3727267,2.9992368,2.6634734,2.493705,2.5804756,2.9086938,2.8181508,2.674791,2.7125173,3.006782,3.0558262,3.1576872,3.3236825,3.500996,3.5839937,3.3425457,3.5387223,4.0178456,4.4894238,4.5007415,4.4403796,4.3347464,3.9914372,3.4896781,3.1727777,3.1614597,3.259548,3.338773,3.350091,3.3274553,3.361409,3.3350005,3.2331395,3.0897799,3.006782,2.7879698,2.7238352,2.71629,2.6634734,2.4559789,2.372981,2.2484846,2.1692593,2.1843498,2.3201644,3.0030096,3.7952607,4.496969,5.0553174,5.553304,5.553304,5.142088,4.5007415,3.9348478,3.8593953,4.1272516,4.5912848,5.1760416,5.666483,5.692891,5.300538,5.2288585,5.2250857,4.908185,3.783943,3.8820312,3.531177,3.048281,2.6106565,2.2447119,1.780679,1.5241405,1.3355093,1.1544232,1.0072908,0.83752275,0.6187105,0.39989826,0.21503963,0.090543,0.090543,0.15467763,0.241448,0.32444575,0.3961256,0.6790725,1.177059,1.7693611,2.2862108,2.516341,2.0787163,1.6222287,1.1732863,0.9318384,1.237421,2.1994405,3.3123648,3.561358,2.595566,0.70170826,0.33576363,0.26408374,0.1659955,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,17.591751,15.045229,13.487134,12.506252,11.827179,11.314102,10.853842,9.378746,7.4811153,5.7872066,4.957229,4.5950575,3.9159849,3.0331905,2.1654868,1.629774,1.6335466,1.5165952,1.0299267,0.3772625,0.21881226,0.16976812,0.090543,0.08299775,0.13204187,0.12826926,0.090543,0.049044125,0.02263575,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.0150905,0.026408374,0.026408374,0.02263575,0.011317875,0.003772625,0.003772625,0.00754525,0.018863125,0.0452715,0.08299775,0.11317875,0.094315626,0.060362,0.03772625,0.033953626,0.033953626,0.02263575,0.018863125,0.02263575,0.0452715,0.06790725,0.11317875,0.17354076,0.2867195,0.5357128,0.77716076,0.8601585,0.6752999,0.34330887,0.2263575,0.23013012,0.29803738,0.3961256,0.5017591,0.5998474,0.7696155,1.1544232,1.6109109,1.9429018,1.8787673,1.7014539,1.4637785,1.4298248,1.6524098,2.003264,2.4974778,2.9728284,3.7235808,4.6327834,5.172269,4.991183,4.9119577,4.727099,4.4215164,4.195159,4.7044635,5.119452,5.342037,5.2175403,4.534695,4.398881,4.6856003,5.081726,5.353355,5.3646727,5.5570765,5.1873593,4.5309224,3.8895764,3.5689032,3.7990334,3.7877154,3.3312278,2.6634734,2.4484336,2.795515,2.9200118,2.6106565,1.9429018,1.2713746,1.0487897,1.0638802,1.2562841,1.388326,1.056335,0.8865669,0.935611,1.1016065,1.3091009,1.5165952,1.4864142,1.146878,0.7809334,0.5281675,0.4074435,0.41498876,0.47157812,0.48666862,0.43007925,0.362172,0.32067314,0.24899325,0.17731337,0.1358145,0.15467763,0.24899325,0.2867195,0.2867195,0.26031113,0.23013012,0.23013012,0.4640329,0.7054809,0.814887,0.7394345,0.58475685,0.69793564,1.0450171,1.569412,2.1881225,1.7919968,1.4109617,1.1053791,1.0186088,1.3505998,2.2975287,3.4632697,4.772371,5.764571,5.587258,5.7306175,5.915476,5.670255,4.776143,3.2557755,1.8523588,0.77338815,0.30181,0.32444575,0.35085413,0.3055826,0.19240387,0.13204187,0.14713238,0.13958712,0.15845025,0.16222288,0.19240387,0.24522063,0.26408374,0.181086,0.13204187,0.08299775,0.033953626,0.0,0.0,0.02263575,0.241448,0.7054809,1.3355093,1.116697,1.0299267,1.1053791,1.358145,1.8146327,1.0223814,0.60362,0.46026024,0.41121614,0.1659955,0.033953626,0.0,0.0,0.0,0.0,0.0,0.026408374,0.06790725,0.090543,0.041498873,0.041498873,0.181086,0.27540162,0.271629,0.21881226,0.150905,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.049044125,0.08299775,0.10186087,0.10940613,0.12826926,0.12826926,0.10940613,0.0754525,0.056589376,0.071679875,0.090543,0.094315626,0.060362,0.041498873,0.030181,0.033953626,0.041498873,0.0452715,0.033953626,0.030181,0.030181,0.033953626,0.03772625,0.1056335,0.17731337,0.1659955,0.124496624,0.2263575,0.4640329,0.5470306,0.5470306,0.48666862,0.32821837,0.19994913,0.17354076,0.25276586,0.32067314,0.13958712,0.056589376,0.14335975,0.23390275,0.24899325,0.19994913,0.13958712,0.1358145,0.13958712,0.120724,0.08677038,0.060362,0.0452715,0.041498873,0.03772625,0.02263575,0.030181,0.02263575,0.02263575,0.0452715,0.094315626,0.090543,0.08299775,0.06413463,0.05281675,0.090543,0.29803738,0.70170826,1.1544232,1.478869,1.4373702,1.3694628,1.4109617,1.2525115,0.935611,0.8526133,0.814887,0.845068,1.1280149,1.9202662,3.5462675,4.5837393,4.3800178,3.3048196,2.1277604,2.04099,2.6597006,3.663219,4.8365054,5.379763,3.8820312,2.3503454,1.4411428,0.9695646,0.724344,0.5017591,0.3734899,0.30935526,0.2678564,0.24522063,0.26408374,0.32444575,0.23767537,0.13204187,0.06790725,0.056589376,0.0754525,0.094315626,0.13204187,0.19994913,0.28294688,0.30181,0.3055826,0.2867195,0.25276586,0.21881226,0.19994913,0.19240387,0.19240387,0.22258487,0.29803738,0.30181,0.35462674,0.4376245,0.51684964,0.56589377,0.55080324,0.55080324,0.5772116,0.6073926,0.60362,0.6752999,0.83752275,1.146878,1.4713237,1.4977322,1.2487389,1.0186088,1.0110635,1.2826926,1.7316349,1.931584,2.173032,2.7615614,3.7009451,4.696918,5.481624,6.319147,6.643593,6.296511,5.5382137,4.7006907,4.244203,4.032936,3.9763467,4.032936,4.2064767,4.504514,4.817642,5.062863,5.2137675,5.5759397,5.7381625,5.7570257,5.7306175,5.7909794,6.1305156,6.688864,7.356619,7.9753294,8.326183,8.820397,9.318384,9.688101,9.903141,10.020092,9.778644,9.635284,9.703192,9.88805,9.87296,9.978593,10.106862,10.065364,9.820143,9.507015,9.239159,9.039209,8.903395,8.831716,8.809079,8.503497,7.8734684,7.3188925,6.9491754,6.541732,6.2323766,5.9796104,5.7570257,5.5759397,5.4703064,5.4250345,5.281675,5.05909,4.821415,4.6818275,4.659192,4.5799665,4.436607,4.2404304,4.0404816,4.06689,4.115934,4.214022,4.3385186,4.436607,3.9574835,3.712263,3.5387223,3.3425457,3.1161883,3.0218725,3.0822346,3.1425967,3.1727777,3.2520027,2.9464202,2.595566,2.3428001,2.263575,2.3578906,2.6785638,2.957738,3.1237335,3.2520027,3.5538127,3.682082,3.731126,3.742444,3.7537618,3.8292143,3.8292143,4.115934,4.6214657,5.119452,5.2099953,4.8440504,4.3686996,4.0103,3.85185,3.8556228,3.874486,3.7877154,3.7273536,3.7462165,3.8405323,3.8858037,3.7273536,3.4745877,3.240685,3.1652324,2.9728284,2.7728794,2.6182017,2.5427492,2.5427492,2.6219745,2.6521554,2.7087448,2.8709676,3.2105038,4.1197066,4.719554,5.0779533,5.240176,5.2137675,5.221313,5.194905,4.825187,4.293247,4.2517486,4.696918,4.908185,5.0213637,5.1873593,5.594803,6.0512905,5.7419353,5.251494,4.847823,4.466788,4.183841,3.591539,3.0407357,2.6446102,2.2673476,1.901403,1.7391801,1.5203679,1.1921495,0.90920264,0.69039035,0.694163,0.7092535,0.6488915,0.55457586,0.35085413,0.20749438,0.14713238,0.16976812,0.26408374,0.59230214,1.0751982,1.4637785,1.5845025,1.358145,1.0638802,0.8337501,0.663982,0.6149379,0.8337501,1.2411937,1.6033657,1.5279131,0.9695646,0.23767537,0.1056335,0.1358145,0.23013012,0.26408374,0.09808825,0.018863125,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,16.731592,16.052519,13.920986,11.781908,10.33322,9.510788,9.137298,8.273367,7.250985,6.349328,5.802297,5.3344917,4.5988297,3.6368105,2.6031113,1.7580433,1.7693611,1.50905,1.0035182,0.47157812,0.33576363,0.19994913,0.1056335,0.08299775,0.10940613,0.1056335,0.08299775,0.060362,0.049044125,0.041498873,0.00754525,0.02263575,0.03772625,0.033953626,0.018863125,0.0150905,0.011317875,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.018863125,0.056589376,0.094315626,0.10940613,0.090543,0.056589376,0.030181,0.02263575,0.02263575,0.02263575,0.026408374,0.03772625,0.0452715,0.07922512,0.124496624,0.18485862,0.271629,0.422534,0.58098423,0.633801,0.5470306,0.3772625,0.2678564,0.21881226,0.23013012,0.32067314,0.482896,0.7205714,0.7054809,0.7167987,0.80356914,0.90920264,0.87147635,1.8372684,2.957738,3.7537618,3.9008942,3.2218218,3.5123138,4.142342,4.406426,4.466788,5.372218,5.775889,5.6287565,5.342037,5.0553174,4.666737,4.3913355,4.3347464,4.376245,4.3913355,4.221567,4.085753,4.195159,4.3422914,4.395108,4.2894745,4.247976,4.3007927,4.0895257,3.5990841,3.1576872,3.7386713,3.7688525,3.4745877,3.0445085,2.6634734,2.6823363,2.6597006,2.4899325,2.1202152,1.5543215,1.4750963,1.5128226,1.6335466,1.6637276,1.2713746,0.97710985,0.9016574,0.97333723,1.2110126,1.7429527,1.8900851,1.6788181,1.2789198,0.875249,0.66020936,0.59230214,0.6073926,0.56212115,0.43007925,0.31312788,0.2263575,0.1659955,0.12826926,0.10940613,0.124496624,0.181086,0.20372175,0.20749438,0.1961765,0.18485862,0.16976812,0.452715,0.7205714,0.80734175,0.67152727,0.7922512,1.4109617,2.0975795,2.4974778,2.335255,1.8825399,1.569412,1.4071891,1.4637785,1.871222,3.150142,4.346064,5.323174,5.7004366,4.8666863,5.0515447,5.3156285,5.1156793,4.2706113,2.938875,1.6976813,0.7054809,0.23390275,0.22258487,0.27917424,0.26408374,0.116951376,0.030181,0.05281675,0.071679875,0.11317875,0.1659955,0.19240387,0.18863125,0.181086,0.14713238,0.16976812,0.16222288,0.094315626,0.0,0.0452715,0.15845025,0.3734899,0.68661773,1.0450171,0.8865669,0.7582976,0.84129536,1.2449663,2.033445,1.0450171,0.49421388,0.27540162,0.2263575,0.13958712,0.08677038,0.056589376,0.026408374,0.0,0.0,0.0,0.0,0.026408374,0.07922512,0.1358145,0.116951376,0.1056335,0.10940613,0.120724,0.10940613,0.0754525,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.0150905,0.0150905,0.018863125,0.03772625,0.08299775,0.08299775,0.08677038,0.08299775,0.0754525,0.090543,0.0754525,0.06790725,0.08299775,0.116951376,0.13204187,0.09808825,0.056589376,0.033953626,0.041498873,0.056589376,0.124496624,0.24522063,0.24899325,0.1358145,0.0754525,0.08677038,0.11317875,0.120724,0.124496624,0.20372175,0.2867195,0.35085413,0.39989826,0.41498876,0.38103512,0.38103512,0.3055826,0.25276586,0.23390275,0.18863125,0.181086,0.1961765,0.32067314,0.5319401,0.7054809,0.39989826,0.26031113,0.21881226,0.19240387,0.11317875,0.060362,0.026408374,0.003772625,0.0,0.00754525,0.026408374,0.02263575,0.018863125,0.116951376,0.49044126,4.4101987,8.944894,7.6584287,1.7467253,0.02263575,0.10940613,0.32821837,0.5885295,0.84129536,1.0940613,1.8259505,3.4594972,3.9008942,2.8219235,1.6637276,0.8941121,0.5583485,0.6187105,1.177059,2.4823873,4.3724723,4.402653,3.4368613,2.3126192,1.8297231,2.516341,3.240685,3.9273026,4.266839,3.731126,2.5389767,1.7467253,1.267602,0.98465514,0.7432071,0.9016574,0.8941121,0.65643674,0.331991,0.2867195,0.34330887,0.32444575,0.271629,0.20749438,0.12826926,0.08677038,0.0754525,0.10186087,0.1659955,0.27540162,0.35839936,0.43007925,0.46026024,0.45648763,0.45648763,0.46026024,0.4678055,0.44139713,0.38480774,0.32821837,0.24899325,0.21881226,0.23390275,0.28294688,0.34330887,0.39989826,0.46026024,0.513077,0.5281675,0.5017591,0.5357128,0.70170826,1.0110635,1.3845534,1.6788181,1.5845025,1.4826416,1.4750963,1.6410918,2.0258996,2.4371157,2.8294687,3.3651814,3.9574835,4.304565,4.7421894,5.247721,5.5080323,5.5193505,5.594803,5.0251365,4.3121104,3.863168,3.7952607,3.9386206,4.315883,4.8855495,5.451443,5.9418845,6.398372,6.749226,6.6020937,6.2097406,5.802297,5.59103,5.8098426,6.319147,6.9755836,7.6697464,8.296002,9.009028,9.95973,10.808571,11.385782,11.68382,11.506506,11.299012,11.227332,11.332966,11.52537,11.4838705,11.400873,11.242422,11.038701,10.899114,10.27663,9.650374,9.118435,8.707218,8.36391,7.914967,7.3868,7.009537,6.7567716,6.3832817,6.085244,5.8211603,5.583485,5.3759904,5.1760416,4.983638,4.776143,4.4441524,4.0404816,3.7914882,3.772625,3.85185,3.9801195,4.1008434,4.1310244,4.1310244,4.2027044,4.402653,4.6931453,4.9459114,4.5497856,4.255521,3.92353,3.4859054,2.9615107,2.8709676,2.957738,3.059599,3.1312788,3.2482302,2.6634734,2.282438,2.1353056,2.1881225,2.3503454,2.7540162,3.1539145,3.4444065,3.6481283,3.9310753,4.063117,4.2102494,4.478106,4.738417,4.640329,4.9949555,5.666483,6.221059,6.349328,5.8702044,5.270357,4.938366,4.772371,4.708236,4.7044635,4.61392,4.436607,4.398881,4.538468,4.689373,4.666737,4.2404304,3.783943,3.4934506,3.361409,3.2067313,3.029418,2.916239,2.9049213,2.9841464,2.916239,2.8596497,2.938875,3.2520027,3.863168,4.8440504,5.3609,5.5382137,5.511805,5.409944,5.6589375,5.783434,5.6287565,5.6815734,7.0510364,7.092535,6.530414,5.7306175,5.1873593,5.534441,6.0362,6.0776987,5.9192486,5.6363015,5.0968165,4.315883,3.4255435,2.7125173,2.2220762,1.7316349,1.3392819,1.1280149,0.935611,0.724344,0.573439,0.5093044,0.52062225,0.56212115,0.6111652,0.67152727,0.70170826,0.452715,0.211267,0.124496624,0.19240387,0.3961256,0.7394345,1.0186088,1.0676528,0.784706,0.62248313,0.6488915,0.73566186,0.73566186,0.48666862,0.9016574,1.3543724,1.6146835,1.4298248,0.543258,0.20749438,0.090543,0.1056335,0.13958712,0.049044125,0.011317875,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,11.249968,12.808062,12.3893,11.23865,10.155907,9.457971,9.159933,8.699674,8.080963,7.2472124,6.092789,5.2779026,4.738417,3.9461658,2.8709676,1.9579924,1.8070874,1.4298248,0.9695646,0.5696664,0.38480774,0.241448,0.15845025,0.120724,0.10940613,0.1056335,0.090543,0.071679875,0.06413463,0.05281675,0.0150905,0.0452715,0.06790725,0.06413463,0.03772625,0.0150905,0.00754525,0.011317875,0.011317875,0.00754525,0.011317875,0.011317875,0.018863125,0.0452715,0.07922512,0.094315626,0.09808825,0.08677038,0.060362,0.033953626,0.026408374,0.026408374,0.033953626,0.041498873,0.05281675,0.06413463,0.10186087,0.14335975,0.18863125,0.24899325,0.35839936,0.5055317,0.56589377,0.5394854,0.452715,0.32821837,0.24899325,0.2678564,0.3470815,0.47912338,0.694163,0.62625575,0.573439,0.55457586,0.59607476,0.72811663,2.9200118,4.45547,5.1534057,4.927048,3.7914882,4.074435,4.6742826,4.6629643,4.398881,5.534441,6.530414,6.628502,6.1078796,5.2779026,4.4705606,3.8556228,3.640583,3.682082,3.7801702,3.6707642,3.4670424,3.4179983,3.591539,3.8443048,3.8292143,3.6141748,3.7877154,3.7084904,3.2105038,2.6144292,3.2105038,3.6858547,3.9273026,3.8971217,3.62172,2.9426475,2.5389767,2.3390274,2.2560298,2.1881225,2.252257,2.082489,1.841041,1.6524098,1.6109109,1.2751472,1.0601076,0.995973,1.2034674,1.8636768,1.9806281,1.7995421,1.4071891,0.97710985,0.77338815,0.663982,0.6073926,0.5093044,0.35839936,0.23767537,0.16222288,0.12826926,0.120724,0.124496624,0.13204187,0.13958712,0.13958712,0.1358145,0.1358145,0.1358145,0.12826926,0.32444575,0.5357128,0.66020936,0.6828451,0.8978847,1.5165952,2.142851,2.4522061,2.2069857,1.871222,1.7354075,1.7995421,2.0862615,2.6521554,3.682082,4.406426,4.7535076,4.617693,3.8782585,3.8782585,3.9386206,3.6934,3.0633714,2.2296214,1.3543724,0.59230214,0.1961765,0.17354076,0.27917424,0.23767537,0.116951376,0.06790725,0.10940613,0.12826926,0.10940613,0.1659955,0.19994913,0.1961765,0.241448,0.24899325,0.22258487,0.2565385,0.32444575,0.26408374,0.38103512,0.694163,0.965792,1.0827434,1.0751982,1.1846043,1.0223814,0.88279426,0.97710985,1.4222796,0.95447415,0.5998474,0.34330887,0.17731337,0.090543,0.0754525,0.056589376,0.026408374,0.0,0.0,0.0,0.0,0.026408374,0.07922512,0.1358145,0.116951376,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.011317875,0.003772625,0.0,0.011317875,0.05281675,0.0452715,0.033953626,0.026408374,0.033953626,0.071679875,0.0754525,0.05281675,0.060362,0.1056335,0.150905,0.14713238,0.09808825,0.06790725,0.08299775,0.13958712,0.32444575,0.39989826,0.3169005,0.150905,0.0754525,0.05281675,0.049044125,0.08299775,0.14713238,0.21503963,0.19240387,0.19240387,0.20749438,0.23767537,0.29426476,0.4376245,0.44894236,0.3961256,0.33576363,0.32444575,0.32821837,0.31312788,0.5696664,0.95447415,0.91297525,0.44516975,0.28294688,0.24522063,0.21881226,0.14335975,0.090543,0.041498873,0.011317875,0.00754525,0.02263575,0.03772625,0.030181,0.018863125,0.124496624,0.55080324,4.666737,9.242931,8.299775,3.1312788,2.3126192,0.98842776,0.4074435,0.26408374,0.41498876,0.8903395,1.991946,4.274384,5.5797124,5.2137675,3.9499383,2.3201644,1.2789198,0.8563859,1.116697,2.1805773,4.395108,4.8063245,3.802806,2.2711203,1.6109109,2.1503963,2.8219235,3.5274043,3.9612563,3.62172,2.6710186,1.9391292,1.4411428,1.1431054,0.9242931,1.1280149,1.1921495,0.95447415,0.5357128,0.36594462,0.27540162,0.29049212,0.32821837,0.33953625,0.29803738,0.15845025,0.10186087,0.09808825,0.1358145,0.21503963,0.3169005,0.41498876,0.482896,0.5394854,0.6375736,0.6752999,0.69039035,0.66775465,0.60362,0.5017591,0.44894236,0.4376245,0.422534,0.39989826,0.392353,0.5319401,0.7394345,0.8111144,0.7205714,0.5998474,0.5357128,0.6073926,0.8299775,1.20724,1.7655885,2.1353056,2.3956168,2.4899325,2.4974778,2.6182017,2.7841973,3.029418,3.3878171,3.7575345,3.904667,4.0291634,4.1762958,4.323428,4.5535583,5.040227,4.776143,4.214022,3.8782585,3.9499383,4.266839,4.817642,5.5570765,6.33801,6.9680386,7.2170315,7.1264887,6.7152724,6.2399216,5.855114,5.621211,5.7494807,6.1305156,6.7756343,7.6508837,8.661947,9.563604,10.518079,11.336739,11.910177,12.2270775,12.219532,12.174261,12.200669,12.355347,12.649611,12.468526,12.204442,11.932813,11.68382,11.449917,10.514306,9.623966,8.903395,8.367682,7.914967,7.4471617,7.0812173,6.8133607,6.587003,6.255012,6.013564,5.753253,5.492942,5.2137675,4.881777,4.6026025,4.346064,4.002755,3.610402,3.361409,3.350091,3.5123138,3.8254418,4.217795,4.564876,4.659192,4.715781,4.8629136,5.0779533,5.2137675,4.8968673,4.515832,3.9989824,3.3953626,2.867195,3.0256453,3.0709167,3.0407357,2.9803739,2.938875,2.5314314,2.372981,2.444661,2.6785638,2.9615107,3.2935016,3.5689032,3.7688525,3.942393,4.191386,4.285702,4.4894238,4.930821,5.5683947,6.187105,6.5643673,6.990674,7.1566696,6.9567204,6.48137,6.175787,6.175787,6.1833324,6.175787,6.3719635,6.4210076,6.3531003,6.2663302,6.1795597,6.0286546,5.7004366,5.1571784,4.6818275,4.349837,4.036709,3.663219,3.470815,3.429316,3.5085413,3.6481283,3.5424948,3.591539,3.8593953,4.3875628,5.2137675,6.058836,6.2889657,6.149379,5.8890676,5.7419353,6.0362,6.1644692,6.138061,6.417235,7.8734684,7.647111,6.9189944,5.9418845,5.1835866,5.342037,5.621211,5.7494807,5.5193505,4.949684,4.274384,3.5123138,2.795515,2.1164427,1.4977322,0.995973,0.724344,0.56589377,0.44516975,0.33953625,0.29426476,0.3169005,0.32067314,0.35462674,0.44516975,0.58475685,0.784706,0.6149379,0.36594462,0.20749438,0.16222288,0.211267,0.38480774,0.56212115,0.6375736,0.5093044,0.47912338,0.56589377,0.6451189,0.58475685,0.24899325,0.55457586,1.0186088,1.4713237,1.5279131,0.5998474,0.20749438,0.049044125,0.00754525,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.666737,6.515323,8.213005,9.333474,9.895596,10.370946,10.627484,10.397354,9.567377,8.058327,5.8211603,4.708236,4.3875628,3.8141239,2.7992878,2.022127,1.4977322,1.1695137,0.9016574,0.6488915,0.45648763,0.4376245,0.42630664,0.35085413,0.22258487,0.15467763,0.124496624,0.09808825,0.0754525,0.06413463,0.0452715,0.08299775,0.09808825,0.08677038,0.06413463,0.030181,0.0452715,0.0452715,0.033953626,0.02263575,0.033953626,0.049044125,0.06413463,0.07922512,0.090543,0.07922512,0.08677038,0.08299775,0.071679875,0.056589376,0.05281675,0.0452715,0.049044125,0.060362,0.08677038,0.124496624,0.150905,0.17354076,0.19994913,0.26031113,0.4074435,0.59230214,0.66020936,0.6111652,0.482896,0.362172,0.30935526,0.35085413,0.41498876,0.47912338,0.5470306,0.55457586,0.5885295,0.7469798,1.0601076,1.5052774,4.032936,4.870459,4.745962,4.195159,3.5538127,4.1083884,4.4139714,4.5007415,4.745962,5.8702044,6.8397694,7.1981683,6.56814,5.2628117,4.266839,3.8367596,3.5990841,3.3840446,3.1161883,2.8143783,2.565385,2.5389767,2.9841464,3.6971724,4.002755,3.8367596,3.5990841,3.0445085,2.2975287,1.8561316,2.0636258,2.886058,3.7801702,4.3649273,4.436607,3.3425457,2.5616124,2.214531,2.305074,2.6974268,2.7238352,2.2371666,1.6410918,1.3392819,1.7391801,1.50905,1.2864652,1.1996948,1.3619176,1.8825399,1.7693611,1.4939595,1.1393328,0.814887,0.6828451,0.573439,0.4640329,0.362172,0.271629,0.16976812,0.1358145,0.124496624,0.13204187,0.150905,0.150905,0.124496624,0.10186087,0.090543,0.094315626,0.09808825,0.1056335,0.16976812,0.32444575,0.543258,0.754525,0.8563859,1.0601076,1.3732355,1.7467253,2.0749438,1.8221779,1.8334957,2.0787163,2.5578396,3.2859564,3.7688525,3.874486,3.6745367,3.3123648,2.9841464,2.6219745,2.3013012,2.0485353,1.8259505,1.5316857,1.0940613,0.56589377,0.211267,0.14713238,0.33576363,0.241448,0.15845025,0.150905,0.20372175,0.23013012,0.16222288,0.14713238,0.14713238,0.181086,0.3169005,0.33953625,0.21503963,0.2867195,0.55457586,0.69039035,1.0487897,1.3958713,1.5505489,1.4637785,1.237421,1.750498,1.6033657,1.1921495,0.8111144,0.6488915,0.724344,0.633801,0.44516975,0.2263575,0.041498873,0.00754525,0.0,0.026408374,0.060362,0.03772625,0.02263575,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.02263575,0.0150905,0.011317875,0.02263575,0.0452715,0.060362,0.041498873,0.0452715,0.07922512,0.11317875,0.15845025,0.15467763,0.15845025,0.20372175,0.31312788,0.513077,0.38858038,0.18863125,0.06413463,0.03772625,0.030181,0.026408374,0.056589376,0.12826926,0.2263575,0.1961765,0.16976812,0.14713238,0.1358145,0.150905,0.30181,0.44139713,0.513077,0.52062225,0.5470306,0.47157812,0.46026024,0.84129536,1.297783,0.87902164,0.46026024,0.27917424,0.211267,0.17354076,0.15467763,0.120724,0.060362,0.026408374,0.026408374,0.041498873,0.06790725,0.060362,0.03772625,0.060362,0.21503963,0.754525,0.9808825,1.8372684,3.783943,6.7944975,3.5085413,1.2449663,0.29426476,0.44139713,0.94315624,1.7014539,3.150142,4.9647746,6.4021444,6.3342376,4.5007415,2.7502437,1.6863633,1.6863633,2.9351022,5.194905,6.1795597,5.010046,2.5729303,1.5618668,1.7542707,2.41448,3.4557245,4.376245,4.2706113,3.0671442,2.1390784,1.5279131,1.1883769,0.965792,0.90543,0.9507015,0.8941121,0.69039035,0.47157812,0.21881226,0.181086,0.24522063,0.33576363,0.40367088,0.21881226,0.1358145,0.10186087,0.094315626,0.10940613,0.16222288,0.2263575,0.29426476,0.38858038,0.55457586,0.6149379,0.63002837,0.633801,0.63002837,0.60362,0.66775465,0.73566186,0.7394345,0.66775465,0.5772116,0.73566186,1.0751982,1.2261031,1.1317875,1.0450171,0.87147635,0.7997965,0.87902164,1.1657411,1.7165444,2.4861598,2.9652832,3.0445085,2.8143783,2.595566,2.5276587,2.5917933,2.8898308,3.4029078,3.9725742,4.032936,4.063117,4.1498876,4.293247,4.3913355,4.2064767,4.093298,4.093298,4.2819295,4.7836885,5.4967146,6.221059,7.001992,7.541477,7.2358947,6.6247296,6.19465,6.0022464,5.9720654,5.9003854,5.9418845,6.221059,6.900131,7.9941926,9.348565,10.378491,10.963248,11.302785,11.544232,11.778135,11.989402,12.30253,12.672247,13.000465,13.151371,12.864652,12.472299,12.068627,11.642321,11.068882,10.0465,9.114662,8.401636,7.91874,7.564113,7.2698483,7.020855,6.7756343,6.515323,6.270103,6.096562,5.80607,5.4401255,5.0251365,4.587512,4.2781568,4.002755,3.7499893,3.5160866,3.3123648,3.3576362,3.5689032,3.9725742,4.5233774,5.119452,5.353355,5.330719,5.198677,5.028909,4.7836885,4.4630156,4.025391,3.4859054,2.987919,2.8143783,3.2972744,3.2859564,3.0369632,2.746471,2.5540671,2.757789,2.9992368,3.2972744,3.6292653,3.942393,4.0517993,4.1083884,4.142342,4.2102494,4.406426,4.4894238,4.7648253,5.2665844,6.1531515,7.707473,7.858378,7.6282477,7.303802,7.1000805,7.194396,7.4584794,7.7187905,7.8734684,8.069645,8.710991,9.06939,9.14107,8.854351,8.280911,7.643338,6.9680386,6.4549613,6.1041074,5.794752,5.304311,4.6327834,4.3347464,4.2630663,4.327201,4.5233774,4.715781,5.0741806,5.59103,6.25124,7.0472636,7.466025,7.1868505,6.6322746,6.1305156,5.9117036,6.092789,6.1078796,6.1041074,6.205968,6.5002327,6.40969,6.138061,5.6023483,5.040227,4.979865,4.9760923,4.696918,3.904667,2.8822856,2.4295704,2.093807,1.8448136,1.4034165,0.814887,0.4376245,0.39989826,0.392353,0.331991,0.2263575,0.16222288,0.15467763,0.19240387,0.24522063,0.32067314,0.4640329,0.66020936,0.6375736,0.51684964,0.35839936,0.1961765,0.124496624,0.16222288,0.26408374,0.39989826,0.55080324,0.6111652,0.58098423,0.44894236,0.271629,0.1358145,0.2263575,0.5470306,0.90543,0.98842776,0.362172,0.11317875,0.018863125,0.0,0.0,0.0,0.011317875,0.0150905,0.018863125,0.018863125,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.9464202,2.969056,3.7990334,5.198677,6.828451,8.269594,9.016574,9.0543,8.541223,7.496206,5.798525,4.9685473,4.221567,3.4934506,2.8030603,2.2447119,1.50905,1.0789708,0.9393836,0.94692886,0.8224323,1.0676528,1.2487389,1.0601076,0.58098423,0.29049212,0.19240387,0.1659955,0.16222288,0.15467763,0.1659955,0.20372175,0.20372175,0.16222288,0.1056335,0.090543,0.1659955,0.12826926,0.06790725,0.033953626,0.0452715,0.120724,0.120724,0.10186087,0.090543,0.090543,0.07922512,0.08677038,0.09808825,0.10186087,0.0754525,0.05281675,0.06413463,0.10186087,0.16222288,0.26031113,0.23390275,0.211267,0.19994913,0.21503963,0.27540162,0.31312788,0.32821837,0.32444575,0.31312788,0.35085413,0.3734899,0.3169005,0.3055826,0.38858038,0.5357128,0.66775465,0.80356914,1.4449154,2.6408374,3.983892,5.4967146,5.243949,4.5950575,4.247976,4.2102494,4.798779,5.2175403,5.5306683,5.783434,6.0286546,5.7570257,5.7570257,5.956975,6.1229706,5.828706,5.7306175,5.1571784,4.032936,2.8634224,2.71629,2.546522,2.4672968,2.5012503,2.686109,3.0520537,3.187868,2.9464202,2.4182527,1.8297231,1.5241405,1.539231,1.7429527,2.4220252,3.4255435,4.1800685,4.1310244,3.0746894,2.203213,1.9051756,1.7693611,1.5505489,1.267602,1.0714256,1.0450171,1.1883769,1.3619176,1.3505998,1.2940104,1.3091009,1.478869,1.297783,1.1581959,1.0374719,0.87902164,0.6111652,0.5017591,0.42630664,0.36594462,0.27917424,0.120724,0.049044125,0.041498873,0.06413463,0.090543,0.090543,0.090543,0.090543,0.090543,0.09808825,0.120724,0.15845025,0.23013012,0.38480774,0.59607476,0.77716076,0.9016574,1.2336484,1.750498,2.3201644,2.686109,2.052308,1.7919968,1.8523588,2.1994405,2.8219235,3.7273536,4.0895257,3.92353,3.240685,2.0447628,1.8485862,1.7014539,1.50905,1.2638294,1.0072908,1.0676528,0.73566186,0.35839936,0.19994913,0.45648763,0.32444575,0.2263575,0.18863125,0.20749438,0.24522063,0.23013012,0.090543,0.0,0.0,0.0,0.011317875,0.060362,0.14713238,0.3470815,0.8224323,1.8863125,1.5731846,1.0186088,0.7997965,0.94692886,1.3015556,1.1959221,0.97710985,0.8563859,0.9318384,0.56589377,0.33576363,0.2263575,0.19994913,0.21503963,0.041498873,0.0,0.1358145,0.3055826,0.18485862,0.120724,0.07922512,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.08677038,0.18485862,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.049044125,0.060362,0.060362,0.05281675,0.041498873,0.033953626,0.0452715,0.02263575,0.0150905,0.026408374,0.05281675,0.0754525,0.10186087,0.18863125,0.3055826,0.422534,0.5357128,0.41121614,0.26408374,0.1358145,0.060362,0.060362,0.03772625,0.011317875,0.011317875,0.056589376,0.150905,0.24899325,0.32821837,0.2867195,0.150905,0.090543,0.150905,0.32444575,0.55080324,0.7432071,0.77716076,0.6451189,0.47157812,0.6375736,1.0978339,1.4034165,1.2562841,0.67152727,0.24899325,0.1659955,0.1659955,0.14335975,0.10186087,0.071679875,0.06413463,0.0754525,0.124496624,0.12826926,0.090543,0.041498873,0.030181,0.77338815,1.539231,2.5502944,5.0025005,11.031156,7.91874,2.9766011,0.18485862,0.211267,0.38103512,0.7130261,1.1242423,2.293756,4.06689,5.43258,5.6287565,4.1762958,2.8256962,2.6898816,4.2404304,7.964011,9.288202,7.7942433,4.4441524,1.5882751,1.7089992,2.4974778,3.7273536,5.0666356,6.1041074,3.942393,2.4974778,1.6184561,1.1242423,0.80734175,0.73566186,0.663982,0.5696664,0.4979865,0.5357128,0.38858038,0.24899325,0.15845025,0.120724,0.120724,0.08677038,0.06790725,0.049044125,0.03772625,0.060362,0.08677038,0.120724,0.1358145,0.13958712,0.150905,0.19994913,0.22258487,0.21503963,0.19994913,0.21503963,0.23767537,0.29049212,0.32821837,0.331991,0.32067314,0.331991,0.59230214,1.0072908,1.4977322,1.9994912,1.7655885,1.599593,1.478869,1.4373702,1.5731846,1.9881734,2.1805773,2.1277604,1.961765,1.9994912,2.1805773,2.5314314,3.127506,3.85185,4.3649273,4.3649273,4.146115,4.0480266,4.074435,3.8895764,3.8895764,4.074435,4.2894745,4.587512,5.2326307,6.2097406,6.6020937,6.752999,6.820906,6.760544,6.428553,6.4021444,6.541732,6.7152724,6.790725,6.752999,7.066127,7.7376537,8.797762,10.299266,11.249968,11.664956,11.7555,11.763044,11.947904,12.128989,12.340257,12.574159,12.796744,12.955194,12.7477,12.3289385,11.876224,11.41219,10.789707,9.835234,8.884532,8.114917,7.6018395,7.3075747,7.1981683,7.1076255,7.0170827,6.9265394,6.8661776,6.696409,6.221059,5.6061206,4.991183,4.5007415,4.221567,4.0480266,3.8782585,3.6669915,3.4481792,3.6669915,4.025391,4.5497856,5.1798143,5.753253,5.9117036,5.9682927,5.7117543,5.100589,4.255521,3.6330378,3.1312788,2.8181508,2.71629,2.776652,2.9464202,2.9539654,2.9313297,2.9954643,3.2482302,3.7273536,4.1008434,4.3196554,4.395108,4.395108,4.395108,4.4403796,4.4818783,4.52715,4.640329,4.859141,5.5193505,6.3908267,7.183078,7.537705,7.7942433,7.884786,8.058327,8.296002,8.329956,8.477088,8.714764,9.190115,9.918231,10.770844,11.065109,10.853842,10.31813,9.631512,8.971302,8.43559,7.798016,7.424526,7.281166,6.9265394,6.5002327,6.156924,5.80607,5.560849,5.7079816,6.571913,7.0284004,7.3868,7.752744,8.009283,7.5716586,6.858632,6.1606965,5.726845,5.753253,6.1305156,5.915476,5.80607,6.1342883,6.8661776,7.145352,6.8435416,5.987156,4.9685473,4.515832,4.0517993,3.2784111,2.4974778,1.9542197,1.8297231,1.478869,1.0676528,0.8186596,0.7092535,0.48666862,0.4376245,0.39989826,0.29426476,0.150905,0.0754525,0.08677038,0.10186087,0.124496624,0.21881226,0.48666862,0.7809334,0.69039035,0.5357128,0.452715,0.36594462,0.15845025,0.16222288,0.331991,0.67152727,1.2223305,1.2449663,1.1883769,1.0299267,0.7092535,0.1358145,0.5772116,1.3807807,1.8825399,1.7052265,0.77716076,0.35085413,0.09808825,0.0,0.0,0.0,0.011317875,0.0150905,0.026408374,0.0452715,0.0452715,0.02263575,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.6144292,2.71629,2.7992878,3.1840954,3.7914882,4.1083884,4.217795,4.466788,4.617693,4.478106,3.893349,3.31991,3.108643,3.1840954,3.2859564,2.987919,1.5128226,0.9280658,0.8262049,0.9205205,1.0450171,1.0336993,1.0186088,0.9808825,0.9620194,1.0601076,0.8639311,0.6187105,0.41498876,0.3055826,0.27917424,0.27540162,0.23767537,0.20372175,0.18485862,0.150905,0.15845025,0.13204187,0.1056335,0.09808825,0.120724,0.19240387,0.27917424,0.331991,0.32444575,0.2867195,0.2565385,0.21881226,0.18485862,0.150905,0.124496624,0.150905,0.21881226,0.29803738,0.3734899,0.44139713,0.47535074,0.5696664,0.6790725,0.754525,0.7394345,0.65643674,0.55080324,0.43007925,0.31312788,0.25276586,0.27917424,0.30935526,0.362172,0.45648763,0.59607476,0.66020936,0.7130261,1.1544232,1.9164935,2.4672968,2.987919,3.451952,4.025391,4.5912848,4.749735,4.8855495,5.1647234,5.5797124,5.956975,5.9796104,5.1345425,4.678055,4.293247,3.874486,3.5349495,3.904667,4.032936,3.9273026,3.6594462,3.3764994,2.8634224,2.4559789,2.2183034,2.161714,2.2447119,2.516341,2.8294687,3.0822346,3.1425967,2.8558772,2.4672968,2.2560298,2.6710186,3.4255435,3.5085413,3.187868,2.3993895,1.780679,1.5052774,1.2826926,1.0638802,0.8941121,0.90543,1.0714256,1.237421,1.1846043,1.0601076,0.97333723,0.9922004,1.1129243,1.0676528,1.0072908,0.91674787,0.7582976,0.5017591,0.39989826,0.31312788,0.24899325,0.211267,0.20749438,0.14335975,0.08677038,0.056589376,0.056589376,0.056589376,0.06413463,0.08299775,0.09808825,0.1056335,0.10940613,0.20372175,0.3961256,0.47157812,0.46026024,0.63002837,1.0374719,1.7052265,2.4559789,3.0709167,3.270866,2.4786146,1.9051756,1.7919968,2.214531,3.0407357,3.8858037,4.044254,3.6707642,2.8294687,1.50905,1.3619176,1.267602,1.1695137,1.0110635,0.7130261,0.6790725,0.452715,0.25276586,0.1961765,0.2867195,0.24899325,0.19994913,0.26031113,0.36594462,0.2565385,0.17731337,0.06413463,0.06413463,0.14713238,0.10940613,0.02263575,0.026408374,0.150905,0.7130261,2.3013012,5.873977,4.870459,2.8747404,1.6750455,1.2638294,1.7542707,1.6863633,1.3807807,0.98842776,0.4678055,0.6375736,0.7205714,0.70170826,0.6073926,0.482896,0.39989826,0.33576363,0.27917424,0.1961765,0.03772625,0.02263575,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.03772625,0.06790725,0.1056335,0.14713238,0.08677038,0.049044125,0.026408374,0.02263575,0.033953626,0.018863125,0.02263575,0.033953626,0.0452715,0.041498873,0.0452715,0.06413463,0.10186087,0.181086,0.33953625,0.29426476,0.18863125,0.11317875,0.09808825,0.09808825,0.08299775,0.05281675,0.06790725,0.13958712,0.2263575,0.2565385,0.271629,0.24522063,0.181086,0.13958712,0.16222288,0.23390275,0.35462674,0.4979865,0.63002837,0.47912338,0.45648763,0.6073926,0.87147635,1.0978339,0.8639311,0.6149379,0.43385187,0.32444575,0.21503963,0.15467763,0.116951376,0.09808825,0.10186087,0.11317875,0.16222288,0.21503963,0.18863125,0.090543,0.030181,0.3169005,0.76584285,1.1996948,2.3503454,5.881522,8.314865,4.7421894,1.2940104,0.32444575,0.4074435,0.5093044,0.83752275,1.4901869,2.4672968,3.651901,6.598321,6.398372,4.5912848,2.806833,2.7653341,5.6098933,6.677546,5.956975,3.9876647,1.8561316,1.6071383,2.1805773,3.3878171,4.5950575,4.7233267,3.6179473,2.3918443,1.5354583,1.146878,0.91674787,0.8563859,0.9318384,0.8526133,0.62625575,0.5357128,0.47535074,0.5055317,0.452715,0.30181,0.1961765,0.2263575,0.21881226,0.17731337,0.1056335,0.02263575,0.030181,0.049044125,0.06790725,0.0754525,0.07922512,0.13958712,0.18485862,0.241448,0.331991,0.47157812,0.49421388,0.47157812,0.4074435,0.32067314,0.26031113,0.28294688,0.42630664,0.72811663,1.1581959,1.6071383,1.9240388,2.2862108,2.493705,2.4672968,2.2786655,2.0787163,2.0485353,1.9768555,1.871222,1.9240388,2.4295704,3.006782,3.5424948,3.8707132,3.7763977,3.6707642,3.451952,3.31991,3.3840446,3.6594462,4.0404816,4.4630156,4.715781,4.7006907,4.4403796,4.9987283,5.5985756,6.1342883,6.6813188,7.4811153,7.8621507,7.9828744,8.031919,8.039464,7.888559,7.8017883,8.160188,8.975075,10.140816,11.446144,12.291212,12.815607,13.189097,13.505998,13.777626,13.373956,12.626976,11.98563,11.706455,11.857361,11.981857,11.710228,11.1631975,10.457717,9.737145,9.291975,8.843033,8.401636,7.986647,7.6131573,7.4471617,7.281166,7.1264887,6.964266,6.7567716,6.5643673,6.3455553,6.043745,5.66271,5.221313,4.8025517,4.4894238,4.3422914,4.327201,4.304565,4.395108,4.587512,4.938366,5.4438977,6.043745,6.6322746,6.3229194,5.621211,4.9685473,4.719554,4.0593443,3.7877154,3.7047176,3.731126,3.9008942,3.7877154,3.6292653,3.6443558,3.8367596,3.99521,4.1498876,4.134797,4.115934,4.1197066,4.0517993,4.112161,4.2894745,4.4403796,4.515832,4.5761943,4.798779,5.2590394,5.8136153,6.387054,6.964266,7.5905213,8.126234,8.394091,8.446907,8.563859,8.503497,8.793989,9.129752,9.382519,9.612649,9.778644,9.87296,9.65792,9.144843,8.59404,8.145098,7.6093845,7.1604424,6.8359966,6.549277,6.307829,6.126743,6.017337,5.975838,5.975838,6.560595,7.0812173,7.2962565,7.1679873,6.888813,6.458734,5.96452,5.534441,5.1873593,4.847823,4.8968673,5.0666356,5.481624,6.205968,7.232122,6.9680386,5.938112,4.961002,4.3611546,3.9688015,3.270866,2.6710186,2.2258487,1.9278114,1.7089992,1.8334957,1.6033657,1.3128735,1.026154,0.573439,0.30935526,0.181086,0.094315626,0.033953626,0.026408374,0.041498873,0.060362,0.07922512,0.11317875,0.20749438,0.33576363,0.31312788,0.2263575,0.16976812,0.23013012,0.21881226,0.15467763,0.18485862,0.34330887,0.55080324,0.58475685,0.56589377,0.56212115,0.5319401,0.32067314,0.29049212,0.6488915,1.0336993,1.177059,0.91297525,0.41498876,0.13204187,0.0150905,0.0,0.0,0.003772625,0.003772625,0.0150905,0.033953626,0.033953626,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.595566,2.505023,2.5238862,2.7653341,3.1010978,3.1312788,2.9954643,2.8936033,2.704972,2.425798,2.173032,1.9391292,2.0070364,2.474842,2.938875,2.4786146,1.358145,0.9205205,0.87902164,1.0299267,1.237421,1.2713746,1.1808317,1.0789708,1.0487897,1.1431054,1.2525115,1.2034674,1.0110635,0.724344,0.41498876,0.482896,0.48666862,0.47535074,0.45648763,0.3961256,0.28294688,0.2565385,0.30181,0.38858038,0.48666862,0.5583485,0.6413463,0.6790725,0.6413463,0.5281675,0.44894236,0.3734899,0.32067314,0.29803738,0.31312788,0.35462674,0.45648763,0.513077,0.513077,0.51684964,0.5583485,0.72811663,0.8563859,0.87902164,0.83752275,0.7997965,0.7394345,0.6451189,0.52439487,0.40367088,0.3169005,0.331991,0.40367088,0.4979865,0.56589377,0.7167987,0.91674787,1.3355093,2.022127,2.897376,3.4368613,3.9612563,4.3611546,4.6026025,4.745962,4.485651,4.1197066,3.8405323,3.6783094,3.5047686,3.0860074,2.8822856,2.8634224,2.9539654,3.0256453,3.0935526,3.1765501,3.3048196,3.4368613,3.4481792,3.0558262,2.6408374,2.3314822,2.1881225,2.1994405,1.991946,2.0145817,2.161714,2.263575,2.0636258,1.9127209,2.0560806,2.7389257,3.5387223,3.3425457,2.776652,2.033445,1.4675511,1.1996948,1.1242423,1.0336993,0.8526133,0.7922512,0.87902164,0.9507015,0.8978847,0.80734175,0.7582976,0.77338815,0.80356914,0.73188925,0.7054809,0.66020936,0.56212115,0.4074435,0.33953625,0.27540162,0.21503963,0.1659955,0.1358145,0.09808825,0.060362,0.041498873,0.03772625,0.0452715,0.056589376,0.0754525,0.090543,0.1056335,0.1056335,0.150905,0.2565385,0.32067314,0.38103512,0.59607476,1.0412445,1.6976813,2.293756,2.6634734,2.7389257,2.2748928,1.7957695,1.7391801,2.1881225,2.8407867,2.9916916,3.0746894,2.969056,2.595566,1.9240388,1.6939086,1.4750963,1.267602,1.056335,0.8337501,0.5394854,0.2867195,0.1659955,0.1659955,0.16222288,0.2678564,0.29049212,0.3055826,0.30181,0.17731337,0.116951376,0.1056335,0.21881226,0.3734899,0.3470815,0.23767537,0.23390275,0.271629,0.8186596,2.8634224,7.624475,6.851087,5.119452,4.447925,4.2706113,2.203213,1.4222796,1.177059,0.91674787,0.29426476,0.6451189,0.7167987,0.58475685,0.40367088,0.422534,0.35839936,0.29049212,0.18485862,0.06790725,0.0,0.0,0.033953626,0.033953626,0.0,0.0,0.0,0.02263575,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.011317875,0.003772625,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.0,0.003772625,0.02263575,0.0452715,0.071679875,0.120724,0.08677038,0.060362,0.056589376,0.06413463,0.049044125,0.0150905,0.011317875,0.026408374,0.049044125,0.056589376,0.071679875,0.0754525,0.08299775,0.10940613,0.16976812,0.16222288,0.23013012,0.28294688,0.271629,0.18863125,0.09808825,0.090543,0.15845025,0.27917424,0.4074435,0.29803738,0.241448,0.21881226,0.2263575,0.26408374,0.27540162,0.29426476,0.3470815,0.43007925,0.5319401,0.46026024,0.4640329,0.5772116,0.7582976,0.8941121,0.9318384,1.1732863,1.2185578,0.90543,0.33953625,0.18485862,0.124496624,0.09808825,0.090543,0.094315626,0.150905,0.21881226,0.23013012,0.15845025,0.049044125,0.10186087,0.45648763,0.9695646,1.7693611,3.2482302,6.349328,5.036454,2.2786655,0.23013012,0.211267,0.29049212,0.5470306,0.9997456,1.6524098,2.516341,4.1762958,4.4818783,3.5877664,2.4672968,2.9086938,5.100589,5.149633,4.3007927,3.2067313,1.9504471,1.3656902,1.6373192,2.5389767,3.5575855,3.8858037,3.3727267,2.4107075,1.6146835,1.2449663,1.1846043,0.9620194,0.8601585,0.7394345,0.5772116,0.47157812,0.4979865,0.5394854,0.47912338,0.331991,0.24899325,0.241448,0.20749438,0.17731337,0.13958712,0.041498873,0.026408374,0.03772625,0.056589376,0.0754525,0.08677038,0.1358145,0.19240387,0.31312788,0.52062225,0.7997965,1.146878,1.297783,1.20724,0.935611,0.63002837,0.4979865,0.4979865,0.6111652,0.7997965,1.026154,1.3958713,1.8334957,2.1805773,2.3163917,2.1654868,1.9202662,1.7882242,1.7127718,1.7089992,1.8523588,2.4371157,3.0935526,3.561358,3.682082,3.3651814,3.127506,2.9766011,3.0369632,3.3576362,3.904667,4.5422406,5.1269975,5.2552667,4.859141,4.195159,4.3686996,4.9685473,5.674028,6.4021444,7.322665,8.469543,8.7751255,8.635539,8.3525915,8.099826,8.190369,8.718536,9.58624,10.559577,11.268831,11.646093,12.0233555,12.540206,13.13628,13.539951,13.026875,12.00072,11.012292,10.487898,10.684074,11.09529,11.140562,10.774617,10.133271,9.522105,9.22784,8.971302,8.631766,8.160188,7.5792036,7.220804,7.183078,7.2472124,7.273621,7.1793056,6.9227667,6.7341356,6.5568223,6.3455553,6.0512905,5.828706,5.5759397,5.372218,5.2175403,5.0666356,4.9647746,4.9534564,5.0477724,5.311856,5.824933,5.926794,5.3382645,4.7044635,4.3913355,4.508287,4.3121104,4.5912848,4.7535076,4.568649,4.172523,3.9650288,3.9348478,3.9876647,4.0291634,3.942393,3.9876647,3.9574835,3.9273026,3.9122121,3.8858037,4.1197066,4.357382,4.5460134,4.666737,4.745962,5.0515447,5.5570765,6.2021956,6.8850408,7.4509344,7.564113,7.605612,7.5490227,7.488661,7.624475,7.914967,8.669493,9.352338,9.665465,9.57115,9.171251,8.669493,8.099826,7.5226145,7.0359454,6.688864,6.258785,5.8966126,5.66271,5.511805,5.3609,5.311856,5.3571277,5.4778514,5.666483,6.1229706,6.488915,6.579458,6.3455553,5.855114,5.4288073,5.1798143,5.081726,5.05909,4.9987283,5.070408,5.2590394,5.5570765,5.87775,6.0701537,5.617439,4.98741,4.29702,3.651901,3.180323,2.5389767,1.8976303,1.659955,1.8334957,2.0372176,2.0296721,1.8749946,1.569412,1.1053791,0.47535074,0.20372175,0.07922512,0.026408374,0.011317875,0.02263575,0.030181,0.03772625,0.0452715,0.05281675,0.071679875,0.10186087,0.094315626,0.06413463,0.041498873,0.07922512,0.13958712,0.16976812,0.17731337,0.1659955,0.181086,0.20372175,0.19994913,0.211267,0.22258487,0.17354076,0.10940613,0.21503963,0.36594462,0.44894236,0.3961256,0.18485862,0.060362,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.02263575,0.02263575,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.9615107,2.6936543,2.757789,2.886058,2.9426475,2.9426475,3.1576872,2.9803739,2.516341,1.9504471,1.5430037,1.81086,1.9127209,2.1390784,2.3428001,1.9051756,1.3770081,1.1657411,1.1883769,1.3430545,1.4977322,1.5505489,1.4335974,1.2411937,1.0827434,1.0638802,1.2449663,1.3128735,1.237421,1.0412445,0.7922512,0.8865669,0.8903395,0.7997965,0.66020936,0.55080324,0.47912338,0.482896,0.5394854,0.633801,0.7469798,0.94692886,1.0374719,1.0714256,1.0940613,1.1242423,0.95824677,0.76584285,0.5885295,0.47912338,0.49421388,0.52439487,0.6111652,0.66775465,0.70170826,0.79602385,0.8526133,0.94315624,0.9242931,0.8186596,0.7997965,0.84129536,0.84129536,0.79602385,0.73566186,0.7507524,0.8299775,0.7167987,0.62625575,0.63002837,0.6752999,0.98842776,1.4637785,2.323937,3.7537618,5.9230213,6.1342883,5.621211,4.67051,3.9008942,4.2819295,4.3083377,3.8858037,3.138824,2.2975287,1.7014539,1.5165952,1.5165952,1.7618159,2.142851,2.3956168,2.2673476,2.1579416,2.2673476,2.5502944,2.727608,2.505023,2.2975287,2.293756,2.5012503,2.7615614,2.2711203,2.0145817,1.8863125,1.7693611,1.5316857,1.569412,1.8523588,2.4786146,3.199186,3.440634,2.625747,1.8334957,1.3128735,1.1317875,1.20724,1.146878,0.9205205,0.7809334,0.754525,0.6790725,0.6526641,0.6790725,0.66775465,0.5998474,0.5281675,0.42630664,0.42630664,0.42630664,0.392353,0.32821837,0.27540162,0.23390275,0.18485862,0.124496624,0.056589376,0.041498873,0.030181,0.030181,0.041498873,0.05281675,0.049044125,0.049044125,0.060362,0.07922512,0.08299775,0.1056335,0.15467763,0.25276586,0.44894236,0.80734175,1.3543724,2.033445,2.372981,2.293756,2.123988,1.8259505,1.4335974,1.4411428,1.8863125,2.335255,2.123988,2.263575,2.425798,2.4295704,2.2409391,1.7655885,1.4600059,1.2336484,1.026154,0.80356914,0.41876137,0.181086,0.09808825,0.10940613,0.11317875,0.33953625,0.4678055,0.3961256,0.22258487,0.21503963,0.181086,0.15467763,0.33576363,0.6790725,0.86770374,0.8262049,0.5357128,0.4678055,1.1355602,3.1010978,7.164215,7.5226145,7.405663,7.9753294,8.318638,4.1612053,2.1315331,1.2525115,0.875249,0.694163,0.66775465,0.513077,0.29049212,0.120724,0.19994913,0.18485862,0.15845025,0.120724,0.06790725,0.0,0.0,0.033953626,0.033953626,0.0,0.0,0.0,0.02263575,0.0452715,0.060362,0.060362,0.011317875,0.03772625,0.05281675,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.011317875,0.011317875,0.003772625,0.0,0.0,0.003772625,0.011317875,0.018863125,0.030181,0.056589376,0.05281675,0.049044125,0.060362,0.06790725,0.041498873,0.0150905,0.018863125,0.03772625,0.060362,0.06413463,0.0754525,0.0754525,0.08299775,0.10186087,0.120724,0.13204187,0.2565385,0.34330887,0.331991,0.2263575,0.11317875,0.12826926,0.23390275,0.38858038,0.543258,0.392353,0.2565385,0.19240387,0.20372175,0.24899325,0.27540162,0.32444575,0.41121614,0.5319401,0.67152727,0.7696155,0.7469798,0.8224323,0.9997456,1.0940613,0.97710985,1.9466745,2.6332922,2.3126192,0.91297525,0.34330887,0.1659955,0.1358145,0.116951376,0.08299775,0.11317875,0.15845025,0.18863125,0.1659955,0.056589376,0.033953626,0.28294688,0.845068,1.539231,1.9768555,4.4101987,6.1833324,4.817642,1.3166461,0.1659955,0.12826926,0.25276586,0.55457586,1.0186088,1.5731846,1.9391292,2.2107582,2.0900342,2.0070364,3.1237335,7.413208,7.0887623,4.859141,2.6597006,1.6524098,1.0714256,1.327964,2.2598023,3.5953116,4.927048,4.3422914,3.0369632,1.9693103,1.5316857,1.5241405,1.2336484,0.875249,0.63002837,0.52439487,0.422534,0.44516975,0.4640329,0.422534,0.3470815,0.31312788,0.29049212,0.211267,0.14335975,0.10186087,0.03772625,0.030181,0.041498873,0.060362,0.090543,0.124496624,0.181086,0.23767537,0.3470815,0.52439487,0.77338815,1.2449663,1.5203679,1.5015048,1.2562841,1.0148361,0.7922512,0.56212115,0.452715,0.48666862,0.58475685,0.87902164,1.2638294,1.659955,1.9504471,1.9994912,1.8749946,2.052308,2.1503963,2.0447628,1.8599042,2.2786655,2.7238352,3.0331905,3.138824,3.0369632,2.8143783,2.7200627,2.837014,3.2142766,3.8405323,4.3875628,4.881777,5.062863,4.878004,4.478106,4.6290107,5.20245,5.938112,6.6322746,7.1302614,7.9828744,8.284684,8.194141,7.9300575,7.7942433,8.009283,8.529905,9.205205,9.827688,10.125726,10.148361,10.431308,10.978339,11.646093,12.162943,11.887542,11.133017,10.287949,9.695646,9.676784,10.050273,10.227587,10.091772,9.733373,9.446653,9.310839,9.163706,8.801534,8.216777,7.594294,7.254758,7.394345,7.594294,7.6810646,7.7225633,7.665974,7.6093845,7.5905213,7.598067,7.541477,7.4773426,7.141579,6.6624556,6.119198,5.5495315,5.2854476,5.0779533,4.9421387,4.9421387,5.2099953,5.2137675,4.8063245,4.293247,4.055572,4.52715,4.5460134,4.7421894,4.8138695,4.606375,4.112161,3.9989824,4.112161,4.2102494,4.164978,3.9348478,3.8178966,3.8443048,3.874486,3.874486,3.9159849,4.2781568,4.5761943,4.8402777,5.0854983,5.330719,5.8437963,6.3153744,6.8171334,7.3188925,7.7037,7.4207535,7.1038527,6.8661776,6.790725,6.9227667,7.5527954,8.477088,9.137298,9.273112,8.922258,8.29223,7.6131573,6.903904,6.2399216,5.745708,5.4250345,5.070408,4.7874613,4.6214657,4.561104,4.5988297,4.7044635,4.8855495,5.160951,5.5495315,5.8928404,5.9230213,5.723072,5.3684454,4.9232755,5.081726,5.2892203,5.462761,5.5193505,5.3759904,5.4174895,5.511805,5.6098933,5.523123,4.9157305,4.3121104,3.9461658,3.5085413,2.9728284,2.6068838,2.1654868,1.4449154,1.0978339,1.2751472,1.6146835,1.6939086,1.5882751,1.3128735,0.8978847,0.3772625,0.16222288,0.071679875,0.041498873,0.03772625,0.03772625,0.026408374,0.02263575,0.018863125,0.018863125,0.02263575,0.018863125,0.0150905,0.011317875,0.003772625,0.0,0.049044125,0.124496624,0.15467763,0.13204187,0.094315626,0.08677038,0.071679875,0.06790725,0.08299775,0.08299775,0.0452715,0.03772625,0.03772625,0.033953626,0.02263575,0.018863125,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.783943,3.4066803,3.3236825,3.150142,2.8747404,2.867195,3.4217708,3.3878171,3.0030096,2.4408884,1.8259505,2.3767538,2.444661,2.2220762,1.9164935,1.7542707,1.5882751,1.5354583,1.5769572,1.6637276,1.7127718,1.6675003,1.5882751,1.4335974,1.2298758,1.0978339,1.116697,1.1317875,1.1581959,1.2147852,1.2902378,1.3204187,1.2751472,1.1053791,0.875249,0.7507524,0.8224323,0.845068,0.83752275,0.8224323,0.84884065,1.1581959,1.2789198,1.3430545,1.4637785,1.7316349,1.5618668,1.2902378,0.995973,0.76584285,0.73566186,0.69039035,0.7432071,0.845068,0.98842776,1.2110126,1.2449663,1.1544232,0.9507015,0.73566186,0.7205714,0.784706,0.79602385,0.7696155,0.784706,1.0072908,1.3694628,1.177059,0.9393836,0.87902164,0.935611,1.3091009,1.9806281,3.361409,5.6551647,8.846806,8.669493,7.0963078,4.9119577,3.259548,3.6179473,4.0517993,3.9650288,3.2935016,2.2899833,1.5316857,1.1506506,1.0714256,1.1393328,1.237421,1.297783,1.2713746,1.1280149,1.2110126,1.4901869,1.5769572,1.4600059,1.5128226,1.8749946,2.4672968,2.9803739,2.674791,2.4899325,2.3163917,2.1088974,1.8787673,1.9994912,2.0070364,2.1466236,2.6031113,3.4972234,2.4786146,1.7014539,1.3053282,1.2525115,1.3468271,1.1883769,0.965792,0.8262049,0.754525,0.59230214,0.543258,0.6375736,0.6187105,0.452715,0.35462674,0.31312788,0.35462674,0.3734899,0.33576363,0.29426476,0.23013012,0.19240387,0.150905,0.09808825,0.041498873,0.033953626,0.026408374,0.033953626,0.05281675,0.06413463,0.05281675,0.03772625,0.033953626,0.041498873,0.056589376,0.10940613,0.18863125,0.3169005,0.56589377,1.0374719,1.7240896,2.493705,2.674791,2.2409391,1.8070874,1.4071891,0.9922004,1.0186088,1.4675511,1.8297231,1.780679,1.9429018,2.1051247,2.1390784,2.003264,1.3241913,1.0412445,0.91297525,0.754525,0.45648763,0.23390275,0.10186087,0.0452715,0.05281675,0.09808825,0.392353,0.60362,0.4979865,0.23013012,0.33576363,0.331991,0.23767537,0.38480774,0.7997965,1.1996948,1.3015556,0.8111144,0.9242931,2.0372176,3.7462165,6.096562,7.805561,9.371201,10.695392,11.0613365,6.63982,3.5802212,1.6863633,0.875249,1.1959221,0.68661773,0.3470815,0.1358145,0.0452715,0.08677038,0.13958712,0.16222288,0.181086,0.15467763,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049044125,0.120724,0.120724,0.02263575,0.071679875,0.1056335,0.06790725,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.018863125,0.00754525,0.00754525,0.030181,0.030181,0.033953626,0.03772625,0.030181,0.026408374,0.026408374,0.026408374,0.026408374,0.0150905,0.011317875,0.041498873,0.06413463,0.071679875,0.05281675,0.03772625,0.030181,0.0452715,0.090543,0.150905,0.18863125,0.23013012,0.2565385,0.26031113,0.23390275,0.21881226,0.271629,0.36594462,0.47912338,0.58098423,0.49421388,0.30181,0.16976812,0.14335975,0.14713238,0.1961765,0.29049212,0.43007925,0.6187105,0.8337501,1.0940613,1.0827434,1.1393328,1.327964,1.4524606,0.9280658,2.3578906,3.8367596,3.9574835,1.7957695,0.66775465,0.30935526,0.23767537,0.19240387,0.1056335,0.090543,0.090543,0.10940613,0.11317875,0.0452715,0.033953626,0.12826926,0.5394854,1.2223305,1.901403,4.919503,8.254503,7.484888,3.4972234,2.505023,1.1317875,0.33953625,0.150905,0.41121614,0.7507524,1.1053791,1.1393328,1.1431054,1.5430037,2.8785129,9.5183325,9.699419,6.417235,2.655928,1.3807807,0.94692886,1.2789198,2.3993895,4.1800685,6.356873,5.6325293,3.8367596,2.3880715,1.7995421,1.6373192,1.4411428,1.0072908,0.6828451,0.55080324,0.42630664,0.38858038,0.41498876,0.452715,0.44139713,0.35839936,0.34330887,0.2263575,0.11317875,0.049044125,0.0150905,0.026408374,0.033953626,0.060362,0.10940613,0.1659955,0.2565385,0.3169005,0.362172,0.41121614,0.4979865,0.7696155,1.0299267,1.1242423,1.086516,1.1204696,0.91674787,0.52439487,0.2867195,0.29803738,0.41121614,0.68661773,1.0714256,1.50905,1.9051756,2.1466236,2.1088974,2.6332922,2.8747404,2.546522,1.9089483,2.0108092,2.071171,2.173032,2.3654358,2.6446102,2.6144292,2.5917933,2.674791,2.969056,3.591539,3.832987,4.1008434,4.466788,4.8365054,4.9421387,5.2665844,5.80607,6.485142,7.069899,7.183078,6.9944468,7.0472636,7.073672,7.0585814,7.201941,7.4773426,7.911195,8.29223,8.563859,8.778898,8.82417,9.239159,9.80128,10.378491,10.921749,10.974566,10.702937,10.231359,9.7069645,9.307066,9.34102,9.352338,9.273112,9.156161,9.156161,9.144843,8.99771,8.548768,7.9262853,7.5565677,7.5527954,7.8923316,8.13378,8.156415,8.156415,8.326183,8.401636,8.518587,8.707218,8.888305,8.880759,8.397863,7.647111,6.760544,5.794752,5.4740787,5.142088,4.889322,4.7535076,4.7044635,5.040227,5.0741806,4.610148,4.0782075,4.5422406,4.5007415,4.214022,4.0103,3.9763467,3.9348478,3.9914372,4.146115,4.2819295,4.315883,4.191386,3.9348478,3.9084394,3.9348478,3.9612563,4.08198,4.485651,4.82896,5.160951,5.5306683,5.9909286,6.6850915,6.94163,6.9869013,6.9982195,7.115171,6.9454026,6.779407,6.670001,6.651138,6.760544,7.3490734,7.9489207,8.171506,7.9300575,7.4509344,7.0246277,6.700182,6.187105,5.523123,5.040227,4.696918,4.4139714,4.1989317,4.06689,4.06689,4.376245,4.5988297,4.847823,5.168496,5.515578,5.670255,5.402399,4.9459114,4.5196047,4.327201,5.1798143,5.772116,6.047518,5.9607477,5.485397,5.3986263,5.3948536,5.3646727,5.1043615,4.2894745,3.5500402,3.0181,2.704972,2.5616124,2.4710693,2.2183034,1.5052774,0.94315624,0.7696155,0.8601585,1.1619685,1.0186088,0.76584285,0.55457586,0.35085413,0.21503963,0.14713238,0.11317875,0.090543,0.071679875,0.033953626,0.0150905,0.003772625,0.003772625,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.003772625,0.011317875,0.030181,0.07922512,0.13958712,0.14335975,0.124496624,0.10186087,0.10940613,0.13958712,0.12826926,0.056589376,0.018863125,0.003772625,0.00754525,0.026408374,0.033953626,0.030181,0.02263575,0.011317875,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,5.1269975,4.5535583,4.0706625,3.8405323,3.8556228,3.9688015,3.4179983,2.7879698,2.3390274,2.082489,1.7391801,1.5203679,1.8485862,2.033445,1.901403,1.8146327,1.7165444,1.6675003,1.6033657,1.5430037,1.5430037,1.4675511,1.5882751,1.6788181,1.599593,1.2826926,1.5241405,1.6222287,1.599593,1.50905,1.448688,1.3996439,1.3807807,1.4147344,1.4939595,1.5580941,1.5203679,1.4373702,1.3166461,1.177059,1.0676528,1.056335,1.1544232,1.2336484,1.2713746,1.3430545,1.5015048,1.5128226,1.4713237,1.4071891,1.297783,1.0789708,1.1581959,1.3015556,1.358145,1.297783,1.1242423,0.9922004,0.8639311,0.7205714,0.55080324,0.52439487,0.5357128,0.543258,0.55457586,0.6413463,0.70170826,0.7997965,0.9695646,1.1431054,1.1280149,1.1883769,1.6524098,2.6068838,3.9876647,5.5985756,6.907676,6.8397694,5.9418845,4.6290107,3.187868,2.384299,1.5316857,1.1053791,1.2525115,1.7995421,1.5580941,1.3505998,1.1732863,1.0299267,0.9318384,0.8563859,0.8111144,0.8224323,0.88279426,0.9318384,1.0299267,1.1619685,1.1695137,1.0751982,1.0978339,1.1846043,1.2525115,1.3656902,1.5882751,1.9542197,2.5993385,2.4974778,2.4107075,2.6672459,3.1425967,2.1051247,1.5807298,1.3732355,1.3091009,1.237421,1.0902886,0.94315624,0.814887,0.7130261,0.6413463,0.59230214,0.5357128,0.422534,0.32821837,0.42630664,0.573439,0.6752999,0.6375736,0.48666862,0.36594462,0.29426476,0.23767537,0.18485862,0.124496624,0.0754525,0.041498873,0.041498873,0.05281675,0.06413463,0.0754525,0.11317875,0.1056335,0.07922512,0.06790725,0.090543,0.12826926,0.19994913,0.31312788,0.4640329,0.67152727,1.2223305,1.8146327,2.04099,1.8448136,1.5241405,1.1846043,0.84129536,0.95824677,1.4750963,1.8146327,1.8636768,1.7014539,1.539231,1.4411428,1.3430545,0.9280658,0.7054809,0.52062225,0.29803738,0.030181,0.030181,0.02263575,0.0150905,0.011317875,0.0,0.29426476,0.47535074,0.47157812,0.33576363,0.27540162,0.35839936,0.49044126,0.422534,0.22258487,0.26031113,0.5281675,0.9808825,2.0787163,3.8103511,5.6778007,7.605612,9.514561,10.642575,10.623712,9.476834,6.156924,3.5877664,1.7542707,0.7205714,0.6111652,0.6111652,0.49044126,0.32067314,0.23013012,0.42630664,0.5017591,0.4640329,0.3055826,0.09808825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.041498873,0.049044125,0.033953626,0.0452715,0.094315626,0.09808825,0.10940613,0.13958712,0.150905,0.07922512,0.033953626,0.0150905,0.0150905,0.0150905,0.003772625,0.026408374,0.056589376,0.0754525,0.0754525,0.05281675,0.026408374,0.033953626,0.06790725,0.090543,0.1659955,0.23767537,0.26408374,0.271629,0.38103512,0.55080324,0.7130261,0.7507524,0.663982,0.58098423,0.49421388,0.3169005,0.1961765,0.18485862,0.24522063,0.3055826,0.31312788,0.31312788,0.331991,0.38103512,0.6149379,0.76207024,0.86770374,0.97710985,1.1581959,1.1242423,1.6637276,3.1048703,4.2404304,2.335255,1.1393328,0.63002837,0.40367088,0.25276586,0.1659955,0.13204187,0.11317875,0.1056335,0.094315626,0.0452715,0.033953626,0.08677038,0.52062225,1.6561824,3.8292143,10.336992,9.042982,5.7419353,5.2288585,11.306557,5.4212623,1.5807298,0.018863125,0.116951376,0.3961256,0.56589377,0.6187105,0.59607476,0.97333723,2.6710186,4.3686996,5.0213637,4.508287,3.2482302,2.2107582,1.3468271,1.1091517,1.5807298,2.6106565,3.8292143,4.3196554,3.451952,2.3277097,1.5015048,0.97710985,0.9280658,0.87147635,0.784706,0.66020936,0.48666862,0.48666862,0.5696664,0.694163,0.69793564,0.32067314,0.16222288,0.094315626,0.08677038,0.10186087,0.0754525,0.041498873,0.011317875,0.041498873,0.12826926,0.21503963,0.32444575,0.44139713,0.52062225,0.5583485,0.59607476,0.6451189,0.83752275,0.97333723,0.9507015,0.77716076,0.59607476,0.44894236,0.35839936,0.33953625,0.41121614,0.754525,1.2147852,1.7655885,2.2786655,2.546522,2.5616124,2.444661,2.2447119,2.0183544,1.8448136,1.6750455,1.5505489,1.5807298,1.7655885,1.9844007,2.2296214,2.4069347,2.7992878,3.4444065,4.164978,4.38379,4.715781,4.991183,5.0854983,4.927048,4.9534564,5.3080835,5.836251,6.462507,7.17176,6.964266,6.590776,6.2021956,6.0286546,6.40969,6.9567204,7.699928,8.13378,8.216777,8.375228,8.888305,9.688101,10.450171,11.031156,11.457462,11.521597,11.370691,11.083972,10.710483,10.284176,10.016319,9.654147,9.273112,8.91094,8.605357,8.2507305,7.7414265,7.1566696,6.7379084,6.8963585,7.4207535,8.039464,8.582722,8.816625,8.439363,8.058327,7.7716074,7.6508837,7.7150183,7.9338303,8.09228,7.9300575,7.4811153,6.820906,6.089017,5.8437963,5.5193505,5.383536,5.402399,5.2175403,5.0854983,5.0515447,4.7346444,4.0404816,3.1727777,3.5160866,3.7462165,3.7348988,3.5689032,3.5538127,3.640583,3.7801702,3.9084394,4.044254,4.2894745,4.323428,4.0970707,3.92353,3.9725742,4.2404304,4.6931453,4.9534564,5.142088,5.3910813,5.8437963,6.379509,6.349328,6.1116524,5.8928404,5.783434,6.013564,6.156924,6.2361493,6.2851934,6.3342376,6.356873,6.428553,6.530414,6.5832305,6.4247804,6.058836,5.5268955,4.9044123,4.3422914,4.074435,3.8292143,3.7047176,3.7160356,3.8480775,4.044254,4.4705606,4.5950575,4.6516466,4.6856003,4.561104,4.4177437,4.2781568,4.2102494,4.2781568,4.5460134,4.6554193,4.7950063,4.9044123,4.9949555,5.142088,5.20245,5.0439997,4.6856003,4.191386,3.6934,3.1048703,2.6672459,2.595566,2.776652,2.776652,2.5314314,2.0145817,1.7089992,1.7278622,1.7995421,1.4939595,1.026154,0.6451189,0.44894236,0.35085413,0.362172,0.30181,0.23013012,0.181086,0.1659955,0.08299775,0.041498873,0.02263575,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.026408374,0.0150905,0.0150905,0.0150905,0.0150905,0.02263575,0.0452715,0.094315626,0.16976812,0.18863125,0.13958712,0.090543,0.030181,0.0150905,0.0150905,0.026408374,0.0754525,0.11317875,0.094315626,0.071679875,0.049044125,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.011317875,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.0286546,5.670255,5.198677,4.6554193,4.0782075,3.5047686,3.2746384,2.9539654,2.6446102,2.3578906,1.9957186,2.2560298,2.3314822,2.1088974,1.780679,1.841041,1.7240896,1.5505489,1.3920987,1.3053282,1.3355093,1.3694628,1.388326,1.4071891,1.3996439,1.3166461,1.297783,1.3091009,1.3091009,1.2902378,1.2789198,1.5015048,1.6825907,1.780679,1.7844516,1.690136,1.5467763,1.4449154,1.3958713,1.3619176,1.2525115,1.4034165,1.5505489,1.5920477,1.5279131,1.4637785,1.4864142,1.4637785,1.5430037,1.690136,1.6863633,1.4298248,1.1808317,1.0751982,1.0978339,1.0638802,0.875249,0.7922512,0.7922512,0.8262049,0.84129536,0.58475685,0.5885295,0.73188925,0.90920264,1.0450171,1.0072908,1.0374719,1.1695137,1.3091009,1.2261031,1.4260522,1.9240388,2.41448,2.927557,3.8178966,4.6856003,4.647874,3.8971217,2.8219235,2.003264,1.8749946,1.7995421,1.780679,1.8146327,1.8863125,1.9051756,1.7769064,1.539231,1.2034674,0.784706,0.7092535,0.7092535,0.7809334,0.88279426,0.94315624,0.9997456,1.0525624,1.0412445,0.995973,1.0487897,1.1053791,1.1355602,1.2713746,1.4864142,1.599593,1.720317,1.7014539,1.7316349,1.841041,1.9353566,1.5430037,1.2525115,1.0827434,1.026154,1.0412445,1.237421,1.297783,1.2261031,1.0148361,0.6790725,0.63002837,0.56212115,0.41876137,0.26031113,0.2678564,0.3470815,0.4376245,0.543258,0.62625575,0.62248313,0.5998474,0.5319401,0.46026024,0.3772625,0.26031113,0.08677038,0.03772625,0.041498873,0.056589376,0.08677038,0.094315626,0.094315626,0.090543,0.09808825,0.150905,0.16976812,0.21503963,0.29049212,0.40367088,0.573439,1.056335,1.4637785,1.5543215,1.3053282,0.9280658,0.86770374,1.0601076,1.2147852,1.2940104,1.4977322,1.6637276,1.4864142,1.1996948,0.9393836,0.73188925,0.58098423,0.43007925,0.2867195,0.150905,0.018863125,0.018863125,0.00754525,0.003772625,0.14713238,0.73188925,0.6149379,0.52062225,0.5093044,0.5583485,0.55457586,0.62248313,0.66020936,0.47912338,0.21503963,0.32067314,0.5093044,0.62248313,2.2899833,5.1873593,7.0057645,7.383027,8.567632,8.899622,7.884786,6.1795597,4.938366,3.270866,1.7467253,0.754525,0.48666862,0.362172,0.24899325,0.15467763,0.1056335,0.1358145,0.1961765,0.24522063,0.24899325,0.20372175,0.1358145,0.1056335,0.1056335,0.1358145,0.16222288,0.120724,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0452715,0.0452715,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.02263575,0.02263575,0.033953626,0.033953626,0.03772625,0.060362,0.094315626,0.116951376,0.181086,0.18863125,0.16222288,0.11317875,0.06413463,0.033953626,0.030181,0.030181,0.026408374,0.026408374,0.033953626,0.0452715,0.07922512,0.13204187,0.17731337,0.19994913,0.23390275,0.22258487,0.181086,0.17354076,0.23767537,0.29803738,0.33953625,0.36971724,0.422534,0.3961256,0.31312788,0.23767537,0.2263575,0.3169005,0.30935526,0.271629,0.211267,0.17731337,0.23390275,0.45648763,0.73566186,0.845068,0.84129536,1.0638802,1.1996948,1.0902886,2.0598533,3.6783094,3.7386713,1.6033657,0.62625575,0.2678564,0.1659955,0.120724,0.120724,0.12826926,0.13204187,0.120724,0.071679875,0.056589376,0.27917424,0.88279426,1.690136,2.1805773,3.199186,2.7313805,1.9844007,2.5993385,6.670001,5.1798143,2.0673985,0.1659955,0.06790725,0.150905,0.2565385,0.362172,0.49421388,0.9507015,2.3163917,4.4705606,4.346064,3.482133,2.6823363,2.0183544,1.5128226,1.418507,1.7240896,2.3767538,3.2935016,3.6934,3.5575855,3.1048703,2.4333432,1.539231,1.2826926,1.2562841,1.2147852,1.0751982,0.9016574,0.72811663,0.56212115,0.5055317,0.52439487,0.41876137,0.2678564,0.15467763,0.10186087,0.11317875,0.1358145,0.150905,0.1056335,0.0754525,0.1056335,0.19994913,0.241448,0.29426476,0.35839936,0.4376245,0.5357128,0.63002837,0.7884786,0.94692886,1.0412445,0.9997456,0.94315624,0.8337501,0.73188925,0.6790725,0.7054809,0.8903395,1.2600567,1.8938577,2.6672459,3.2670932,3.0445085,2.6144292,2.1051247,1.6788181,1.5165952,1.6184561,1.6561824,1.7165444,1.8448136,2.0447628,2.3465726,2.7992878,3.3651814,3.9197574,4.2404304,4.3800178,4.447925,4.4705606,4.4139714,4.195159,4.2291126,4.727099,5.4778514,6.3116016,7.0849895,7.2887115,6.990674,6.515323,6.168242,6.2135134,6.802043,7.3717093,7.7678347,7.9828744,8.122461,8.495952,9.148616,9.940866,10.665211,11.031156,11.102836,11.027383,10.955703,10.887795,10.676529,10.650121,10.593531,10.393582,10.0276375,9.559832,8.714764,7.726336,6.9152217,6.515323,6.651138,7.062354,7.435844,7.6282477,7.6018395,7.435844,7.4697976,7.2057137,7.0170827,7.039718,7.141579,6.937857,6.964266,7.2660756,7.6320205,7.6018395,7.6320205,7.5490227,7.1906233,6.688864,6.488915,6.537959,6.096562,5.409944,4.6252384,3.8103511,3.3878171,3.1463692,3.048281,3.0860074,3.2520027,3.3651814,3.4179983,3.4444065,3.519859,3.7613072,3.9461658,3.9725742,3.9914372,4.123479,4.447925,4.617693,4.6026025,4.376245,4.1272516,4.255521,4.5422406,4.3422914,4.1800685,4.214022,4.2819295,4.4630156,4.6742826,4.908185,5.13077,5.247721,5.2326307,5.20245,5.172269,5.0968165,4.8968673,4.4743333,4.236658,3.9499383,3.62172,3.4896781,3.5651307,3.5274043,3.500996,3.531177,3.5802212,3.7235808,3.874486,3.99521,4.085753,4.146115,4.3121104,4.349837,4.466788,4.6856003,4.8138695,4.798779,4.8365054,4.8365054,4.7120085,4.4101987,4.1272516,3.7386713,3.199186,2.5691576,2.0070364,1.8334957,1.7240896,1.7014539,1.7618159,1.8485862,1.750498,1.3128735,0.90920264,0.73566186,0.7997965,0.7205714,0.4678055,0.30935526,0.27917424,0.181086,0.16222288,0.16222288,0.16222288,0.15467763,0.13204187,0.1056335,0.08677038,0.06413463,0.033953626,0.0150905,0.003772625,0.011317875,0.011317875,0.003772625,0.003772625,0.003772625,0.003772625,0.00754525,0.0150905,0.02263575,0.030181,0.0452715,0.056589376,0.05281675,0.041498873,0.041498873,0.033953626,0.033953626,0.03772625,0.026408374,0.026408374,0.026408374,0.026408374,0.02263575,0.011317875,0.003772625,0.0,0.00754525,0.011317875,0.0,0.011317875,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,7.1000805,6.8661776,6.3116016,5.5382137,4.738417,4.183841,4.014073,3.6971724,3.3651814,3.059599,2.7389257,2.4484336,2.252257,2.003264,1.720317,1.5543215,1.5618668,1.4562333,1.327964,1.2751472,1.3996439,1.4260522,1.418507,1.4562333,1.5203679,1.5015048,1.4373702,1.4260522,1.4939595,1.6146835,1.6939086,1.8900851,1.9768555,1.961765,1.8749946,1.7316349,1.629774,1.5052774,1.4524606,1.4901869,1.5618668,1.6184561,1.7919968,1.9089483,1.8372684,1.4675511,1.418507,1.358145,1.3128735,1.3430545,1.5203679,1.4562333,1.3355093,1.2864652,1.2713746,1.0714256,0.8186596,0.7507524,0.76207024,0.77716076,0.77716076,0.67152727,0.8224323,1.0827434,1.3468271,1.5279131,1.1732863,1.146878,1.2600567,1.4034165,1.5165952,1.7693611,1.9051756,1.7919968,1.629774,1.9429018,2.305074,2.4408884,2.2107582,1.8372684,1.9089483,2.1956677,2.3503454,2.4597516,2.5389767,2.5201135,2.4295704,2.2409391,1.9164935,1.4750963,1.0035182,0.98842776,1.0186088,1.0676528,1.1016065,1.0751982,1.0714256,1.0902886,1.0940613,1.0714256,1.0374719,1.0940613,1.1732863,1.3317367,1.5241405,1.6033657,1.6712729,1.750498,1.7127718,1.5430037,1.3656902,1.1355602,0.94692886,0.8563859,0.8526133,0.8526133,0.8186596,0.8299775,0.8262049,0.7809334,0.68661773,0.6526641,0.573439,0.43385187,0.30181,0.31312788,0.26408374,0.241448,0.27917424,0.362172,0.4376245,0.44139713,0.422534,0.3961256,0.35085413,0.26031113,0.13204187,0.06790725,0.05281675,0.056589376,0.06413463,0.06413463,0.060362,0.060362,0.0754525,0.120724,0.14713238,0.18863125,0.25276586,0.36971724,0.5583485,0.875249,1.0751982,1.0902886,0.91674787,0.6149379,0.7432071,1.1016065,1.2713746,1.2185578,1.2713746,1.3128735,1.1544232,0.8639311,0.5394854,0.31312788,0.29426476,0.21881226,0.1358145,0.06790725,0.00754525,0.0150905,0.02263575,0.094315626,0.3470815,0.9620194,0.9016574,0.845068,0.8224323,0.7582976,0.47157812,0.5885295,0.7469798,0.6488915,0.3772625,0.392353,0.51684964,0.65643674,2.795515,6.349328,8.152642,7.907422,8.59404,8.484633,7.0849895,5.1534057,4.08198,2.8709676,1.7542707,0.8941121,0.3734899,0.26031113,0.181086,0.124496624,0.09808825,0.1056335,0.181086,0.2565385,0.30935526,0.32067314,0.26031113,0.23013012,0.23767537,0.2263575,0.18485862,0.1358145,0.094315626,0.13204187,0.13958712,0.08677038,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.030181,0.011317875,0.0150905,0.03772625,0.060362,0.060362,0.10186087,0.120724,0.12826926,0.12826926,0.13958712,0.15467763,0.120724,0.0754525,0.03772625,0.02263575,0.03772625,0.06413463,0.1056335,0.16222288,0.2263575,0.20749438,0.21881226,0.21503963,0.181086,0.13204187,0.13204187,0.15845025,0.22258487,0.3055826,0.35462674,0.34330887,0.31312788,0.30935526,0.331991,0.33576363,0.2678564,0.19240387,0.14713238,0.1358145,0.150905,0.2263575,0.3961256,0.52062225,0.6187105,0.87147635,1.1053791,0.84129536,1.4826416,3.6141748,6.983129,3.7877154,1.6939086,0.52439487,0.0754525,0.08677038,0.10186087,0.11317875,0.124496624,0.13204187,0.1056335,0.08299775,0.181086,0.87902164,1.9240388,2.3277097,1.3166461,0.814887,0.7469798,1.2940104,2.916239,2.6597006,1.6976813,1.0978339,0.90920264,0.18485862,0.14335975,0.22258487,0.422534,0.8601585,1.7618159,3.1161883,3.4142256,3.4896781,3.4066803,2.444661,1.6486372,1.4335974,1.6863633,2.1994405,2.6823363,2.9728284,2.9501927,2.5691576,1.9089483,1.1846043,1.1657411,1.2751472,1.4298248,1.5656394,1.629774,1.1242423,0.7507524,0.5394854,0.47157812,0.51684964,0.55080324,0.5319401,0.41498876,0.26408374,0.23390275,0.19240387,0.13204187,0.090543,0.08299775,0.116951376,0.124496624,0.13958712,0.181086,0.26408374,0.3734899,0.513077,0.66020936,0.814887,0.9507015,1.0336993,1.1204696,1.1280149,1.1053791,1.0789708,1.0525624,1.2223305,1.5203679,1.991946,2.595566,3.1916409,3.0369632,2.6936543,2.3578906,2.1994405,2.3880715,2.7615614,2.8143783,2.5729303,2.1956677,1.9957186,2.2560298,2.8747404,3.4029078,3.5877664,3.3689542,3.2142766,3.1463692,3.1840954,3.2972744,3.4179983,3.7613072,4.4743333,5.406172,6.3531003,7.073672,7.145352,6.7567716,6.1305156,5.6061206,5.643847,6.066381,6.4021444,6.5455046,6.5266414,6.5266414,6.809588,7.364164,8.114917,8.89585,9.424017,9.65792,9.680555,9.7220545,9.839006,9.929549,10.325675,10.536942,10.540714,10.431308,10.438853,9.759781,8.83926,7.884786,7.149124,6.930312,6.9793563,7.149124,7.2094865,7.1302614,7.0849895,7.2660756,7.1679873,6.9755836,6.8133607,6.779407,6.673774,6.3531003,6.205968,6.3455553,6.587003,7.33021,7.466025,7.2094865,6.9189944,7.1076255,7.394345,7.145352,6.5455046,5.8513412,5.3948536,4.7912335,4.036709,3.350091,2.9464202,3.0445085,3.1954134,3.097325,3.0331905,3.1199608,3.3123648,3.4594972,3.5349495,3.7990334,4.2630663,4.7308717,4.9232755,4.5761943,4.0103,3.5424948,3.4594972,3.3915899,3.0935526,2.897376,2.9237845,3.0633714,3.2218218,3.4029078,3.5953116,3.7650797,3.874486,3.9386206,3.9688015,3.9386206,3.8405323,3.682082,3.4557245,3.3350005,3.229367,3.138824,3.150142,3.2218218,3.2444575,3.3161373,3.4594972,3.6179473,3.7084904,3.8593953,4.002755,4.112161,4.236658,4.3121104,4.327201,4.425289,4.538468,4.3875628,4.45547,4.5233774,4.3385186,3.8669407,3.2746384,2.7691069,2.4069347,2.033445,1.6146835,1.2298758,1.478869,1.7618159,1.7919968,1.5354583,1.20724,0.87902164,0.60362,0.422534,0.33576363,0.29426476,0.25276586,0.1659955,0.150905,0.211267,0.24899325,0.19994913,0.16222288,0.150905,0.1659955,0.18485862,0.20372175,0.21503963,0.18863125,0.124496624,0.071679875,0.03772625,0.018863125,0.00754525,0.0,0.0,0.00754525,0.003772625,0.003772625,0.00754525,0.0150905,0.02263575,0.033953626,0.049044125,0.056589376,0.056589376,0.049044125,0.03772625,0.030181,0.026408374,0.0150905,0.018863125,0.02263575,0.02263575,0.018863125,0.02263575,0.011317875,0.00754525,0.011317875,0.0150905,0.00754525,0.0150905,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,7.816879,7.6584287,7.118943,6.3342376,5.541986,5.0553174,4.7120085,4.304565,3.9989824,3.7688525,3.410453,2.9011486,2.7841973,2.6068838,2.2484846,1.901403,1.9240388,1.9881734,1.991946,1.9466745,1.961765,1.7919968,1.7693611,1.8334957,1.9051756,1.8749946,1.7089992,1.720317,1.9089483,2.1503963,2.2107582,2.2899833,2.2560298,2.1390784,1.9579924,1.7655885,1.6637276,1.5731846,1.5430037,1.569412,1.6184561,1.5015048,1.6146835,1.7240896,1.6486372,1.2600567,1.1393328,1.0789708,1.0035182,0.9620194,1.1280149,1.0902886,1.0676528,1.0940613,1.0978339,0.90543,0.7167987,0.6752999,0.69793564,0.72811663,0.73566186,0.90543,1.3053282,1.6675003,1.8448136,1.8221779,1.20724,1.0412445,1.0601076,1.1695137,1.4298248,1.9278114,1.8825399,1.4864142,1.0638802,1.0525624,1.1959221,1.4713237,1.7014539,2.04099,3.0105548,3.3048196,3.4255435,3.5538127,3.6368105,3.380272,2.9313297,2.4408884,1.9844007,1.6033657,1.3317367,1.4750963,1.7618159,1.8938577,1.7731338,1.5128226,1.237421,1.1317875,1.1016065,1.0789708,1.0186088,1.0902886,1.20724,1.3619176,1.5052774,1.5543215,1.6675003,1.7580433,1.6410918,1.3317367,1.0751982,0.875249,0.7394345,0.68661773,0.68661773,0.663982,0.52062225,0.45648763,0.47157812,0.543258,0.63002837,0.6187105,0.55457586,0.452715,0.35839936,0.32821837,0.20749438,0.1358145,0.120724,0.14713238,0.18863125,0.1961765,0.20749438,0.20749438,0.1961765,0.181086,0.13958712,0.094315626,0.06413463,0.056589376,0.0452715,0.03772625,0.026408374,0.033953626,0.056589376,0.090543,0.116951376,0.16222288,0.23390275,0.33953625,0.4979865,0.72811663,0.80734175,0.77338815,0.66775465,0.55080324,0.7809334,1.0978339,1.2261031,1.146878,1.0902886,0.97333723,0.7809334,0.52439487,0.2678564,0.11317875,0.116951376,0.08299775,0.049044125,0.02263575,0.0,0.00754525,0.026408374,0.15467763,0.45648763,0.97333723,0.875249,1.0110635,1.1544232,1.0827434,0.573439,0.5772116,0.68661773,0.66775465,0.52439487,0.48666862,0.55080324,0.694163,2.938875,6.7039547,8.782671,8.83926,8.518587,7.647111,6.296511,4.7950063,3.8254418,2.746471,1.7240896,0.875249,0.27917424,0.15845025,0.1056335,0.07922512,0.094315626,0.21503963,0.30181,0.36594462,0.4074435,0.42630664,0.43007925,0.46026024,0.51684964,0.4979865,0.392353,0.2867195,0.19240387,0.1659955,0.13958712,0.08677038,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.00754525,0.018863125,0.033953626,0.041498873,0.018863125,0.011317875,0.05281675,0.120724,0.12826926,0.094315626,0.071679875,0.06790725,0.094315626,0.14713238,0.1961765,0.15845025,0.10186087,0.06413463,0.049044125,0.0754525,0.1358145,0.21503963,0.271629,0.23767537,0.181086,0.15467763,0.15467763,0.1659955,0.1659955,0.17354076,0.17354076,0.29049212,0.47912338,0.52439487,0.44894236,0.36971724,0.35839936,0.40367088,0.3961256,0.271629,0.17354076,0.13204187,0.1358145,0.12826926,0.11317875,0.16222288,0.26408374,0.4376245,0.7507524,0.9016574,0.6790725,0.88279426,2.293756,5.6778007,3.5462675,1.7919968,0.62625575,0.10186087,0.10186087,0.124496624,0.1358145,0.14713238,0.14335975,0.116951376,0.090543,0.071679875,1.0072908,3.1199608,5.915476,2.9351022,1.20724,0.56589377,0.70170826,1.1581959,1.2562841,1.5241405,1.569412,1.1657411,0.27917424,0.1358145,0.14713238,0.392353,0.8337501,1.3468271,1.841041,2.4182527,3.1237335,3.5651307,2.8898308,1.599593,1.1996948,1.3166461,1.5882751,1.6524098,1.8184053,1.8938577,1.7957695,1.5128226,1.1091517,1.0714256,1.0940613,1.2525115,1.5203679,1.7391801,1.3505998,1.0072908,0.7167987,0.52062225,0.5093044,0.6149379,0.6790725,0.60362,0.42630664,0.33953625,0.22258487,0.15467763,0.11317875,0.090543,0.071679875,0.060362,0.05281675,0.06790725,0.120724,0.20749438,0.331991,0.45648763,0.5885295,0.72811663,0.8526133,0.9808825,1.0525624,1.116697,1.1808317,1.2110126,1.3845534,1.6410918,1.9579924,2.3201644,2.71629,2.6710186,2.6597006,2.7804246,3.1312788,3.7914882,4.3649273,4.274384,3.5990841,2.7011995,2.233394,2.4974778,3.0671442,3.3764994,3.2105038,2.7238352,2.4031622,2.3088465,2.4484336,2.7728794,3.169005,3.6594462,4.2027044,4.8365054,5.485397,5.9494295,5.987156,5.7494807,5.311856,4.90064,4.8666863,5.13077,5.3344917,5.409944,5.4288073,5.643847,6.1116524,6.647365,7.152897,7.541477,7.7338815,7.835742,7.937603,8.107371,8.371455,8.714764,9.371201,9.895596,10.159679,10.246449,10.450171,10.321902,9.963503,9.348565,8.601585,7.9753294,7.360391,7.0585814,6.881268,6.722818,6.560595,6.700182,6.7152724,6.5040054,6.1644692,6.013564,5.987156,5.59103,5.240176,5.168496,5.4363527,6.2851934,6.511551,6.5530496,6.696409,7.0585814,6.930312,6.983129,6.779407,6.224831,5.5683947,5.2326307,4.5007415,3.6368105,2.9652832,2.8936033,2.9615107,2.8294687,2.7313805,2.8332415,3.2557755,3.4896781,3.5123138,3.5764484,3.7763977,4.0291634,4.244203,3.9650288,3.519859,3.1463692,3.006782,2.9539654,2.7238352,2.5276587,2.4899325,2.625747,2.6483827,2.7238352,2.8294687,2.927557,2.9652832,3.078462,3.1916409,3.259548,3.2670932,3.2369123,3.240685,3.2444575,3.289729,3.380272,3.4783602,3.5123138,3.531177,3.6141748,3.7688525,3.9348478,3.9763467,4.06689,4.142342,4.168751,4.1574326,4.183841,4.2027044,4.2404304,4.1083884,3.399135,3.2670932,3.1954134,2.916239,2.3993895,1.8448136,1.4109617,1.1883769,1.0751982,1.0223814,1.0525624,1.5467763,1.8523588,1.7882242,1.3807807,0.8563859,0.44516975,0.2867195,0.24899325,0.21503963,0.090543,0.06790725,0.0754525,0.124496624,0.21503963,0.32821837,0.2565385,0.1659955,0.116951376,0.12826926,0.16222288,0.19240387,0.21881226,0.19994913,0.13958712,0.094315626,0.0754525,0.060362,0.041498873,0.026408374,0.018863125,0.026408374,0.0150905,0.003772625,0.0,0.00754525,0.02263575,0.033953626,0.05281675,0.06413463,0.06413463,0.0452715,0.030181,0.02263575,0.0150905,0.0150905,0.026408374,0.026408374,0.02263575,0.018863125,0.02263575,0.011317875,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,8.073418,7.997965,7.699928,7.1378064,6.4210076,5.824933,5.3910813,5.0251365,4.82896,4.67051,4.183841,4.036709,4.172523,4.006528,3.5349495,3.3236825,3.2142766,3.289729,3.229367,2.9728284,2.6974268,2.3277097,2.3126192,2.3503454,2.3163917,2.2484846,2.0258996,2.1692593,2.4861598,2.746471,2.6634734,2.5276587,2.4672968,2.372981,2.191895,1.9579924,1.7655885,1.6863633,1.659955,1.6184561,1.5128226,1.358145,1.3694628,1.3091009,1.1431054,1.0072908,0.845068,0.784706,0.7696155,0.76584285,0.77338815,0.65643674,0.6413463,0.66020936,0.6488915,0.5583485,0.5281675,0.5281675,0.60362,0.73188925,0.84129536,1.1393328,1.6524098,2.0145817,2.0560806,1.7769064,1.1921495,0.8941121,0.84129536,0.9997456,1.3166461,2.093807,2.2560298,2.052308,1.7655885,1.7165444,2.0975795,2.3428001,2.6219745,3.2218218,4.561104,4.6856003,4.715781,4.7535076,4.6327834,3.904667,3.108643,2.323937,1.81086,1.6863633,1.9051756,2.595566,3.6707642,4.0517993,3.5085413,2.6710186,1.7467253,1.3204187,1.1431054,1.0676528,1.0450171,1.1204696,1.2223305,1.327964,1.4071891,1.3996439,1.448688,1.4562333,1.3355093,1.1053791,0.91674787,0.77338815,0.663982,0.573439,0.5055317,0.48666862,0.48666862,0.4376245,0.422534,0.46026024,0.5093044,0.513077,0.5017591,0.45648763,0.38103512,0.27540162,0.16976812,0.124496624,0.116951376,0.10940613,0.056589376,0.056589376,0.060362,0.05281675,0.0452715,0.08677038,0.10186087,0.08299775,0.060362,0.049044125,0.041498873,0.018863125,0.018863125,0.033953626,0.060362,0.10186087,0.12826926,0.19240387,0.27917424,0.3734899,0.47912338,0.6828451,0.724344,0.6451189,0.55457586,0.59607476,0.8224323,1.0223814,1.0940613,1.026154,0.91674787,0.73566186,0.49044126,0.271629,0.13204187,0.0754525,0.060362,0.030181,0.00754525,0.0,0.0,0.0,0.060362,0.21503963,0.49421388,0.8941121,0.56589377,0.814887,1.1695137,1.2600567,0.8299775,0.6413463,0.55457586,0.5470306,0.56212115,0.513077,0.6413463,0.9318384,2.9615107,6.368191,8.846806,9.74469,7.9526935,5.987156,4.8855495,4.195159,3.6443558,2.637065,1.5618668,0.70170826,0.20749438,0.041498873,0.0,0.00754525,0.071679875,0.29426476,0.3772625,0.42630664,0.44139713,0.452715,0.5319401,0.63002837,0.7507524,0.754525,0.62625575,0.452715,0.24899325,0.1056335,0.03772625,0.02263575,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.026408374,0.02263575,0.011317875,0.003772625,0.003772625,0.0150905,0.041498873,0.06413463,0.060362,0.049044125,0.02263575,0.07922512,0.1961765,0.23013012,0.20749438,0.15845025,0.120724,0.1056335,0.10940613,0.12826926,0.1056335,0.07922512,0.06413463,0.071679875,0.10940613,0.19240387,0.3169005,0.392353,0.24899325,0.17354076,0.124496624,0.13204187,0.1961765,0.271629,0.24522063,0.19994913,0.34330887,0.6149379,0.6790725,0.56589377,0.43007925,0.35462674,0.3734899,0.43007925,0.28294688,0.1961765,0.15467763,0.13958712,0.13958712,0.1358145,0.13958712,0.18485862,0.32821837,0.67152727,0.68661773,0.52062225,0.2867195,0.22258487,0.7092535,0.98465514,0.90543,0.66775465,0.3961256,0.124496624,0.181086,0.20372175,0.19240387,0.16222288,0.11317875,0.090543,0.06413463,1.0601076,3.9461658,9.439108,5.455216,2.3692086,0.7394345,0.5017591,0.9808825,1.4034165,1.5203679,1.20724,0.6413463,0.31312788,0.14713238,0.11317875,0.36971724,0.83752275,1.1959221,1.3468271,1.6939086,2.2296214,2.7502437,2.8407867,1.5505489,1.1732863,1.1355602,1.0525624,0.7469798,0.6752999,0.875249,1.2336484,1.5241405,1.388326,1.0601076,0.86770374,0.875249,1.0487897,1.2525115,1.3505998,1.2261031,0.9620194,0.66775465,0.4640329,0.47535074,0.55457586,0.6073926,0.59607476,0.5357128,0.3961256,0.30181,0.22258487,0.15467763,0.1056335,0.06790725,0.041498873,0.03772625,0.049044125,0.08677038,0.14713238,0.21881226,0.32821837,0.44894236,0.543258,0.6451189,0.7432071,0.8865669,1.056335,1.1921495,1.3091009,1.5015048,1.7278622,1.9579924,2.1579416,2.2258487,2.5540671,3.1237335,3.9084394,4.8402777,5.413717,5.172269,4.304565,3.2784111,2.8521044,3.1463692,3.470815,3.4783602,3.1237335,2.637065,2.354118,2.3088465,2.5502944,3.006782,3.4972234,3.893349,4.002755,4.025391,4.0706625,4.1612053,4.327201,4.4101987,4.425289,4.3686996,4.22534,4.406426,4.6327834,4.90064,5.2779026,5.9003854,6.537959,6.9491754,7.020855,6.752999,6.255012,5.975838,6.089017,6.398372,6.820906,7.364164,8.099826,8.941121,9.567377,9.842778,9.812597,10.148361,10.540714,10.623712,10.246449,9.476834,8.428044,7.5716586,6.94163,6.436098,5.8098426,5.885295,5.915476,5.704209,5.330719,5.142088,5.040227,4.9345937,4.8629136,4.881777,5.032682,5.3684454,5.5985756,5.904158,6.2436943,6.3644185,5.523123,5.6476197,5.7494807,5.2892203,4.1762958,4.3007927,4.044254,3.5424948,3.0256453,2.8181508,2.6483827,2.5578396,2.474842,2.5616124,3.2029586,3.572676,3.5424948,3.180323,2.7238352,2.5616124,2.7389257,2.9049213,2.9501927,2.8747404,2.7804246,2.9426475,2.8785129,2.8030603,2.8407867,3.0105548,2.848332,2.7691069,2.7841973,2.837014,2.8030603,2.9351022,3.1161883,3.31991,3.531177,3.7462165,3.92353,4.08198,4.221567,4.3196554,4.346064,4.346064,4.3422914,4.3347464,4.315883,4.29702,4.195159,4.142342,4.0480266,3.8593953,3.5424948,3.5877664,3.5877664,3.5387223,3.199186,2.1088974,1.6373192,1.3543724,1.1317875,0.8941121,0.6187105,0.44516975,0.362172,0.41498876,0.6375736,1.0450171,1.5015048,1.5052774,1.2789198,0.97710985,0.6526641,0.41498876,0.30181,0.241448,0.17354076,0.060362,0.060362,0.08677038,0.1358145,0.1961765,0.27917424,0.20749438,0.10940613,0.049044125,0.041498873,0.049044125,0.06790725,0.08677038,0.08299775,0.06790725,0.07922512,0.120724,0.14713238,0.14335975,0.1056335,0.056589376,0.041498873,0.02263575,0.00754525,0.003772625,0.00754525,0.0150905,0.0150905,0.02263575,0.041498873,0.041498873,0.030181,0.02263575,0.018863125,0.018863125,0.018863125,0.026408374,0.02263575,0.0150905,0.018863125,0.018863125,0.00754525,0.003772625,0.003772625,0.003772625,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,8.13378,8.243186,8.488406,8.265821,7.533932,6.851087,7.020855,7.066127,6.911449,6.537959,5.96452,5.915476,5.7306175,5.485397,5.3873086,5.753253,5.5570765,5.0515447,4.164978,3.187868,2.746471,2.6106565,2.6974268,2.595566,2.2975287,2.2107582,2.4672968,2.9728284,3.3463185,3.410453,3.187868,2.5540671,2.4861598,2.6144292,2.6898816,2.595566,2.252257,1.9579924,1.7429527,1.6712729,1.8297231,1.9768555,2.003264,1.6939086,1.2147852,1.1280149,1.0940613,0.8903395,0.69039035,0.5885295,0.62625575,0.87147635,1.1242423,1.1431054,0.8639311,0.41121614,0.41121614,0.44894236,0.5470306,0.7205714,0.97710985,0.98842776,1.0299267,1.1431054,1.3015556,1.3732355,1.2864652,1.1581959,1.3694628,1.9240388,2.425798,2.9501927,3.5500402,3.8480775,3.8669407,4.014073,5.0741806,5.0025005,4.659192,4.587512,4.991183,5.3571277,5.372218,5.062863,4.395108,3.2972744,2.5767028,2.0673985,1.8523588,2.1353056,3.2331395,5.4212623,8.182823,8.907167,7.2585306,5.172269,3.0860074,2.0787163,1.6071383,1.3656902,1.267602,1.2902378,1.3053282,1.3317367,1.3770081,1.448688,1.2902378,1.20724,1.1581959,1.0978339,0.97710985,0.8526133,0.7130261,0.55080324,0.39989826,0.35085413,0.35085413,0.35839936,0.35839936,0.35085413,0.35085413,0.3772625,0.41876137,0.41876137,0.35839936,0.27540162,0.23767537,0.17354076,0.1056335,0.056589376,0.030181,0.030181,0.02263575,0.00754525,0.003772625,0.0150905,0.026408374,0.030181,0.02263575,0.0150905,0.0150905,0.0150905,0.033953626,0.056589376,0.08677038,0.1358145,0.22258487,0.3169005,0.452715,0.62625575,0.80734175,0.8563859,0.80734175,0.694163,0.5696664,0.47157812,0.58475685,0.7092535,0.8224323,0.8563859,0.73188925,0.6111652,0.46026024,0.27917424,0.11317875,0.0754525,0.08677038,0.0452715,0.00754525,0.0,0.0,0.0,0.21881226,0.47157812,0.6375736,0.68661773,0.32067314,0.27540162,0.42630664,0.6111652,0.6111652,0.58475685,0.5696664,0.56589377,0.5017591,0.24522063,0.84129536,2.173032,3.9914372,6.149379,8.590267,10.103089,7.213259,4.466788,3.5236318,3.1576872,2.2560298,1.6373192,1.1280149,0.6451189,0.18485862,0.03772625,0.0,0.030181,0.08677038,0.1358145,0.19994913,0.26031113,0.28294688,0.27540162,0.27540162,0.32444575,0.41876137,0.3772625,0.20749438,0.120724,0.1358145,0.18485862,0.18485862,0.10940613,0.0,0.0,0.0,0.0,0.026408374,0.1358145,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.026408374,0.030181,0.02263575,0.0150905,0.0150905,0.0150905,0.00754525,0.011317875,0.03772625,0.060362,0.09808825,0.071679875,0.033953626,0.02263575,0.060362,0.27917424,0.3734899,0.3772625,0.3169005,0.18485862,0.08677038,0.033953626,0.0150905,0.02263575,0.0452715,0.0452715,0.056589376,0.13958712,0.271629,0.32067314,0.29426476,0.30935526,0.39989826,0.51684964,0.5017591,0.17354076,0.08299775,0.094315626,0.12826926,0.150905,0.2867195,0.31312788,0.2678564,0.211267,0.19994913,0.150905,0.1358145,0.14335975,0.150905,0.150905,0.12826926,0.11317875,0.1358145,0.23013012,0.42630664,0.5998474,0.422534,0.21881226,0.15845025,0.24522063,0.4640329,1.0412445,1.3958713,1.1393328,0.0754525,0.211267,0.24522063,0.2263575,0.18485862,0.1358145,0.124496624,0.094315626,0.11317875,0.9808825,4.22534,5.3986263,3.3312278,1.3317367,0.6488915,0.44139713,0.56589377,0.5772116,0.51684964,0.39989826,0.23013012,0.120724,0.1358145,0.30181,0.6451189,1.2223305,1.478869,1.7052265,1.901403,1.9994912,1.8787673,2.0108092,2.2560298,2.354118,2.1164427,1.418507,0.7582976,0.58475685,0.7092535,0.91297525,0.9620194,0.72811663,0.7432071,0.8601585,0.9997456,1.1431054,1.3392819,1.3317367,1.1921495,0.9507015,0.6111652,0.573439,0.6187105,0.73566186,0.8865669,1.0223814,0.97333723,0.80734175,0.55457586,0.30181,0.1659955,0.120724,0.071679875,0.033953626,0.011317875,0.0,0.011317875,0.05281675,0.120724,0.21503963,0.33576363,0.5055317,0.73188925,0.9695646,1.1695137,1.267602,1.2185578,1.20724,1.2902378,1.4864142,1.7542707,2.0975795,2.4823873,3.1010978,3.863168,4.425289,4.606375,4.515832,4.2291126,3.874486,3.6330378,3.802806,3.8443048,3.6669915,3.2482302,2.625747,2.3428001,2.3918443,2.7351532,3.289729,3.9386206,4.304565,4.4215164,4.2630663,3.953711,3.7688525,3.7198083,3.7801702,3.9273026,4.104616,4.22534,4.349837,4.689373,5.1534057,5.6589375,6.1342883,6.096562,5.832478,5.458988,5.0251365,4.485651,4.1083884,4.123479,4.459243,5.0553174,5.873977,6.828451,7.8244243,8.922258,9.80128,9.767326,9.767326,10.589758,11.0613365,10.868933,10.589758,10.453944,9.661693,8.473316,7.066127,5.553304,5.772116,5.855114,5.80607,5.6778007,5.5683947,5.5080323,5.3646727,5.119452,4.8629136,4.776143,4.9949555,5.3080835,5.485397,5.413717,5.0968165,4.644101,4.447925,4.1008434,3.5877664,3.2972744,3.6745367,3.5764484,3.31991,3.0897799,2.9313297,2.4182527,2.1503963,2.0862615,2.1051247,2.0447628,2.1315331,2.1881225,2.071171,1.8523588,1.8146327,2.071171,2.565385,2.938875,3.048281,2.9766011,2.7691069,2.7351532,2.9464202,3.361409,3.8141239,3.6443558,3.4368613,3.270866,3.1916409,3.2029586,3.4745877,3.7688525,4.08198,4.478106,5.111907,5.4665337,5.6551647,5.6363015,5.4212623,5.0666356,4.821415,4.8968673,4.8968673,4.7006907,4.45547,4.13857,3.8858037,3.519859,2.9803739,2.335255,2.0673985,1.7354075,1.4298248,1.1695137,0.9016574,0.7432071,0.6488915,0.6111652,0.58475685,0.47157812,0.38858038,0.3470815,0.36594462,0.46026024,0.65643674,0.7922512,0.694163,0.52439487,0.3734899,0.27540162,0.21503963,0.14335975,0.10186087,0.09808825,0.120724,0.071679875,0.05281675,0.041498873,0.033953626,0.0452715,0.033953626,0.030181,0.02263575,0.011317875,0.0,0.0,0.0,0.00754525,0.030181,0.090543,0.19994913,0.31312788,0.32821837,0.241448,0.1056335,0.033953626,0.00754525,0.00754525,0.02263575,0.0452715,0.033953626,0.011317875,0.00754525,0.0150905,0.0150905,0.0150905,0.02263575,0.030181,0.030181,0.030181,0.030181,0.02263575,0.02263575,0.030181,0.030181,0.018863125,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,9.49947,9.4127,9.216523,8.631766,7.858378,7.594294,7.3679366,6.9265394,6.6662283,6.571913,6.221059,5.5985756,5.5382137,5.6891184,5.8664317,6.043745,6.066381,5.8890676,5.4363527,4.7836885,4.187614,3.7801702,3.4444065,3.1010978,2.8558772,2.9954643,3.4632697,3.9650288,3.9801195,3.5802212,3.410453,3.2218218,3.1652324,3.0369632,2.7804246,2.4974778,2.3126192,2.425798,2.584248,2.6974268,2.8558772,2.7087448,2.41448,1.9881734,1.5203679,1.1883769,0.995973,0.8299775,0.69039035,0.6073926,0.6149379,0.67152727,0.70170826,0.6526641,0.543258,0.46026024,0.5583485,0.6488915,0.784706,0.97333723,1.1732863,1.0751982,1.0827434,1.1393328,1.1996948,1.2147852,1.267602,1.4826416,1.991946,2.686109,3.2557755,3.7990334,4.346064,4.927048,5.6023483,6.4436436,7.220804,7.2170315,7.1981683,7.4169807,7.624475,7.5037513,6.477597,5.240176,4.142342,3.199186,2.8294687,2.8181508,3.1124156,3.7650797,4.9421387,7.8810134,10.114408,10.208723,8.190369,5.5268955,3.5160866,2.4710693,2.0598533,1.991946,2.0108092,2.0749438,2.0636258,1.9655377,1.7844516,1.5354583,1.2902378,1.1431054,1.056335,0.9808825,0.87902164,0.68661773,0.573439,0.5093044,0.44516975,0.32821837,0.3055826,0.331991,0.35839936,0.35462674,0.32821837,0.31312788,0.32444575,0.33576363,0.35462674,0.3961256,0.48666862,0.3961256,0.24899325,0.120724,0.018863125,0.018863125,0.0150905,0.0150905,0.011317875,0.0150905,0.00754525,0.0150905,0.030181,0.0452715,0.026408374,0.03772625,0.049044125,0.1056335,0.20749438,0.34330887,0.51684964,0.62625575,0.7469798,0.88279426,0.965792,0.76207024,0.6187105,0.52062225,0.47157812,0.47157812,0.60362,0.7130261,0.80734175,0.8337501,0.67152727,0.452715,0.24899325,0.10940613,0.0452715,0.041498873,0.041498873,0.018863125,0.0,0.02263575,0.120724,0.33576363,0.36971724,0.47912338,0.73566186,1.0299267,0.67152727,0.67152727,0.7997965,0.814887,0.4640329,0.5281675,0.5281675,0.36971724,0.16976812,0.24522063,1.5354583,3.6556737,5.873977,7.6282477,8.518587,8.088508,5.311856,3.1463692,2.516341,2.3163917,1.4034165,0.9507015,0.68661773,0.46026024,0.23013012,0.0452715,0.0,0.033953626,0.10940613,0.18485862,0.34330887,0.47535074,0.4979865,0.422534,0.32444575,0.26408374,0.2678564,0.23013012,0.14713238,0.10940613,0.0452715,0.071679875,0.071679875,0.02263575,0.0,0.0,0.0,0.0,0.003772625,0.026408374,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.05281675,0.06413463,0.05281675,0.030181,0.0150905,0.0150905,0.003772625,0.00754525,0.0150905,0.02263575,0.03772625,0.071679875,0.060362,0.030181,0.00754525,0.02263575,0.1056335,0.181086,0.26408374,0.30935526,0.1961765,0.116951376,0.1056335,0.1358145,0.16976812,0.15467763,0.056589376,0.033953626,0.05281675,0.08299775,0.10186087,0.14335975,0.1659955,0.18863125,0.1961765,0.124496624,0.116951376,0.15845025,0.23390275,0.30181,0.2867195,0.3734899,0.45648763,0.40367088,0.241448,0.16222288,0.124496624,0.12826926,0.14335975,0.150905,0.150905,0.13958712,0.15467763,0.17354076,0.181086,0.16976812,0.36971724,0.3470815,0.25276586,0.25276586,0.513077,0.47912338,0.56589377,0.87147635,1.0676528,0.4074435,0.13958712,0.14713238,0.19240387,0.18485862,0.17354076,0.16222288,0.08677038,0.17354076,0.6752999,1.871222,2.4069347,1.629774,0.7922512,0.45648763,0.49044126,0.4979865,0.5093044,0.5319401,0.49044126,0.241448,0.181086,0.21881226,0.3772625,0.6828451,1.1581959,1.991946,3.4934506,4.4743333,4.478106,3.7801702,2.372981,1.901403,1.6976813,1.3619176,0.77338815,0.44516975,0.44139713,0.5885295,0.7092535,0.63002837,0.56589377,0.5998474,0.70170826,0.8563859,1.0714256,1.3920987,1.7618159,2.0183544,2.0108092,1.599593,1.2487389,0.9695646,0.8224323,0.7997965,0.8262049,0.77716076,0.76584285,0.6790725,0.47912338,0.181086,0.16222288,0.15467763,0.14335975,0.1056335,0.03772625,0.011317875,0.018863125,0.071679875,0.17354076,0.33576363,0.573439,0.8186596,1.0525624,1.2261031,1.2525115,1.0676528,0.8978847,0.8601585,1.0110635,1.327964,1.7957695,2.2371666,2.6936543,3.1350515,3.4745877,3.6858547,3.8443048,3.9574835,4.0404816,4.1083884,4.074435,3.8593953,3.7273536,3.6896272,3.5274043,3.187868,2.9237845,2.8898308,3.0709167,3.2784111,3.5764484,3.6934,3.6443558,3.4896781,3.3048196,3.3651814,3.500996,3.712263,3.99521,4.3611546,4.7648253,5.149633,5.300538,5.2175403,5.0968165,4.8930945,4.696918,4.5460134,4.429062,4.2894745,4.1762958,4.1612053,4.349837,4.745962,5.251494,5.8437963,6.485142,7.17176,7.8319697,8.360137,9.046755,9.748463,10.012547,9.955957,10.272858,10.148361,9.5183325,8.782671,8.099826,7.3981175,7.069899,7.0812173,7.01331,6.696409,6.217286,5.794752,5.4438977,5.3156285,5.3194013,5.119452,4.821415,4.678055,4.6742826,4.6856003,4.485651,4.1498876,3.904667,3.9386206,4.2027044,4.406426,4.187614,4.002755,3.6896272,3.2444575,2.7841973,3.0520537,3.2444575,3.4481792,3.7273536,4.1574326,3.4330888,2.4974778,1.8674494,1.7391801,1.9881734,2.252257,2.7200627,2.9954643,2.9728284,2.8407867,2.7917426,2.8521044,2.9652832,3.0860074,3.218049,3.240685,3.3010468,3.3236825,3.308592,3.350091,3.7273536,4.0480266,4.323428,4.52715,4.636556,4.666737,4.6516466,4.5950575,4.447925,4.112161,3.6858547,3.3915899,3.2255943,3.108643,2.9049213,2.637065,2.4899325,2.3918443,2.2371666,1.8825399,1.388326,1.0148361,0.7507524,0.573439,0.46026024,0.4376245,0.46026024,0.5055317,0.543258,0.5093044,0.44516975,0.39989826,0.40367088,0.4678055,0.59607476,0.67152727,0.70170826,0.6413463,0.4979865,0.32444575,0.1659955,0.09808825,0.0754525,0.071679875,0.08677038,0.124496624,0.16222288,0.18863125,0.18863125,0.14335975,0.090543,0.094315626,0.150905,0.22258487,0.21881226,0.19994913,0.1961765,0.20749438,0.25276586,0.3734899,0.49044126,0.4376245,0.38480774,0.36594462,0.241448,0.12826926,0.060362,0.049044125,0.07922512,0.13204187,0.090543,0.03772625,0.00754525,0.003772625,0.003772625,0.003772625,0.011317875,0.02263575,0.030181,0.030181,0.030181,0.03772625,0.041498873,0.041498873,0.041498873,0.041498873,0.033953626,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,9.631512,9.5032425,9.582467,9.529651,9.2995205,9.125979,8.329956,7.4735703,6.9152217,6.722818,6.670001,6.398372,6.228604,6.2021956,6.3342376,6.587003,6.7454534,6.752999,6.5266414,6.092789,5.59103,5.1571784,4.8930945,4.6214657,4.3121104,4.104616,4.5799665,4.919503,4.908185,4.647874,4.5724216,4.666737,4.636556,4.2064767,3.5764484,3.4255435,3.0633714,2.6219745,2.4408884,2.5502944,2.6634734,2.5767028,2.1202152,1.6222287,1.2562841,1.0487897,0.84884065,0.72811663,0.6451189,0.573439,0.49044126,0.5319401,0.543258,0.51684964,0.482896,0.52062225,0.6187105,0.7432071,0.94315624,1.1883769,1.3958713,1.448688,1.4449154,1.4222796,1.4071891,1.4147344,1.4750963,1.7165444,2.0900342,2.493705,2.757789,3.1916409,3.7462165,4.4894238,5.4665337,6.730363,7.4735703,7.835742,8.024373,8.07719,7.854605,7.3188925,6.149379,5.0251365,4.2781568,3.8782585,4.146115,4.4403796,5.240176,6.7341356,8.82417,10.789707,11.336739,10.295494,8.080963,5.7079816,4.0895257,3.0897799,2.757789,2.8219235,2.6634734,2.474842,2.263575,2.0447628,1.81086,1.5580941,1.3392819,1.1808317,1.0487897,0.91674787,0.7809334,0.6828451,0.5998474,0.543258,0.5055317,0.4678055,0.41876137,0.38480774,0.36594462,0.35085413,0.32821837,0.3055826,0.29049212,0.32067314,0.38858038,0.45648763,0.5093044,0.4074435,0.26031113,0.13204187,0.02263575,0.018863125,0.011317875,0.00754525,0.00754525,0.00754525,0.0,0.0150905,0.033953626,0.05281675,0.056589376,0.12826926,0.27540162,0.6187105,1.0186088,1.0827434,0.9997456,0.8299775,0.76207024,0.8262049,0.8865669,0.80356914,0.5998474,0.45648763,0.452715,0.56589377,0.76584285,0.814887,0.784706,0.70170826,0.58475685,0.3470815,0.15467763,0.060362,0.06413463,0.094315626,0.094315626,0.03772625,0.06413463,0.1961765,0.35462674,0.543258,0.5281675,0.58475685,0.784706,1.0223814,0.80734175,0.9808825,1.1242423,0.97333723,0.41876137,0.3734899,0.392353,0.43007925,0.4678055,0.5093044,1.8485862,3.8669407,5.20245,5.4665337,5.221313,4.6931453,3.742444,3.0935526,2.9011486,2.727608,1.9655377,1.4901869,1.1016065,0.68661773,0.20749438,0.041498873,0.0,0.1056335,0.271629,0.29803738,0.44516975,0.5772116,0.5772116,0.4678055,0.41876137,0.33953625,0.18485862,0.0754525,0.05281675,0.041498873,0.03772625,0.033953626,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.033953626,0.060362,0.049044125,0.026408374,0.018863125,0.02263575,0.018863125,0.02263575,0.026408374,0.033953626,0.041498873,0.0452715,0.03772625,0.018863125,0.011317875,0.02263575,0.05281675,0.0754525,0.1056335,0.12826926,0.09808825,0.11317875,0.14713238,0.16976812,0.1659955,0.120724,0.071679875,0.06413463,0.06413463,0.056589376,0.0452715,0.1056335,0.16976812,0.19994913,0.18485862,0.120724,0.12826926,0.14335975,0.1961765,0.2678564,0.2565385,0.29426476,0.38858038,0.38858038,0.28294688,0.20749438,0.16222288,0.15467763,0.150905,0.13204187,0.08677038,0.090543,0.120724,0.15845025,0.17354076,0.1056335,0.17354076,0.19240387,0.1961765,0.2678564,0.55080324,0.6828451,0.7205714,0.90920264,1.0751982,0.6451189,0.15467763,0.07922512,0.116951376,0.13204187,0.15467763,0.150905,0.10940613,0.1659955,0.5055317,1.3656902,1.6675003,1.3430545,0.8337501,0.44516975,0.3734899,0.32067314,0.32821837,0.41121614,0.5093044,0.49044126,0.42630664,0.3961256,0.482896,0.7205714,1.0714256,1.7089992,3.3425457,4.9044123,5.6287565,5.036454,3.92353,3.3123648,3.108643,2.8407867,1.6260014,0.5998474,0.3169005,0.35085413,0.41876137,0.3734899,0.3734899,0.46026024,0.59230214,0.7469798,0.94315624,1.2449663,1.569412,1.8334957,1.9429018,1.7995421,1.4600059,1.086516,0.77716076,0.59607476,0.5583485,0.51684964,0.48666862,0.44516975,0.38103512,0.30181,0.39989826,0.47157812,0.4678055,0.3772625,0.211267,0.071679875,0.033953626,0.08677038,0.211267,0.38103512,0.5281675,0.6488915,0.754525,0.84884065,0.9016574,0.83752275,0.7809334,0.7809334,0.8639311,1.0450171,1.3204187,1.5958204,1.8938577,2.2107582,2.5125682,2.8332415,3.187868,3.5538127,3.893349,4.172523,4.2102494,4.112161,4.08198,4.1800685,4.3196554,4.0480266,3.651901,3.2557755,2.9237845,2.6634734,2.6219745,2.6483827,2.8256962,3.169005,3.591539,4.22534,4.538468,4.6742826,4.738417,4.8063245,5.1156793,5.300538,5.1873593,4.776143,4.2517486,3.9914372,3.9122121,4.0178456,4.2404304,4.4630156,4.5007415,4.5007415,4.4818783,4.5007415,4.647874,5.0025005,5.4891696,6.0701537,6.7114997,7.360391,7.9451485,8.379,8.560086,8.631766,8.993938,9.405154,9.363655,9.114662,8.771353,8.307321,7.888559,7.699928,7.488661,7.0887623,6.4436436,5.7683434,5.342037,5.1232247,4.991183,4.745962,4.7950063,4.8855495,4.878004,4.727099,4.496969,4.4931965,4.5007415,4.719554,5.1760416,5.7192993,5.704209,5.492942,5.062863,4.617693,4.587512,4.7572803,4.6629643,4.4139714,4.187614,4.2102494,3.9159849,3.500996,3.1954134,3.0671442,3.0181,3.1463692,3.4896781,3.6669915,3.5236318,3.138824,2.8521044,2.7653341,2.795515,2.8822856,2.9652832,3.0633714,3.138824,3.169005,3.1765501,3.240685,3.519859,3.7499893,3.893349,3.92353,3.8480775,3.7763977,3.7198083,3.6443558,3.4896781,3.187868,2.806833,2.5238862,2.372981,2.3013012,2.1805773,1.9391292,1.7844516,1.6712729,1.5279131,1.2487389,0.845068,0.55080324,0.38858038,0.331991,0.331991,0.41121614,0.5093044,0.573439,0.5772116,0.5281675,0.44516975,0.4074435,0.41876137,0.47535074,0.56212115,0.55080324,0.5055317,0.43385187,0.33953625,0.21503963,0.17354076,0.18863125,0.18485862,0.15467763,0.15845025,0.17731337,0.2678564,0.3470815,0.38480774,0.4074435,0.271629,0.18485862,0.1659955,0.19240387,0.19240387,0.18863125,0.20749438,0.23767537,0.29803738,0.43385187,0.55457586,0.55080324,0.48666862,0.392353,0.2565385,0.17731337,0.16222288,0.15845025,0.14713238,0.14335975,0.10186087,0.05281675,0.0150905,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.02263575,0.030181,0.041498873,0.0452715,0.0452715,0.0452715,0.0452715,0.03772625,0.02263575,0.011317875,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,9.733373,9.933322,10.34831,10.642575,10.601076,10.140816,8.903395,8.152642,7.654656,7.3000293,7.122716,7.2962565,7.1566696,7.020855,7.0887623,7.4471617,7.6810646,7.7414265,7.575431,7.2698483,7.0548086,6.8171334,6.670001,6.5002327,6.2889657,6.1078796,6.5455046,6.3832817,6.1229706,6.0286546,6.138061,6.5266414,6.19465,5.292993,4.3347464,4.1762958,3.7462165,3.0897799,2.71629,2.6446102,2.4031622,2.1881225,1.720317,1.3355093,1.1544232,1.0676528,0.90543,0.7997965,0.694163,0.5696664,0.422534,0.47535074,0.5470306,0.5998474,0.6187105,0.5998474,0.66775465,0.7884786,0.97333723,1.237421,1.5769572,1.7844516,1.8334957,1.8146327,1.7919968,1.8146327,1.8561316,1.9806281,2.1768045,2.3993895,2.5993385,3.097325,3.7952607,4.7610526,6.043745,7.7037,7.809334,7.8508325,7.752744,7.405663,6.6662283,6.0248823,5.2590394,4.6214657,4.3007927,4.4403796,5.198677,6.1116524,7.798016,10.227587,12.721292,13.528633,12.294985,10.054046,7.586749,5.4212623,4.4101987,3.7084904,3.470815,3.4557245,3.048281,2.7653341,2.3465726,1.9957186,1.7844516,1.629774,1.4562333,1.2449663,1.0601076,0.9205205,0.7884786,0.72811663,0.6073926,0.5017591,0.452715,0.46026024,0.4640329,0.41876137,0.36971724,0.331991,0.3055826,0.30935526,0.31312788,0.33953625,0.3772625,0.39989826,0.3772625,0.28294688,0.181086,0.090543,0.018863125,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0150905,0.03772625,0.0754525,0.150905,0.36594462,0.6828451,1.1846043,1.6373192,1.478869,1.2034674,0.9242931,0.784706,0.814887,0.9507015,1.116697,0.90920264,0.6828451,0.5998474,0.6488915,0.84884065,0.8262049,0.69039035,0.55080324,0.49044126,0.27540162,0.116951376,0.060362,0.12826926,0.31312788,0.33953625,0.241448,0.2678564,0.42630664,0.4640329,0.46026024,0.5998474,0.724344,0.7696155,0.7469798,0.5583485,0.6828451,0.79602385,0.72811663,0.47157812,0.3470815,0.31312788,0.38480774,0.68661773,1.4298248,2.2183034,3.0671442,3.3425457,2.9954643,2.5238862,2.4295704,2.8558772,3.1312788,3.0633714,2.9351022,2.9501927,2.7804246,2.305074,1.4411428,0.150905,0.211267,0.24522063,0.3055826,0.3734899,0.34330887,0.48666862,0.6451189,0.6488915,0.482896,0.28294688,0.241448,0.090543,0.0,0.0,0.0,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.041498873,0.0452715,0.033953626,0.018863125,0.011317875,0.02263575,0.02263575,0.02263575,0.0452715,0.071679875,0.056589376,0.041498873,0.02263575,0.0150905,0.018863125,0.030181,0.056589376,0.0452715,0.02263575,0.011317875,0.030181,0.10940613,0.15467763,0.16222288,0.14713238,0.120724,0.1056335,0.10186087,0.10186087,0.08677038,0.06413463,0.094315626,0.17731337,0.23390275,0.241448,0.20749438,0.150905,0.124496624,0.15845025,0.23767537,0.2867195,0.271629,0.32067314,0.34330887,0.31312788,0.29426476,0.23767537,0.19994913,0.16976812,0.1358145,0.06413463,0.05281675,0.06790725,0.13958712,0.21503963,0.18485862,0.1358145,0.120724,0.150905,0.271629,0.5357128,1.0035182,1.0902886,1.0336993,0.8941121,0.52062225,0.14335975,0.049044125,0.06413463,0.094315626,0.13204187,0.13204187,0.116951376,0.124496624,0.3055826,0.9507015,1.1808317,1.086516,0.7809334,0.42630664,0.23013012,0.21881226,0.33576363,0.52439487,0.69793564,0.7432071,0.6488915,0.55457586,0.59230214,0.8337501,1.2864652,1.9051756,3.4217708,5.304311,6.771862,6.7944975,6.405917,6.0776987,5.802297,5.198677,3.4896781,1.599593,0.73188925,0.38858038,0.26031113,0.241448,0.2565385,0.34330887,0.4640329,0.59607476,0.7432071,0.965792,1.1846043,1.3732355,1.5015048,1.5203679,1.2940104,0.97710985,0.68661773,0.4979865,0.44139713,0.3961256,0.41876137,0.513077,0.69039035,0.9507015,1.1393328,1.2411937,1.2298758,1.0336993,0.5394854,0.24522063,0.116951376,0.11317875,0.18485862,0.28294688,0.32821837,0.36594462,0.38858038,0.42630664,0.52439487,0.6526641,0.79602385,0.9016574,0.95824677,0.97333723,0.95447415,1.0072908,1.1431054,1.3505998,1.6146835,2.0183544,2.4974778,3.0256453,3.5349495,3.9197574,4.134797,4.266839,4.3309736,4.3800178,4.4743333,4.2328854,3.8178966,3.2935016,2.7540162,2.293756,2.093807,2.11267,2.463524,3.2142766,4.398881,5.5683947,6.1418333,6.115425,5.692891,5.2779026,5.1345425,4.9421387,4.5988297,4.112161,3.591539,3.440634,3.5953116,3.9084394,4.247976,4.515832,4.466788,4.376245,4.2291126,4.1008434,4.142342,4.376245,4.821415,5.4363527,6.126743,6.700182,7.062354,7.2623034,7.4207535,7.605612,7.835742,8.36391,8.7600355,8.903395,8.797762,8.567632,8.280911,7.960239,7.647111,7.284939,6.730363,6.1720147,5.7117543,5.2967653,5.0251365,5.1534057,5.621211,5.9305663,5.802297,5.323174,4.930821,4.979865,5.172269,5.564622,6.047518,6.360646,5.934339,5.674028,5.455216,5.406172,5.915476,5.6287565,5.2250857,4.7950063,4.508287,4.617693,4.9534564,5.1835866,5.1458607,4.8063245,4.2706113,3.9197574,3.7386713,3.6066296,3.4066803,3.0105548,2.6144292,2.5087957,2.5616124,2.6597006,2.71629,2.806833,2.8709676,2.927557,2.9954643,3.0897799,3.1463692,3.1840954,3.1840954,3.1312788,3.0105548,2.8822856,2.7653341,2.6483827,2.5012503,2.2786655,2.0372176,1.8787673,1.7919968,1.7467253,1.6976813,1.5279131,1.4222796,1.3317367,1.1959221,0.91674787,0.573439,0.33576363,0.241448,0.28294688,0.41876137,0.5394854,0.6149379,0.63002837,0.5885295,0.51684964,0.4376245,0.422534,0.47157812,0.55457586,0.62248313,0.5093044,0.35462674,0.23767537,0.17731337,0.150905,0.20372175,0.3055826,0.38480774,0.40367088,0.33576363,0.271629,0.30935526,0.48666862,0.73188925,0.8563859,0.6752999,0.4640329,0.30181,0.211267,0.16222288,0.20372175,0.241448,0.30181,0.38858038,0.48666862,0.69793564,0.7696155,0.67152727,0.47912338,0.36594462,0.49421388,0.7054809,0.7507524,0.573439,0.32067314,0.1659955,0.07922512,0.03772625,0.018863125,0.02263575,0.0150905,0.003772625,0.003772625,0.00754525,0.00754525,0.0150905,0.026408374,0.041498873,0.05281675,0.056589376,0.056589376,0.049044125,0.033953626,0.018863125,0.00754525,0.00754525,0.011317875,0.011317875,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,9.971047,10.676529,11.306557,11.672502,11.510279,10.47658,9.0957985,8.707218,8.60913,8.356364,7.752744,7.884786,7.911195,7.9451485,8.107371,8.526133,8.816625,8.843033,8.66572,8.480861,8.620448,8.756263,8.684583,8.560086,8.529905,8.748717,9.099571,8.465771,7.805561,7.5905213,7.8131065,8.27714,7.4018903,6.156924,5.20245,4.9119577,4.538468,4.172523,3.8593953,3.470815,2.6898816,2.04099,1.5958204,1.4109617,1.4071891,1.3656902,1.2411937,1.1091517,0.9242931,0.7054809,0.543258,0.5470306,0.6375736,0.7469798,0.7997965,0.7092535,0.7432071,0.845068,1.0035182,1.2789198,1.8259505,2.173032,2.3918443,2.5238862,2.5804756,2.5616124,2.5616124,2.5691576,2.6634734,2.9049213,3.338773,4.0706625,5.0175915,6.1342883,7.4509344,9.084481,8.443134,7.726336,7.069899,6.3908267,5.3873086,4.847823,4.5988297,4.459243,4.4630156,4.8629136,5.8173876,7.496206,10.250222,13.43809,15.437581,15.373446,12.808062,9.680555,7.020855,4.919503,4.561104,4.22534,3.9725742,3.7160356,3.2142766,2.916239,2.384299,1.9881734,1.8523588,1.8297231,1.6486372,1.3204187,1.0601076,0.9280658,0.8262049,0.73566186,0.56589377,0.422534,0.3470815,0.32821837,0.392353,0.3961256,0.36971724,0.331991,0.29803738,0.3169005,0.34330887,0.331991,0.29049212,0.24899325,0.18485862,0.124496624,0.0754525,0.033953626,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.06413463,0.16976812,0.35839936,0.68661773,1.0374719,1.388326,1.5656394,1.2562841,1.0336993,0.90543,0.8299775,0.8262049,0.9997456,1.2789198,1.1431054,0.9205205,0.77338815,0.68661773,0.77338815,0.7054809,0.60362,0.5470306,0.5998474,0.3055826,0.120724,0.06413463,0.181086,0.5357128,0.5696664,0.44516975,0.43385187,0.51684964,0.3772625,0.211267,0.513077,0.7469798,0.7130261,0.5093044,0.24522063,0.15467763,0.16976812,0.26408374,0.452715,0.362172,0.32067314,0.35462674,0.83752275,2.4786146,2.4484336,1.8297231,1.5165952,1.659955,1.6524098,1.8033148,2.3088465,2.505023,2.3277097,2.3428001,3.3123648,3.8556228,3.6330378,2.4220252,0.1358145,0.45648763,0.573439,0.5017591,0.34330887,0.28294688,0.422534,0.58475685,0.6187105,0.4376245,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.033953626,0.071679875,0.041498873,0.02263575,0.00754525,0.003772625,0.018863125,0.02263575,0.018863125,0.05281675,0.1056335,0.07922512,0.05281675,0.030181,0.0150905,0.0150905,0.026408374,0.06790725,0.056589376,0.0452715,0.0452715,0.03772625,0.10186087,0.12826926,0.150905,0.17731337,0.1961765,0.15467763,0.13958712,0.13958712,0.13958712,0.116951376,0.08677038,0.15845025,0.23390275,0.24899325,0.20372175,0.15467763,0.14335975,0.18485862,0.271629,0.36594462,0.33576363,0.34330887,0.331991,0.30935526,0.34330887,0.31312788,0.26031113,0.21503963,0.16976812,0.08677038,0.03772625,0.03772625,0.11317875,0.23013012,0.26408374,0.19994913,0.150905,0.17354076,0.2867195,0.47157812,1.0714256,1.1619685,1.0336993,0.7884786,0.35085413,0.120724,0.05281675,0.06413463,0.10186087,0.13204187,0.124496624,0.10186087,0.094315626,0.13958712,0.27540162,0.52439487,0.6451189,0.58475685,0.38858038,0.18485862,0.26031113,0.52439487,0.7997965,1.0035182,1.1431054,1.2261031,1.0638802,0.95824677,1.1091517,1.629774,2.4220252,4.0216184,6.0248823,7.8206515,8.567632,8.624221,8.812852,8.627994,7.5603404,5.1043615,2.8709676,1.6825907,1.0072908,0.5885295,0.46026024,0.41121614,0.3734899,0.38480774,0.43385187,0.5017591,0.62248313,0.7997965,1.0299267,1.2864652,1.5430037,1.1619685,0.8262049,0.63002837,0.5696664,0.5470306,0.5885295,0.8639311,1.3996439,1.9730829,2.1353056,1.9542197,1.9051756,1.8863125,1.6939086,1.0299267,0.73188925,0.44139713,0.23013012,0.124496624,0.08677038,0.08677038,0.11317875,0.13204187,0.16222288,0.2867195,0.52062225,0.76584285,0.94692886,1.0186088,0.97333723,0.7997965,0.7092535,0.7054809,0.7922512,0.9620194,1.3505998,1.841041,2.4182527,2.9916916,3.4179983,3.7990334,4.1008434,4.2404304,4.1989317,4.032936,3.7763977,3.4142256,3.006782,2.6182017,2.2899833,2.2183034,2.323937,2.6936543,3.500996,4.98741,6.330465,7.2283497,7.2396674,6.470052,5.583485,4.870459,4.2592936,3.731126,3.3123648,3.0935526,3.1463692,3.5236318,3.9122121,4.146115,4.2102494,3.9763467,3.7537618,3.6141748,3.6028569,3.7575345,3.983892,4.376245,4.927048,5.523123,5.9192486,6.258785,6.356873,6.4511886,6.6662283,7.020855,7.326438,7.854605,8.197914,8.27714,8.348819,8.213005,7.8621507,7.598067,7.462252,7.250985,6.990674,6.579458,6.119198,5.938112,6.579458,6.9491754,7.039718,6.617184,5.87775,5.4212623,5.379763,5.6513925,6.1078796,6.405917,5.9720654,4.647874,4.315883,4.447925,4.798779,5.4212623,4.878004,4.5535583,4.4403796,4.610148,5.198677,5.847569,6.277648,6.2323766,5.643847,4.6554193,3.7877154,3.0407357,2.584248,2.4031622,2.2748928,2.052308,2.0900342,2.233394,2.354118,2.354118,2.3126192,2.3578906,2.474842,2.6219745,2.7389257,2.5917933,2.444661,2.3654358,2.3277097,2.2447119,2.093807,1.9127209,1.7618159,1.6448646,1.5430037,1.4637785,1.4637785,1.4373702,1.3770081,1.3543724,1.3807807,1.6146835,1.7618159,1.5958204,0.965792,0.5772116,0.33576363,0.23767537,0.29426476,0.51684964,0.62625575,0.6375736,0.6413463,0.6375736,0.56589377,0.49044126,0.49044126,0.55457586,0.6451189,0.6790725,0.482896,0.32444575,0.2263575,0.20749438,0.26408374,0.26408374,0.35839936,0.5017591,0.59230214,0.47912338,0.38858038,0.35839936,0.6111652,1.056335,1.2826926,1.1581959,0.8526133,0.56212115,0.3772625,0.29426476,0.422534,0.5093044,0.59607476,0.6752999,0.6752999,0.91297525,0.965792,0.8337501,0.68661773,0.8563859,1.4147344,1.9768555,1.9240388,1.267602,0.60362,0.24899325,0.13204187,0.10186087,0.08299775,0.07922512,0.041498873,0.018863125,0.0150905,0.026408374,0.026408374,0.0150905,0.0150905,0.033953626,0.06413463,0.07922512,0.07922512,0.06790725,0.05281675,0.033953626,0.02263575,0.018863125,0.0150905,0.0150905,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,9.446653,10.250222,11.283921,12.377983,12.770335,11.125471,9.940866,9.167479,9.235386,9.669238,9.110889,8.390318,8.299775,8.59404,9.061845,9.552286,9.978593,9.929549,9.827688,9.914458,10.269085,10.902886,11.155652,11.080199,10.899114,10.970794,10.970794,10.842525,10.340765,9.680555,9.522105,9.205205,8.088508,7.352846,7.254758,7.1566696,6.5568223,6.006019,5.3759904,4.5912848,3.6179473,2.5314314,1.8938577,1.6524098,1.6939086,1.8146327,1.7429527,1.5882751,1.3619176,1.116697,0.94692886,0.8111144,0.7507524,0.76207024,0.8224323,0.87147635,0.8337501,1.0072908,1.3317367,1.7882242,2.4107075,3.1312788,3.712263,4.142342,4.3196554,4.0895257,3.9801195,3.9159849,3.8707132,3.9612563,4.425289,5.2552667,6.4247804,7.1679873,7.352846,7.462252,7.816879,7.4018903,6.752999,6.168242,5.692891,5.0062733,4.881777,5.2250857,5.7570257,6.013564,7.0246277,8.7600355,11.955449,15.546988,16.693865,15.509261,12.083718,8.688355,6.3832817,5.0062733,5.1269975,4.6554193,4.074435,3.651901,3.4330888,2.5917933,2.0862615,1.9164935,2.003264,2.1956677,1.9164935,1.4600059,1.0412445,0.76584285,0.65643674,0.6451189,0.60362,0.543258,0.47157812,0.41121614,0.35085413,0.35462674,0.38480774,0.422534,0.45648763,0.35839936,0.27917424,0.21503963,0.150905,0.0754525,0.05281675,0.0452715,0.041498873,0.030181,0.030181,0.018863125,0.00754525,0.0,0.0,0.0,0.011317875,0.05281675,0.1659955,0.392353,0.7469798,0.88279426,0.8978847,0.8186596,0.7205714,0.73188925,0.7809334,0.77338815,0.6526641,0.46026024,0.35085413,0.29049212,0.30181,0.41121614,0.5772116,0.68661773,0.5885295,0.59230214,0.70170826,0.9318384,1.297783,0.5998474,0.19994913,0.06413463,0.14713238,0.36594462,0.29426476,0.14713238,0.090543,0.14335975,0.1659955,0.181086,0.23767537,0.422534,0.6790725,0.83752275,0.694163,0.6752999,0.5772116,0.32821837,0.0,0.0,0.32821837,0.9393836,1.659955,2.1956677,1.7089992,1.0450171,0.80734175,1.0412445,1.237421,1.3204187,1.0789708,0.8941121,0.9507015,1.2223305,1.9655377,3.259548,3.821669,2.897376,0.26031113,0.392353,0.41876137,0.35085413,0.24899325,0.19994913,0.16222288,0.1358145,0.15845025,0.19240387,0.1056335,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.0452715,0.018863125,0.0,0.00754525,0.030181,0.041498873,0.026408374,0.033953626,0.06790725,0.090543,0.056589376,0.03772625,0.018863125,0.003772625,0.0150905,0.026408374,0.06790725,0.12826926,0.15845025,0.060362,0.03772625,0.049044125,0.13958712,0.2565385,0.24522063,0.18485862,0.18485862,0.21503963,0.23767537,0.21503963,0.116951376,0.19994913,0.27540162,0.23013012,0.0452715,0.13204187,0.19994913,0.241448,0.2565385,0.24522063,0.34330887,0.43007925,0.36971724,0.22258487,0.26031113,0.34330887,0.36594462,0.3055826,0.18485862,0.060362,0.02263575,0.02263575,0.041498873,0.06790725,0.090543,0.12826926,0.18485862,0.26408374,0.31312788,0.23013012,0.19240387,0.32821837,0.9280658,1.5467763,1.0223814,0.21503963,0.060362,0.120724,0.1659955,0.1659955,0.13204187,0.094315626,0.16222288,0.31312788,0.3961256,0.8601585,0.97710985,0.80734175,0.513077,0.36594462,0.41498876,0.5470306,0.7054809,1.1091517,2.2447119,3.1350515,2.7804246,2.1277604,1.6675003,1.4335974,1.690136,3.5500402,5.666483,7.2887115,8.239413,8.424272,9.156161,10.084227,9.525878,4.4705606,2.8709676,2.6182017,2.4295704,1.8900851,1.448688,1.0940613,0.7884786,0.56212115,0.41876137,0.32067314,0.271629,0.38858038,0.845068,1.750498,3.1425967,1.81086,1.0148361,0.694163,0.7054809,0.77716076,1.2298758,2.0183544,3.4745877,4.6742826,3.4783602,1.6976813,1.1242423,1.146878,1.3807807,1.6637276,1.8825399,1.3317367,0.6488915,0.19994913,0.0754525,0.06413463,0.060362,0.056589376,0.07922512,0.21503963,0.31312788,0.392353,0.48666862,0.6073926,0.7167987,0.77716076,0.72811663,0.68661773,0.7167987,0.83752275,1.0714256,1.4147344,1.8033148,2.2220762,2.686109,3.1727777,3.5236318,3.731126,3.7763977,3.6179473,3.410453,3.1840954,2.9464202,2.7540162,2.7313805,2.8030603,2.9237845,3.1425967,3.519859,4.1197066,5.119452,6.398372,7.1604424,6.952948,5.6476197,4.6554193,3.832987,3.187868,2.776652,2.71629,2.8747404,3.1350515,3.3915899,3.5538127,3.5387223,3.440634,3.3350005,3.2859564,3.3312278,3.4632697,3.7688525,3.9461658,4.0480266,4.112161,4.134797,4.67051,4.7874613,4.6252384,4.7006907,5.9192486,6.7756343,7.383027,7.6584287,7.677292,7.6886096,7.54525,7.1302614,7.1264887,7.567886,7.8734684,7.4584794,7.3377557,7.4094353,7.6282477,7.9941926,7.360391,6.6624556,5.9494295,5.4212623,5.43258,5.9192486,6.4549613,6.515323,5.9003854,4.715781,3.6669915,3.3576362,3.2029586,2.9803739,2.806833,2.8332415,3.059599,3.259548,3.3048196,3.1576872,3.8669407,4.2894745,4.395108,3.9688015,2.6408374,2.0183544,1.6976813,1.5015048,1.3807807,1.418507,1.478869,1.4939595,1.6524098,1.9127209,1.9994912,1.5467763,1.4335974,1.478869,1.5656394,1.6637276,1.5165952,1.4147344,1.3732355,1.4034165,1.5241405,1.5505489,1.539231,1.4298248,1.2864652,1.297783,1.4449154,1.7278622,1.7769064,1.5882751,1.5241405,1.9542197,3.1124156,3.7462165,3.1237335,1.0374719,0.7205714,0.49421388,0.35462674,0.29426476,0.32067314,0.38103512,0.47157812,0.694163,0.94315624,0.87147635,0.69793564,0.63002837,0.58475685,0.5319401,0.45648763,0.27540162,0.28294688,0.38858038,0.52062225,0.65643674,0.41121614,0.2678564,0.19994913,0.211267,0.32067314,0.45648763,0.5885295,0.72811663,0.91674787,1.2223305,1.3430545,1.0148361,0.7054809,0.6149379,0.68661773,0.9808825,1.20724,1.3128735,1.2600567,1.0525624,0.88279426,0.7582976,0.7092535,0.9922004,2.0900342,3.3236825,4.1536603,3.4896781,1.7014539,0.6413463,0.18863125,0.18485862,0.25276586,0.2263575,0.150905,0.06790725,0.03772625,0.049044125,0.08677038,0.1358145,0.0754525,0.041498873,0.03772625,0.056589376,0.090543,0.090543,0.071679875,0.060362,0.056589376,0.0452715,0.033953626,0.02263575,0.00754525,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,8.00551,8.850578,9.314611,9.710737,10.001229,9.81637,9.178797,9.027891,9.265567,9.691874,10.001229,9.574923,9.623966,10.20495,10.967021,11.1631975,11.570641,11.883769,11.959221,11.898859,12.038446,12.204442,12.559069,12.808062,12.875969,12.913695,12.932558,12.66093,12.200669,11.593277,10.827434,9.680555,8.835487,8.541223,8.6732645,8.729855,8.688355,8.401636,8.050782,7.7414265,7.484888,7.0246277,6.0362,4.8138695,3.5538127,2.3767538,2.1088974,1.8825399,1.690136,1.5316857,1.4109617,1.267602,1.1355602,1.086516,1.1129243,1.1506506,1.2223305,1.4147344,1.7240896,2.1768045,2.837014,3.8405323,4.568649,5.0251365,5.198677,5.0666356,5.160951,5.142088,5.0477724,5.070408,5.534441,6.375736,7.2962565,7.635793,7.4773426,7.6584287,7.8244243,7.541477,7.2283497,7.020855,6.741681,6.273875,6.2814207,6.56814,6.9982195,7.488661,8.677037,10.699164,13.5663595,16.195879,16.437326,14.441608,11.208468,8.269594,6.2927384,5.0779533,4.6327834,4.0782075,3.640583,3.3689542,3.138824,2.5238862,2.2862108,2.2862108,2.4333432,2.686109,2.082489,1.5618668,1.2223305,1.0299267,0.80356914,0.70170826,0.663982,0.694163,0.7432071,0.694163,0.5357128,0.46026024,0.4074435,0.3470815,0.2867195,0.20749438,0.14713238,0.10940613,0.090543,0.0754525,0.060362,0.041498873,0.026408374,0.0150905,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.030181,0.14335975,0.30181,0.482896,0.663982,0.543258,0.45648763,0.4074435,0.41121614,0.5017591,0.5093044,0.48666862,0.43007925,0.34330887,0.25276586,0.42630664,0.87147635,0.97710985,0.68661773,0.5017591,0.47535074,0.5017591,0.543258,0.58098423,0.62625575,0.29049212,0.20749438,0.29049212,0.482896,0.73188925,0.5319401,0.2867195,0.20372175,0.31312788,0.47157812,0.6413463,0.84884065,0.9280658,0.8337501,0.63002837,0.241448,0.13958712,0.116951376,0.06790725,0.011317875,0.23767537,0.36594462,0.47912338,0.76584285,1.5241405,1.2336484,0.7205714,0.5017591,0.6488915,0.79602385,0.8337501,0.77338815,0.814887,1.0186088,1.3053282,1.7278622,2.516341,2.806833,2.0862615,0.211267,0.49044126,0.6187105,0.6149379,0.573439,0.663982,0.5772116,0.41876137,0.21503963,0.03772625,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.026408374,0.033953626,0.02263575,0.02263575,0.018863125,0.011317875,0.00754525,0.00754525,0.018863125,0.03772625,0.049044125,0.056589376,0.026408374,0.011317875,0.00754525,0.0150905,0.026408374,0.041498873,0.071679875,0.09808825,0.1056335,0.08677038,0.10186087,0.120724,0.14713238,0.15845025,0.14713238,0.15467763,0.1659955,0.17731337,0.17354076,0.13958712,0.08299775,0.18485862,0.44139713,0.7130261,0.7167987,0.6187105,0.45648763,0.31312788,0.21881226,0.14713238,0.14713238,0.1659955,0.15467763,0.124496624,0.150905,0.2263575,0.23767537,0.20372175,0.14713238,0.08677038,0.049044125,0.06413463,0.116951376,0.15467763,0.090543,0.07922512,0.11317875,0.331991,0.63002837,0.6790725,0.59607476,0.55080324,0.62625575,0.73566186,0.6187105,0.28294688,0.16976812,0.120724,0.094315626,0.19240387,0.14713238,0.090543,0.094315626,0.24899325,0.663982,1.0110635,0.98842776,0.8865669,0.8337501,0.7922512,0.73566186,0.7507524,1.0751982,1.7354075,2.546522,2.5012503,2.2069857,1.750498,1.3543724,1.3845534,2.2484846,3.5839937,4.9119577,5.945657,6.6058664,7.5301595,9.046755,8.846806,6.4247804,3.078462,1.8599042,2.2598023,2.7540162,2.505023,1.3505998,1.2223305,1.0638802,0.94315624,0.8639311,0.784706,0.7167987,0.68661773,0.7507524,0.9620194,1.3845534,1.237421,1.1053791,1.0035182,0.94315624,0.935611,1.1846043,1.4373702,1.8146327,2.161714,2.0862615,1.9768555,1.81086,1.4411428,1.026154,1.0525624,0.88279426,0.6149379,0.3772625,0.21881226,0.124496624,0.0754525,0.060362,0.06790725,0.09808825,0.150905,0.17354076,0.150905,0.16222288,0.23013012,0.35085413,0.52062225,0.6375736,0.7092535,0.7809334,0.91297525,1.1053791,1.3430545,1.8561316,2.5540671,3.0256453,3.1652324,3.2218218,3.1124156,2.8596497,2.6031113,2.727608,2.7917426,2.7992878,2.7917426,2.8030603,2.9766011,3.1124156,3.199186,3.2859564,3.4745877,3.9461658,4.5837393,5.1835866,5.5080323,5.304311,4.9119577,4.395108,3.9008942,3.5047686,3.229367,3.1237335,3.0256453,2.9049213,2.776652,2.686109,2.7351532,2.8256962,2.957738,3.1161883,3.2670932,3.3689542,3.361409,3.3312278,3.289729,3.1954134,3.1765501,3.350091,3.6254926,3.9989824,4.564876,5.1269975,5.8136153,6.4247804,6.790725,6.7643166,6.820906,6.930312,7.2472124,7.677292,7.8734684,7.967784,8.578949,8.846806,8.465771,7.6886096,6.7039547,6.1606965,6.1003346,6.4511886,7.032173,6.319147,6.8661776,8.013056,8.2507305,5.240176,3.731126,3.1765501,2.9652832,2.7691069,2.5389767,2.4861598,2.493705,2.5087957,2.5502944,2.7087448,3.0143273,2.9124665,2.637065,2.3013012,1.9202662,1.6976813,1.5580941,1.4411428,1.3392819,1.3091009,1.3015556,1.3204187,1.3619176,1.4071891,1.4260522,1.2940104,1.1846043,1.1280149,1.1393328,1.1883769,1.1883769,1.297783,1.4675511,1.6373192,1.7580433,1.7127718,1.6976813,1.7731338,1.8787673,1.8334957,1.8523588,1.931584,2.0258996,2.0975795,2.0749438,2.1692593,2.7917426,2.9313297,2.2069857,0.8903395,0.70170826,0.66020936,0.67152727,0.633801,0.44139713,0.3772625,0.43385187,0.68661773,1.0186088,1.1016065,0.98842776,0.8601585,0.7092535,0.5394854,0.3470815,0.19240387,0.211267,0.2867195,0.35085413,0.38858038,0.33953625,0.29426476,0.2678564,0.2867195,0.4074435,0.46026024,0.46026024,0.4376245,0.482896,0.7205714,1.026154,1.2034674,1.1544232,0.97333723,0.9318384,1.056335,1.2902378,1.4373702,1.3505998,0.91674787,0.94315624,1.4600059,2.4220252,3.6971724,5.070408,5.5495315,4.749735,3.0671442,1.418507,1.2147852,1.8561316,2.2220762,2.5125682,2.795515,2.9954643,2.0145817,1.3694628,0.94692886,0.633801,0.32067314,0.0754525,0.00754525,0.00754525,0.0150905,0.030181,0.041498873,0.0452715,0.049044125,0.049044125,0.056589376,0.0452715,0.041498873,0.030181,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.7643166,7.8319697,8.812852,9.359882,9.488152,9.582467,9.220296,9.265567,9.752235,10.487898,11.027383,11.129244,11.223559,11.638548,12.347801,12.966512,13.59654,13.947394,13.924759,13.626721,13.332457,13.185325,13.177779,13.298503,13.434318,13.377728,13.189097,13.045737,12.717519,12.132762,11.400873,10.872705,10.005001,9.175024,8.575176,8.216777,8.469543,8.605357,8.59404,8.741172,9.680555,10.231359,10.095545,9.424017,8.356364,7.032173,5.8136153,4.82896,3.8556228,2.8936033,2.1315331,1.8448136,1.7014539,1.690136,1.7618159,1.8334957,1.9693103,2.214531,2.6295197,3.289729,4.2894745,5.372218,6.198423,6.56814,6.5266414,6.3455553,6.307829,6.1531515,6.039973,6.1078796,6.5002327,7.326438,8.114917,8.480861,8.492179,8.66572,8.409182,7.8998766,7.7716074,8.016829,7.9828744,7.6131573,7.4509344,7.5905213,8.065872,8.865668,10.552032,13.087236,15.403628,16.505234,15.482853,12.90615,9.986138,7.4169807,5.583485,4.5761943,4.085753,3.7273536,3.4632697,3.2331395,2.957738,2.5502944,2.5012503,2.4786146,2.354118,2.2107582,1.8863125,1.4939595,1.1506506,0.91674787,0.7922512,0.7432071,0.7167987,0.7167987,0.73188925,0.72811663,0.63002837,0.5394854,0.452715,0.36594462,0.27917424,0.17731337,0.116951376,0.07922512,0.056589376,0.056589376,0.0452715,0.030181,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.06413463,0.1659955,0.27540162,0.36971724,0.43007925,0.29803738,0.271629,0.30181,0.36594462,0.47157812,0.41876137,0.36594462,0.3169005,0.27540162,0.24899325,0.392353,0.69039035,0.76207024,0.5772116,0.4678055,0.4678055,0.5055317,0.47912338,0.3734899,0.24899325,0.1358145,0.35462674,0.6752999,0.88279426,0.79602385,0.513077,0.3470815,0.44516975,0.6488915,0.49421388,0.4678055,0.6187105,0.7054809,0.66020936,0.6073926,0.543258,0.38103512,0.21503963,0.094315626,0.033953626,0.31312788,0.39989826,0.3961256,0.5017591,1.0299267,0.8224323,0.49044126,0.38103512,0.5394854,0.694163,0.8224323,0.9393836,1.1355602,1.4562333,1.8938577,2.5427492,2.4597516,1.9693103,1.2411937,0.27917424,0.44516975,0.5357128,0.5583485,0.5357128,0.513077,0.422534,0.30181,0.13958712,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.026408374,0.018863125,0.011317875,0.00754525,0.0150905,0.018863125,0.011317875,0.0,0.0,0.011317875,0.026408374,0.03772625,0.0452715,0.02263575,0.011317875,0.0150905,0.026408374,0.030181,0.033953626,0.049044125,0.060362,0.06413463,0.06413463,0.08677038,0.10186087,0.10186087,0.090543,0.094315626,0.11317875,0.124496624,0.13958712,0.14335975,0.120724,0.094315626,0.14713238,0.33576363,0.58098423,0.663982,0.56212115,0.36594462,0.22258487,0.19240387,0.22258487,0.2565385,0.241448,0.18863125,0.124496624,0.1056335,0.19240387,0.26031113,0.2565385,0.18485862,0.10186087,0.056589376,0.05281675,0.094315626,0.150905,0.14713238,0.10186087,0.11317875,0.24522063,0.42630664,0.49044126,0.452715,0.422534,0.3961256,0.362172,0.29803738,0.211267,0.21503963,0.16976812,0.07922512,0.1056335,0.08677038,0.08677038,0.10940613,0.21881226,0.52062225,0.845068,1.2185578,1.5769572,1.8561316,1.9994912,2.0447628,2.0447628,2.0447628,2.0598533,2.0749438,1.9353566,1.9278114,2.0787163,2.3126192,2.4899325,2.5729303,3.3764994,4.4630156,5.458988,6.0211096,6.8473144,7.6622014,7.2887115,5.3759904,2.4031622,1.4034165,1.6825907,2.3993895,2.7011995,1.720317,1.448688,1.2638294,1.1657411,1.1431054,1.1581959,1.3317367,1.4222796,1.5354583,1.7316349,2.0636258,2.2447119,2.252257,2.0900342,1.8146327,1.5241405,1.5015048,1.4977322,1.4939595,1.4939595,1.50905,1.5241405,1.3619176,1.0902886,0.8224323,0.72811663,0.5319401,0.44139713,0.36971724,0.26031113,0.10940613,0.056589376,0.060362,0.09808825,0.1659955,0.28294688,0.25276586,0.16222288,0.124496624,0.16976812,0.241448,0.3470815,0.4979865,0.65643674,0.8224323,1.0223814,1.2487389,1.4449154,1.720317,2.033445,2.1881225,2.191895,2.1994405,2.173032,2.123988,2.1202152,2.3578906,2.625747,2.8219235,2.9200118,2.9501927,2.9351022,2.8558772,2.8106055,2.8256962,2.8898308,2.9916916,3.2482302,3.5802212,3.904667,4.13857,4.2819295,4.293247,4.187614,4.002755,3.8065786,3.5689032,3.2482302,2.867195,2.4861598,2.2069857,2.1466236,2.1994405,2.305074,2.4182527,2.5314314,2.6898816,2.7313805,2.7087448,2.686109,2.7313805,2.8936033,3.1539145,3.5160866,3.9273026,4.2706113,4.4441524,5.1647234,5.824933,6.066381,5.7419353,6.066381,6.587003,7.062354,7.375482,7.564113,7.8621507,8.299775,8.537451,8.341274,7.594294,7.3415284,7.3905725,7.273621,6.9454026,6.809588,6.379509,6.40969,6.9944468,7.333983,5.7192993,3.8480775,3.0407357,2.8030603,2.8332415,3.0218725,2.5616124,2.191895,2.0108092,2.0296721,2.1805773,2.263575,2.1541688,2.0183544,1.9164935,1.8221779,1.8033148,1.7165444,1.5731846,1.4034165,1.2713746,1.2411937,1.2261031,1.2223305,1.2298758,1.2713746,1.20724,1.1129243,1.0638802,1.0827434,1.1506506,1.2449663,1.3920987,1.5543215,1.6863633,1.7316349,1.7731338,1.8674494,2.0258996,2.191895,2.2258487,2.1692593,2.1805773,2.2748928,2.3390274,2.1654868,2.4408884,3.0860074,3.259548,2.6144292,1.2864652,0.8563859,0.8978847,1.1317875,1.3656902,1.4901869,1.1129243,1.0336993,1.3619176,1.8259505,1.7731338,1.3468271,1.0412445,0.8639311,0.7582976,0.6413463,0.56589377,0.73566186,0.9318384,1.0186088,0.94315624,0.5998474,0.52062225,0.5998474,0.72811663,0.8224323,0.9016574,0.9695646,0.9620194,0.91297525,0.935611,1.2940104,1.4373702,1.4147344,1.3392819,1.3770081,2.082489,2.5540671,2.4710693,1.8749946,1.1581959,1.6222287,2.6597006,3.9725742,5.1571784,5.7117543,5.2892203,3.85185,2.252257,1.2298758,1.4034165,2.8030603,3.9650288,4.255521,3.5764484,2.335255,1.237421,0.724344,0.47912338,0.30935526,0.14713238,0.030181,0.0,0.0,0.0,0.00754525,0.011317875,0.0150905,0.02263575,0.030181,0.033953626,0.03772625,0.03772625,0.030181,0.02263575,0.02263575,0.011317875,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.719554,5.9720654,7.303802,8.22055,8.771353,9.563604,10.016319,10.250222,10.431308,10.70671,11.204697,11.695138,11.868678,12.396846,13.422999,14.539697,15.286676,16.022339,16.350557,16.150608,15.562078,14.988639,14.622695,14.505743,14.471789,14.154889,13.936077,13.962485,13.72481,13.102326,12.336484,11.864905,10.891568,9.9257765,9.231613,8.835487,8.929804,9.016574,8.933576,8.971302,9.876732,10.589758,10.993429,11.0613365,10.819888,10.344538,9.016574,7.6131573,5.9909286,4.3083377,3.0445085,2.584248,2.3805263,2.3578906,2.4522061,2.6031113,2.8558772,3.240685,3.8065786,4.6327834,5.8211603,6.8699503,7.6848373,7.986647,7.805561,7.5112963,7.2887115,7.1076255,7.066127,7.224577,7.586749,8.182823,8.654402,8.922258,9.012801,9.016574,8.726082,8.318638,8.262049,8.473316,8.307321,7.8998766,7.598067,7.779153,8.5563135,9.774872,11.774363,14.596286,16.286423,15.992157,14.000212,11.295239,8.778898,6.63982,5.093044,4.3800178,3.9461658,3.6556737,3.4142256,3.2218218,3.1652324,3.0407357,2.916239,2.6068838,2.123988,1.6750455,1.5279131,1.2487389,0.9620194,0.7809334,0.7922512,0.88279426,0.90543,0.87902164,0.8262049,0.7809334,0.70170826,0.5998474,0.49044126,0.392353,0.3055826,0.211267,0.13958712,0.08677038,0.060362,0.05281675,0.030181,0.0150905,0.003772625,0.0,0.0,0.0,0.003772625,0.00754525,0.018863125,0.049044125,0.094315626,0.14713238,0.19994913,0.23390275,0.24899325,0.18863125,0.21881226,0.29426476,0.392353,0.5017591,0.40367088,0.331991,0.271629,0.2263575,0.22258487,0.31312788,0.44894236,0.5583485,0.5885295,0.5281675,0.48666862,0.513077,0.452715,0.28294688,0.124496624,0.150905,0.5470306,0.98842776,1.2034674,0.97333723,0.62248313,0.4678055,0.5885295,0.79602385,0.63002837,0.49044126,0.4376245,0.392353,0.362172,0.4376245,0.6111652,0.43385187,0.21503963,0.14335975,0.28294688,0.331991,0.36971724,0.422534,0.4979865,0.6073926,0.513077,0.40367088,0.38858038,0.5093044,0.7092535,0.94692886,1.1883769,1.4600059,1.7919968,2.2183034,2.8143783,2.3767538,1.6222287,0.9393836,0.3961256,0.39989826,0.38858038,0.3470815,0.29049212,0.27917424,0.23767537,0.19240387,0.10186087,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.018863125,0.00754525,0.0,0.0,0.00754525,0.0150905,0.0150905,0.00754525,0.011317875,0.02263575,0.030181,0.033953626,0.041498873,0.041498873,0.026408374,0.018863125,0.02263575,0.02263575,0.03772625,0.041498873,0.0452715,0.056589376,0.0754525,0.094315626,0.094315626,0.0754525,0.060362,0.0754525,0.094315626,0.10186087,0.1056335,0.1056335,0.1056335,0.13958712,0.18863125,0.271629,0.35462674,0.3734899,0.362172,0.30181,0.27540162,0.29803738,0.32821837,0.362172,0.33576363,0.24899325,0.14713238,0.09808825,0.15467763,0.24899325,0.2678564,0.18863125,0.094315626,0.060362,0.049044125,0.071679875,0.120724,0.15845025,0.181086,0.20749438,0.25276586,0.30935526,0.331991,0.3470815,0.38858038,0.35462674,0.23767537,0.13958712,0.150905,0.18863125,0.17354076,0.1056335,0.08299775,0.08299775,0.120724,0.17731337,0.27540162,0.45648763,0.6073926,0.97333723,1.3958713,1.7467253,1.9391292,2.033445,2.033445,1.8523588,1.5241405,1.1921495,1.1016065,1.237421,1.690136,2.3465726,2.8747404,3.500996,4.3611546,4.6327834,4.4630156,4.9534564,6.277648,7.654656,7.8508325,6.488915,4.044254,3.2784111,3.0218725,3.1010978,3.1199608,2.4522061,1.7127718,1.3392819,1.2185578,1.2638294,1.3958713,1.8146327,2.263575,2.6483827,3.0935526,3.9348478,4.5724216,5.100589,5.062863,4.4139714,3.519859,2.7200627,2.2711203,1.9730829,1.7354075,1.5769572,1.3468271,1.086516,0.8941121,0.7696155,0.63002837,0.51684964,0.48666862,0.44894236,0.35085413,0.18485862,0.07922512,0.0754525,0.1358145,0.24899325,0.422534,0.482896,0.38480774,0.30181,0.31312788,0.392353,0.331991,0.3772625,0.5093044,0.70170826,0.935611,1.1544232,1.3053282,1.3807807,1.3920987,1.3770081,1.4071891,1.5467763,1.7429527,1.9466745,2.1202152,2.3805263,2.7426984,3.0709167,3.2935016,3.4029078,3.127506,2.7615614,2.4786146,2.3390274,2.3088465,2.2447119,2.2598023,2.3428001,2.4974778,2.7540162,3.048281,3.3538637,3.5538127,3.62172,3.6330378,3.4859054,3.2444575,2.9313297,2.565385,2.1768045,1.9542197,1.8448136,1.7957695,1.7882242,1.8297231,1.9881734,2.0560806,2.0787163,2.142851,2.3578906,2.8294687,3.218049,3.5538127,3.8065786,3.8895764,4.1989317,4.8025517,5.070408,4.8629136,4.5460134,5.010046,5.7796617,6.330465,6.5756855,6.8774953,7.364164,7.4697976,7.484888,7.4094353,6.960493,7.2585306,7.5527954,7.24344,6.379509,5.66271,5.5759397,5.4778514,5.66271,5.945657,5.6513925,4.508287,4.123479,3.874486,3.5274043,3.2784111,2.625747,2.0560806,1.7127718,1.6184561,1.6524098,1.659955,1.6373192,1.6260014,1.6222287,1.5731846,1.6071383,1.5618668,1.448688,1.2940104,1.1695137,1.1355602,1.1393328,1.1355602,1.1280149,1.1695137,1.116697,1.0902886,1.1242423,1.2336484,1.4071891,1.5807298,1.7240896,1.8259505,1.8599042,1.81086,1.8787673,2.052308,2.2711203,2.463524,2.5238862,2.4031622,2.3314822,2.3126192,2.2975287,2.1805773,2.5238862,3.0143273,2.9916916,2.2975287,1.267602,0.97333723,1.2525115,1.7580433,2.1805773,2.2296214,2.0900342,2.1202152,2.293756,2.4559789,2.3088465,2.1202152,2.003264,1.81086,1.4713237,0.9808825,1.0601076,1.3543724,1.6335466,1.7693611,1.7354075,1.237421,0.9393836,0.8601585,0.8903395,0.8262049,0.83752275,0.97710985,1.20724,1.5128226,1.9051756,2.0560806,1.8070874,1.5203679,1.3996439,1.478869,2.4220252,2.9803739,2.7917426,2.0145817,1.3128735,1.8372684,3.0105548,4.304565,5.2175403,5.27413,4.3422914,2.7804246,1.4750963,0.90543,1.1431054,2.7804246,4.187614,4.508287,3.5236318,1.6373192,0.62248313,0.2678564,0.24899325,0.33953625,0.4074435,0.35462674,0.3169005,0.33576363,0.3470815,0.1659955,0.060362,0.018863125,0.033953626,0.0754525,0.071679875,0.030181,0.02263575,0.02263575,0.026408374,0.030181,0.02263575,0.02263575,0.0150905,0.003772625,0.0,0.003772625,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.8332415,3.9612563,4.8968673,5.904158,7.213259,9.039209,10.567122,11.174516,10.974566,10.570895,11.038701,11.578186,11.891314,12.792972,14.298248,15.645076,16.33924,17.523844,18.546225,18.912169,18.316093,17.214487,16.905132,16.803272,16.51278,15.833707,15.679029,15.731846,15.554533,14.962231,14.030393,13.011784,12.15917,11.7555,11.763044,11.7894535,11.506506,11.117926,10.608622,10.121953,9.940866,10.057818,10.269085,10.536942,10.846297,11.212241,10.559577,9.235386,7.364164,5.3910813,4.0895257,3.5085413,3.218049,3.1765501,3.3236825,3.5990841,3.983892,4.429062,5.032682,5.8702044,6.9944468,7.911195,8.560086,8.793989,8.654402,8.36391,8.209232,8.284684,8.582722,8.9788475,9.224068,9.246704,9.107117,9.06939,9.122208,8.967529,8.684583,8.646856,8.695901,8.624221,8.197914,7.865923,7.7112455,8.141325,9.318384,11.151879,13.04951,15.358356,16.056292,14.683057,12.37421,10.140816,8.013056,6.258785,5.081726,4.6290107,4.3724723,3.9688015,3.519859,3.259548,3.5424948,3.7801702,3.5802212,2.9351022,2.082489,1.5165952,1.2336484,1.0110635,0.87902164,0.8563859,0.94692886,1.1921495,1.3392819,1.3807807,1.3204187,1.1657411,0.87147635,0.6413463,0.47912338,0.36594462,0.28294688,0.23390275,0.15467763,0.10186087,0.07922512,0.056589376,0.026408374,0.00754525,0.003772625,0.003772625,0.0,0.0,0.011317875,0.02263575,0.041498873,0.0754525,0.1056335,0.1056335,0.120724,0.15467763,0.17354076,0.18485862,0.21503963,0.28294688,0.38103512,0.482896,0.3961256,0.36594462,0.34330887,0.29049212,0.181086,0.25276586,0.3734899,0.5357128,0.6526641,0.5583485,0.45648763,0.44139713,0.392353,0.2867195,0.20372175,0.30181,0.6375736,0.965792,1.1242423,1.026154,0.7394345,0.55457586,0.5055317,0.5885295,0.7432071,0.69039035,0.47157812,0.24522063,0.124496624,0.19994913,0.38103512,0.20749438,0.0452715,0.120724,0.52439487,0.32821837,0.271629,0.3470815,0.41876137,0.24522063,0.2867195,0.3734899,0.41498876,0.47157812,0.7205714,1.0638802,1.4713237,1.7769064,1.9542197,2.1088974,2.2560298,2.0296721,1.6033657,1.056335,0.392353,0.36594462,0.29049212,0.14713238,0.05281675,0.2678564,0.29426476,0.2565385,0.1358145,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.011317875,0.0150905,0.030181,0.03772625,0.03772625,0.030181,0.033953626,0.06790725,0.041498873,0.018863125,0.0150905,0.018863125,0.0452715,0.05281675,0.056589376,0.06413463,0.1056335,0.10940613,0.10186087,0.08677038,0.07922512,0.1056335,0.124496624,0.11317875,0.094315626,0.08677038,0.124496624,0.20372175,0.2678564,0.28294688,0.23390275,0.1358145,0.25276586,0.4074435,0.49044126,0.46026024,0.3470815,0.3169005,0.32067314,0.27540162,0.181086,0.120724,0.116951376,0.18485862,0.211267,0.16222288,0.071679875,0.060362,0.071679875,0.11317875,0.15467763,0.1659955,0.271629,0.32821837,0.3734899,0.41121614,0.392353,0.38103512,0.47157812,0.45648763,0.3470815,0.35839936,0.33953625,0.29049212,0.25276586,0.24522063,0.24899325,0.25276586,0.28294688,0.33576363,0.42630664,0.55457586,0.43007925,0.35839936,0.43007925,0.59607476,0.7167987,0.7884786,0.77716076,0.69039035,0.56212115,0.47535074,0.42630664,0.543258,0.7922512,1.2110126,1.931584,3.874486,5.0741806,4.644101,3.451952,4.104616,6.145606,8.99771,9.906913,8.439363,6.4926877,6.043745,5.7683434,5.6325293,5.243949,3.8405323,2.3163917,1.5316857,1.2713746,1.327964,1.4713237,1.8825399,2.595566,3.2972744,4.1083884,5.613666,6.7756343,8.073418,8.533678,7.907422,6.696409,5.311856,4.3649273,3.4972234,2.7011995,2.3088465,1.9089483,1.4864142,1.1393328,0.8978847,0.73188925,0.62625575,0.6073926,0.6149379,0.59230214,0.5093044,0.26408374,0.1659955,0.18485862,0.29803738,0.47535074,0.66775465,0.62248313,0.5281675,0.5093044,0.62248313,0.41498876,0.32821837,0.35839936,0.482896,0.6752999,0.7997965,0.875249,0.8978847,0.8941121,0.9205205,1.0299267,1.3392819,1.7278622,2.0749438,2.2711203,2.5087957,2.7804246,3.1237335,3.4934506,3.7499893,3.3915899,2.8785129,2.3918443,2.0598533,1.9542197,1.8372684,1.7089992,1.6260014,1.6260014,1.690136,1.7769064,2.0258996,2.323937,2.6031113,2.8332415,2.957738,3.097325,3.1954134,3.1727777,2.9237845,2.5389767,2.191895,1.9127209,1.7278622,1.6863633,1.7240896,1.7165444,1.7240896,1.8259505,2.0975795,2.625747,3.0709167,3.3689542,3.451952,3.2670932,3.9386206,4.236658,3.9574835,3.410453,3.429316,3.9197574,4.7120085,5.281675,5.6023483,6.1305156,6.820906,6.9227667,6.8058157,6.6134114,6.247467,6.2851934,6.432326,6.2021956,5.534441,4.7836885,4.7572803,4.9949555,5.353355,5.617439,5.462761,5.7494807,6.2135134,5.847569,4.5535583,3.1350515,2.4899325,1.9806281,1.6033657,1.3656902,1.2826926,1.2826926,1.2638294,1.2298758,1.1846043,1.1619685,1.1619685,1.1657411,1.1544232,1.1355602,1.1355602,1.116697,1.1355602,1.1280149,1.1016065,1.1053791,1.1129243,1.1808317,1.297783,1.4713237,1.720317,1.9353566,2.0749438,2.1315331,2.1013522,1.9994912,2.0070364,2.1843498,2.4974778,2.7879698,2.7615614,2.5804756,2.4597516,2.3390274,2.2409391,2.2711203,2.2711203,2.2560298,1.81086,1.0827434,0.7922512,1.3128735,2.0975795,2.795515,3.1463692,2.969056,3.2444575,3.1312788,2.8256962,2.5502944,2.5804756,3.1048703,3.2972744,3.0633714,2.4371157,1.5920477,1.6712729,1.8523588,2.022127,2.1051247,2.093807,1.720317,1.237421,0.8978847,0.7205714,0.482896,0.36971724,0.58475685,1.146878,1.9881734,2.9464202,2.595566,1.9051756,1.3166461,1.0714256,1.2223305,1.8787673,2.2673476,2.0900342,1.4977322,1.0902886,1.3015556,2.203213,3.2369123,3.9914372,4.1989317,3.4217708,2.0749438,0.97333723,0.513077,0.6790725,2.2711203,3.289729,3.5839937,3.108643,1.8863125,0.97710985,0.5772116,0.58475685,0.8186596,1.0223814,0.9922004,0.8601585,0.875249,0.95447415,0.68661773,0.32444575,0.13204187,0.10186087,0.14713238,0.1358145,0.030181,0.00754525,0.011317875,0.0150905,0.02263575,0.026408374,0.026408374,0.02263575,0.0150905,0.003772625,0.011317875,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.0291634,4.406426,4.2894745,4.749735,5.9984736,7.4169807,8.892077,10.03141,11.019837,11.891314,12.528888,12.736382,13.20796,13.947394,14.950912,16.218515,16.905132,17.37671,18.493408,19.768555,19.379974,17.912424,18.444365,18.987621,18.689585,17.82188,17.248442,17.05981,17.022083,16.852316,16.203424,15.935568,15.841252,15.939341,16.146835,16.28265,16.03743,15.445127,14.766054,14.211478,13.932304,14.124708,14.109617,13.909668,13.505998,12.849561,11.981857,10.499215,8.390318,6.224831,5.1873593,4.6252384,4.38379,4.538468,4.9760923,5.4174895,5.783434,5.8211603,6.1003346,6.8359966,7.8734684,8.495952,8.771353,8.820397,8.805306,8.926031,9.42779,10.110635,11.257513,12.336484,11.993175,11.042474,10.069136,9.88805,10.382264,10.529396,8.918486,8.7600355,9.193887,9.623966,9.733373,10.076681,10.574668,11.216014,12.457208,15.226315,16.65614,16.969267,15.588487,13.094781,11.216014,10.103089,8.197914,6.432326,5.2779026,4.715781,5.1798143,4.847823,4.002755,3.2255943,3.3727267,3.9688015,4.395108,3.85185,2.5540671,1.7240896,1.2864652,1.1921495,1.2185578,1.2638294,1.3732355,1.7278622,2.0900342,2.3465726,2.4107075,2.2258487,1.3505998,0.67152727,0.33576363,0.271629,0.19994913,0.1358145,0.094315626,0.071679875,0.056589376,0.0452715,0.033953626,0.02263575,0.0150905,0.011317875,0.0,0.0,0.018863125,0.03772625,0.05281675,0.0754525,0.0754525,0.049044125,0.049044125,0.08677038,0.1358145,0.18485862,0.23390275,0.28294688,0.32444575,0.33576363,0.33576363,0.5281675,0.7092535,0.6790725,0.23013012,0.20372175,0.23390275,0.26408374,0.29049212,0.35085413,0.32821837,0.23013012,0.22258487,0.32821837,0.41121614,0.5093044,0.44139713,0.30935526,0.16976812,0.060362,0.24522063,0.271629,0.181086,0.08677038,0.18485862,0.20749438,0.17731337,0.10940613,0.116951376,0.3961256,0.7130261,0.5017591,0.2263575,0.09808825,0.060362,0.29426476,0.13958712,0.0,0.0,0.0,0.071679875,0.1659955,0.2867195,0.4640329,0.73188925,1.2336484,2.0900342,2.4672968,2.2447119,1.9994912,1.901403,1.6675003,1.2826926,0.73188925,0.0,0.21881226,0.2565385,0.14713238,0.10940613,0.55080324,0.573439,0.4074435,0.17354076,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.03772625,0.030181,0.033953626,0.0452715,0.071679875,0.056589376,0.033953626,0.018863125,0.030181,0.018863125,0.02263575,0.030181,0.030181,0.030181,0.018863125,0.033953626,0.10186087,0.19240387,0.23013012,0.23013012,0.14713238,0.10940613,0.17354076,0.32067314,0.271629,0.1961765,0.116951376,0.06413463,0.0754525,0.32067314,0.5998474,0.6187105,0.38480774,0.21503963,0.150905,0.27540162,0.3470815,0.29049212,0.1659955,0.15467763,0.20749438,0.24522063,0.20749438,0.060362,0.03772625,0.08677038,0.23013012,0.38480774,0.33576363,0.27540162,0.3055826,0.3734899,0.41498876,0.36594462,0.16976812,0.26031113,0.5093044,0.8601585,1.3128735,1.116697,0.91297525,0.754525,0.6752999,0.68661773,0.724344,0.7130261,0.694163,0.6526641,0.52062225,0.32444575,0.27540162,0.32444575,0.4376245,0.59607476,0.80356914,0.7922512,0.68661773,0.62248313,0.73188925,1.0601076,1.3996439,1.2185578,0.6149379,0.32067314,0.55080324,1.1506506,2.6446102,4.7648253,6.4247804,7.2057137,8.967529,9.748463,8.503497,5.111907,5.0138187,6.7756343,9.820143,11.393328,6.560595,3.92353,2.3767538,1.7014539,1.5316857,1.3732355,1.2751472,1.5354583,2.4220252,3.8820312,5.553304,6.2361493,7.3792543,8.616675,9.525878,9.612649,9.684328,8.926031,7.1302614,4.957229,3.904667,3.138824,2.2409391,1.599593,1.2826926,1.0374719,0.7432071,0.8262049,1.0299267,1.1921495,1.267602,0.76584285,0.422534,0.2565385,0.2678564,0.42630664,0.513077,0.5357128,0.55080324,0.573439,0.55080324,0.4376245,0.38480774,0.38480774,0.43007925,0.5017591,0.49044126,0.452715,0.392353,0.32444575,0.27540162,0.38480774,0.6413463,1.086516,1.6109109,1.9542197,2.0636258,1.9429018,2.0787163,2.5314314,2.9464202,2.957738,2.704972,2.4220252,2.2711203,2.3201644,2.0372176,1.8938577,1.7655885,1.6033657,1.4335974,1.3241913,1.3807807,1.6524098,2.0749438,2.4408884,2.8822856,3.519859,4.1800685,4.719554,5.036454,4.3875628,3.742444,3.138824,2.6898816,2.5804756,2.565385,2.4710693,2.323937,2.2296214,2.3654358,2.5729303,2.7615614,2.9766011,3.180323,3.2670932,3.3010468,3.0897799,2.867195,2.795515,2.9916916,3.5764484,4.1083884,4.6214657,5.20245,5.9984736,6.7039547,7.3377557,7.7187905,7.6886096,7.1264887,6.089017,6.4134626,6.7643166,6.4926877,5.6778007,6.175787,6.4134626,6.5341864,6.587003,6.5002327,7.145352,7.7037,6.9265394,4.9421387,3.218049,2.1956677,1.8448136,1.7014539,1.5241405,1.3430545,1.2449663,1.2487389,1.2864652,1.3204187,1.358145,1.297783,1.2713746,1.3204187,1.4411428,1.5882751,1.599593,1.4562333,1.3505998,1.3619176,1.4335974,1.5807298,1.6712729,1.720317,1.7467253,1.7693611,1.9051756,1.9730829,1.9881734,1.961765,1.9391292,1.9730829,2.1315331,2.5804756,3.078462,2.9464202,2.7238352,2.8822856,2.9351022,2.7238352,2.3805263,1.6486372,1.1431054,0.8224323,0.67152727,0.73188925,2.5993385,4.146115,4.7346444,4.738417,5.5683947,4.9459114,3.078462,2.022127,2.3013012,2.897376,3.5085413,3.2142766,2.8709676,2.897376,3.2670932,2.727608,2.3088465,2.0485353,1.7995421,1.2525115,0.94692886,0.79602385,0.7582976,0.7507524,0.6413463,0.6149379,1.1242423,1.8372684,2.444661,2.6408374,1.5769572,0.8262049,0.44139713,0.5017591,1.1129243,1.7127718,1.8448136,1.3656902,0.6149379,0.38103512,0.51684964,0.94315624,1.448688,1.8787673,2.1353056,2.161714,1.4901869,0.7884786,0.44516975,0.58098423,2.4823873,3.2821836,3.0860074,2.2899833,1.5580941,1.0072908,0.63002837,0.52062225,0.6790725,1.0223814,1.3996439,1.146878,1.026154,1.3091009,1.7844516,0.9922004,0.482896,0.1961765,0.071679875,0.060362,0.02263575,0.00754525,0.0,0.0,0.0,0.011317875,0.0150905,0.02263575,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.293756,3.5538127,4.3724723,4.9685473,5.560849,6.3908267,7.816879,9.529651,10.842525,11.68382,12.611885,13.249459,13.645585,13.834216,13.909668,14.034165,14.856597,16.278877,17.972786,19.836462,22.013268,21.45869,20.640032,19.97605,19.57615,19.28566,19.08571,18.980076,18.97253,19.029121,19.08571,19.413929,19.911915,20.48158,21.047476,21.590733,21.013521,20.383493,19.983595,20.089228,20.960705,21.537916,21.368149,20.375948,18.761265,16.999449,15.124454,13.600313,12.140307,10.748209,9.691874,8.318638,7.2887115,6.6134114,6.330465,6.515323,6.851087,7.2094865,7.598067,8.141325,9.0807085,10.125726,10.3634,10.38981,10.487898,10.646348,11.0613365,11.363147,11.61214,11.763044,11.676274,11.574413,11.476325,11.457462,11.608367,12.015811,12.181807,12.58925,13.245687,14.136025,15.203679,16.493916,18.406637,20.070366,20.8098,20.1345,18.5085,16.788181,15.0376835,13.241914,11.314102,9.646602,8.088508,6.651138,5.4250345,4.5799665,4.459243,4.214022,3.99521,3.9574835,4.2517486,3.8254418,3.4142256,2.8558772,2.2409391,1.9089483,1.81086,1.9202662,2.335255,2.9841464,3.6330378,4.2781568,4.708236,4.7421894,4.3196554,3.4745877,1.6750455,0.7167987,0.3772625,0.34330887,0.22258487,0.14335975,0.08677038,0.05281675,0.03772625,0.033953626,0.030181,0.0150905,0.003772625,0.003772625,0.0,0.0,0.011317875,0.02263575,0.041498873,0.06413463,0.0754525,0.07922512,0.094315626,0.124496624,0.16222288,0.19240387,0.2263575,0.25276586,0.25276586,0.2263575,0.21503963,0.29049212,0.35085413,0.331991,0.19240387,0.20749438,0.23390275,0.25276586,0.271629,0.31312788,0.32067314,0.32444575,0.5772116,0.9205205,0.7922512,0.31312788,0.38480774,0.46026024,0.31312788,0.03772625,0.08299775,0.23013012,0.41121614,0.5470306,0.5357128,0.35462674,0.19240387,0.24522063,0.452715,0.52062225,0.543258,0.5055317,0.38103512,0.19994913,0.03772625,0.06413463,0.026408374,0.0,0.0150905,0.071679875,0.17731337,0.25276586,0.38103512,0.5885295,0.86770374,1.4260522,2.3201644,2.6106565,2.2748928,2.2069857,2.7238352,2.3956168,1.7731338,1.1544232,0.55080324,0.15467763,0.05281675,0.06790725,0.13204187,0.2678564,0.24522063,0.12826926,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.018863125,0.0150905,0.00754525,0.00754525,0.02263575,0.02263575,0.018863125,0.0150905,0.018863125,0.026408374,0.030181,0.026408374,0.02263575,0.030181,0.026408374,0.03772625,0.056589376,0.071679875,0.071679875,0.07922512,0.06413463,0.06413463,0.10186087,0.19994913,0.150905,0.07922512,0.0452715,0.071679875,0.16222288,0.3169005,0.4074435,0.40367088,0.331991,0.2867195,0.3734899,0.36971724,0.2867195,0.1961765,0.241448,0.36594462,0.4376245,0.3470815,0.14713238,0.049044125,0.06413463,0.12826926,0.20749438,0.25276586,0.21503963,0.124496624,0.24899325,0.44894236,0.62248313,0.7205714,0.56212115,0.6187105,0.9205205,1.4222796,1.9730829,2.0673985,1.9957186,1.8372684,1.7052265,1.7354075,1.9579924,1.7240896,1.4222796,1.2411937,1.1657411,0.8941121,0.8601585,1.056335,1.448688,1.9881734,1.7240896,0.9808825,0.5394854,0.5998474,0.7696155,1.0789708,1.6260014,2.6634734,4.22534,6.119198,3.127506,1.5354583,1.0789708,1.388326,1.991946,2.7728794,3.874486,5.036454,6.590776,9.457971,11.59705,9.537196,6.820906,4.7836885,2.546522,2.191895,1.8561316,1.6524098,1.5882751,1.5580941,1.8184053,2.1202152,2.4484336,2.776652,3.0520537,3.4029078,4.1310244,5.1043615,6.1795597,7.220804,8.152642,7.250985,5.824933,4.6742826,4.0517993,3.85185,3.5990841,3.4142256,3.1161883,2.2447119,1.5920477,1.1808317,0.9922004,0.9507015,0.9242931,0.79602385,0.7130261,0.6149379,0.5017591,0.41498876,0.62625575,0.68661773,0.68661773,0.7432071,0.9997456,1.0676528,1.0714256,1.0110635,0.91297525,0.8224323,0.7394345,0.6828451,0.65643674,0.6488915,0.63002837,0.58098423,0.69793564,0.91297525,1.1619685,1.3656902,1.4675511,1.5279131,1.6675003,2.0070364,2.674791,3.1576872,3.4330888,3.3651814,2.9992368,2.5502944,1.9881734,1.8334957,1.9655377,2.3880715,3.1916409,2.535204,2.1013522,1.8448136,1.7542707,1.8561316,2.3163917,3.0407357,4.0895257,5.2665844,6.1078796,6.3116016,5.745708,4.957229,4.266839,3.7763977,3.6745367,3.4481792,3.180323,2.957738,2.867195,2.837014,2.867195,2.8709676,2.8256962,2.7653341,2.7238352,2.5729303,2.686109,3.1124156,3.6028569,3.6707642,3.9008942,4.3913355,5.2250857,6.4964604,7.7414265,8.688355,9.159933,9.329701,9.714509,9.631512,9.386291,9.831461,10.759526,10.887795,10.197406,10.11818,10.314357,10.529396,10.601076,9.461743,8.16396,6.3531003,4.3649273,3.218049,2.6936543,2.4823873,2.2899833,2.0372176,1.8938577,1.8636768,1.780679,1.7580433,1.8448136,2.0296721,2.0258996,2.11267,2.2748928,2.4786146,2.686109,2.425798,2.0447628,1.8070874,1.8259505,2.0447628,2.3277097,2.5125682,2.4333432,2.142851,1.8938577,2.123988,2.4107075,2.6446102,2.7540162,2.6710186,2.5012503,2.5238862,2.8558772,3.218049,2.957738,2.9728284,3.229367,3.0520537,2.4069347,1.9278114,1.6939086,2.4295704,3.3010468,3.8707132,4.0895257,5.1458607,5.624984,5.27413,4.266839,3.2029586,2.1692593,1.4449154,1.2525115,1.7127718,2.837014,3.8593953,3.6443558,3.3161373,3.380272,3.7160356,3.610402,2.9766011,2.1088974,1.2940104,0.8111144,0.663982,0.7507524,1.1053791,1.4373702,1.1431054,0.8941121,1.3807807,1.931584,2.1654868,1.9693103,1.0336993,0.49044126,0.33576363,0.5885295,1.297783,1.5543215,1.4071891,0.88279426,0.30935526,0.331991,0.4979865,0.66775465,0.8563859,1.056335,1.2336484,1.4034165,1.0902886,0.7997965,0.8299775,1.2751472,2.0258996,2.1202152,1.6448646,1.0110635,0.935611,1.4109617,2.1541688,2.2899833,1.871222,1.901403,2.2899833,2.0372176,1.6071383,1.3091009,1.297783,1.8787673,2.1013522,2.093807,1.9164935,1.5618668,0.90920264,0.32067314,0.026408374,0.011317875,0.011317875,0.0150905,0.0150905,0.0150905,0.018863125,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.0258996,2.8219235,3.7801702,4.5988297,5.1835866,5.6476197,6.809588,8.050782,8.952439,9.635284,10.767072,11.510279,12.113899,12.766563,13.358865,13.472044,13.849306,15.531898,17.286167,18.693357,20.157135,20.421219,20.798481,21.273832,21.553007,21.05502,20.549488,20.055275,19.70442,19.572378,19.696875,20.093,20.862616,21.639776,22.296213,22.963968,23.477045,23.171463,22.643295,22.307531,22.428255,23.443092,24.118391,23.967487,22.733839,20.37972,18.225552,16.863634,15.999702,15.335721,14.554788,13.068373,11.072655,9.26934,8.080963,7.6320205,8.013056,8.582722,9.235386,9.95973,10.838752,11.61214,11.846043,11.944131,12.113899,12.351574,12.668475,12.46098,12.264804,12.362892,12.777881,13.13628,13.472044,13.845533,14.351066,15.135772,16.180788,17.354074,18.391546,19.342249,20.57967,22.201899,24.167437,25.001186,24.125937,21.892544,20.541943,18.893307,17.105082,15.207452,13.068373,11.129244,9.261794,7.5565677,6.175787,5.3269467,4.9157305,4.6818275,4.640329,4.7120085,4.727099,3.8367596,3.199186,2.7615614,2.5427492,2.6483827,3.048281,3.5839937,4.327201,5.138315,5.715527,6.0776987,6.1041074,5.6061206,4.6026025,3.3161373,1.5845025,0.73188925,0.40367088,0.30935526,0.24899325,0.16976812,0.1056335,0.06790725,0.05281675,0.0754525,0.06790725,0.033953626,0.011317875,0.0150905,0.00754525,0.0150905,0.02263575,0.033953626,0.056589376,0.08677038,0.07922512,0.07922512,0.09808825,0.13958712,0.21503963,0.23013012,0.22258487,0.2263575,0.23767537,0.20749438,0.18863125,0.18485862,0.181086,0.17354076,0.1659955,0.21881226,0.26031113,0.29049212,0.3055826,0.31312788,0.28294688,0.29803738,0.6073926,1.0035182,0.8111144,0.31312788,0.34330887,0.38480774,0.23767537,0.02263575,0.041498873,0.10940613,0.211267,0.30935526,0.35839936,0.22258487,0.116951376,0.17354076,0.35085413,0.43007925,0.40367088,0.30935526,0.24899325,0.21503963,0.08677038,0.018863125,0.09808825,0.19240387,0.22258487,0.1659955,0.24522063,0.331991,0.47157812,0.6828451,0.95447415,1.5279131,2.4107075,2.625747,2.1881225,2.1202152,2.7540162,2.6898816,2.4559789,2.3314822,2.335255,1.5656394,0.98465514,0.4979865,0.15467763,0.14335975,0.07922512,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.003772625,0.0,0.0,0.00754525,0.02263575,0.0150905,0.003772625,0.0,0.0,0.018863125,0.02263575,0.0150905,0.0,0.00754525,0.0150905,0.0150905,0.011317875,0.00754525,0.0150905,0.018863125,0.02263575,0.02263575,0.026408374,0.030181,0.030181,0.0452715,0.060362,0.06790725,0.0754525,0.094315626,0.094315626,0.090543,0.090543,0.1056335,0.06413463,0.056589376,0.071679875,0.10940613,0.17354076,0.32444575,0.4074435,0.44894236,0.46026024,0.43385187,0.46026024,0.43007925,0.33953625,0.2565385,0.3055826,0.3772625,0.35462674,0.23767537,0.090543,0.026408374,0.06790725,0.150905,0.22258487,0.23390275,0.14713238,0.10186087,0.23013012,0.4979865,0.8224323,1.0638802,1.2638294,1.6260014,1.8561316,1.8674494,1.7882242,2.0183544,2.161714,2.1579416,2.033445,1.9164935,2.4182527,2.5276587,2.1013522,1.4449154,1.3166461,1.3166461,1.5882751,1.7316349,1.690136,1.7316349,1.6071383,1.7391801,2.04099,2.3390274,2.354118,2.9086938,3.0633714,2.886058,2.8445592,3.8065786,4.6026025,5.1269975,3.7198083,1.1657411,0.694163,0.9016574,1.3543724,2.2069857,3.6745367,6.047518,7.7150183,6.485142,4.5007415,2.8709676,1.6410918,1.4524606,1.3505998,1.2902378,1.2600567,1.2826926,1.6561824,2.3013012,2.686109,2.6898816,2.6106565,2.505023,2.776652,3.2670932,3.8556228,4.4705606,4.8063245,4.2592936,3.5160866,2.9652832,2.71629,2.7125173,2.6710186,2.6182017,2.4597516,1.9994912,1.5543215,1.2487389,1.0940613,1.0827434,1.1959221,1.0940613,0.94315624,0.79602385,0.69793564,0.7054809,0.875249,0.86770374,0.77338815,0.724344,0.8865669,1.0902886,1.237421,1.3015556,1.2864652,1.2110126,1.1129243,1.0676528,1.0940613,1.177059,1.2751472,1.3015556,1.3505998,1.4562333,1.5958204,1.7240896,1.8070874,1.7995421,1.8184053,1.9881734,2.4371157,3.078462,3.4330888,3.519859,3.3161373,2.7540162,2.2899833,2.0258996,2.04099,2.293756,2.595566,2.1768045,2.071171,2.0862615,2.1579416,2.3390274,2.5125682,2.757789,3.1765501,3.8178966,4.6931453,5.0213637,4.749735,4.3724723,4.168751,4.2102494,4.432834,4.2819295,4.063117,3.953711,3.9876647,4.187614,3.9197574,3.3010468,2.584248,2.1353056,2.0900342,2.0070364,2.1353056,2.5502944,3.1765501,3.3274553,3.380272,3.6934,4.429062,5.5495315,6.937857,8.367682,9.58624,10.653893,11.936585,12.7477,12.917468,12.838243,12.642066,12.208215,11.1631975,10.910432,11.068882,11.197151,10.79348,8.6732645,6.5756855,4.8930945,3.8065786,3.2746384,2.9728284,2.8521044,2.7728794,2.6974268,2.6785638,2.704972,2.7691069,2.8596497,2.9652832,3.0671442,3.0369632,3.0822346,3.1916409,3.3312278,3.4632697,3.3915899,3.108643,2.8407867,2.727608,2.837014,2.9803739,3.0218725,2.867195,2.5540671,2.252257,2.5238862,2.546522,2.4295704,2.252257,2.0749438,2.161714,2.1466236,2.1956677,2.3163917,2.384299,2.2899833,2.4408884,2.3956168,2.0258996,1.5430037,1.4977322,2.1881225,3.1199608,3.9122121,4.304565,4.4630156,4.134797,3.3953626,2.4333432,1.5467763,1.3053282,1.4373702,1.9202662,2.7691069,4.014073,4.8365054,4.7120085,4.164978,3.5500402,3.097325,2.9351022,2.335255,1.6524098,1.146878,0.97710985,1.0940613,1.5279131,1.8976303,1.9127209,1.3656902,1.1581959,1.4260522,1.7014539,1.6788181,1.2336484,0.6752999,0.39989826,0.43385187,0.8299775,1.6825907,1.5882751,1.0638802,0.5055317,0.19994913,0.29426476,0.38480774,0.41876137,0.482896,0.5885295,0.7054809,0.8111144,0.72811663,0.5772116,0.51684964,0.73566186,1.146878,1.2751472,1.1016065,0.80734175,0.7696155,1.4147344,2.1956677,2.3163917,1.8485862,1.7542707,2.1315331,2.5540671,2.969056,3.3576362,3.7273536,3.85185,3.3651814,2.6634734,2.1768045,2.3692086,1.5128226,0.62248313,0.13204187,0.060362,0.02263575,0.011317875,0.00754525,0.011317875,0.02263575,0.05281675,0.0452715,0.056589376,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.3088465,2.565385,3.1199608,3.6896272,4.142342,4.508287,5.458988,6.6247296,7.5829763,8.318638,9.224068,9.763554,10.4049,11.329193,12.464753,13.52486,13.660675,14.7321005,15.935568,16.920223,17.795471,18.632996,19.896824,21.247423,22.228306,22.269806,22.084948,21.41342,20.53817,19.666695,18.968758,19.247932,20.070366,20.915434,21.613369,22.330168,23.477045,23.69963,23.673222,23.69963,23.665676,24.639013,25.525581,25.834936,25.12191,22.97906,21.221016,20.213724,19.74592,19.455427,18.821627,17.320122,14.928277,12.521342,10.642575,9.49947,9.695646,10.329447,11.185833,12.140307,13.166461,13.547497,13.656902,13.70972,13.804035,13.924759,14.094527,13.920986,13.973803,14.449154,15.17727,15.871433,16.625957,17.47857,18.433046,19.421474,20.06282,21.07011,22.077402,23.073374,24.401339,25.808527,27.117628,27.268534,26.091475,24.314568,23.861853,23.00924,21.375692,18.851807,15.596032,13.008011,10.450171,8.080963,6.304056,5.80607,5.523123,5.383536,5.349582,5.304311,5.0553174,4.2328854,3.8103511,3.663219,3.7462165,4.112161,4.7233267,5.4174895,6.1908774,6.964266,7.6131573,7.4999785,6.828451,5.6061206,4.0480266,2.5729303,1.1996948,0.6375736,0.422534,0.31312788,0.271629,0.19994913,0.15467763,0.13204187,0.120724,0.120724,0.10186087,0.071679875,0.0452715,0.033953626,0.02263575,0.030181,0.0452715,0.06790725,0.090543,0.120724,0.07922512,0.0754525,0.090543,0.1358145,0.20749438,0.21503963,0.19994913,0.2263575,0.27917424,0.24522063,0.1961765,0.14713238,0.124496624,0.1358145,0.15845025,0.211267,0.2565385,0.28294688,0.2867195,0.241448,0.4640329,0.67152727,0.8941121,1.0148361,0.7809334,0.41876137,0.2867195,0.20372175,0.1056335,0.0452715,0.13958712,0.11317875,0.06413463,0.06413463,0.150905,0.12826926,0.10186087,0.10940613,0.15467763,0.23013012,0.21503963,0.11317875,0.124496624,0.21503963,0.1056335,0.02263575,0.22258487,0.43007925,0.47535074,0.29426476,0.43385187,0.58098423,0.7394345,0.90920264,1.0827434,1.5807298,2.3767538,2.5767028,2.142851,1.9202662,2.1013522,2.1202152,2.1956677,2.4408884,2.8596497,1.9693103,1.1959221,0.5394854,0.10186087,0.06413463,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.018863125,0.0150905,0.011317875,0.00754525,0.00754525,0.030181,0.02263575,0.00754525,0.0,0.0,0.0150905,0.02263575,0.018863125,0.00754525,0.02263575,0.02263575,0.0150905,0.003772625,0.0,0.00754525,0.0150905,0.018863125,0.030181,0.041498873,0.030181,0.030181,0.0452715,0.060362,0.0754525,0.10186087,0.124496624,0.13204187,0.13204187,0.116951376,0.090543,0.056589376,0.071679875,0.094315626,0.10186087,0.11317875,0.20749438,0.29049212,0.3734899,0.4376245,0.43385187,0.44516975,0.4640329,0.45648763,0.43007925,0.4376245,0.33576363,0.22258487,0.12826926,0.060362,0.02263575,0.0754525,0.14713238,0.18485862,0.16976812,0.09808825,0.124496624,0.271629,0.4979865,0.76207024,1.0223814,1.4600059,1.8599042,1.9542197,1.7655885,1.599593,1.9504471,2.282438,2.595566,2.806833,2.7879698,3.31991,3.772625,3.3463185,2.3314822,2.082489,2.6182017,3.240685,3.5877664,3.6141748,3.5651307,3.1425967,3.1652324,3.7990334,4.557331,4.3007927,4.5233774,4.3007927,3.3840446,2.2711203,2.2107582,3.9008942,4.9459114,3.772625,1.2336484,0.63002837,0.4979865,0.6149379,1.1016065,1.9730829,3.1312788,3.9989824,3.893349,3.5047686,3.0105548,2.0447628,1.2487389,1.0827434,1.1393328,1.2034674,1.2147852,1.3845534,1.9579924,2.3993895,2.6483827,3.1350515,2.8332415,2.6483827,2.6446102,2.8219235,3.108643,3.4745877,3.1916409,2.5729303,1.9278114,1.5882751,1.5128226,1.4675511,1.4373702,1.3996439,1.3355093,1.1544232,1.0110635,0.9318384,0.9393836,1.086516,1.0336993,0.9318384,0.84129536,0.8224323,0.935611,1.418507,1.4901869,1.2940104,1.0035182,0.8224323,0.95447415,1.1355602,1.2562841,1.3053282,1.3468271,1.388326,1.5618668,1.7919968,2.0372176,2.2447119,2.4371157,2.5012503,2.505023,2.5201135,2.6332922,2.6219745,2.5502944,2.5389767,2.637065,2.8181508,3.229367,3.451952,3.5877664,3.5990841,3.3236825,2.9011486,2.5276587,2.3465726,2.323937,2.2296214,2.2484846,2.637065,3.3161373,4.1083884,4.715781,4.90064,4.5761943,4.093298,3.7273536,3.6745367,3.561358,3.3274553,3.218049,3.3840446,3.874486,4.1762958,4.1612053,4.2328854,4.504514,4.817642,5.2779026,5.100589,4.236658,3.006782,2.11267,1.8448136,1.7467253,1.8485862,2.1805773,2.7502437,2.8785129,2.806833,2.9426475,3.4632697,4.293247,5.406172,6.7039547,8.073418,9.582467,11.45369,12.909923,13.264549,12.774108,11.864905,11.159425,10.378491,10.163452,10.299266,10.310584,9.457971,7.364164,5.406172,4.214022,3.8103511,3.6179473,3.3048196,3.127506,3.0860074,3.150142,3.270866,3.3463185,3.4972234,3.7235808,3.9612563,4.1272516,3.9084394,3.7613072,3.7537618,3.8593953,3.9461658,3.8669407,3.62172,3.4066803,3.3236825,3.380272,3.289729,3.2105038,3.0935526,2.927557,2.7540162,2.8219235,2.4974778,1.9994912,1.5543215,1.3656902,1.6410918,1.8259505,1.9655377,2.123988,2.3880715,1.9655377,1.7127718,1.5769572,1.4713237,1.267602,1.3920987,1.7354075,2.1994405,2.6219745,2.7992878,2.5427492,2.0296721,1.4600059,1.0035182,0.8224323,1.1732863,1.7089992,2.5125682,3.6179473,4.9949555,5.379763,4.961002,4.093298,3.187868,2.7200627,2.9539654,2.8256962,2.3578906,1.7391801,1.3241913,1.5354583,1.9051756,2.04099,1.7957695,1.2713746,1.3053282,1.6071383,1.9579924,1.991946,1.2336484,0.66020936,0.4678055,0.663982,1.20724,2.003264,1.4222796,0.7130261,0.24899325,0.14335975,0.2263575,0.40367088,0.41121614,0.35462674,0.3169005,0.362172,0.40367088,0.44894236,0.36971724,0.211267,0.17354076,0.41498876,0.6111652,0.7054809,0.7130261,0.7092535,1.1883769,1.6373192,1.7240896,1.4826416,1.327964,1.659955,2.1881225,2.8256962,3.5274043,4.285702,4.557331,4.0291634,3.150142,2.4107075,2.3201644,1.901403,1.3770081,0.9922004,0.7884786,0.60362,0.29803738,0.14335975,0.06413463,0.030181,0.0452715,0.0452715,0.0754525,0.06790725,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.5578396,2.7011995,2.7502437,2.7502437,2.8558772,3.3463185,4.1800685,5.66271,7.0510364,7.967784,8.401636,8.669493,9.163706,9.982366,11.317875,13.445636,13.766309,13.951167,14.4114275,15.282904,16.444872,17.467255,18.470772,19.60256,20.8513,22.03213,22.88097,22.737612,21.813318,20.387266,18.821627,18.863125,19.57615,20.462717,21.23988,21.83218,22.567842,23.145054,23.98635,25.057775,25.850027,26.453646,26.823364,26.834682,26.291424,24.940825,23.703403,23.205416,23.129965,23.073374,22.515026,20.964478,18.836716,16.4826,14.290704,12.657157,12.31762,12.736382,13.528633,14.520834,15.735619,16.090246,16.078928,15.988385,15.916705,15.799753,15.90916,16.343012,17.222033,18.30855,19.006485,19.84778,20.975796,22.03213,22.873425,23.563816,23.337458,23.405365,23.846762,24.710693,26.02734,27.113855,27.872154,28.204145,28.181509,28.057013,27.974014,27.574116,25.702894,22.054766,17.154125,13.483362,10.416218,7.7301087,5.881522,5.987156,6.1003346,6.1531515,6.115425,5.938112,5.5683947,5.1043615,5.0779533,5.2665844,5.553304,5.934339,6.3531003,6.94163,7.643338,8.492179,9.623966,9.114662,7.673519,5.515578,3.229367,1.8070874,0.80734175,0.52062225,0.44894236,0.362172,0.271629,0.211267,0.20749438,0.21503963,0.1961765,0.13958712,0.13204187,0.124496624,0.090543,0.041498873,0.041498873,0.0452715,0.07922512,0.1056335,0.116951376,0.120724,0.071679875,0.0754525,0.09808825,0.120724,0.14335975,0.15467763,0.16976812,0.23767537,0.3169005,0.26408374,0.18485862,0.12826926,0.120724,0.14713238,0.1659955,0.17731337,0.1961765,0.211267,0.19994913,0.120724,0.66020936,1.086516,1.1619685,0.94315624,0.77716076,0.55457586,0.23767537,0.041498873,0.0150905,0.071679875,0.23013012,0.1961765,0.11317875,0.06413463,0.09808825,0.14335975,0.14335975,0.09808825,0.03772625,0.03772625,0.026408374,0.011317875,0.08299775,0.181086,0.071679875,0.041498873,0.30935526,0.55457586,0.5998474,0.40367088,0.6752999,0.8903395,1.0412445,1.1393328,1.1959221,1.5580941,2.1994405,2.4031622,2.0598533,1.6675003,1.2261031,1.1016065,1.177059,1.388326,1.7316349,0.94315624,0.422534,0.124496624,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.02263575,0.02263575,0.02263575,0.02263575,0.018863125,0.011317875,0.0,0.011317875,0.0150905,0.00754525,0.0,0.003772625,0.003772625,0.00754525,0.0150905,0.02263575,0.03772625,0.030181,0.011317875,0.0,0.0,0.003772625,0.0150905,0.026408374,0.03772625,0.049044125,0.03772625,0.041498873,0.049044125,0.05281675,0.06413463,0.07922512,0.1056335,0.13204187,0.14335975,0.13958712,0.12826926,0.10186087,0.10186087,0.094315626,0.071679875,0.049044125,0.0452715,0.06790725,0.1358145,0.22258487,0.271629,0.34330887,0.41121614,0.47157812,0.513077,0.5055317,0.3169005,0.2263575,0.15845025,0.090543,0.0452715,0.07922512,0.10940613,0.09808825,0.060362,0.056589376,0.13204187,0.29803738,0.41876137,0.4979865,0.6752999,1.0827434,1.2223305,1.1959221,1.2223305,1.599593,2.0598533,2.372981,2.9200118,3.6443558,4.06689,4.617693,5.1760416,4.90064,3.9763467,3.6254926,4.195159,4.7421894,5.485397,6.270103,6.5568223,5.5382137,4.45547,5.0138187,6.696409,6.752999,5.7381625,5.05909,4.376245,3.783943,3.7952607,2.3503454,1.5430037,1.2638294,1.2449663,1.0940613,0.8526133,0.8299775,1.1619685,1.9579924,3.289729,4.006528,3.712263,3.361409,3.1124156,2.323937,1.3430545,1.1959221,1.3204187,1.4260522,1.4826416,1.4109617,1.5165952,1.8448136,2.505023,3.6707642,3.3010468,2.7313805,2.3767538,2.425798,2.848332,3.85185,3.7499893,3.2029586,2.5087957,1.599593,1.1506506,0.9507015,0.9016574,0.90920264,0.9016574,0.8563859,0.76207024,0.6752999,0.633801,0.663982,0.784706,0.9620194,1.1091517,1.2600567,1.5958204,2.4031622,2.4107075,1.9806281,1.3996439,0.9016574,0.8639311,0.9808825,1.0751982,1.116697,1.2298758,1.4750963,1.9579924,2.5238862,3.0256453,3.31991,3.5953116,3.651901,3.561358,3.4896781,3.6745367,3.6556737,3.5538127,3.5123138,3.5538127,3.5764484,3.6556737,3.7160356,3.8065786,3.9461658,4.1272516,3.572676,3.180323,2.9766011,2.9426475,3.0256453,3.2369123,4.014073,5.323174,6.8171334,7.84706,8.179051,7.6207023,6.7567716,5.772116,4.4403796,3.5651307,2.8785129,2.5880208,2.7351532,3.187868,3.229367,3.2746384,3.6330378,4.2706113,4.8402777,5.7419353,6.058836,5.2967653,3.783943,2.674791,2.1466236,1.9994912,2.11267,2.3880715,2.7238352,2.6408374,2.5012503,2.5389767,2.8634224,3.4783602,4.025391,4.610148,5.3910813,6.617184,8.643084,10.265312,10.435081,9.967276,9.378746,8.922258,8.409182,8.284684,8.409182,8.394091,7.598067,6.432326,5.2967653,4.5761943,4.29702,4.112161,3.712263,3.4066803,3.3048196,3.399135,3.5802212,3.6292653,3.6971724,3.9122121,4.255521,4.5535583,4.085753,3.731126,3.6254926,3.7160356,3.7650797,3.4783602,3.1954134,3.097325,3.187868,3.270866,3.0331905,2.9237845,2.8709676,2.8407867,2.8332415,2.6483827,2.2069857,1.6524098,1.1846043,1.0751982,1.2940104,1.7354075,2.2296214,2.6295197,2.8256962,2.1805773,1.5505489,1.2185578,1.2298758,1.3807807,1.4939595,1.5769572,1.5920477,1.5052774,1.3015556,1.1393328,0.88279426,0.6752999,0.6526641,0.935611,1.4750963,2.1277604,2.916239,3.893349,5.1760416,5.13077,4.304565,3.3274553,2.7653341,3.0935526,4.1083884,4.719554,4.221567,2.8181508,1.6109109,1.6260014,1.750498,1.7882242,1.6675003,1.448688,1.8485862,2.2409391,2.6219745,2.7011995,1.8749946,0.9997456,0.6488915,0.8639311,1.4411428,1.9391292,1.0676528,0.4678055,0.19240387,0.17731337,0.24522063,0.49421388,0.49421388,0.32444575,0.13958712,0.12826926,0.18863125,0.2867195,0.29426476,0.1961765,0.094315626,0.116951376,0.19240387,0.32067314,0.47912338,0.63002837,0.814887,0.935611,1.0186088,1.0299267,0.86770374,1.1393328,1.1959221,1.2562841,1.5241405,2.214531,3.338773,3.7084904,3.4670424,2.7615614,1.720317,1.9278114,2.2748928,2.4220252,2.214531,1.7052265,1.2185578,0.9620194,0.5885295,0.13204187,0.018863125,0.0150905,0.049044125,0.06413463,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.5314314,2.71629,2.7540162,2.746471,2.916239,3.6028569,4.2102494,4.949684,5.7419353,6.462507,6.911449,7.326438,7.8696957,9.084481,10.917976,12.725064,13.347548,13.743673,14.181297,14.713238,15.150862,15.82239,16.603323,17.40312,18.274595,19.410156,20.862616,22.239624,22.888515,22.703657,22.141537,21.617142,22.115128,23.111101,23.94485,23.835445,23.809036,24.005213,24.457928,25.144547,25.985842,26.755457,27.313805,27.502436,27.24967,26.566826,24.918188,25.016277,25.872662,26.642279,26.642279,25.32186,23.548725,21.38701,19.164934,17.455936,16.28265,15.946886,16.233604,16.94286,17.882242,18.968758,19.232841,19.15739,19.032892,18.934805,19.398838,20.402355,22.228306,24.193844,24.657877,25.061548,26.049976,26.404602,25.921707,25.419947,25.850027,25.687803,25.329405,25.174726,25.650078,27.125174,28.430502,29.20389,29.667923,30.607307,30.780848,29.724512,26.238607,20.719257,15.150862,10.525623,7.914967,6.6020937,6.255012,6.9265394,7.3415284,7.537705,7.488661,7.194396,6.6662283,6.436098,6.617184,6.8737226,7.0548086,7.201941,7.250985,7.960239,9.0957985,10.552032,12.359119,11.664956,9.684328,6.205968,2.5012503,1.3430545,0.8299775,0.63002837,0.482896,0.30935526,0.19994913,0.18485862,0.211267,0.21503963,0.18863125,0.150905,0.19994913,0.1961765,0.120724,0.041498873,0.0754525,0.10186087,0.124496624,0.120724,0.08677038,0.060362,0.060362,0.09808825,0.12826926,0.13204187,0.1056335,0.15467763,0.1961765,0.23013012,0.23767537,0.150905,0.1056335,0.10186087,0.124496624,0.150905,0.150905,0.116951376,0.116951376,0.120724,0.120724,0.120724,0.23013012,0.2867195,0.27540162,0.31312788,0.65643674,0.65643674,0.27917424,0.018863125,0.0,0.0,0.0,0.08299775,0.14335975,0.1358145,0.060362,0.08677038,0.08299775,0.0452715,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0452715,0.15467763,0.29426476,0.3961256,0.42630664,0.36594462,0.694163,0.8601585,0.91674787,0.9507015,1.0978339,1.3920987,1.8033148,1.8938577,1.6184561,1.3128735,0.95824677,0.8865669,0.875249,0.80356914,0.65643674,0.13204187,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.003772625,0.0150905,0.0150905,0.00754525,0.011317875,0.03772625,0.060362,0.02263575,0.0150905,0.00754525,0.003772625,0.0150905,0.026408374,0.030181,0.02263575,0.02263575,0.060362,0.08677038,0.08299775,0.06413463,0.041498873,0.030181,0.06790725,0.094315626,0.1056335,0.1056335,0.090543,0.1056335,0.1358145,0.14713238,0.1358145,0.120724,0.09808825,0.071679875,0.06790725,0.08677038,0.1358145,0.150905,0.14335975,0.13204187,0.12826926,0.150905,0.32444575,0.44894236,0.4074435,0.23013012,0.1056335,0.033953626,0.041498873,0.060362,0.056589376,0.0452715,0.071679875,0.13204187,0.22258487,0.35839936,0.56589377,0.79602385,0.9280658,0.8865669,0.86770374,1.3430545,1.7316349,1.5920477,1.8146327,2.6295197,3.6179473,4.9949555,5.5495315,5.6363015,5.481624,5.1873593,3.832987,3.1727777,3.9197574,5.2967653,5.0666356,4.52715,3.9084394,5.485397,8.903395,11.185833,8.20546,6.1795597,4.798779,4.13857,4.640329,3.663219,2.987919,3.0407357,3.3538637,2.546522,1.6222287,1.1431054,1.4222796,2.3616633,3.4481792,4.2064767,3.5538127,2.4823873,1.6675003,1.4335974,1.690136,1.7731338,1.5543215,1.3015556,1.6788181,1.9466745,1.9504471,2.2748928,2.938875,3.4029078,2.4371157,1.6750455,1.2110126,1.1016065,1.358145,1.5052774,2.1088974,3.451952,4.504514,2.9313297,1.659955,1.0601076,0.8563859,0.86770374,0.97710985,1.086516,1.1053791,1.086516,1.0638802,1.0525624,1.3204187,1.7995421,2.2598023,2.8294687,4.014073,3.9386206,2.9237845,1.81086,1.0487897,0.67152727,0.7696155,0.9507015,1.1506506,1.2789198,1.20724,1.3996439,1.9089483,2.7426984,3.6368105,4.0291634,4.0782075,3.92353,3.85185,4.002755,4.395108,4.847823,4.5761943,4.123479,3.783943,3.6028569,3.942393,3.9386206,3.9499383,4.1498876,4.515832,3.8443048,3.6141748,3.7650797,4.0970707,4.255521,4.0970707,5.292993,6.760544,7.907422,8.650629,8.322411,8.2507305,8.345046,8.16396,6.881268,5.243949,3.6179473,2.8332415,2.8936033,2.9916916,2.9049213,2.8181508,2.916239,3.289729,3.9386206,6.205968,6.8925858,5.764571,3.772625,3.0520537,2.8558772,2.8332415,2.8521044,2.8558772,2.867195,2.9426475,2.8521044,2.8634224,3.0897799,3.4783602,3.429316,3.610402,4.0178456,4.870459,6.590776,7.61693,8.213005,8.107371,7.356619,6.3342376,5.089271,4.6931453,4.6818275,4.768598,4.851596,5.070408,5.0439997,4.8440504,4.5535583,4.2706113,3.9688015,3.7160356,3.6669915,3.7877154,3.8593953,3.6783094,3.5387223,3.440634,3.380272,3.3576362,2.8822856,2.595566,2.4522061,2.3503454,2.1654868,2.093807,2.0862615,2.1390784,2.1956677,2.1353056,2.0145817,1.8448136,1.6561824,1.5015048,1.4637785,1.5128226,1.4713237,1.3053282,1.0978339,1.0374719,1.1581959,1.4109617,1.750498,2.082489,2.2296214,1.9730829,1.7693611,1.9466745,2.3578906,2.3956168,1.6863633,1.418507,1.4864142,1.7165444,1.8749946,1.7919968,1.4939595,1.1242423,0.97333723,1.50905,2.7804246,3.7575345,4.4139714,4.749735,4.7610526,4.432834,4.0480266,3.6443558,3.4594972,3.9348478,5.05909,6.138061,5.5759397,3.5047686,1.7693611,1.3543724,2.0485353,2.7691069,3.0746894,3.1576872,3.9386206,3.6028569,2.7389257,2.0108092,2.1805773,1.5580941,0.95447415,0.784706,0.9997456,1.0827434,0.935611,0.633801,0.47535074,0.52439487,0.6111652,0.3055826,0.15467763,0.0754525,0.030181,0.030181,0.12826926,0.24522063,0.33576363,0.362172,0.29049212,0.25276586,0.30935526,0.4376245,0.58475685,0.65643674,0.30181,0.150905,0.1056335,0.10940613,0.120724,0.36594462,0.59230214,0.6828451,0.69039035,0.8224323,1.2147852,1.8636768,2.1805773,1.9542197,1.3430545,1.1959221,2.2409391,3.3878171,3.7575345,2.6710186,3.169005,3.3878171,2.3126192,0.5055317,0.090543,0.06790725,0.060362,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6524098,1.8184053,1.871222,2.0787163,2.5767028,3.3689542,4.478106,5.8098426,7.0812173,8.024373,8.390318,7.956466,8.080963,9.510788,11.502733,11.834724,11.830952,12.487389,13.864397,15.596032,16.886269,16.365646,16.731592,17.4333,18.063328,18.346275,19.440336,20.602304,21.541689,22.107582,22.299986,22.60557,23.552498,24.586197,25.385994,25.872662,26.189562,27.196854,28.22678,28.562544,27.415667,27.811792,28.539907,29.354795,29.95087,29.958416,29.10203,27.626932,26.993132,27.476028,28.181509,28.158873,27.849518,27.359077,26.823364,26.404602,25.808527,25.416174,25.412401,25.706667,25.914162,26.140518,26.24238,25.959433,25.370903,24.891779,25.816072,26.40083,26.97804,27.740112,28.720995,28.1966,27.63825,27.62316,28.057013,28.132465,28.215462,28.317324,27.974014,27.17799,26.34424,26.310287,26.766775,27.5213,28.596497,30.230043,28.683268,25.646305,21.013521,15.697892,11.623458,8.91094,7.9715567,7.6131573,7.3453007,7.3905725,8.684583,8.959985,8.601585,8.058327,7.877241,7.877241,8.0206,8.201687,8.465771,9.031664,9.812597,10.86516,12.298758,14.015302,15.716756,14.592513,11.065109,6.085244,1.6750455,0.91674787,0.5998474,0.47535074,0.35462674,0.19240387,0.11317875,0.10940613,0.14335975,0.1659955,0.15845025,0.13958712,0.20749438,0.19994913,0.14335975,0.09808825,0.17354076,0.19994913,0.21503963,0.20372175,0.16976812,0.1358145,0.11317875,0.13204187,0.14713238,0.13958712,0.1056335,0.15467763,0.181086,0.18863125,0.17354076,0.116951376,0.09808825,0.12826926,0.30935526,0.52439487,0.44516975,0.14713238,0.2263575,0.35462674,0.3772625,0.3169005,0.33953625,0.28294688,0.16976812,0.07922512,0.15467763,0.14713238,0.060362,0.003772625,0.0,0.0,0.0,0.0150905,0.030181,0.026408374,0.011317875,0.08677038,0.10186087,0.060362,0.0,0.0,0.0,0.0,0.0,0.07922512,0.39989826,0.995973,0.8978847,0.67152727,0.59230214,0.66020936,1.1544232,1.3015556,1.1280149,0.86770374,0.965792,0.9242931,0.91674787,0.88279426,0.814887,0.76207024,0.7130261,0.754525,0.73188925,0.5696664,0.26408374,0.05281675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.003772625,0.0150905,0.033953626,0.03772625,0.03772625,0.03772625,0.02263575,0.018863125,0.0150905,0.0150905,0.0150905,0.026408374,0.041498873,0.033953626,0.030181,0.033953626,0.060362,0.08677038,0.0754525,0.056589376,0.06413463,0.12826926,0.14713238,0.15467763,0.120724,0.06790725,0.056589376,0.0754525,0.094315626,0.116951376,0.14335975,0.16976812,0.1358145,0.10186087,0.071679875,0.060362,0.08677038,0.12826926,0.15467763,0.124496624,0.07922512,0.1056335,0.18863125,0.3055826,0.3169005,0.1961765,0.0452715,0.02263575,0.026408374,0.03772625,0.03772625,0.0452715,0.049044125,0.071679875,0.1358145,0.29049212,0.5772116,0.90543,0.98842776,1.0336993,1.1808317,1.4901869,1.9089483,1.8938577,1.7693611,1.7769064,2.04099,3.832987,5.5382137,5.8400235,4.7421894,3.5538127,2.3918443,2.3465726,3.451952,5.270357,6.8850408,6.319147,5.062863,4.014073,3.9499383,5.5193505,5.617439,5.715527,5.775889,5.753253,5.59103,5.032682,5.4250345,5.926794,6.047518,5.613666,4.779916,4.466788,4.6742826,5.4401255,6.828451,6.4247804,5.0138187,3.6934,3.0445085,3.1048703,3.6254926,3.4029078,2.8747404,2.3465726,1.9730829,2.1051247,2.203213,2.3956168,2.6785638,2.938875,2.6106565,2.173032,1.7354075,1.4071891,1.3204187,1.3505998,1.3996439,1.5580941,1.6561824,1.2336484,1.1355602,0.98842776,0.7884786,0.6187105,0.66020936,0.80734175,0.995973,1.146878,1.2034674,1.1506506,1.0487897,1.0751982,1.1317875,1.2223305,1.448688,1.5505489,1.50905,1.4675511,1.3920987,1.0601076,1.1581959,1.4939595,1.9240388,2.1994405,1.9504471,1.267602,1.2298758,1.5316857,1.9429018,2.3314822,2.6332922,2.9916916,3.4557245,4.093298,4.979865,4.9044123,4.032936,3.2482302,2.8634224,2.6106565,2.5729303,2.282438,2.0145817,1.901403,1.9051756,2.1503963,2.6182017,3.2784111,4.0404816,4.745962,4.957229,5.1345425,5.621211,6.25124,6.3342376,5.534441,5.723072,5.8513412,5.2967653,3.8782585,3.1425967,2.6785638,2.6597006,3.2670932,4.6629643,4.5988297,3.3236825,2.4182527,2.4220252,2.8256962,4.0216184,3.99521,3.500996,3.1727777,3.5274043,3.9386206,4.244203,4.4101987,4.4931965,4.6629643,5.372218,6.477597,6.25124,4.6856003,3.5160866,3.0746894,3.1425967,3.5462675,4.2517486,5.3571277,5.1345425,4.8100967,4.3800178,3.9197574,3.5990841,3.2331395,3.0445085,3.2784111,3.772625,3.9386206,3.4255435,3.6896272,4.2781568,4.9534564,5.6891184,4.6214657,3.783943,3.429316,3.470815,3.5047686,3.380272,3.150142,2.897376,2.6634734,2.4522061,2.1843498,2.1277604,2.1202152,2.0598533,1.8863125,1.9504471,2.0900342,2.3126192,2.4484336,2.173032,1.8561316,1.5656394,1.5845025,1.8636768,2.003264,1.7278622,1.6637276,1.6109109,1.4637785,1.20724,1.4977322,1.7731338,1.9353566,1.9957186,2.093807,1.991946,1.720317,2.022127,2.7728794,3.006782,1.5958204,1.1204696,1.1393328,1.358145,1.6335466,1.5656394,1.478869,1.4713237,1.7240896,2.535204,3.7160356,4.98741,5.613666,5.492942,5.1647234,4.949684,4.5460134,3.9650288,3.240685,2.3993895,2.867195,3.4896781,3.7613072,3.429316,2.4672968,2.003264,2.5201135,3.0671442,3.2255943,3.1463692,2.9124665,2.2560298,1.6373192,1.5731846,2.6332922,1.961765,1.2298758,0.9507015,1.2638294,1.9240388,2.1202152,1.1883769,0.3961256,0.211267,0.2678564,0.3055826,0.241448,0.1358145,0.06413463,0.090543,0.24899325,0.38480774,0.41876137,0.35085413,0.27917424,0.241448,0.25276586,0.271629,0.2867195,0.29049212,0.23013012,0.23013012,0.2565385,0.2565385,0.16976812,0.27917424,0.3734899,0.35085413,0.24899325,0.27540162,0.47157812,0.84129536,1.3732355,1.9278114,2.233394,1.3355093,2.0975795,3.3312278,3.6783094,1.5958204,1.4034165,1.5203679,1.1129243,0.27917424,0.030181,0.056589376,0.06790725,0.06413463,0.03772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.599593,1.5241405,1.5128226,1.7052265,2.1051247,2.5880208,3.3727267,4.395108,5.6287565,6.820906,7.4773426,7.2170315,7.5905213,8.737399,10.178542,10.77839,11.46878,12.325166,13.43809,14.769827,16.146835,16.493916,17.282394,17.991648,18.368912,18.448135,19.089483,19.753464,20.432537,21.19838,22.183035,23.126192,24.239115,25.33695,26.261242,26.857317,27.260988,27.88347,28.32487,28.29846,27.634478,28.438047,29.415157,30.305496,30.860073,30.844982,30.154593,28.905853,28.230553,28.32487,28.472,28.472,28.434275,28.777584,29.566063,30.516764,30.562035,30.73935,31.067568,31.297697,30.890253,30.192318,29.434021,28.464457,27.53639,27.298714,28.049467,28.445593,28.524818,28.430502,28.411638,28.5135,28.358822,28.464457,28.834173,28.981306,28.358822,27.626932,27.540163,27.902334,27.555252,27.008223,27.487347,27.864609,27.619389,26.842226,23.265778,19.534653,15.663939,12.181807,10.148361,8.944894,8.643084,8.816625,9.031664,8.835487,8.801534,8.98262,9.039209,8.952439,8.993938,8.892077,8.956212,9.167479,9.578695,10.27663,11.344283,12.706201,14.369928,15.973294,16.803272,15.041456,10.582213,5.492942,1.6486372,0.72811663,0.4640329,0.331991,0.23767537,0.15845025,0.1358145,0.12826926,0.116951376,0.15467763,0.23390275,0.27540162,0.23013012,0.1961765,0.181086,0.20372175,0.32821837,0.32821837,0.30181,0.2565385,0.20749438,0.181086,0.15467763,0.13958712,0.13204187,0.124496624,0.124496624,0.17354076,0.17731337,0.16222288,0.12826926,0.07922512,0.08299775,0.12826926,0.2678564,0.42630664,0.41876137,0.32444575,0.52439487,0.73188925,0.7997965,0.7432071,0.513077,0.41876137,0.362172,0.271629,0.08677038,0.08677038,0.13958712,0.16976812,0.15467763,0.10940613,0.06413463,0.09808825,0.27917424,0.60362,1.0072908,1.297783,1.2110126,0.87147635,0.44516975,0.14713238,0.62248313,1.3694628,1.7467253,1.6788181,1.6222287,1.6109109,1.2713746,0.9318384,0.7696155,0.77716076,1.2411937,1.3241913,1.0638802,0.7167987,0.7205714,0.65643674,0.60362,0.55457586,0.52439487,0.543258,0.60362,0.5885295,0.5017591,0.32821837,0.06790725,0.07922512,0.08299775,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.011317875,0.0150905,0.00754525,0.00754525,0.003772625,0.0,0.0,0.00754525,0.02263575,0.033953626,0.0452715,0.049044125,0.02263575,0.018863125,0.0150905,0.0150905,0.0150905,0.02263575,0.033953626,0.049044125,0.056589376,0.056589376,0.05281675,0.05281675,0.05281675,0.05281675,0.06790725,0.124496624,0.150905,0.14713238,0.1358145,0.13204187,0.1659955,0.20372175,0.17354076,0.116951376,0.07922512,0.10940613,0.13204187,0.14713238,0.14713238,0.1358145,0.13204187,0.120724,0.09808825,0.071679875,0.056589376,0.071679875,0.09808825,0.14335975,0.15845025,0.116951376,0.041498873,0.018863125,0.018863125,0.030181,0.041498873,0.0452715,0.0452715,0.056589376,0.13204187,0.30181,0.56212115,0.8639311,1.2110126,1.6335466,2.0070364,2.0485353,2.1881225,2.2484846,1.9881734,1.6486372,1.931584,3.4444065,5.0553174,5.50426,4.5535583,2.9954643,1.9240388,1.8259505,2.5729303,4.055572,6.156924,6.5228686,5.945657,4.825187,3.874486,4.123479,4.6516466,5.6589375,6.56814,7.043491,6.990674,5.564622,5.243949,5.824933,6.5756855,6.2135134,5.5193505,5.281675,5.881522,7.0170827,7.7225633,6.168242,5.1081343,4.5497856,4.395108,4.4403796,5.1571784,5.2854476,4.7950063,4.0291634,3.712263,3.5651307,3.1048703,3.0860074,3.7084904,4.5988297,5.5570765,5.8513412,5.541986,4.689373,3.3538637,2.637065,2.1390784,1.780679,1.5618668,1.569412,1.6675003,1.418507,1.0978339,0.875249,0.8186596,0.8903395,1.116697,1.3845534,1.5958204,1.659955,1.50905,1.3958713,1.3732355,1.3996439,1.3656902,1.3656902,1.448688,1.5165952,1.4901869,1.297783,1.3053282,1.4750963,1.7618159,2.0636258,2.2183034,1.6222287,1.4411428,1.3958713,1.4071891,1.5882751,1.8636768,2.2899833,2.9841464,3.9310753,4.979865,5.1458607,4.881777,4.6214657,4.45547,4.1498876,3.7084904,3.0143273,2.425798,2.1654868,2.3126192,3.0520537,3.2444575,3.2972744,3.4179983,3.5839937,3.99521,3.92353,3.863168,4.002755,4.2328854,4.044254,4.5120597,4.727099,4.244203,3.0897799,2.263575,1.9881734,2.2183034,2.8936033,3.953711,3.85185,3.1954134,2.7615614,2.8558772,3.3350005,3.7877154,3.5274043,3.2821836,3.3840446,3.7575345,4.085753,4.4403796,4.715781,4.9232755,5.20245,6.530414,7.635793,7.4207535,5.9230213,4.304565,3.399135,3.1237335,3.180323,3.3878171,3.6481283,3.150142,2.686109,2.3390274,2.161714,2.191895,2.052308,1.9768555,2.2447119,2.6936543,2.746471,2.3956168,2.8030603,3.5953116,4.496969,5.3458095,4.3686996,3.4481792,2.8747404,2.6936543,2.6936543,3.0746894,3.3425457,3.2255943,2.7691069,2.3277097,1.8900851,1.7919968,1.8448136,1.9202662,1.9164935,1.961765,1.8976303,1.8976303,2.003264,2.1277604,1.8787673,1.6524098,1.6184561,1.7618159,1.8787673,1.780679,1.8787673,1.9730829,1.931584,1.7014539,1.6637276,1.7618159,1.9806281,2.305074,2.7200627,2.6521554,2.4861598,2.3616633,2.3013012,2.2258487,1.5769572,1.3166461,1.4524606,1.9089483,2.5427492,2.5767028,2.969056,3.832987,4.983638,5.915476,6.5756855,6.6586833,6.175787,5.455216,5.1269975,5.7872066,5.987156,5.7419353,4.98741,3.5877664,2.9351022,3.4142256,4.7874613,5.8664317,4.534695,2.9954643,2.214531,2.2748928,2.9086938,3.482133,3.380272,3.2482302,3.3123648,3.6858547,4.376245,3.31991,2.0485353,1.237421,1.1996948,1.8900851,2.1768045,1.5769572,0.8941121,0.48666862,0.2565385,0.23013012,0.29049212,0.331991,0.31312788,0.25276586,0.5281675,0.8601585,1.1280149,1.1393328,0.6488915,0.2263575,0.124496624,0.14335975,0.17731337,0.21503963,0.21503963,0.23013012,0.24522063,0.23767537,0.15467763,0.17731337,0.23390275,0.31312788,0.38480774,0.38480774,0.38480774,0.5998474,1.1091517,1.7618159,2.173032,1.8863125,2.4786146,3.3350005,3.7575345,2.957738,2.757789,2.535204,1.8070874,0.7507524,0.20749438,0.060362,0.026408374,0.041498873,0.056589376,0.0452715,0.03772625,0.018863125,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4298248,1.3619176,1.3996439,1.5958204,1.9089483,2.2107582,2.71629,3.4255435,4.4101987,5.5457587,6.5002327,6.760544,7.3415284,8.171506,9.175024,10.246449,11.608367,12.419481,13.000465,13.611631,14.456699,15.437581,16.520325,17.467255,18.1086,18.368912,18.829172,19.251705,19.719511,20.417446,21.62846,22.862108,24.250433,25.529354,26.359331,26.34424,27.2044,27.872154,27.747658,27.083675,26.966724,27.811792,28.532362,29.154846,29.656605,29.977278,30.03764,29.796192,29.69056,29.758467,29.667923,29.80751,29.913143,30.07914,30.52431,31.599506,32.199356,32.731293,33.346233,33.90458,33.97249,33.372643,32.701115,31.931498,31.165655,30.637487,30.573353,30.309269,29.818829,29.215208,28.75872,29.554745,29.758467,29.90937,30.282862,30.863846,29.932007,28.74363,28.290915,28.404093,27.78161,26.819592,26.815819,26.381968,24.872917,22.367893,18.059555,14.875461,12.449662,10.699164,9.8239155,9.35611,9.208978,9.510788,10.005001,10.054046,9.529651,9.635284,9.774872,9.718282,9.578695,9.386291,9.242931,9.171251,9.190115,9.314611,10.665211,12.427027,14.358611,15.769572,15.516807,13.189097,8.820397,4.606375,1.7919968,0.663982,0.3734899,0.20749438,0.12826926,0.116951376,0.14335975,0.16976812,0.16976812,0.19240387,0.241448,0.27917424,0.23013012,0.24899325,0.29049212,0.34330887,0.43007925,0.40367088,0.3470815,0.27917424,0.2263575,0.211267,0.18485862,0.13958712,0.10940613,0.120724,0.14335975,0.17731337,0.17354076,0.150905,0.10940613,0.056589376,0.10186087,0.1659955,0.24522063,0.30935526,0.30935526,0.35085413,0.5055317,0.724344,0.9280658,0.9922004,0.6828451,0.5017591,0.38858038,0.27917424,0.1056335,0.14713238,0.22258487,0.25276586,0.22258487,0.1659955,0.15845025,0.33576363,0.7696155,1.4411428,2.2220762,2.7653341,2.7426984,2.4484336,2.082489,1.7391801,2.5087957,3.561358,4.0480266,3.712263,2.8822856,1.8938577,1.2902378,0.965792,0.83752275,0.8865669,1.20724,1.1808317,0.8865669,0.5357128,0.48666862,0.4640329,0.46026024,0.452715,0.452715,0.5017591,0.5998474,0.49044126,0.32067314,0.16222288,0.0,0.06413463,0.08299775,0.049044125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.041498873,0.041498873,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.011317875,0.0150905,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.00754525,0.0150905,0.026408374,0.033953626,0.018863125,0.011317875,0.00754525,0.011317875,0.0150905,0.00754525,0.026408374,0.056589376,0.090543,0.1056335,0.08299775,0.071679875,0.071679875,0.071679875,0.06790725,0.0754525,0.094315626,0.09808825,0.124496624,0.18863125,0.2867195,0.2867195,0.22258487,0.14713238,0.09808825,0.1056335,0.124496624,0.16222288,0.181086,0.17354076,0.14335975,0.094315626,0.05281675,0.033953626,0.041498873,0.049044125,0.0452715,0.03772625,0.041498873,0.041498873,0.026408374,0.018863125,0.026408374,0.041498873,0.05281675,0.041498873,0.033953626,0.03772625,0.094315626,0.23013012,0.45648763,0.72811663,1.2034674,1.7127718,2.071171,2.0787163,2.1994405,2.2711203,2.0296721,1.6712729,1.8334957,2.848332,3.9989824,4.6327834,4.4177437,3.3576362,2.5767028,2.1579416,2.3578906,3.2142766,4.5724216,5.413717,5.9796104,5.9305663,5.43258,5.160951,5.7079816,6.5945487,7.383027,7.6395655,6.9491754,5.3759904,5.1571784,5.8437963,6.5455046,5.9003854,5.2892203,5.0477724,5.5495315,6.5530496,7.232122,5.987156,5.7117543,6.0022464,6.3342376,6.0814714,6.1305156,6.0550632,5.621211,5.1043615,5.2779026,5.1534057,4.504514,4.3800178,5.3759904,7.624475,9.129752,9.333474,8.43559,6.7454534,4.67051,3.4179983,2.9011486,2.6408374,2.4295704,2.3314822,2.305074,1.9655377,1.5656394,1.2789198,1.1846043,1.2147852,1.3807807,1.6788181,2.0636258,2.4672968,2.7200627,2.6597006,2.5880208,2.5880208,2.546522,2.41448,2.3692086,2.2975287,2.161714,1.9730829,1.8221779,1.7165444,1.7278622,1.8938577,2.2107582,2.1088974,1.9693103,1.7354075,1.4713237,1.3619176,1.4637785,1.7240896,2.305074,3.1539145,3.9914372,4.564876,5.1760416,5.855114,6.5756855,7.250985,7.4471617,6.730363,5.6778007,4.7572803,4.346064,4.5497856,4.2328854,3.62172,2.957738,2.5238862,2.7200627,2.7238352,2.6785638,2.757789,3.1539145,3.229367,3.591539,3.7914882,3.591539,2.9803739,2.1088974,1.6561824,1.7089992,2.1843498,2.8181508,2.9992368,3.1124156,3.270866,3.5953116,4.2404304,4.7233267,4.557331,4.2894745,4.191386,4.2404304,4.376245,4.644101,4.927048,5.149633,5.2628117,6.0362,6.507778,6.379509,5.624984,4.496969,3.7273536,3.4066803,3.308592,3.2482302,3.059599,2.6597006,2.1994405,1.9391292,1.9278114,1.9881734,1.7127718,1.6637276,1.8221779,2.0070364,1.8599042,1.6825907,2.04099,2.6974268,3.3538637,3.651901,3.0520537,2.4786146,2.093807,1.9730829,2.0787163,2.6332922,3.1312788,3.2142766,2.8747404,2.4522061,2.0145817,1.8636768,1.8825399,1.991946,2.1353056,2.2371666,2.2371666,2.1541688,2.0862615,2.1994405,2.0447628,2.003264,2.0636258,2.1843498,2.3088465,2.3993895,2.6182017,2.727608,2.5993385,2.1994405,1.9693103,1.8976303,1.9806281,2.2258487,2.6521554,2.8558772,2.9615107,2.8106055,2.4597516,2.1805773,2.093807,2.0862615,2.444661,3.218049,4.214022,4.647874,5.2590394,6.398372,7.854605,8.812852,8.409182,7.2698483,5.802297,4.568649,4.266839,5.541986,6.7341356,7.062354,6.2097406,4.3196554,3.2369123,3.6745367,5.2062225,6.462507,5.1081343,3.0822346,1.7693611,1.7278622,2.795515,4.093298,4.817642,5.1081343,4.82896,4.236658,3.9688015,3.2029586,2.233394,1.4901869,1.237421,1.5656394,1.7844516,1.5580941,1.1355602,0.69039035,0.29803738,0.15845025,0.26031113,0.4074435,0.47912338,0.43007925,0.6149379,0.91674787,1.20724,1.2638294,0.7469798,0.21503963,0.06413463,0.08677038,0.1659955,0.25276586,0.2867195,0.26031113,0.19994913,0.1358145,0.08677038,0.08677038,0.1358145,0.26408374,0.41121614,0.4376245,0.4640329,0.84884065,1.3204187,1.6637276,1.6863633,1.8636768,2.4823873,3.2520027,3.9197574,4.2630663,4.1498876,3.3312278,2.11267,0.9242931,0.33576363,0.21503963,0.10940613,0.05281675,0.041498873,0.056589376,0.06413463,0.0452715,0.026408374,0.0150905,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9997456,1.1619685,1.3317367,1.5958204,1.9466745,2.293756,2.7804246,3.4217708,4.1197066,4.889322,5.847569,6.571913,7.213259,7.9715567,8.922258,10.005001,11.314102,11.932813,12.427027,12.955194,13.29473,13.747445,14.543469,15.682802,16.886269,17.591751,18.312323,19.025349,19.711966,20.43631,21.34174,22.481071,23.92976,25.204908,25.823618,25.291677,26.536644,27.528845,27.23458,26.02734,25.691576,25.872662,25.880207,26.178246,26.951633,28.102283,29.524563,30.437538,30.980797,31.286379,31.456148,32.195583,32.618114,32.154083,31.22979,31.248653,31.912636,32.26349,32.98029,34.251663,35.764484,36.60201,37.145267,37.375397,37.073586,35.82485,34.655334,33.440548,32.414394,31.742867,31.508965,32.131447,32.116356,32.10881,32.489845,33.35755,32.489845,31.429739,30.131956,28.64177,27.064812,25.518036,24.30325,22.718748,20.564579,18.153872,14.901869,13.12119,12.095036,11.3669195,10.733118,10.061591,9.763554,9.842778,10.220041,10.736891,10.93684,10.933067,10.63503,10.106862,9.57115,9.352338,8.812852,8.088508,7.281166,6.436098,8.213005,10.359629,12.510024,13.717264,12.449662,9.891823,6.5530496,3.7273536,1.9051756,0.7809334,0.35839936,0.15467763,0.08677038,0.08677038,0.13204187,0.2263575,0.3055826,0.27917424,0.19994913,0.24899325,0.3470815,0.4074435,0.4376245,0.44516975,0.43385187,0.392353,0.33576363,0.2678564,0.20749438,0.19994913,0.17731337,0.120724,0.10186087,0.12826926,0.14713238,0.15845025,0.1659955,0.15467763,0.11317875,0.060362,0.1358145,0.2263575,0.31312788,0.36594462,0.32067314,0.30935526,0.3055826,0.47912338,0.7922512,1.0299267,0.9507015,0.6752999,0.3734899,0.16222288,0.120724,0.17354076,0.19994913,0.18485862,0.14713238,0.13204187,0.24522063,0.5885295,1.177059,1.9542197,2.8181508,3.5651307,3.942393,4.217795,4.4177437,4.3083377,4.719554,5.149633,5.221313,4.6554193,3.270866,1.7542707,1.0412445,0.80734175,0.84129536,1.0487897,1.1204696,0.98465514,0.7092535,0.43385187,0.38480774,0.35462674,0.35462674,0.3772625,0.42630664,0.48666862,0.5772116,0.41876137,0.2263575,0.090543,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.03772625,0.08677038,0.08677038,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.00754525,0.011317875,0.003772625,0.02263575,0.05281675,0.10940613,0.16222288,0.150905,0.14713238,0.13204187,0.10186087,0.06413463,0.033953626,0.02263575,0.049044125,0.10186087,0.18485862,0.31312788,0.2565385,0.211267,0.1961765,0.19240387,0.15845025,0.11317875,0.116951376,0.12826926,0.124496624,0.090543,0.049044125,0.033953626,0.030181,0.026408374,0.026408374,0.018863125,0.00754525,0.003772625,0.003772625,0.0,0.011317875,0.041498873,0.071679875,0.07922512,0.049044125,0.033953626,0.02263575,0.026408374,0.090543,0.2867195,0.543258,0.94692886,1.2525115,1.3996439,1.5128226,1.8900851,1.9579924,1.8334957,1.6260014,1.4147344,2.0145817,2.897376,3.772625,4.293247,4.0480266,3.4972234,2.9049213,2.7841973,3.1161883,3.3425457,4.112161,5.3873086,6.1305156,6.19465,6.3153744,7.383027,8.201687,8.43559,7.8508325,6.2851934,6.56814,7.3981175,7.798016,7.352846,6.19465,5.715527,5.4212623,5.1458607,5.1760416,6.25124,6.3342376,6.790725,7.7640624,8.7751255,8.710991,6.990674,5.9305663,5.5683947,5.7570257,6.1795597,6.0512905,5.613666,5.6476197,6.858632,9.87296,10.770844,10.182315,8.484633,6.2851934,4.4101987,3.2633207,3.0520537,3.029418,2.8332415,2.4974778,2.3880715,2.173032,1.8599042,1.5920477,1.6071383,1.629774,1.6146835,1.7542707,2.173032,2.9124665,3.712263,3.9273026,3.9725742,4.006528,3.9348478,3.6934,3.5236318,3.338773,3.0822346,2.7351532,2.5502944,2.3767538,2.2975287,2.323937,2.3993895,2.6483827,2.5993385,2.3163917,1.9127209,1.5580941,1.50905,1.6939086,2.11267,2.6144292,2.9049213,3.4670424,4.349837,5.553304,7.1264887,9.190115,10.604849,10.427535,9.190115,7.4811153,5.9117036,4.8629136,4.22534,3.4670424,2.5729303,2.04099,1.8863125,2.0258996,2.3692086,2.7728794,3.0746894,2.867195,2.8558772,2.9313297,2.9652832,2.806833,2.1541688,1.5882751,1.3694628,1.5920477,2.214531,2.806833,3.1954134,3.5839937,4.0895257,4.7346444,5.594803,5.7306175,5.4665337,5.0854983,4.821415,4.7233267,4.7535076,4.8553686,4.930821,4.8327327,4.561104,4.6026025,4.696918,4.6856003,4.52715,4.2630663,4.025391,3.85185,3.7198083,3.5387223,3.187868,2.6332922,2.3163917,2.2975287,2.2673476,1.8221779,1.6788181,1.6448646,1.5656394,1.3015556,1.0902886,1.2940104,1.6788181,1.9202662,1.5920477,1.3505998,1.2713746,1.3430545,1.5430037,1.8146327,2.0975795,2.3918443,2.6219745,2.704972,2.5729303,2.372981,2.252257,2.2183034,2.2899833,2.5201135,2.7389257,3.0181,3.0671442,2.8558772,2.5917933,2.505023,2.6182017,2.837014,3.0520537,3.1652324,3.2520027,3.440634,3.470815,3.1954134,2.565385,2.4031622,2.263575,2.0673985,1.8938577,1.991946,2.595566,3.0369632,3.3953626,3.6443558,3.663219,3.7235808,4.0593443,4.696918,5.534441,6.326692,6.952948,7.284939,7.8395147,8.68081,9.420244,8.186596,6.6322746,4.919503,3.482133,3.0256453,4.1800685,6.047518,6.900131,6.085244,4.0178456,3.2067313,3.410453,4.0593443,4.45547,3.7763977,2.3163917,1.6373192,1.8900851,2.9313297,4.3422914,5.613666,5.8513412,4.6327834,2.6446102,1.6675003,1.6939086,1.6335466,1.4411428,1.1921495,1.0714256,1.1695137,1.056335,0.8299775,0.56589377,0.28294688,0.15845025,0.22258487,0.36594462,0.4979865,0.5281675,0.44516975,0.47912338,0.5319401,0.5281675,0.41498876,0.17731337,0.094315626,0.124496624,0.21503963,0.30181,0.35462674,0.29049212,0.16222288,0.033953626,0.0150905,0.026408374,0.071679875,0.13204187,0.19994913,0.27917424,0.5017591,1.1204696,1.5052774,1.4335974,1.0789708,1.2449663,1.9957186,3.0746894,4.0970707,4.5724216,4.2102494,2.886058,1.6373192,0.97333723,0.9016574,0.845068,0.55080324,0.24899325,0.06413463,0.026408374,0.05281675,0.06790725,0.06413463,0.05281675,0.030181,0.026408374,0.02263575,0.0150905,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.97710985,1.0487897,1.1695137,1.4071891,1.7316349,2.0145817,2.293756,2.7313805,3.1463692,3.5160866,3.9688015,5.0062733,6.0248823,7.062354,8.062099,8.880759,9.367428,10.050273,11.393328,13.098554,14.0983,13.29473,13.275867,13.890805,14.992412,16.433554,17.836971,19.38752,20.89657,22.14531,22.903606,23.673222,23.854307,24.284388,25.159636,26.061293,26.121656,25.770802,25.235088,24.639013,24.016531,23.322369,22.847017,23.137508,24.291933,25.940569,28.234325,30.147047,31.207153,31.384468,31.067568,32.127674,32.587936,32.350258,31.614597,30.867619,30.429993,30.256453,31.286379,33.580135,36.300198,39.472977,41.09143,41.5781,41.231018,40.204865,38.363823,36.99436,36.485058,36.31906,35.11182,34.315796,34.4667,34.36107,33.640495,32.761475,31.4901,30.067822,28.619133,27.442074,26.97804,25.061548,22.862108,20.010002,16.954176,14.954685,13.928532,13.717264,13.815352,13.917213,13.932304,12.185578,11.208468,10.823661,10.917976,11.442371,11.321648,10.868933,10.310584,9.767326,9.276885,8.873214,7.6923823,6.300284,5.0062733,3.8593953,6.047518,8.231868,10.250222,11.09529,8.91094,6.700182,4.7836885,3.308592,2.2220762,1.2826926,0.5357128,0.2678564,0.20749438,0.20372175,0.23013012,0.362172,0.452715,0.40367088,0.3470815,0.6413463,0.87147635,0.7205714,0.513077,0.3961256,0.33576363,0.32444575,0.27540162,0.19994913,0.124496624,0.0754525,0.06413463,0.071679875,0.094315626,0.120724,0.120724,0.1358145,0.1659955,0.16976812,0.14713238,0.120724,0.10940613,0.19994913,0.36971724,0.55080324,0.62625575,0.6752999,0.7130261,0.7884786,0.9318384,1.1732863,1.6146835,1.4298248,1.0412445,0.66020936,0.3055826,0.21881226,0.150905,0.07922512,0.033953626,0.1056335,0.29049212,0.59230214,0.95824677,1.3920987,1.9542197,2.806833,3.9650288,5.0553174,5.726845,5.613666,4.7346444,3.802806,3.0897799,2.5502944,1.8297231,1.1355602,0.79602385,0.77338815,0.965792,1.2223305,0.8903395,0.69793564,0.6073926,0.56589377,0.52062225,0.47157812,0.41121614,0.38858038,0.392353,0.36594462,0.3169005,0.22258487,0.13204187,0.060362,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.033953626,0.08677038,0.1659955,0.21503963,0.2263575,0.1659955,0.09808825,0.056589376,0.0452715,0.0452715,0.071679875,0.116951376,0.150905,0.150905,0.17731337,0.24899325,0.26031113,0.1961765,0.120724,0.03772625,0.0150905,0.026408374,0.041498873,0.030181,0.018863125,0.02263575,0.02263575,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.011317875,0.0,0.0,0.03772625,0.08677038,0.120724,0.120724,0.09808825,0.056589376,0.030181,0.056589376,0.150905,0.35839936,0.8337501,1.2110126,1.3166461,1.1581959,1.5241405,1.7014539,1.7240896,1.6335466,1.448688,1.8749946,2.927557,3.9989824,4.5497856,4.074435,2.8294687,2.625747,2.7540162,2.916239,3.218049,4.587512,5.20245,5.0138187,4.5233774,4.7912335,6.462507,9.224068,9.944639,8.650629,8.529905,13.230596,13.72481,12.2119875,10.212496,8.575176,8.575176,8.254503,7.118943,5.6778007,5.4476705,5.5570765,6.417235,8.333729,10.910432,13.045737,8.786444,6.730363,6.7454534,7.6093845,7.0359454,5.8136153,5.0062733,5.613666,7.1868505,7.798016,7.5037513,6.907676,6.043745,4.9345937,3.6179473,3.2633207,2.7804246,2.2183034,1.7391801,1.6184561,1.569412,1.5203679,1.5316857,1.6825907,2.0598533,1.9240388,1.5354583,1.2110126,1.2261031,1.7995421,2.5314314,3.410453,4.2894745,4.8629136,4.67051,4.1800685,3.821669,3.3576362,2.7728794,2.2598023,2.5616124,2.9501927,3.3538637,3.6179473,3.5085413,3.4368613,3.4444065,3.2746384,2.8747404,2.4107075,2.4597516,3.1048703,3.9273026,4.406426,3.904667,3.4896781,3.2218218,3.270866,3.904667,5.4778514,6.700182,7.488661,7.322665,6.119198,4.22534,2.444661,1.7354075,1.4826416,1.3694628,1.358145,1.4562333,1.7655885,2.3428001,2.9803739,3.1727777,3.1124156,3.1161883,3.127506,3.0256453,2.625747,1.8561316,1.5165952,1.4562333,1.629774,2.1051247,2.4710693,2.9954643,3.62172,4.1989317,4.45547,4.689373,5.2665844,5.5193505,5.2364035,4.7006907,3.8556228,3.3463185,2.9539654,2.757789,3.1124156,3.8443048,4.7610526,5.523123,6.0626082,6.5756855,6.1003346,5.1835866,4.244203,3.5877664,3.4179983,2.7691069,2.1881225,1.780679,1.6071383,1.6939086,1.4260522,1.0110635,0.724344,0.6149379,0.52062225,0.543258,0.68661773,0.80734175,0.83752275,0.76207024,0.77338815,0.8601585,1.056335,1.327964,1.5731846,1.6561824,1.8523588,2.1654868,2.5125682,2.7313805,2.5616124,2.5012503,2.565385,2.776652,3.1425967,3.3010468,3.3312278,3.3463185,3.3953626,3.4934506,3.6028569,3.6141748,3.4745877,3.2255943,3.006782,2.957738,2.9615107,3.0445085,3.078462,2.8219235,2.6408374,2.5012503,2.3993895,2.3465726,2.3956168,2.9200118,3.591539,4.3309736,5.138315,6.1041074,7.152897,8.412953,9.333474,9.49947,8.620448,7.997965,7.6131573,7.3075747,7.0510364,6.94163,6.771862,5.8588867,4.67051,3.5387223,2.6710186,3.0256453,4.093298,5.111907,5.4703064,4.7006907,3.7235808,3.169005,2.8747404,2.71629,2.595566,2.082489,2.0636258,2.3390274,2.7200627,3.0369632,3.097325,3.0030096,2.5502944,1.8787673,1.448688,1.3770081,1.1393328,0.7167987,0.25276586,0.0452715,0.1056335,0.150905,0.19994913,0.24899325,0.26031113,0.32067314,0.362172,0.44894236,0.5281675,0.44139713,0.22258487,0.150905,0.094315626,0.02263575,0.0,0.03772625,0.10940613,0.23013012,0.35085413,0.35085413,0.23013012,0.14335975,0.071679875,0.0150905,0.0150905,0.026408374,0.056589376,0.11317875,0.19240387,0.29049212,0.58475685,0.7922512,0.7205714,0.47157812,0.45648763,0.935611,1.6863633,2.9237845,4.217795,4.485651,3.3123648,2.2786655,1.8825399,2.2598023,3.1727777,2.4899325,1.659955,0.87902164,0.29426476,0.0150905,0.003772625,0.06413463,0.1056335,0.1056335,0.090543,0.06790725,0.041498873,0.030181,0.026408374,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.9016574,1.056335,1.1657411,1.2751472,1.4147344,1.5882751,1.8485862,2.214531,2.6823363,3.1916409,3.6254926,4.0970707,5.451443,6.7567716,7.5112963,7.635793,8.903395,10.125726,11.389555,12.623203,13.573905,13.385274,12.683565,12.642066,13.517315,14.664193,16.06761,18.312323,20.839981,23.23937,25.246407,26.034885,26.683777,27.78161,28.819082,28.1966,26.842226,25.382221,23.97126,22.703657,21.613369,21.11161,20.692848,20.549488,21.53037,25.12191,28.023058,30.331905,30.92798,30.048958,29.32084,29.260479,29.701876,30.214954,30.629942,31.041159,30.735577,30.92798,31.954134,33.670677,35.432495,37.164127,38.446823,39.46543,40.17091,40.318043,39.197575,37.760204,36.334152,35.06278,33.915897,32.07486,30.331905,28.924715,27.800474,26.608324,25.261497,23.933533,22.986605,22.503708,22.315077,20.398582,18.814081,17.41821,16.4411,16.478827,16.263786,15.852571,15.116908,14.200161,13.528633,12.90615,12.121444,11.348056,10.665211,10.076681,9.484379,8.89585,8.360137,7.907422,7.5565677,7.0057645,5.907931,4.647874,3.5462675,2.848332,4.0178456,5.3344917,6.477597,6.862405,5.6023483,4.4101987,3.259548,2.0447628,0.94692886,0.42630664,0.36594462,0.4376245,0.4979865,0.47912338,0.3734899,0.3055826,0.35462674,0.4979865,0.62625575,0.56589377,0.60362,0.63002837,0.5394854,0.35462674,0.21503963,0.181086,0.14335975,0.1056335,0.0754525,0.0754525,0.08299775,0.10186087,0.11317875,0.11317875,0.1358145,0.1358145,0.120724,0.18485862,0.33953625,0.5017591,0.51684964,0.55457586,0.5998474,0.60362,0.49044126,0.724344,1.0299267,1.1091517,0.9393836,0.784706,0.66775465,0.58098423,0.4678055,0.30935526,0.10940613,0.11317875,0.10940613,0.09808825,0.11317875,0.26408374,0.36971724,0.41876137,0.452715,0.56589377,0.8903395,1.6071383,2.535204,3.2746384,3.5123138,2.9916916,2.191895,1.4864142,1.0487897,0.8978847,0.9280658,0.94315624,0.84884065,0.8111144,0.8865669,1.026154,0.9507015,0.80734175,0.6375736,0.52062225,0.58098423,0.49044126,0.35839936,0.32067314,0.35839936,0.3055826,0.18863125,0.120724,0.071679875,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.00754525,0.0,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.00754525,0.003772625,0.003772625,0.003772625,0.003772625,0.02263575,0.05281675,0.090543,0.13958712,0.124496624,0.1056335,0.094315626,0.07922512,0.0452715,0.0452715,0.071679875,0.1358145,0.20749438,0.23767537,0.21503963,0.18485862,0.14335975,0.094315626,0.049044125,0.02263575,0.02263575,0.041498873,0.05281675,0.030181,0.026408374,0.02263575,0.011317875,0.003772625,0.003772625,0.003772625,0.011317875,0.0150905,0.011317875,0.0,0.0,0.0150905,0.06790725,0.14335975,0.18485862,0.14713238,0.090543,0.060362,0.08299775,0.13958712,0.271629,0.52439487,0.845068,1.2902378,2.052308,2.5616124,2.625747,2.474842,2.2748928,2.1202152,2.2748928,3.2105038,4.055572,4.1272516,2.927557,2.6182017,2.4899325,2.1805773,2.0372176,3.1350515,4.979865,7.152897,7.8508325,6.858632,5.534441,5.8702044,6.722818,7.281166,7.0887623,6.039973,6.4926877,6.387054,6.0324273,5.6815734,5.5495315,5.987156,5.1835866,4.1083884,3.429316,3.519859,3.783943,4.719554,6.5341864,8.488406,8.89585,7.752744,6.9755836,7.069899,7.635793,7.375482,5.8437963,5.6815734,5.9984736,5.9192486,4.5761943,4.6629643,4.776143,4.5233774,3.8782585,3.2255943,2.746471,2.1503963,1.8863125,2.1051247,2.6672459,3.1954134,3.4670424,3.6443558,3.99521,4.878004,4.9421387,4.3347464,3.097325,1.7089992,1.0940613,1.4034165,1.9429018,2.5616124,3.1576872,3.7047176,3.5085413,3.3161373,3.0671442,2.776652,2.5389767,2.6785638,3.1350515,3.4255435,3.4217708,3.350091,3.4444065,3.4783602,3.3764994,3.0445085,2.372981,2.2296214,2.3314822,2.4786146,3.0218725,4.8930945,6.6850915,5.240176,3.4783602,2.7691069,2.927557,3.8858037,4.776143,5.3646727,5.2250857,3.7613072,2.674791,2.1051247,1.8900851,1.841041,1.7618159,1.5845025,1.6335466,2.263575,3.6481283,5.7872066,5.5985756,4.8742313,3.572676,2.3163917,2.3918443,2.5502944,2.5012503,2.2899833,2.0183544,1.8485862,2.0108092,2.4069347,2.9728284,3.6368105,4.3196554,4.749735,5.142088,5.3344917,5.3156285,5.2364035,5.0779533,4.7950063,4.349837,3.772625,3.1614597,2.7502437,3.1916409,4.315883,5.6476197,6.405917,5.8702044,4.538468,3.4594972,2.9313297,2.4672968,1.7882242,1.3468271,1.0601076,0.8941121,0.8639311,0.73188925,0.5998474,0.513077,0.47157812,0.43385187,0.41876137,0.4640329,0.49421388,0.482896,0.47157812,0.5017591,0.6451189,0.8639311,1.1091517,1.3015556,1.5052774,1.7467253,1.961765,2.1088974,2.1315331,1.9542197,1.8221779,1.8033148,1.9127209,2.142851,2.3314822,2.4861598,2.6634734,2.867195,3.0445085,3.259548,3.5538127,3.519859,3.1463692,2.7992878,2.7200627,2.9086938,3.180323,3.3689542,3.3350005,2.9954643,2.7389257,2.6710186,2.7917426,3.0181,3.4632697,4.074435,4.644101,5.2288585,6.115425,8.065872,9.122208,9.49947,9.420244,9.144843,8.2507305,7.2170315,6.507778,6.349328,6.749226,7.454707,7.8244243,7.443389,6.1606965,4.074435,2.9426475,2.9313297,3.8405323,4.938366,4.930821,4.285702,3.361409,2.9464202,3.1765501,3.5349495,3.7160356,3.5538127,3.2784111,3.0822346,3.1463692,3.470815,3.6707642,3.500996,2.9200118,2.071171,1.4034165,0.84129536,0.4376245,0.20749438,0.1056335,0.09808825,0.17731337,0.3169005,0.4678055,0.5394854,0.72811663,0.8903395,0.754525,0.392353,0.211267,0.28294688,0.25276586,0.18485862,0.13204187,0.14713238,0.62248313,1.1204696,1.6561824,2.1051247,2.1956677,1.6712729,0.7092535,0.1056335,0.033953626,0.06413463,0.08677038,0.11317875,0.14335975,0.17354076,0.20372175,0.46026024,0.66775465,0.6073926,0.36594462,0.33576363,0.8601585,2.2447119,3.7914882,4.9760923,5.4363527,3.7386713,2.8219235,2.6446102,2.927557,3.150142,2.444661,1.3996439,0.7205714,0.52439487,0.32067314,0.0754525,0.018863125,0.03772625,0.06790725,0.1056335,0.12826926,0.116951376,0.08299775,0.049044125,0.026408374,0.0150905,0.011317875,0.00754525,0.0,0.0,0.65643674,0.8639311,1.0638802,1.237421,1.388326,1.5354583,1.6373192,1.9542197,2.425798,2.9501927,3.3463185,3.7575345,4.6290107,5.515578,6.2361493,6.8774953,8.273367,9.95973,11.627231,13.155144,14.588741,13.52486,12.645839,12.706201,13.611631,14.422746,15.350811,16.807045,19.1008,21.998177,24.699375,26.193335,27.970242,29.784874,30.716713,29.188799,27.596752,26.148064,24.69183,23.156372,21.560553,20.406128,20.606077,21.171972,22.062311,24.17498,26.721502,28.573862,29.264252,29.256706,29.928234,30.275316,30.577126,30.8148,31.007204,31.22979,31.08643,30.607307,30.505445,31.161882,32.606796,33.565044,34.444065,35.406086,36.156837,35.96821,35.191048,34.991096,34.210163,32.572845,30.71294,29.294434,27.800474,26.491373,25.54067,25.02382,23.409138,21.273832,20.002459,19.76101,19.500698,18.376457,17.520071,16.82968,16.316603,16.120426,15.901614,15.448899,14.690601,13.713491,12.770335,12.00072,11.117926,10.367173,9.8239155,9.367428,8.967529,8.601585,8.235641,7.7829256,7.1076255,6.3229194,5.3873086,4.610148,4.044254,3.4745877,3.3350005,3.3727267,3.3840446,3.1312788,2.3390274,1.841041,1.388326,0.9205205,0.513077,0.36971724,0.42630664,0.47912338,0.4979865,0.47912338,0.40367088,0.30935526,0.34330887,0.48666862,0.67152727,0.7884786,0.694163,0.573439,0.4074435,0.2263575,0.10940613,0.08677038,0.071679875,0.06413463,0.06790725,0.1056335,0.13204187,0.16222288,0.19240387,0.271629,0.48666862,0.47157812,0.26408374,0.16976812,0.2678564,0.392353,0.47535074,0.4678055,0.41876137,0.362172,0.29426476,0.47912338,0.70170826,0.7922512,0.73188925,0.6488915,0.52439487,0.39989826,0.2867195,0.181086,0.08677038,0.23013012,0.2678564,0.23013012,0.18485862,0.2678564,0.29426476,0.26408374,0.21503963,0.21503963,0.35839936,0.7582976,1.2562841,1.6524098,1.7995421,1.5920477,1.146878,0.7884786,0.58475685,0.56589377,0.7092535,0.95824677,1.2600567,1.3920987,1.3128735,1.1959221,1.1053791,0.995973,0.8865669,0.8111144,0.814887,0.66775465,0.4678055,0.3470815,0.31312788,0.24522063,0.15467763,0.071679875,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.00754525,0.00754525,0.00754525,0.00754525,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0150905,0.030181,0.049044125,0.06790725,0.094315626,0.09808825,0.094315626,0.07922512,0.060362,0.03772625,0.060362,0.07922512,0.11317875,0.1659955,0.22258487,0.16976812,0.116951376,0.0754525,0.041498873,0.02263575,0.0150905,0.018863125,0.026408374,0.030181,0.02263575,0.0150905,0.00754525,0.003772625,0.003772625,0.018863125,0.011317875,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0150905,0.05281675,0.10186087,0.1358145,0.1056335,0.0754525,0.08299775,0.116951376,0.12826926,0.181086,0.29426476,0.46026024,0.73566186,1.2562841,1.6448646,1.7580433,1.750498,1.7052265,1.6486372,1.720317,2.1353056,2.5314314,2.6332922,2.2748928,2.3918443,2.2183034,2.0636258,2.2673476,3.187868,3.9876647,5.855114,7.7187905,8.45068,6.8737226,7.3679366,9.1976595,9.846551,8.646856,6.809588,5.3194013,5.6853456,6.3832817,6.470052,5.587258,6.326692,6.1531515,5.142088,3.9914372,4.006528,4.2027044,4.195159,4.949684,6.3153744,7.062354,6.752999,6.971811,7.6131573,7.8131065,5.934339,4.6214657,4.4931965,4.395108,3.893349,3.2935016,3.9310753,4.0291634,3.7537618,3.2859564,2.8332415,2.4672968,2.1579416,2.123988,2.516341,3.4255435,4.315883,5.0213637,6.33801,8.284684,10.125726,9.208978,7.062354,4.349837,2.1164427,1.7957695,1.6712729,1.5015048,1.4373702,1.569412,1.9089483,2.033445,2.535204,2.9313297,3.0218725,2.8558772,2.7426984,2.957738,3.2859564,3.5500402,3.62172,3.7650797,3.9084394,4.1310244,4.357382,4.3611546,4.4516973,4.4743333,4.4403796,4.666737,5.783434,6.458734,5.27413,3.651901,2.5616124,2.5012503,3.500996,5.0741806,6.221059,6.379509,5.413717,4.878004,4.7346444,4.927048,5.070408,4.4630156,3.7914882,3.2142766,3.0935526,3.531177,4.3686996,3.9386206,3.4142256,2.7351532,2.2220762,2.5729303,3.2859564,3.5990841,3.3538637,2.7653341,2.4371157,2.4371157,2.625747,2.9728284,3.451952,4.032936,4.7950063,5.0968165,5.0666356,4.98741,5.3269467,5.4250345,5.2779026,4.957229,4.496969,3.8707132,3.2670932,3.470815,4.1272516,4.7950063,4.927048,4.727099,3.953711,3.0256453,2.263575,1.8900851,1.5279131,1.2751472,1.056335,0.8526133,0.70170826,0.69039035,0.8601585,1.0601076,1.0902886,0.724344,0.5394854,0.4640329,0.47535074,0.58098423,0.845068,1.2034674,1.0299267,0.79602385,0.724344,0.7582976,0.88279426,1.0374719,1.2110126,1.3694628,1.4713237,1.5354583,1.7316349,1.7278622,1.50905,1.3958713,1.5505489,1.7618159,2.0598533,2.4220252,2.8030603,2.8181508,2.9124665,3.0897799,3.2520027,3.1576872,3.1161883,3.2972744,3.7047176,4.2517486,4.7346444,4.425289,4.044254,3.6858547,3.5764484,4.0706625,4.7044635,5.4363527,5.383536,4.7308717,4.719554,6.115425,6.94163,7.356619,7.5263867,7.647111,7.424526,7.1000805,6.937857,7.1868505,8.099826,8.967529,8.990166,8.514814,7.6282477,6.138061,4.247976,3.4972234,3.6707642,4.183841,4.112161,3.5802212,2.848332,2.6332922,3.0445085,3.5839937,4.0706625,3.9574835,3.4066803,2.6144292,1.81086,2.3692086,2.8143783,2.8785129,2.3126192,0.8903395,0.56212115,0.35085413,0.24899325,0.23390275,0.241448,0.22258487,0.392353,0.66775465,0.8865669,0.80356914,1.1317875,1.4826416,1.3505998,0.7884786,0.42630664,0.35462674,0.33576363,0.33576363,0.362172,0.4678055,0.9205205,1.3015556,1.5958204,1.7278622,1.5279131,1.0223814,0.41121614,0.08677038,0.11317875,0.22258487,0.35839936,0.34330887,0.26031113,0.181086,0.1659955,0.29803738,0.45648763,0.482896,0.38858038,0.35085413,0.6828451,1.6033657,2.595566,3.31991,3.6330378,2.4484336,2.04099,2.384299,3.2520027,4.22534,3.712263,2.0787163,0.91674787,0.6375736,0.46026024,0.3734899,0.23013012,0.09808825,0.030181,0.041498873,0.071679875,0.08677038,0.08677038,0.0754525,0.06790725,0.049044125,0.041498873,0.030181,0.00754525,0.0,0.46026024,0.6526641,0.91297525,1.2298758,1.5279131,1.7014539,1.7957695,2.1994405,2.6672459,3.0935526,3.5047686,4.1612053,4.52715,4.859141,5.3986263,6.379509,7.537705,9.012801,10.484125,11.849815,13.257004,12.483616,12.0724,12.396846,13.340002,14.313339,14.592513,15.237633,16.705183,19.119663,22.273579,24.797464,27.189308,28.954897,29.524563,28.26828,26.812046,26.125427,25.555761,24.574879,22.737612,21.794455,22.296213,22.933788,23.314823,23.978804,25.808527,26.853544,27.366621,27.785383,28.751175,29.59247,30.060276,30.241362,30.094229,29.464201,28.871899,28.030603,27.589207,27.88347,28.95867,29.388748,29.913143,30.629942,31.33165,31.50142,31.120384,31.38824,31.188292,30.188545,28.788902,28.106056,26.93277,25.66894,24.650331,24.17498,22.40562,20.326904,19.119663,18.829172,18.357594,17.772837,17.30503,16.791954,16.15438,15.380992,14.913187,14.5132885,14.068119,13.472044,12.642066,11.823407,10.993429,10.212496,9.593785,9.288202,9.178797,9.020347,8.850578,8.601585,8.126234,7.3717093,6.6850915,6.255012,5.904158,5.0666356,3.9461658,2.916239,2.033445,1.2902378,0.6187105,0.45648763,0.41876137,0.5093044,0.65643674,0.7469798,0.77716076,0.7696155,0.73566186,0.68661773,0.62248313,0.543258,0.52062225,0.5281675,0.56589377,0.6526641,0.5470306,0.3772625,0.21881226,0.11317875,0.071679875,0.071679875,0.06790725,0.09808825,0.1659955,0.23767537,0.20749438,0.20372175,0.23013012,0.32067314,0.5470306,0.6187105,0.52062225,0.41121614,0.35462674,0.35085413,0.43007925,0.3734899,0.2867195,0.2263575,0.21503963,0.29049212,0.36594462,0.41876137,0.44516975,0.4376245,0.38858038,0.29426476,0.19240387,0.124496624,0.10186087,0.27540162,0.32821837,0.29049212,0.21881226,0.18485862,0.16222288,0.124496624,0.09808825,0.1056335,0.1961765,0.4074435,0.5772116,0.724344,0.845068,0.935611,0.7432071,0.6488915,0.69793564,0.8337501,0.91297525,1.1996948,1.7655885,1.9504471,1.6335466,1.2336484,1.056335,0.9507015,0.9016574,0.90543,0.965792,0.7884786,0.5357128,0.31312788,0.17354076,0.12826926,0.090543,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.003772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.041498873,0.06413463,0.094315626,0.1056335,0.120724,0.09808825,0.060362,0.026408374,0.018863125,0.07922512,0.116951376,0.1358145,0.14335975,0.1659955,0.120724,0.08299775,0.056589376,0.033953626,0.02263575,0.0150905,0.0150905,0.011317875,0.00754525,0.00754525,0.0,0.0,0.0,0.003772625,0.02263575,0.011317875,0.00754525,0.00754525,0.00754525,0.00754525,0.00754525,0.0150905,0.026408374,0.0452715,0.071679875,0.07922512,0.090543,0.10940613,0.124496624,0.116951376,0.15845025,0.241448,0.32821837,0.4074435,0.513077,0.6526641,0.73188925,0.814887,0.91674787,0.9997456,1.1242423,1.3091009,1.4562333,1.539231,1.6222287,1.7316349,1.6448646,1.780679,2.3805263,3.4859054,3.9688015,5.0477724,6.4964604,7.4811153,6.571913,7.383027,9.050528,9.374973,8.186596,7.364164,5.6891184,5.772116,6.4021444,6.5945487,5.587258,6.187105,6.752999,6.217286,4.8327327,4.1762958,5.783434,6.1229706,5.8966126,5.7909794,6.48137,6.56814,7.4094353,8.107371,7.77538,5.515578,4.402653,4.085753,3.8669407,3.5085413,3.2331395,4.0593443,4.617693,4.644101,4.191386,3.6179473,3.1614597,2.8219235,2.71629,2.9652832,3.6934,4.2630663,5.0138187,6.4511886,8.314865,9.590013,8.461998,6.360646,4.006528,2.3013012,2.323937,2.0560806,1.4826416,0.98465514,0.754525,0.784706,0.94692886,1.5467763,2.1692593,2.5767028,2.7087448,2.757789,2.9426475,3.3123648,3.7613072,4.063117,4.7610526,5.342037,5.915476,6.485142,6.9793563,7.1604424,7.122716,7.2170315,7.61693,8.296002,8.52236,7.273621,5.240176,3.3312278,2.6521554,3.429316,4.9987283,6.307829,6.72659,6.0739264,5.6023483,5.9230213,6.7379084,7.484888,7.3415284,6.2889657,5.4778514,5.0515447,4.851596,4.4177437,3.7801702,3.3048196,2.969056,2.8521044,3.1237335,3.731126,4.1083884,3.9801195,3.4481792,2.9652832,2.9124665,3.0030096,3.2331395,3.6254926,4.22534,5.0666356,5.292993,5.142088,4.949684,5.172269,5.1081343,4.859141,4.5460134,4.266839,4.1008434,4.036709,4.406426,4.745962,4.7836885,4.4177437,4.3196554,3.9499383,3.2520027,2.4107075,1.8599042,1.5316857,1.2940104,1.146878,1.0789708,1.0450171,1.146878,1.3392819,1.4675511,1.358145,0.83752275,0.66020936,0.5696664,0.573439,0.6790725,0.91297525,1.1996948,0.9016574,0.5394854,0.35839936,0.32067314,0.38858038,0.4640329,0.573439,0.73188925,0.9205205,1.0789708,1.3317367,1.3543724,1.1317875,0.9695646,1.116697,1.3317367,1.6335466,1.9957186,2.372981,2.2748928,2.2560298,2.5767028,3.1614597,3.6179473,3.863168,4.0103,4.2328854,4.6327834,5.2364035,5.560849,5.715527,5.6778007,5.6061206,5.8211603,5.926794,6.1418333,5.7117543,4.7874613,4.436607,5.062863,5.560849,5.9909286,6.3644185,6.6586833,6.677546,6.771862,6.983129,7.2924843,7.624475,7.726336,7.3717093,7.0284004,6.7152724,6.009792,4.515832,3.8858037,3.8103511,3.942393,3.9348478,3.451952,2.9539654,2.8822856,3.338773,4.0782075,4.82896,4.919503,4.2328854,2.916239,1.358145,1.4034165,1.5203679,1.539231,1.2336484,0.3055826,0.35462674,0.38480774,0.5055317,0.70170826,0.814887,0.48666862,0.47535074,0.66020936,0.84129536,0.7582976,1.1053791,1.4147344,1.3505998,0.91674787,0.48666862,0.2867195,0.3055826,0.35839936,0.38480774,0.41876137,0.6187105,0.7507524,0.7922512,0.7394345,0.62625575,0.44894236,0.38480774,0.35839936,0.32444575,0.271629,0.3470815,0.3055826,0.211267,0.12826926,0.10940613,0.18863125,0.32444575,0.40367088,0.39989826,0.362172,0.48666862,0.8111144,1.2298758,1.6109109,1.8334957,1.4524606,1.6410918,2.372981,3.4330888,4.4177437,3.8556228,2.4786146,1.6561824,1.659955,1.6637276,1.7731338,1.7089992,1.6109109,1.599593,1.780679,1.1091517,0.4074435,0.056589376,0.071679875,0.08677038,0.06413463,0.060362,0.0452715,0.018863125,0.00754525,0.39989826,0.5281675,0.76207024,1.1317875,1.5430037,1.7693611,2.052308,2.5804756,3.0143273,3.3425457,3.8895764,4.908185,5.1798143,5.2628117,5.572167,6.3644185,7.17176,7.937603,8.571404,9.1825695,10.103089,10.868933,11.34051,11.864905,12.653384,13.773854,13.422999,13.660675,14.252977,15.569623,18.602814,21.654867,23.95617,25.502945,26.253696,26.14429,25.042685,25.212452,25.729303,25.66894,24.095757,23.925987,24.061802,23.910898,23.567589,23.824127,24.944597,25.506718,25.789665,25.921707,25.868889,26.668686,27.264761,27.525072,27.238352,26.121656,24.903097,24.337204,24.480564,25.0955,25.63876,25.702894,26.091475,26.570599,27.094994,27.830654,27.796701,27.551481,27.453392,27.59298,27.78161,27.600525,26.366877,25.087955,24.137255,23.258234,21.258741,19.90437,19.112118,18.648085,18.135008,17.599297,17.1164,16.59955,15.98084,15.237633,14.634012,14.237886,13.977575,13.70972,13.185325,12.811834,12.377983,11.710228,10.887795,10.26154,10.065364,9.910686,9.808825,9.767326,9.812597,9.397609,9.035437,8.707218,8.126234,6.730363,5.1534057,3.5689032,2.2447119,1.2713746,0.5583485,0.41498876,0.4678055,0.6828451,0.97710985,1.2261031,1.2487389,1.2487389,1.2336484,1.177059,1.0110635,0.84884065,0.7432071,0.6111652,0.422534,0.20372175,0.150905,0.1056335,0.071679875,0.06413463,0.08677038,0.1056335,0.116951376,0.19240387,0.331991,0.45648763,0.39989826,0.31312788,0.24899325,0.241448,0.29049212,0.452715,0.6451189,0.70170826,0.6149379,0.543258,0.55457586,0.42630664,0.32067314,0.29803738,0.32821837,0.31312788,0.29049212,0.25276586,0.20749438,0.15467763,0.120724,0.12826926,0.12826926,0.10940613,0.124496624,0.241448,0.2678564,0.24522063,0.18863125,0.07922512,0.049044125,0.026408374,0.030181,0.08299775,0.19994913,0.38858038,0.44139713,0.47157812,0.5394854,0.6413463,0.6187105,0.69039035,0.90543,1.1581959,1.20724,1.4600059,1.9881734,2.0447628,1.5203679,0.965792,0.7394345,0.59607476,0.543258,0.60362,0.814887,0.6790725,0.44516975,0.18863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02263575,0.033953626,0.06790725,0.120724,0.1358145,0.12826926,0.08299775,0.033953626,0.00754525,0.00754525,0.090543,0.15467763,0.17354076,0.150905,0.1056335,0.08299775,0.06790725,0.056589376,0.041498873,0.033953626,0.026408374,0.02263575,0.018863125,0.003772625,0.003772625,0.003772625,0.0,0.0,0.003772625,0.011317875,0.003772625,0.011317875,0.018863125,0.018863125,0.0150905,0.011317875,0.003772625,0.0,0.00754525,0.0452715,0.094315626,0.12826926,0.12826926,0.10940613,0.11317875,0.19240387,0.29803738,0.38858038,0.43007925,0.39989826,0.33953625,0.29049212,0.32821837,0.47535074,0.694163,0.8903395,1.1732863,1.3166461,1.2336484,0.9922004,0.8941121,0.9393836,1.1732863,1.81086,3.2482302,4.236658,4.8402777,4.9119577,4.67051,4.719554,5.5193505,5.7079816,5.7570257,6.0324273,6.820906,5.9532022,5.7306175,5.798525,5.7872066,5.3571277,5.3571277,5.8702044,5.696664,4.587512,3.229367,6.4926877,8.348819,8.028146,6.470052,6.3455553,6.7869525,7.5905213,7.745199,6.9755836,5.7381625,4.817642,4.4894238,4.45547,4.2706113,3.350091,3.9008942,5.2779026,6.0626082,5.873977,5.3684454,4.745962,4.146115,3.7914882,3.7160356,3.7801702,3.4972234,3.7537618,4.112161,4.2592936,4.0178456,4.085753,4.104616,3.9008942,3.4179983,2.7200627,2.2786655,1.629774,1.0714256,0.7432071,0.6488915,0.5998474,0.6828451,1.0110635,1.5505489,2.1202152,2.674791,3.1463692,3.561358,4.006528,4.6214657,6.1305156,7.3490734,8.197914,8.741172,9.175024,9.114662,8.952439,9.363655,10.510533,12.053536,13.113645,11.272603,8.013056,4.7535076,2.8521044,2.957738,3.6934,4.6742826,5.2892203,4.727099,4.085753,4.647874,5.8588867,7.194396,8.171506,7.213259,6.692637,6.6322746,6.752999,6.458734,5.938112,5.2779026,4.557331,3.9574835,3.7763977,3.863168,4.044254,4.1008434,3.863168,3.2255943,3.1199608,3.2633207,3.5689032,4.032936,4.708236,5.323174,5.5193505,5.481624,5.3344917,5.1571784,4.798779,4.353609,3.8971217,3.591539,3.6707642,4.266839,4.9723196,5.3873086,5.330719,4.8365054,4.557331,4.2592936,3.8593953,3.2746384,2.4220252,1.7580433,1.3317367,1.1921495,1.3053282,1.5543215,1.8259505,1.9579924,1.8599042,1.5505489,1.1921495,1.0751982,0.90543,0.76207024,0.67152727,0.6111652,0.43385187,0.29049212,0.2263575,0.21503963,0.18485862,0.21503963,0.241448,0.2867195,0.3734899,0.5357128,0.59230214,0.65643674,0.7922512,0.935611,0.9016574,0.94315624,1.0601076,1.2525115,1.478869,1.6788181,1.6825907,1.7882242,2.142851,2.8256962,3.8443048,4.5761943,4.779916,4.5837393,4.3309736,4.561104,5.6325293,6.6134114,7.284939,7.4697976,7.0359454,6.221059,5.6815734,5.409944,5.3382645,5.3382645,5.481624,5.6325293,5.8966126,6.2399216,6.485142,6.2323766,6.0286546,5.983383,5.8513412,5.040227,4.2592936,4.1612053,4.402653,4.5799665,4.2291126,3.6858547,3.6481283,3.9122121,4.3007927,4.6554193,4.247976,3.802806,3.640583,3.953711,4.7836885,5.6551647,5.9305663,5.3344917,3.983892,2.3805263,1.4637785,0.845068,0.56212115,0.58475685,0.84884065,1.0110635,1.026154,1.1581959,1.3770081,1.3619176,0.6488915,0.35839936,0.331991,0.422534,0.49044126,0.724344,0.77716076,0.7582976,0.6752999,0.4376245,0.452715,0.5696664,0.5772116,0.41121614,0.15467763,0.090543,0.06790725,0.056589376,0.10940613,0.35839936,0.5319401,0.72811663,0.73566186,0.5055317,0.1659955,0.06413463,0.049044125,0.07922512,0.12826926,0.18485862,0.2678564,0.331991,0.36594462,0.3734899,0.35839936,0.35462674,0.4074435,0.6073926,0.91297525,1.1732863,1.3392819,1.8636768,2.5880208,3.2142766,3.2784111,2.4861598,2.082489,2.2748928,2.8558772,3.2029586,3.5387223,3.7650797,3.8480775,3.8405323,3.904667,2.3616633,0.8262049,0.0452715,0.03772625,0.06413463,0.056589376,0.056589376,0.0452715,0.026408374,0.018863125,0.41121614,0.52062225,0.63002837,0.77338815,0.97710985,1.2826926,1.7089992,2.1013522,2.4182527,2.8256962,3.6934,5.036454,5.66271,6.1342883,6.730363,7.462252,8.084735,8.578949,8.7600355,8.967529,10.038955,11.151879,12.306303,13.124963,13.396591,13.091009,12.2119875,11.827179,11.921495,12.562841,13.917213,15.746937,18.03692,21.19838,24.28816,25.008732,24.971004,25.174726,25.370903,25.291677,24.657877,23.511,22.767792,22.303759,21.934042,21.409647,21.967995,23.190327,24.514517,25.453901,25.589716,26.016022,25.58217,24.631468,23.778856,23.925987,23.390276,23.043194,23.111101,23.503454,23.820354,23.941078,24.631468,24.87669,24.156118,22.447119,22.043447,21.998177,22.266033,22.82438,23.665676,23.839218,23.322369,23.424229,24.208935,24.491882,21.522825,19.410156,18.078419,17.463482,17.486116,17.108854,16.55428,16.28265,16.286423,16.127972,15.652621,14.992412,14.366156,13.86817,13.487134,13.487134,13.72481,14.18507,14.335975,13.151371,12.128989,11.751727,11.404645,10.876478,10.374719,10.352083,10.355856,10.133271,9.303293,7.3377557,5.617439,3.953711,2.5804756,1.5845025,0.9016574,0.5696664,0.4979865,0.6187105,0.935611,1.4939595,1.4600059,1.4147344,1.5165952,1.6071383,1.20724,0.7432071,0.633801,0.56212115,0.38858038,0.1659955,0.094315626,0.056589376,0.0452715,0.049044125,0.060362,0.10940613,0.1961765,0.3055826,0.44516975,0.6413463,0.8978847,0.694163,0.40367088,0.241448,0.29049212,0.21503963,0.19994913,0.35839936,0.63002837,0.76207024,0.76207024,0.47912338,0.32067314,0.41121614,0.59607476,0.47157812,0.35085413,0.22258487,0.13204187,0.1659955,0.23013012,0.271629,0.26031113,0.22258487,0.26031113,0.4074435,0.35085413,0.21503963,0.090543,0.030181,0.018863125,0.02263575,0.049044125,0.090543,0.150905,0.21503963,0.28294688,0.33953625,0.38480774,0.45648763,0.935611,1.1883769,1.2336484,1.1732863,1.2223305,1.3053282,1.4637785,1.3505998,0.9393836,0.55080324,0.3055826,0.09808825,0.0,0.033953626,0.16976812,0.181086,0.1659955,0.090543,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.018863125,0.049044125,0.060362,0.03772625,0.02263575,0.02263575,0.030181,0.030181,0.06790725,0.094315626,0.094315626,0.071679875,0.0452715,0.02263575,0.0150905,0.02263575,0.033953626,0.0452715,0.056589376,0.060362,0.049044125,0.026408374,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.011317875,0.02263575,0.03772625,0.041498873,0.0150905,0.003772625,0.0,0.0,0.00754525,0.0452715,0.094315626,0.1056335,0.11317875,0.124496624,0.1358145,0.18485862,0.2263575,0.2678564,0.31312788,0.35085413,0.33953625,0.271629,0.32067314,0.52439487,0.7922512,0.8903395,0.98842776,1.0638802,1.0638802,0.9318384,0.784706,0.63002837,0.56589377,0.633801,0.7922512,1.0638802,1.7354075,2.546522,3.2784111,3.7537618,4.534695,5.6363015,7.039718,7.967784,6.881268,6.832224,9.593785,10.868933,9.533423,7.6282477,6.8359966,5.692891,4.3196554,3.0218725,2.2899833,3.2670932,5.2779026,6.307829,6.089017,6.089017,5.80607,5.4250345,5.1760416,4.689373,2.9916916,2.8936033,3.1425967,3.1539145,2.776652,2.2899833,2.3993895,3.5349495,4.851596,5.881522,6.515323,6.3455553,6.126743,5.8098426,5.3080835,4.5007415,3.610402,3.059599,2.746471,2.7125173,3.127506,5.13077,7.424526,8.669493,7.91874,4.6214657,3.059599,2.0296721,1.3694628,0.94315624,0.62625575,0.51684964,0.5357128,0.7167987,1.0827434,1.6335466,2.4031622,3.1614597,3.7952607,4.436607,5.462761,6.903904,8.43559,9.533423,10.054046,10.238904,9.774872,9.740918,10.570895,12.298758,14.558559,14.973549,13.373956,10.057818,6.149379,3.5839937,2.7917426,2.8143783,3.0143273,2.969056,2.4559789,2.2748928,2.546522,3.2029586,4.006528,4.5912848,4.6554193,4.4139714,4.6026025,5.323174,6.043745,6.3719635,6.224831,5.7192993,4.961002,4.0593443,3.9499383,4.1310244,4.2102494,4.032936,3.6783094,3.2369123,3.5047686,4.0216184,4.429062,4.4403796,4.817642,5.168496,5.492942,5.7419353,5.828706,5.643847,5.3269467,4.82896,4.1612053,3.3425457,3.731126,4.29702,4.689373,4.606375,3.7990334,3.6292653,3.8254418,3.9688015,3.863168,3.5085413,2.5804756,1.9579924,1.5241405,1.358145,1.7240896,2.3465726,3.0256453,3.3727267,3.3274553,3.1576872,2.6106565,1.81086,1.146878,0.80734175,0.7922512,0.48666862,0.36594462,0.42630664,0.52439487,0.36594462,0.1358145,0.1056335,0.150905,0.20749438,0.24522063,0.32821837,0.67152727,1.2525115,1.6825907,1.20724,0.6790725,0.5017591,0.55080324,0.72811663,0.94692886,1.1544232,1.3355093,1.750498,2.5276587,3.663219,4.772371,5.198677,4.8138695,4.063117,3.953711,4.478106,5.168496,5.5382137,5.4250345,4.961002,4.459243,4.5535583,4.881777,5.13077,5.0213637,4.7648253,4.7535076,4.979865,5.251494,5.20245,5.3609,4.9421387,4.22534,3.5160866,3.1727777,3.2218218,3.712263,4.3347464,4.779916,4.7308717,4.0706625,3.8065786,4.074435,4.678055,5.081726,4.8138695,4.29702,3.832987,3.6481283,3.8895764,4.195159,4.346064,4.3686996,4.2102494,3.7235808,2.6974268,1.8297231,1.2298758,0.995973,1.1883769,1.5203679,1.7316349,1.7467253,1.4335974,0.58098423,0.24899325,0.26031113,0.36971724,0.44139713,0.44139713,0.5885295,0.47912338,0.45648763,0.6451189,0.97710985,1.720317,2.0447628,1.8184053,1.1808317,0.5357128,0.41121614,0.34330887,0.29049212,0.23767537,0.21503963,0.29803738,0.49421388,0.5017591,0.27917424,0.0452715,0.02263575,0.1358145,0.31312788,0.513077,0.73188925,0.7092535,0.44516975,0.3055826,0.36971724,0.44139713,0.38103512,0.422534,0.6526641,0.98842776,1.1581959,1.2713746,1.4600059,1.7014539,1.8863125,1.8599042,1.2751472,1.0940613,1.2751472,1.750498,2.3956168,3.3463185,4.006528,4.0480266,3.2935016,1.6939086,0.8639311,0.39989826,0.150905,0.026408374,0.0150905,0.026408374,0.041498873,0.041498873,0.030181,0.030181,0.47157812,0.67152727,0.9507015,1.2223305,1.4637785,1.7089992,1.8825399,2.2183034,2.5729303,2.8898308,3.180323,3.742444,4.2102494,4.6516466,5.160951,5.873977,6.809588,8.409182,9.416472,9.4013815,8.744945,10.1294985,11.25374,11.959221,12.189351,11.981857,11.736636,11.8045435,11.838497,11.876224,12.355347,13.754991,16.01102,18.772581,21.394556,22.945105,23.09601,22.941332,22.945105,23.179008,23.314823,23.348776,22.613113,21.613369,20.640032,19.783646,20.677757,21.55678,22.009495,22.243397,23.099783,24.005213,23.839218,23.348776,22.967741,22.790428,21.862362,21.734093,22.164171,22.662159,22.499935,22.009495,21.262514,20.617395,20.096773,19.395065,18.912169,19.176252,20.040184,21.511507,23.752447,23.982576,23.473272,22.65084,21.843498,21.292696,20.443855,20.11941,19.983595,19.889278,19.855326,19.828917,19.685556,19.54597,19.247932,18.33873,17.520071,17.05981,17.237123,17.96524,18.787672,19.372429,18.644312,17.222033,15.558306,13.936077,13.268322,12.925014,12.370438,11.638548,11.351829,11.563096,11.457462,10.86516,9.627739,7.594294,6.2361493,5.0175915,3.983892,3.180323,2.6823363,2.2447119,1.720317,1.7014539,2.282438,3.059599,2.444661,1.9542197,1.6109109,1.3166461,0.8639311,0.60362,0.5696664,0.51684964,0.3772625,0.26408374,0.19240387,0.13204187,0.090543,0.090543,0.16976812,0.27917424,0.4376245,0.76207024,1.1053791,1.056335,0.784706,0.56212115,0.6451189,1.146878,2.0372176,1.1921495,0.6488915,0.47535074,0.5319401,0.47157812,0.56589377,0.87902164,0.95447415,0.7054809,0.41121614,0.22258487,0.23013012,0.3169005,0.3470815,0.181086,0.1056335,0.08299775,0.12826926,0.2263575,0.32067314,0.44894236,0.32821837,0.1659955,0.06413463,0.030181,0.06790725,0.14335975,0.27540162,0.40367088,0.3961256,0.33953625,0.30181,0.28294688,0.28294688,0.2867195,0.392353,0.5696664,0.7884786,0.965792,0.97710985,0.98465514,0.98465514,0.9318384,0.80734175,0.62248313,0.3961256,0.27540162,0.18863125,0.1056335,0.033953626,0.03772625,0.033953626,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.003772625,0.0,0.00754525,0.018863125,0.011317875,0.00754525,0.003772625,0.0150905,0.03772625,0.06790725,0.094315626,0.09808825,0.08677038,0.0754525,0.071679875,0.0452715,0.026408374,0.011317875,0.0150905,0.0452715,0.06790725,0.07922512,0.071679875,0.049044125,0.026408374,0.026408374,0.018863125,0.011317875,0.0150905,0.02263575,0.026408374,0.02263575,0.018863125,0.018863125,0.003772625,0.0,0.00754525,0.011317875,0.0150905,0.033953626,0.06413463,0.09808825,0.15467763,0.21503963,0.24899325,0.2565385,0.21503963,0.18485862,0.1961765,0.241448,0.29803738,0.29049212,0.28294688,0.2867195,0.27917424,0.42630664,0.6526641,0.7507524,0.724344,0.784706,0.95824677,0.98842776,0.94692886,0.8526133,0.67152727,1.780679,2.6521554,2.7087448,2.474842,3.5953116,5.089271,6.326692,7.066127,7.2094865,6.7944975,6.5530496,6.488915,6.4549613,7.413208,11.438599,13.087236,11.714001,8.492179,4.8553686,2.4823873,2.6710186,3.4859054,4.2064767,4.466788,4.2819295,3.5802212,2.8030603,2.5314314,2.625747,2.2107582,2.2975287,3.1954134,3.7273536,3.361409,2.191895,2.3390274,2.5917933,2.6106565,2.584248,3.218049,3.9197574,4.606375,5.081726,5.191132,4.8553686,3.0860074,2.9728284,4.093298,5.80607,7.2660756,7.0510364,6.1342883,5.05909,4.06689,3.0860074,2.957738,2.4408884,1.8523588,1.388326,1.1016065,0.90543,0.80356914,0.935611,1.3807807,2.1956677,3.150142,3.904667,4.3913355,4.6856003,4.98741,6.643593,8.235641,9.6051035,10.231359,9.21275,8.054554,6.934085,7.6697464,10.627484,14.70192,18.176508,16.7995,13.000465,8.827943,5.9418845,4.961002,4.7535076,4.7610526,4.5497856,3.8103511,2.9954643,2.757789,2.927557,3.350091,3.8971217,3.7613072,3.772625,4.266839,5.1156793,5.7494807,6.19465,6.519096,6.647365,6.571913,6.3417826,5.9305663,5.451443,4.825187,4.134797,3.6179473,3.410453,3.5462675,3.6971724,3.7575345,3.8178966,4.3422914,5.081726,5.794752,6.379509,6.8661776,6.8774953,6.643593,6.1795597,5.5004873,4.6214657,4.036709,4.085753,4.285702,4.217795,3.531177,3.1539145,3.3048196,3.8858037,4.7421894,5.6589375,5.794752,5.172269,4.496969,4.2064767,4.447925,5.6363015,7.1793056,8.503497,9.009028,8.07719,6.198423,4.164978,2.4107075,1.2261031,0.7432071,0.90920264,1.7014539,2.2862108,2.2183034,1.4524606,0.8299775,0.4074435,0.20749438,0.18863125,0.2565385,0.32067314,0.40367088,0.6375736,0.9695646,1.1581959,1.0412445,1.0714256,1.297783,1.931584,3.3123648,3.0445085,2.3654358,2.2862108,2.9841464,3.8103511,4.870459,4.719554,3.9084394,2.897376,2.0372176,2.6182017,3.2935016,3.640583,3.572676,3.3236825,2.8898308,2.8634224,3.0331905,3.2255943,3.3123648,3.180323,3.059599,2.9992368,3.0897799,3.4217708,3.832987,4.044254,3.6556737,2.9237845,2.757789,3.7952607,4.9157305,5.8626595,6.3531003,6.1078796,5.674028,5.1156793,4.6214657,4.2894745,4.115934,3.99521,3.772625,3.7235808,3.9688015,4.478106,4.195159,4.0216184,4.0291634,4.063117,3.772625,3.127506,2.214531,1.6071383,1.4562333,1.4939595,1.3091009,1.0601076,0.80734175,0.573439,0.32444575,0.754525,1.3128735,1.478869,1.1921495,0.87147635,0.5583485,0.5583485,0.8526133,1.3996439,2.1466236,2.5917933,2.6031113,2.0862615,1.2449663,0.6073926,0.32067314,0.181086,0.11317875,0.06790725,0.041498873,0.1961765,0.55457586,0.8601585,0.9205205,0.6187105,0.47912338,0.5998474,0.80356914,0.935611,0.84129536,0.47535074,0.31312788,0.28294688,0.30935526,0.28294688,0.30935526,0.32821837,0.40367088,0.5281675,0.6111652,0.67152727,0.6752999,0.76584285,1.0299267,1.4939595,2.1994405,2.565385,2.6634734,2.5427492,2.2107582,3.0369632,4.478106,4.851596,3.8103511,2.3277097,1.3996439,1.6146835,2.4069347,3.0822346,2.848332,1.961765,0.8903395,0.23390275,0.090543,0.07922512,1.0110635,1.0336993,1.1431054,1.297783,1.4826416,1.7165444,1.9730829,2.354118,2.7238352,2.9992368,3.187868,3.429316,3.8858037,4.3649273,4.7572803,5.0213637,5.6891184,6.7454534,7.443389,7.5829763,7.5075235,8.59404,9.390063,10.016319,10.540714,10.970794,11.257513,11.5857315,11.7555,11.876224,12.366665,13.241914,14.354838,15.686575,17.105082,18.402864,19.828917,20.50799,20.82489,20.885252,20.500444,20.60985,20.643805,20.319359,19.662922,19.021576,19.081938,19.625195,20.123182,20.474035,20.994658,21.236107,21.032385,20.95316,21.066338,20.949387,20.37972,20.398582,20.749437,21.134245,21.228561,20.662666,19.866644,19.138527,18.561316,18.03692,17.814335,18.467,19.67424,21.254969,23.16769,23.722265,23.631723,23.114874,22.669704,23.092237,23.220507,23.231825,22.990377,22.582933,22.322622,22.473528,23.273323,23.869398,23.390276,20.949387,20.8513,21.27006,21.405874,21.104065,20.870161,20.394812,18.297232,15.931795,14.064346,12.894833,12.713746,12.604341,12.332711,11.974312,11.917723,12.045992,11.98563,11.246195,9.718282,7.707473,6.1078796,4.8742313,3.9461658,3.3840446,3.3953626,3.531177,3.6858547,3.4859054,3.0218725,2.8256962,2.41448,1.7844516,1.1657411,0.7054809,0.47535074,0.38480774,0.3734899,0.32444575,0.23390275,0.20749438,0.23013012,0.27540162,0.32067314,0.35462674,0.39989826,0.5055317,0.5772116,0.6413463,0.79602385,1.2147852,1.3317367,1.0789708,0.965792,1.1883769,1.6109109,1.0638802,0.6413463,0.38103512,0.30181,0.4074435,0.45648763,0.5394854,0.52439487,0.392353,0.2565385,0.26031113,0.28294688,0.29803738,0.26031113,0.090543,0.049044125,0.060362,0.16222288,0.30181,0.35462674,0.35085413,0.2263575,0.10186087,0.0452715,0.049044125,0.21503963,0.35462674,0.47912338,0.543258,0.4678055,0.36594462,0.30181,0.23767537,0.17354076,0.116951376,0.150905,0.2867195,0.48666862,0.62625575,0.5017591,0.55080324,0.7054809,0.69039035,0.49044126,0.35839936,0.36594462,0.31312788,0.2263575,0.12826926,0.06413463,0.041498873,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.033953626,0.041498873,0.030181,0.02263575,0.0150905,0.00754525,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.003772625,0.0150905,0.030181,0.049044125,0.06413463,0.08299775,0.08677038,0.056589376,0.033953626,0.030181,0.030181,0.030181,0.0452715,0.07922512,0.090543,0.08677038,0.071679875,0.041498873,0.033953626,0.0150905,0.00754525,0.00754525,0.011317875,0.011317875,0.00754525,0.00754525,0.011317875,0.03772625,0.00754525,0.003772625,0.011317875,0.0150905,0.011317875,0.02263575,0.03772625,0.08299775,0.14335975,0.17354076,0.17354076,0.17731337,0.1961765,0.21881226,0.1961765,0.23013012,0.26408374,0.27917424,0.2678564,0.21503963,0.22258487,0.3169005,0.38858038,0.4376245,0.59230214,0.724344,0.7884786,0.8337501,0.8337501,0.694163,1.1883769,1.6788181,1.9466745,2.2862108,3.500996,5.7079816,7.333983,8.262049,8.744945,9.431562,9.74469,9.473062,8.3525915,7.224577,8.050782,9.759781,8.986393,6.952948,5.2175403,5.7004366,5.0968165,3.7575345,3.2746384,3.6858547,3.482133,2.5578396,1.9164935,1.8297231,2.3314822,3.1765501,2.4484336,2.425798,3.3764994,4.4894238,3.9159849,3.6066296,4.3800178,4.647874,3.942393,2.9464202,3.048281,3.2972744,3.591539,3.6971724,3.259548,2.214531,2.1013522,2.7087448,3.682082,4.5460134,4.5837393,4.1574326,3.6707642,3.2821836,2.8936033,2.655928,2.1579416,1.841041,1.7769064,1.6788181,1.4600059,1.4411428,1.6448646,2.1088974,2.8936033,3.9461658,4.715781,4.938366,4.7610526,4.768598,5.6853456,7.1340337,8.926031,10.668983,11.759273,11.578186,10.816116,10.378491,11.317875,14.849052,17.108854,15.7657995,13.04951,10.416218,8.518587,8.0206,7.8508325,7.7376537,7.375482,6.458734,5.27413,4.3083377,3.9725742,4.142342,4.146115,3.5500402,3.519859,3.8895764,4.447925,4.9723196,5.6098933,6.2436943,6.7869525,7.149124,7.250985,7.122716,7.043491,6.5341864,5.50426,4.2592936,3.8858037,3.9801195,4.398881,4.7044635,4.1574326,4.0593443,4.38379,5.191132,6.368191,7.6207023,8.692128,8.812852,8.397863,7.798016,7.2962565,6.488915,5.832478,5.1458607,4.353609,3.4896781,2.9237845,3.1199608,3.9386206,5.311856,7.2094865,8.118689,8.299775,7.986647,7.5829763,7.643338,8.390318,9.635284,10.525623,10.536942,9.473062,7.254758,5.1156793,3.229367,1.8523588,1.327964,1.3355093,1.8146327,2.233394,2.305074,1.9542197,1.358145,1.1393328,1.1129243,1.0148361,0.47912338,0.35839936,0.38103512,0.49421388,0.73188925,1.2185578,1.8297231,2.6068838,3.3689542,4.08198,4.878004,3.591539,2.4031622,2.214531,3.006782,3.8556228,4.5761943,3.9763467,3.0218725,2.1994405,1.539231,2.003264,2.3126192,2.3126192,2.093807,1.9806281,1.8448136,1.9391292,2.1466236,2.384299,2.5917933,2.6898816,2.5767028,2.4220252,2.4220252,2.7841973,3.229367,3.6368105,3.6594462,3.4444065,3.6443558,4.5799665,5.458988,6.149379,6.537959,6.5002327,6.349328,5.9532022,5.270357,4.466788,3.8858037,3.6028569,3.7084904,3.9084394,4.0517993,4.164978,3.4368613,2.7691069,2.1768045,1.8372684,2.0900342,2.052308,1.690136,1.4109617,1.3128735,1.1959221,0.7997965,0.5017591,0.3055826,0.19994913,0.17731337,0.59607476,1.086516,1.3770081,1.3845534,1.2223305,0.8903395,0.6375736,0.58098423,0.76207024,1.1431054,1.4411428,1.4977322,1.2261031,0.7469798,0.3961256,0.19240387,0.10940613,0.071679875,0.041498873,0.056589376,0.452715,1.3770081,2.6597006,3.62172,3.078462,2.4823873,1.9240388,1.5656394,1.358145,1.026154,0.4640329,0.23013012,0.16976812,0.19240387,0.26408374,0.3169005,0.34330887,0.38858038,0.4376245,0.4074435,0.3055826,0.6413463,1.2638294,2.11267,3.2331395,3.470815,3.429316,3.229367,3.0218725,2.9803739,3.6594462,4.859141,5.0553174,3.942393,2.4220252,2.5125682,3.0407357,3.7688525,4.285702,4.014073,3.0558262,1.6939086,0.7054809,0.29049212,0.08299775,1.2411937,1.0412445,0.98842776,1.0601076,1.2336484,1.4939595,1.7995421,2.1541688,2.516341,2.9086938,3.3915899,3.663219,4.006528,4.4177437,4.7912335,4.9345937,5.383536,5.983383,6.579458,7.1793056,7.960239,8.526133,8.880759,9.1825695,9.616421,10.378491,11.351829,11.846043,12.00072,11.974312,11.962994,12.445889,12.815607,13.053283,13.358865,14.143571,15.841252,17.040947,17.765291,17.987877,17.60684,17.765291,18.150099,18.153872,17.731337,17.40312,17.05981,17.248442,17.674747,18.1086,18.387774,18.757492,18.923487,19.191343,19.564833,19.779873,19.74592,19.87419,20.02132,20.16468,20.4099,20.33822,20.447628,20.43631,20.040184,19.017803,18.946123,19.57615,20.572124,21.62846,22.443346,22.677248,22.884743,22.963968,23.092237,23.741129,23.918442,23.775084,23.258234,22.484844,21.73032,21.398329,22.107582,22.631977,22.035902,19.670467,19.67424,20.1345,20.096773,19.372429,18.53868,17.501207,15.497944,13.521088,12.117672,11.3971,11.514051,11.729091,11.955449,12.140307,12.272349,11.91395,11.310329,10.1294985,8.4544525,6.790725,5.523123,4.82896,4.3724723,4.0517993,4.002755,4.478106,5.05909,5.0666356,4.3309736,3.1916409,2.233394,1.3958713,0.7432071,0.35462674,0.32821837,0.32821837,0.30935526,0.25276586,0.20749438,0.3169005,0.51684964,0.7205714,0.8224323,0.8111144,0.754525,0.87147635,0.7809334,0.513077,0.36971724,0.9393836,1.267602,1.0978339,0.8639311,0.7582976,0.7130261,0.59230214,0.41498876,0.25276586,0.24899325,0.6149379,0.59230214,0.41498876,0.28294688,0.2565385,0.24899325,0.30935526,0.30935526,0.26408374,0.18485862,0.08677038,0.090543,0.1358145,0.24522063,0.362172,0.35462674,0.2678564,0.16222288,0.094315626,0.090543,0.1358145,0.30935526,0.43007925,0.4979865,0.4979865,0.38858038,0.28294688,0.20749438,0.14335975,0.0754525,0.030181,0.056589376,0.13204187,0.23390275,0.3055826,0.23013012,0.29426476,0.47912338,0.47912338,0.28294688,0.16222288,0.271629,0.23390275,0.15467763,0.09808825,0.06413463,0.056589376,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.018863125,0.03772625,0.049044125,0.041498873,0.030181,0.02263575,0.0150905,0.00754525,0.0,0.003772625,0.003772625,0.0,0.0,0.003772625,0.00754525,0.011317875,0.018863125,0.00754525,0.00754525,0.011317875,0.011317875,0.011317875,0.011317875,0.033953626,0.06413463,0.094315626,0.11317875,0.094315626,0.08299775,0.08299775,0.0754525,0.056589376,0.033953626,0.07922512,0.1056335,0.120724,0.12826926,0.124496624,0.124496624,0.08677038,0.05281675,0.033953626,0.02263575,0.011317875,0.003772625,0.0,0.00754525,0.03772625,0.00754525,0.0,0.003772625,0.00754525,0.0,0.0,0.003772625,0.030181,0.0754525,0.120724,0.12826926,0.15467763,0.20372175,0.23767537,0.1961765,0.17354076,0.19994913,0.23767537,0.26408374,0.271629,0.17731337,0.13958712,0.16222288,0.241448,0.35839936,0.41876137,0.47912338,0.56212115,0.6375736,0.63002837,0.62248313,0.77338815,1.1695137,1.8900851,2.987919,4.617693,5.7117543,6.5002327,7.3377557,8.703445,10.340765,10.86516,9.861642,7.647111,5.27413,5.5570765,5.0138187,4.214022,4.0404816,5.7004366,5.3194013,4.1498876,3.7009451,4.036709,3.7688525,2.686109,1.8297231,1.5128226,2.033445,3.6707642,4.1083884,3.2218218,3.0935526,3.8292143,3.561358,3.218049,4.06689,4.557331,4.063117,2.8898308,2.6031113,2.2183034,2.0636258,2.1088974,1.9542197,2.1579416,2.2371666,2.2107582,2.142851,2.1164427,2.6483827,3.3123648,3.682082,3.6179473,3.259548,2.7087448,2.2484846,2.123988,2.3390274,2.6672459,2.565385,2.4559789,2.535204,2.927557,3.6858547,4.908185,5.5306683,5.5268955,5.2137675,5.2364035,5.66271,7.1000805,9.854096,13.287186,15.833707,16.222288,15.943113,15.064092,14.547242,16.229834,15.143317,13.008011,11.053791,9.740918,8.744945,8.511042,8.443134,8.812852,9.420244,9.601331,8.050782,6.5530496,5.617439,5.2590394,4.961002,4.217795,3.92353,3.9725742,4.2592936,4.689373,5.462761,6.3417826,7.0812173,7.4735703,7.33021,7.8319697,8.616675,8.699674,7.779153,6.2436943,5.3269467,5.243949,5.594803,5.764571,4.889322,4.3800178,4.2102494,4.5912848,5.5985756,7.1981683,8.8618965,9.544742,9.442881,8.83926,8.096053,7.2585306,6.2927384,5.2326307,4.22534,3.5160866,3.150142,3.4745877,4.3422914,5.692891,7.5301595,8.616675,8.846806,8.390318,7.7716074,7.8508325,8.054554,8.5563135,8.797762,8.484633,7.5565677,5.7494807,4.236658,3.0746894,2.4069347,2.463524,2.1390784,1.9504471,1.9693103,2.2409391,2.7879698,3.1199608,2.9313297,2.5087957,1.8674494,0.76584285,0.55457586,0.5470306,0.5696664,0.62625575,0.91297525,1.7278622,2.9200118,4.093298,4.938366,5.247721,3.7499893,2.746471,2.6446102,3.2859564,3.9348478,4.08198,3.3689542,2.8219235,2.7917426,2.9351022,3.218049,3.1765501,2.8709676,2.4861598,2.3390274,2.2183034,2.1768045,2.1692593,2.214531,2.384299,2.5993385,2.6785638,2.6672459,2.6332922,2.6483827,2.7426984,2.927557,3.0897799,3.3123648,3.893349,4.610148,4.9987283,5.0854983,4.9345937,4.644101,4.5950575,4.496969,4.22534,3.7537618,3.1463692,2.7087448,2.7502437,2.8709676,2.8407867,2.6219745,1.9391292,1.3204187,0.72811663,0.392353,0.8337501,1.0110635,0.95447415,0.87902164,0.84129536,0.7432071,0.46026024,0.30181,0.21881226,0.181086,0.16976812,0.362172,0.6073926,0.8903395,1.1091517,1.0940613,0.8224323,0.47912338,0.241448,0.17731337,0.26408374,0.49044126,0.7092535,0.8978847,0.9695646,0.80734175,0.5281675,0.27917424,0.1056335,0.033953626,0.056589376,0.44139713,1.4826416,3.0445085,4.38379,4.142342,3.3689542,2.2748928,1.448688,1.0374719,0.7432071,0.40367088,0.24899325,0.21881226,0.32067314,0.62248313,0.6488915,0.543258,0.44894236,0.40367088,0.32821837,0.30181,0.8262049,1.6146835,2.5314314,3.6179473,3.218049,2.776652,2.444661,2.4672968,3.1463692,4.255521,5.1232247,5.1873593,4.346064,2.9464202,2.8936033,3.1048703,3.5349495,3.9876647,4.123479,3.742444,2.6144292,1.6750455,1.2525115,1.1016065,1.0299267,0.76207024,0.73188925,0.88279426,1.1431054,1.4335974,1.6825907,1.8523588,2.1541688,2.7087448,3.5839937,3.9989824,4.22534,4.6214657,5.2062225,5.66271,6.085244,6.571913,7.303802,8.265821,9.231613,9.574923,9.752235,9.81637,9.914458,10.306811,11.514051,12.0082655,12.061082,11.744182,10.944386,11.140562,11.3971,11.295239,11.057564,11.544232,12.347801,13.272095,14.200161,14.969776,15.358356,15.739391,15.841252,15.535669,15.01882,14.807553,14.800008,14.754736,14.84528,15.113135,15.482853,16.475054,17.135263,17.591751,17.999193,18.572634,19.074392,19.413929,19.515789,19.515789,19.753464,20.330677,21.304014,22.069857,22.043447,20.65135,20.63626,20.813572,21.058792,21.164427,20.858843,20.251451,20.285404,20.496672,20.598532,20.485353,20.677757,20.749437,20.545715,19.953413,18.900852,17.946377,17.701157,17.327667,16.52787,15.543215,14.852824,14.441608,14.25675,14.109617,13.702174,13.034419,12.336484,11.61214,10.940613,10.457717,10.510533,10.910432,11.438599,11.864905,11.944131,11.208468,9.918231,8.213005,6.4926877,5.4174895,5.062863,5.3269467,5.613666,5.6287565,5.353355,5.7570257,5.926794,5.8588867,5.323174,3.8254418,1.9655377,1.026154,0.573439,0.38103512,0.41876137,0.4678055,0.44894236,0.3734899,0.35839936,0.6149379,0.9318384,1.2034674,1.2789198,1.1657411,1.0412445,1.1883769,0.95824677,0.5319401,0.20749438,0.41876137,0.5583485,0.5772116,0.4640329,0.29426476,0.211267,0.23013012,0.22258487,0.26031113,0.44139713,0.90543,0.875249,0.7167987,0.58098423,0.4979865,0.3961256,0.30181,0.26408374,0.23390275,0.19240387,0.15467763,0.17354076,0.21881226,0.29049212,0.34330887,0.3055826,0.2263575,0.150905,0.124496624,0.16222288,0.23013012,0.29049212,0.32821837,0.34330887,0.331991,0.26408374,0.181086,0.090543,0.03772625,0.030181,0.033953626,0.018863125,0.02263575,0.041498873,0.094315626,0.211267,0.241448,0.25276586,0.24522063,0.20749438,0.12826926,0.16976812,0.10186087,0.049044125,0.03772625,0.0,0.030181,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.026408374,0.033953626,0.02263575,0.018863125,0.0150905,0.011317875,0.003772625,0.00754525,0.00754525,0.0,0.003772625,0.011317875,0.0150905,0.018863125,0.02263575,0.011317875,0.0150905,0.02263575,0.026408374,0.026408374,0.041498873,0.08299775,0.1056335,0.124496624,0.13958712,0.150905,0.17354076,0.150905,0.116951376,0.0754525,0.02263575,0.07922512,0.124496624,0.15845025,0.19994913,0.26031113,0.2867195,0.23767537,0.17354076,0.12826926,0.08677038,0.041498873,0.0150905,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.02263575,0.05281675,0.11317875,0.1358145,0.150905,0.18485862,0.23013012,0.24899325,0.181086,0.16222288,0.17731337,0.21881226,0.29426476,0.23390275,0.16222288,0.13958712,0.16222288,0.17354076,0.24522063,0.30935526,0.36594462,0.41498876,0.44894236,0.5055317,0.56589377,0.7130261,1.0978339,1.9089483,2.1881225,2.1654868,2.3616633,3.0897799,4.4403796,7.2057137,8.541223,8.744945,7.8810134,5.80607,4.304565,3.3010468,2.6106565,2.2711203,2.516341,3.0633714,3.8895764,4.568649,4.851596,4.67051,3.802806,2.4861598,1.5354583,1.5316857,2.8445592,5.3458095,4.515832,2.969056,1.9957186,1.5580941,1.5467763,1.6675003,1.9730829,2.4371157,2.9615107,2.6710186,1.8900851,1.327964,1.3091009,1.7844516,2.8558772,3.399135,3.3651814,2.9086938,2.3956168,2.7238352,3.6179473,4.183841,4.1800685,4.006528,3.4557245,3.0633714,2.8822856,3.0369632,3.6971724,3.8820312,3.663219,3.5575855,3.8669407,4.6554193,6.0701537,6.579458,6.488915,6.19465,6.1720147,6.488915,7.8319697,11.159425,15.482853,17.84829,18.444365,18.889534,18.915941,18.485863,17.810562,13.7700815,10.461489,8.379,7.394345,6.719045,6.4549613,6.4436436,7.3679366,9.178797,11.102836,9.639057,8.27714,7.0963078,6.247467,5.9607477,5.383536,4.8025517,4.5460134,4.719554,5.1873593,6.0362,6.9680386,7.5829763,7.6508837,7.1038527,8.152642,9.699419,10.529396,10.159679,8.873214,7.435844,6.952948,6.8699503,6.7152724,6.096562,5.451443,4.919503,4.5724216,4.7535076,6.0550632,7.54525,8.620448,8.75249,7.8696957,6.3719635,5.485397,4.7950063,4.255521,3.893349,3.8103511,4.0178456,4.4516973,5.1232247,5.9607477,6.828451,7.4094353,6.937857,5.983383,5.1835866,5.251494,5.1534057,5.0477724,5.010046,4.8742313,4.244203,3.2935016,2.6182017,2.354118,2.5578396,3.218049,2.8030603,2.4069347,2.372981,2.9539654,4.274384,5.6098933,5.142088,3.9197574,2.5578396,1.2525115,1.1544232,1.267602,1.267602,1.0110635,0.52062225,0.87147635,1.8599042,3.0746894,4.1008434,4.504514,3.6858547,3.2520027,3.1954134,3.3878171,3.5651307,3.2784111,2.8785129,3.0897799,3.9989824,5.0477724,5.323174,5.172269,4.768598,4.3611546,4.244203,4.074435,3.7575345,3.3538637,2.9766011,2.7841973,2.8332415,3.1840954,3.4594972,3.4330888,3.0407357,2.8143783,2.625747,2.5578396,2.7351532,3.350091,3.9914372,4.1272516,3.731126,2.9237845,1.9579924,1.7316349,1.8334957,2.1956677,2.5125682,2.2258487,1.8070874,1.4713237,1.2562841,1.1016065,0.84884065,0.59607476,0.51684964,0.5357128,0.62248313,0.77716076,0.7054809,0.52439487,0.39989826,0.38858038,0.41876137,0.4074435,0.392353,0.362172,0.3169005,0.27540162,0.33953625,0.41498876,0.55457586,0.694163,0.6752999,0.46026024,0.3055826,0.211267,0.181086,0.22258487,0.41498876,0.7696155,1.2713746,1.6788181,1.4826416,0.9922004,0.49044126,0.14335975,0.00754525,0.00754525,0.1358145,0.694163,1.5543215,2.4031622,2.7502437,2.263575,1.3015556,0.5394854,0.22258487,0.15467763,0.23390275,0.29803738,0.41121614,0.66775465,1.2110126,1.2223305,0.9205205,0.6149379,0.44139713,0.331991,0.5319401,0.95447415,1.4411428,1.9278114,2.4220252,1.9164935,1.4939595,1.2525115,1.4675511,2.584248,4.3121104,5.0968165,5.3344917,5.05909,3.9197574,2.5427492,2.0749438,2.2447119,2.757789,3.2935016,3.6141748,3.059599,2.4974778,2.3088465,2.3918443,0.8865669,0.8978847,1.1016065,1.4675511,1.8749946,2.1051247,2.4107075,2.3126192,2.3692086,2.837014,3.6934,4.0216184,4.52715,5.4703064,6.6247296,7.2472124,7.515069,7.0359454,6.862405,7.3151197,7.9489207,9.024119,9.914458,10.763299,11.257513,10.63503,10.182315,10.26154,10.593531,10.895341,10.895341,10.650121,10.38981,10.125726,10.069136,10.604849,11.106608,11.514051,12.253486,13.219278,13.792717,13.902123,13.856852,13.570132,13.109872,12.694883,12.804289,12.951422,13.200415,13.483362,13.58145,13.155144,13.147598,13.4644985,13.985121,14.558559,15.803526,16.663685,17.120173,17.45971,18.263277,18.802763,19.055529,19.127209,19.078165,18.904623,19.319613,19.08571,18.346275,17.354074,16.463736,15.62244,14.8339615,14.158662,13.7700815,13.977575,15.735619,17.127718,18.184053,18.780127,18.648085,18.463226,18.30855,17.557796,16.22606,14.969776,14.102073,13.290957,12.551523,11.9064045,11.3820095,10.725573,10.174769,10.231359,10.702937,10.725573,10.359629,10.435081,10.506761,10.321902,9.797507,9.929549,9.442881,8.043237,6.296511,5.5985756,5.587258,5.9494295,6.470052,7.1340337,8.14887,8.661947,7.7640624,5.6098933,3.059599,1.6788181,0.87147635,0.633801,0.55080324,0.45648763,0.44139713,0.6375736,0.6488915,0.5696664,0.55457586,0.8224323,0.935611,0.9695646,0.935611,0.87147635,0.87147635,1.0148361,0.7582976,0.422534,0.211267,0.19994913,0.41876137,0.5998474,0.5357128,0.271629,0.1358145,0.1358145,0.33953625,0.5696664,0.7469798,0.87147635,0.90543,0.90543,0.8563859,0.7507524,0.58098423,0.3961256,0.241448,0.1358145,0.094315626,0.1056335,0.15467763,0.18485862,0.21503963,0.23013012,0.18485862,0.1358145,0.094315626,0.094315626,0.13204187,0.1659955,0.19240387,0.18863125,0.16976812,0.17731337,0.27540162,0.26408374,0.1659955,0.094315626,0.071679875,0.0452715,0.02263575,0.0150905,0.02263575,0.05281675,0.1358145,0.1358145,0.10186087,0.056589376,0.030181,0.030181,0.090543,0.05281675,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.03772625,0.02263575,0.011317875,0.0,0.011317875,0.00754525,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.0150905,0.011317875,0.0,0.011317875,0.0150905,0.00754525,0.018863125,0.090543,0.13958712,0.150905,0.14713238,0.12826926,0.090543,0.13958712,0.1358145,0.1056335,0.071679875,0.060362,0.08677038,0.10186087,0.1358145,0.211267,0.32067314,0.4074435,0.39989826,0.362172,0.3055826,0.18485862,0.10940613,0.0452715,0.0150905,0.0150905,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.003772625,0.0150905,0.041498873,0.120724,0.211267,0.29803738,0.3961256,0.3470815,0.29049212,0.23390275,0.22258487,0.32067314,0.34330887,0.3055826,0.26408374,0.23390275,0.19994913,0.26031113,0.32067314,0.36971724,0.38858038,0.35085413,0.35085413,0.35085413,0.33953625,0.3470815,0.45648763,0.9205205,1.0827434,1.1431054,1.4260522,2.3654358,4.123479,5.926794,7.2094865,7.6622014,7.2472124,4.9534564,3.361409,2.293756,1.8599042,2.4559789,2.9803739,3.3425457,3.8292143,4.5007415,5.172269,5.66271,4.719554,3.3764994,2.1843498,1.2223305,1.5128226,1.7882242,2.1654868,2.5616124,2.6710186,2.3163917,2.082489,2.5804756,3.9348478,5.7683434,4.557331,3.361409,2.3277097,1.7844516,2.2107582,3.0181,3.832987,4.0517993,3.6292653,3.0671442,2.8596497,3.3123648,4.191386,5.119452,5.5683947,5.0213637,4.2517486,3.6971724,3.5387223,3.7084904,4.3422914,4.6742826,4.938366,5.3269467,5.9984736,7.364164,8.401636,8.394091,7.488661,6.6850915,6.3644185,6.7454534,8.009283,10.087999,12.649611,15.286676,18.270823,19.908142,19.28566,16.29774,12.608112,9.261794,6.9189944,5.7079816,5.2175403,5.3646727,5.383536,5.311856,5.670255,7.4773426,7.7225633,7.6810646,7.5603404,7.326438,6.730363,6.092789,5.541986,5.168496,5.2137675,6.043745,7.0057645,7.4773426,7.435844,7.1302614,7.0812173,7.9715567,9.688101,11.091517,11.389555,10.133271,8.948667,7.91874,7.91874,8.624221,8.514814,7.145352,6.0739264,5.3948536,5.2854476,5.9796104,7.2887115,7.8998766,7.2585306,5.6287565,4.0895257,3.270866,3.2520027,3.6707642,4.2894745,4.957229,5.692891,6.0022464,6.1078796,6.1418333,6.1795597,5.666483,5.3194013,4.9157305,4.3611546,3.6783094,3.2859564,3.180323,3.180323,3.1840954,3.1576872,3.1463692,2.886058,2.4107075,1.9240388,1.8146327,1.9391292,2.5087957,3.519859,4.825187,6.119198,6.398372,5.828706,4.7610526,3.5123138,2.3654358,2.4974778,3.3274553,3.682082,2.9501927,1.0827434,0.8262049,1.3128735,2.191895,3.0030096,3.1727777,2.795515,2.354118,1.9730829,1.7354075,1.6486372,1.7354075,2.0862615,2.7011995,3.6443558,5.036454,5.87775,5.8966126,5.6023483,5.4778514,5.96452,6.6247296,6.6247296,6.25124,5.5797124,4.45547,3.9197574,4.3875628,4.8327327,4.847823,4.6554193,5.13077,4.957229,4.432834,3.874486,3.6330378,3.9122121,4.3686996,4.3422914,3.640583,2.516341,1.8825399,1.961765,2.4333432,2.9237845,3.0218725,2.8143783,2.3956168,1.8825399,1.4222796,1.1883769,1.2034674,1.297783,1.3958713,1.4260522,1.327964,1.0110635,0.7394345,0.52062225,0.36971724,0.32067314,0.41876137,0.41498876,0.38480774,0.3734899,0.3961256,0.47157812,0.543258,0.62248313,0.69793564,0.7469798,0.79602385,0.7809334,0.6526641,0.41876137,0.1358145,0.36971724,0.7394345,1.0450171,1.116697,0.8224323,0.422534,0.211267,0.094315626,0.033953626,0.0452715,0.094315626,0.14335975,0.14335975,0.10186087,0.0754525,0.090543,0.1358145,0.16222288,0.14335975,0.1056335,0.1056335,0.18863125,0.45648763,0.91674787,1.478869,1.6373192,1.3845534,1.0940613,0.87147635,0.56589377,0.5885295,0.9808825,1.5656394,2.1805773,2.655928,2.372981,2.2862108,2.052308,1.901403,2.6106565,3.731126,4.4441524,5.149633,5.50426,4.395108,2.746471,2.04099,1.6675003,1.3505998,1.1431054,1.4260522,1.659955,1.6863633,1.5241405,1.4034165,1.237421,1.086516,1.116697,1.2449663,1.3958713,1.5203679,1.8636768,2.2069857,2.5276587,2.8634224,3.338773,3.7348988,4.293247,4.7912335,5.040227,4.8930945,5.2967653,5.6325293,6.1720147,7.01331,8.107371,9.250477,9.171251,8.816625,8.597813,8.36391,8.722309,9.035437,9.231613,9.465516,10.087999,10.536942,10.412445,10.110635,9.895596,9.895596,9.978593,10.589758,11.849815,13.189097,13.355092,12.996693,12.736382,13.0646,13.920986,14.698147,14.211478,13.951167,13.81158,13.622949,13.166461,12.717519,12.325166,12.00072,11.827179,11.981857,12.630749,13.245687,14.003984,15.052773,16.531643,17.421982,18.229324,18.323639,17.72002,17.097536,16.588232,16.143063,15.452672,14.305794,12.596795,12.181807,12.162943,12.449662,12.90615,13.317367,14.060574,14.385019,14.70192,15.128226,15.471535,14.252977,13.226823,12.336484,11.498961,10.56335,9.725827,9.359882,9.216523,9.159933,9.175024,9.608876,9.793735,9.737145,9.454198,8.98262,8.733627,8.937348,9.273112,9.533423,9.612649,9.484379,9.009028,8.182823,7.466025,7.798016,8.624221,9.725827,10.253995,9.895596,8.869441,6.0814714,4.3875628,3.1350515,2.0372176,1.1657411,0.7205714,0.55080324,0.47912338,0.452715,0.5281675,0.73188925,0.784706,0.80734175,0.9242931,1.2525115,1.3920987,1.3770081,1.056335,0.6111652,0.55080324,0.845068,0.65643674,0.41121614,0.35085413,0.5017591,0.38103512,0.30935526,0.3169005,0.41121614,0.5885295,0.7922512,1.0676528,1.2487389,1.2789198,1.237421,1.5165952,1.5467763,1.3317367,0.9695646,0.6526641,0.38103512,0.21881226,0.12826926,0.090543,0.094315626,0.181086,0.24522063,0.2867195,0.27917424,0.18485862,0.11317875,0.07922512,0.071679875,0.090543,0.120724,0.13204187,0.12826926,0.124496624,0.17354076,0.35839936,0.32821837,0.17731337,0.0754525,0.056589376,0.033953626,0.00754525,0.003772625,0.018863125,0.08299775,0.24899325,0.24899325,0.24899325,0.15467763,0.018863125,0.018863125,0.02263575,0.033953626,0.02263575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.011317875,0.00754525,0.003772625,0.003772625,0.0,0.003772625,0.0,0.0,0.0,0.003772625,0.003772625,0.003772625,0.003772625,0.011317875,0.03772625,0.060362,0.071679875,0.06413463,0.049044125,0.041498873,0.06413463,0.124496624,0.17731337,0.18485862,0.12826926,0.116951376,0.11317875,0.09808825,0.071679875,0.049044125,0.0452715,0.06790725,0.08677038,0.10186087,0.11317875,0.16976812,0.19994913,0.18863125,0.14335975,0.09808825,0.071679875,0.049044125,0.030181,0.018863125,0.026408374,0.018863125,0.0150905,0.00754525,0.0,0.0,0.003772625,0.0,0.003772625,0.0150905,0.026408374,0.041498873,0.1056335,0.19240387,0.2678564,0.2867195,0.2565385,0.211267,0.18485862,0.1961765,0.23390275,0.211267,0.20372175,0.20749438,0.21881226,0.211267,0.20372175,0.20372175,0.241448,0.3055826,0.33953625,0.3470815,0.29049212,0.23013012,0.21881226,0.29803738,0.5772116,0.8111144,0.9280658,0.9808825,1.1204696,1.5505489,3.7386713,6.1041074,7.598067,7.699928,5.511805,3.8178966,2.535204,1.7693611,1.81086,2.4408884,3.2520027,4.0782075,4.8930945,5.80607,6.089017,5.149633,3.6556737,2.2447119,1.5241405,1.2034674,1.0035182,1.5165952,2.7502437,4.0970707,3.6971724,3.1425967,2.7200627,2.637065,3.0218725,2.8106055,2.8407867,2.686109,2.3201644,2.1013522,2.4974778,3.0407357,3.440634,3.4934506,3.078462,2.655928,2.6446102,3.3123648,4.293247,4.568649,3.9612563,3.8443048,4.036709,4.353609,4.6214657,4.644101,4.8666863,5.4363527,6.2399216,6.900131,7.6622014,8.00551,8.013056,7.8131065,7.5603404,7.654656,7.9526935,8.669493,9.81637,11.208468,13.053283,16.177015,18.821627,20.025093,19.651604,14.803781,10.272858,7.2887115,6.039973,5.6589375,5.745708,5.66271,5.515578,5.4401255,5.5985756,5.6476197,5.7909794,5.9192486,5.9117036,5.6551647,5.4778514,5.194905,5.281675,5.828706,6.541732,6.9491754,7.2962565,7.6093845,8.050782,8.91094,10.31813,11.936585,12.577931,11.932813,10.559577,9.024119,8.258276,8.160188,8.431817,8.575176,7.7640624,6.5228686,5.323174,4.6516466,5.0062733,6.1644692,6.7454534,6.7869525,6.319147,5.3571277,4.647874,4.1197066,4.08198,4.4403796,4.7044635,4.22534,4.3121104,4.534695,4.5799665,4.274384,4.06689,4.006528,4.06689,4.1989317,4.323428,4.3422914,4.2291126,4.0103,3.7462165,3.5236318,3.1425967,2.6785638,2.263575,1.9994912,1.9994912,2.335255,3.4783602,4.908185,6.2135134,7.1076255,6.432326,5.4891696,4.768598,4.315883,3.7462165,4.2291126,4.5912848,3.9989824,2.5276587,1.1581959,1.3505998,1.9994912,2.686109,3.1010978,3.0256453,2.727608,2.3277097,1.9429018,1.6448646,1.4411428,1.3128735,1.5731846,1.9730829,2.3654358,2.704972,3.029418,3.2331395,3.3048196,3.4330888,4.002755,4.8742313,5.27413,5.836251,6.643593,7.201941,6.673774,6.4511886,6.4134626,6.360646,6.009792,5.2364035,4.647874,4.402653,4.5120597,4.8025517,4.851596,4.6516466,3.9876647,2.9426475,1.9089483,1.448688,1.4335974,1.8448136,2.4597516,2.8521044,2.6219745,2.1994405,1.7467253,1.4034165,1.3015556,1.3619176,1.6071383,1.7580433,1.6675003,1.3166461,0.98842776,0.67152727,0.43007925,0.3055826,0.29426476,0.5017591,0.5093044,0.392353,0.23767537,0.1659955,0.23013012,0.38858038,0.543258,0.62248313,0.56589377,0.38858038,0.24522063,0.14713238,0.08299775,0.026408374,0.13204187,0.32444575,0.422534,0.35839936,0.1659955,0.08299775,0.041498873,0.02263575,0.033953626,0.094315626,0.124496624,0.116951376,0.11317875,0.1659955,0.34330887,0.69039035,0.8563859,0.7469798,0.43007925,0.1659955,0.090543,0.07922512,0.150905,0.30181,0.49044126,0.62248313,0.63002837,0.6111652,0.55080324,0.331991,0.27917424,0.3734899,0.56212115,0.8337501,1.2034674,1.7731338,1.8297231,1.4939595,1.1242423,1.3015556,2.2409391,2.8106055,3.097325,3.187868,3.1614597,3.1652324,2.5502944,1.6448646,0.8337501,0.5470306,0.7394345,0.98842776,1.1695137,1.2185578,1.1355602,1.1883769,1.1204696,1.0902886,1.2298758,1.539231,1.8863125,2.4672968,2.6483827,2.5578396,2.4069347,2.5012503,2.8106055,3.259548,4.376245,5.885295,6.692637,6.8246784,6.7944975,6.7567716,6.85486,7.2057137,7.647111,7.5226145,7.5716586,7.9036493,7.9791017,8.050782,8.171506,8.284684,8.492179,9.0543,9.397609,9.435335,9.405154,9.469289,9.703192,10.042727,10.314357,10.982111,12.00072,12.823153,12.30253,12.166716,13.087236,14.592513,15.098045,14.366156,13.607859,13.419228,13.958713,14.966003,14.916959,14.173752,12.6345215,10.891568,10.238904,10.197406,10.676529,11.314102,11.970539,12.736382,14.18507,15.094273,15.169725,14.592513,14.056801,13.547497,13.20796,12.853333,12.351574,11.6008215,11.5857315,11.661184,11.830952,12.08749,12.411936,12.649611,12.664702,12.50248,12.215759,11.823407,10.303039,9.378746,8.827943,8.390318,7.748972,7.364164,7.3490734,7.5792036,7.9489207,8.36391,9.073163,9.733373,10.208723,10.450171,10.495442,10.533169,10.702937,11.099063,11.487643,11.314102,10.329447,9.929549,9.676784,9.465516,9.544742,10.182315,10.638803,10.020092,8.345046,6.5568223,4.1083884,2.7728794,1.9881734,1.4298248,0.9922004,1.0638802,1.146878,1.1204696,1.0148361,1.0148361,1.1280149,1.3920987,1.6788181,1.961765,2.3088465,2.0108092,1.7429527,1.4675511,1.2147852,1.1129243,1.1431054,0.9507015,0.7582976,0.6828451,0.7167987,0.5772116,0.52439487,0.59607476,0.9242931,1.7467253,2.1202152,1.8825399,1.6335466,1.5807298,1.5467763,1.448688,1.2638294,0.98465514,0.6790725,0.47912338,0.30181,0.17354076,0.094315626,0.06413463,0.056589376,0.13204187,0.18863125,0.2263575,0.21503963,0.120724,0.06790725,0.049044125,0.05281675,0.071679875,0.09808825,0.10940613,0.1358145,0.15845025,0.17731337,0.21503963,0.181086,0.10186087,0.06413463,0.06413463,0.049044125,0.011317875,0.003772625,0.030181,0.10186087,0.2565385,0.211267,0.16222288,0.090543,0.026408374,0.033953626,0.041498873,0.030181,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.018863125,0.011317875,0.00754525,0.00754525,0.033953626,0.1358145,0.24899325,0.22258487,0.150905,0.09808825,0.06790725,0.056589376,0.090543,0.1358145,0.16976812,0.17354076,0.1659955,0.124496624,0.094315626,0.08299775,0.08299775,0.049044125,0.041498873,0.056589376,0.0754525,0.041498873,0.06413463,0.07922512,0.08299775,0.0754525,0.06790725,0.049044125,0.03772625,0.026408374,0.0150905,0.02263575,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.02263575,0.049044125,0.08299775,0.11317875,0.11317875,0.116951376,0.124496624,0.150905,0.19240387,0.22258487,0.19994913,0.181086,0.16976812,0.1659955,0.15845025,0.16222288,0.14335975,0.13958712,0.15845025,0.16976812,0.18485862,0.1659955,0.16222288,0.17731337,0.21503963,0.33576363,0.754525,1.146878,1.3317367,1.2864652,1.0751982,1.8787673,3.0860074,4.183841,4.7346444,4.217795,3.2444575,2.655928,2.8634224,3.863168,2.9916916,2.6332922,2.7313805,3.240685,4.0970707,4.425289,3.783943,3.1916409,3.150142,3.6254926,2.9011486,2.1503963,1.6863633,1.7769064,2.6144292,2.9539654,3.5538127,3.8103511,3.6481283,3.4896781,3.289729,3.7952607,4.5761943,5.036454,4.4101987,4.2328854,4.3385186,4.3686996,4.13857,3.6594462,3.4745877,3.2670932,3.2784111,3.5236318,3.7688525,5.2854476,7.835742,7.9036493,5.43258,3.8254418,3.832987,4.3083377,5.05909,5.8136153,6.2361493,7.1906233,8.084735,8.473316,8.431817,8.567632,9.175024,10.386037,11.672502,12.649611,13.083464,14.252977,16.399601,18.859352,20.839981,21.398329,18.859352,14.720782,11.170743,9.22784,8.733627,8.60913,8.424272,8.311093,8.246958,8.0206,7.7640624,7.2170315,6.5568223,5.8966126,5.2854476,5.3873086,5.4288073,5.6551647,6.0211096,6.1908774,6.1078796,6.2927384,6.8473144,7.816879,9.159933,10.578441,11.581959,11.710228,11.057564,10.291721,9.4127,8.831716,8.827943,9.295748,9.718282,8.986393,7.786698,6.405917,5.2288585,4.7421894,5.0025005,5.534441,6.085244,6.360646,6.043745,4.817642,4.08198,3.874486,4.191386,4.9949555,4.7044635,4.3121104,4.195159,4.3422914,4.349837,4.353609,4.187614,4.1197066,4.3686996,5.100589,4.8930945,4.3083377,3.942393,3.9574835,4.08198,4.274384,4.3347464,4.3196554,4.2291126,4.002755,4.036709,4.5196047,5.406172,6.25124,6.2021956,4.9044123,3.9386206,3.5764484,3.8707132,4.666737,5.3873086,5.5080323,4.561104,2.916239,1.780679,1.5279131,2.093807,2.674791,2.8558772,2.6446102,2.4710693,2.11267,1.6033657,1.116697,0.9507015,0.8601585,0.935611,1.3241913,1.9806281,2.6597006,3.6028569,3.953711,3.651901,3.3123648,4.214022,5.0477724,5.6287565,5.9720654,6.115425,6.1418333,6.1720147,5.8928404,5.4401255,5.251494,6.0550632,5.9117036,5.304311,4.930821,4.9685473,5.0515447,4.7836885,4.402653,3.783943,2.9049213,1.8448136,1.4222796,1.3807807,1.6146835,1.9391292,2.1013522,1.7542707,1.3543724,1.0940613,1.177059,1.81086,1.7769064,1.5769572,1.4298248,1.3392819,1.0940613,0.87147635,0.70170826,0.5281675,0.32821837,0.116951376,0.20749438,0.32444575,0.31312788,0.181086,0.09808825,0.07922512,0.16222288,0.241448,0.26408374,0.20749438,0.150905,0.13958712,0.1961765,0.2678564,0.19994913,0.0754525,0.09808825,0.116951376,0.07922512,0.00754525,0.06790725,0.124496624,0.18485862,0.24899325,0.33576363,0.32444575,0.24522063,0.25276586,0.43007925,0.77716076,1.4411428,1.6976813,1.4901869,0.9620194,0.4376245,0.17354076,0.08299775,0.124496624,0.24899325,0.38103512,0.33576363,0.30935526,0.3055826,0.31312788,0.30181,0.30181,0.30181,0.32821837,0.41498876,0.58475685,1.0110635,1.3430545,1.6184561,1.9240388,2.41448,2.505023,1.9957186,1.659955,1.7542707,2.0296721,2.4522061,2.757789,2.8294687,2.4522061,1.3015556,0.83752275,0.7092535,0.72811663,0.754525,0.7092535,0.8978847,0.95824677,1.2185578,1.81086,2.5427492,2.867195,3.350091,3.4632697,3.0671442,2.3993895,2.052308,2.8143783,3.2935016,4.29702,5.8588867,7.224577,7.4094353,7.2358947,6.983129,6.7831798,6.6624556,6.5832305,6.485142,6.688864,7.1378064,7.4018903,7.3188925,7.3905725,7.5603404,7.809334,8.145098,8.273367,8.273367,8.273367,8.431817,8.907167,9.273112,9.224068,9.348565,9.989911,11.25374,11.838497,12.683565,14.04171,15.260268,14.784918,14.147344,13.419228,13.04951,13.347548,14.464244,14.762281,14.053028,12.494934,10.819888,10.329447,9.850324,9.737145,9.590013,9.397609,9.540969,10.95193,11.672502,11.834724,11.676274,11.548005,11.072655,10.736891,10.7557535,11.046246,11.234878,11.446144,11.778135,11.932813,11.823407,11.563096,11.393328,11.140562,10.638803,9.95973,9.405154,8.688355,8.75249,8.831716,8.492179,7.6207023,7.567886,7.7225633,8.107371,8.692128,9.378746,10.159679,11.050018,11.796998,12.279895,12.491161,12.898605,13.347548,14.045483,14.86037,15.350811,14.698147,13.721037,12.709973,11.766817,10.770844,10.280403,9.6201935,8.235641,6.307829,4.7648253,3.3651814,2.323937,1.6410918,1.2940104,1.2223305,1.9278114,2.305074,2.3314822,2.071171,1.6637276,1.5015048,1.7240896,2.04099,2.293756,2.4861598,1.9730829,1.6033657,1.3958713,1.297783,1.1883769,1.1619685,1.1959221,1.3204187,1.4939595,1.6260014,1.5467763,1.418507,1.2902378,1.3958713,2.123988,2.3654358,1.9429018,1.5203679,1.3392819,1.237421,0.97333723,0.7394345,0.5319401,0.36594462,0.28294688,0.19994913,0.120724,0.06413463,0.03772625,0.02263575,0.06413463,0.124496624,0.1659955,0.16222288,0.0754525,0.041498873,0.030181,0.0452715,0.0754525,0.1056335,0.13204187,0.150905,0.15845025,0.14335975,0.094315626,0.06790725,0.056589376,0.05281675,0.056589376,0.041498873,0.00754525,0.018863125,0.05281675,0.09808825,0.15845025,0.10940613,0.049044125,0.018863125,0.018863125,0.026408374,0.041498873,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.02263575,0.018863125,0.018863125,0.018863125,0.03772625,0.120724,0.22258487,0.1961765,0.14713238,0.116951376,0.090543,0.071679875,0.06413463,0.090543,0.14335975,0.19994913,0.2263575,0.1659955,0.10940613,0.090543,0.08677038,0.05281675,0.026408374,0.03772625,0.060362,0.030181,0.026408374,0.02263575,0.033953626,0.049044125,0.049044125,0.033953626,0.041498873,0.033953626,0.0150905,0.0150905,0.011317875,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.018863125,0.018863125,0.011317875,0.011317875,0.0150905,0.05281675,0.11317875,0.17731337,0.23390275,0.24899325,0.19994913,0.16976812,0.14713238,0.13958712,0.13958712,0.1358145,0.1056335,0.08299775,0.06790725,0.06790725,0.06790725,0.08677038,0.120724,0.15467763,0.16976812,0.31312788,0.84884065,1.5543215,2.0598533,1.8221779,1.1883769,1.0450171,1.3204187,1.8825399,2.5314314,3.31991,3.3312278,3.3878171,3.85185,4.61392,3.259548,2.5767028,2.4597516,2.7728794,3.3840446,3.0860074,2.5540671,2.5691576,3.3274553,4.4177437,4.187614,3.8254418,3.0181,1.9806281,1.4675511,2.3201644,3.6443558,4.7308717,5.172269,4.8365054,4.447925,4.772371,5.481624,5.994701,5.455216,5.111907,5.4778514,6.096562,6.1720147,4.5497856,3.8254418,3.4481792,3.0633714,2.7087448,2.7917426,4.957229,7.798016,8.028146,6.009792,5.7419353,5.9909286,5.5570765,5.4288073,5.8136153,6.1531515,7.33021,8.318638,8.741172,8.888305,9.703192,11.136789,13.215506,15.026365,15.916705,15.467763,14.234114,14.984866,16.920223,19.051756,20.202406,19.825144,17.45971,14.811326,13.075918,12.909923,13.441863,12.90615,12.162943,11.717773,11.69891,11.136789,10.03141,8.688355,7.492433,6.9265394,7.496206,7.8017883,7.877241,7.594294,6.6624556,6.0626082,5.956975,6.4926877,7.624475,9.110889,10.54826,10.699164,10.269085,9.827688,9.789962,9.703192,9.616421,10.0276375,10.789707,11.106608,10.412445,9.514561,8.318638,6.907676,5.5306683,4.459243,4.1612053,4.376245,4.949684,5.8211603,5.8513412,5.481624,5.1571784,5.20245,5.794752,5.881522,5.4476705,5.1232247,5.1571784,5.4174895,5.43258,4.8930945,4.406426,4.349837,4.8629136,4.7308717,4.13857,3.6594462,3.5802212,3.893349,4.534695,5.191132,5.873977,6.485142,6.809588,6.330465,5.7909794,5.4438977,5.1835866,4.5724216,3.4859054,2.916239,2.7917426,3.169005,4.2328854,5.270357,5.6061206,5.160951,4.1762958,3.2255943,2.4672968,2.3428001,2.4408884,2.505023,2.4182527,2.444661,2.203213,1.7354075,1.2298758,1.0412445,1.0638802,1.2185578,1.599593,2.142851,2.655928,3.2670932,3.6066296,3.500996,3.3689542,4.191386,4.5912848,4.927048,5.0025005,4.8063245,4.496969,4.6931453,4.564876,4.1498876,3.9159849,4.772371,4.90064,4.3611546,4.104616,4.3422914,4.557331,4.564876,4.395108,3.9914372,3.2859564,2.1692593,1.5958204,1.3317367,1.3166461,1.4335974,1.50905,1.3656902,0.95447415,0.6451189,0.72811663,1.4034165,1.3543724,1.0450171,0.8601585,0.8941121,0.98842776,1.1732863,1.0412445,0.77716076,0.482896,0.19994913,0.150905,0.20749438,0.21503963,0.150905,0.116951376,0.06790725,0.06413463,0.06790725,0.05281675,0.030181,0.09808825,0.16976812,0.25276586,0.32821837,0.36594462,0.30935526,0.17731337,0.0754525,0.0452715,0.06413463,0.16222288,0.32821837,0.573439,0.8111144,0.8526133,0.7167987,0.5055317,0.39989826,0.47535074,0.7167987,1.4675511,1.7731338,1.5882751,1.0601076,0.5055317,0.20749438,0.12826926,0.18863125,0.31312788,0.4376245,0.29803738,0.20372175,0.16222288,0.181086,0.26408374,0.35839936,0.46026024,0.5319401,0.5583485,0.5583485,0.573439,0.8111144,1.2298758,1.8070874,2.5502944,2.6672459,2.3578906,2.1277604,2.123988,2.1390784,2.123988,2.7238352,3.4934506,3.7952607,2.8030603,1.8070874,0.8941121,0.42630664,0.38103512,0.38858038,0.91674787,1.0751982,1.6976813,2.7011995,3.62172,3.6141748,3.7386713,4.044254,3.8367596,3.0746894,2.3692086,3.5538127,4.2517486,4.398881,4.3875628,5.036454,5.6061206,5.8437963,6.0286546,6.2436943,6.3644185,6.3153744,6.119198,5.9230213,5.9003854,6.247467,6.5002327,6.8058157,7.149124,7.4471617,7.537705,7.647111,7.6207023,7.413208,7.1906233,7.333983,7.4207535,7.4811153,7.7640624,8.390318,9.363655,11.246195,13.068373,14.532151,15.16218,14.313339,13.822898,13.460726,12.849561,12.106354,11.84227,12.098808,11.672502,11.1782875,11.012292,11.3669195,10.895341,10.216269,9.4013815,8.726082,8.643084,9.378746,9.944639,10.359629,10.653893,10.868933,10.167224,9.6201935,9.673011,10.223814,10.63503,10.948157,11.691365,12.027128,11.631002,10.676529,10.303039,9.771099,9.092027,8.526133,8.605357,9.020347,9.971047,10.487898,10.1294985,8.967529,8.873214,9.001483,9.371201,9.982366,10.804798,11.61214,12.427027,12.898605,12.951422,12.796744,13.445636,14.517061,15.912932,17.644567,19.821371,20.57967,19.029121,16.837225,14.777372,12.702429,10.585986,8.669493,6.9189944,5.4476705,4.5309224,3.5575855,2.4861598,1.7919968,1.6222287,1.81086,2.938875,3.4066803,3.429316,3.1199608,2.474842,2.1466236,2.1390784,2.2258487,2.2598023,2.1692593,1.750498,1.3732355,1.0676528,0.875249,0.8186596,1.0902886,1.5165952,1.9881734,2.41448,2.7200627,2.6446102,2.305074,1.8485862,1.4826416,1.4750963,1.3996439,1.2600567,1.0638802,0.8337501,0.5998474,0.46026024,0.36594462,0.2867195,0.21881226,0.16222288,0.1056335,0.06413463,0.03772625,0.02263575,0.02263575,0.0452715,0.094315626,0.13204187,0.13204187,0.071679875,0.03772625,0.033953626,0.05281675,0.09808825,0.15467763,0.2263575,0.18863125,0.12826926,0.090543,0.071679875,0.060362,0.056589376,0.0452715,0.02263575,0.011317875,0.003772625,0.033953626,0.06413463,0.071679875,0.033953626,0.018863125,0.00754525,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.02263575,0.02263575,0.0150905,0.00754525,0.02263575,0.056589376,0.08677038,0.094315626,0.071679875,0.06413463,0.05281675,0.0754525,0.1358145,0.19994913,0.26031113,0.20749438,0.12826926,0.0754525,0.056589376,0.060362,0.041498873,0.033953626,0.041498873,0.041498873,0.026408374,0.018863125,0.018863125,0.02263575,0.02263575,0.030181,0.060362,0.060362,0.030181,0.011317875,0.003772625,0.0,0.003772625,0.011317875,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.030181,0.02263575,0.011317875,0.00754525,0.02263575,0.08677038,0.15467763,0.21881226,0.26408374,0.241448,0.15467763,0.124496624,0.124496624,0.13958712,0.15845025,0.11317875,0.07922512,0.06413463,0.06790725,0.07922512,0.06790725,0.07922512,0.094315626,0.116951376,0.15467763,0.41121614,0.9016574,1.690136,2.335255,1.9051756,1.1091517,1.0186088,1.2525115,1.5958204,1.9881734,3.0558262,4.08198,4.6252384,4.515832,3.8971217,3.1539145,2.9954643,3.0935526,3.338773,3.8178966,2.8596497,2.1881225,2.0787163,2.5691576,3.4368613,4.38379,5.142088,5.05909,3.9801195,2.263575,2.6898816,3.6179473,4.8440504,5.824933,5.670255,5.572167,5.4476705,5.191132,4.8365054,4.5422406,4.3875628,5.3571277,6.9491754,7.673519,5.05909,3.610402,3.2972744,3.1199608,2.8558772,3.0671442,3.9386206,4.1536603,4.3422914,5.342037,8.201687,8.850578,7.462252,6.462507,6.6549106,7.220804,8.126234,8.314865,8.390318,8.933576,10.529396,12.619431,14.826416,16.546734,17.101309,15.724301,11.898859,11.514051,12.67602,14.237886,15.773345,16.614641,16.4826,15.690348,14.958458,15.437581,16.878725,16.124199,14.728328,13.849306,14.2077055,13.943622,12.932558,11.514051,10.336992,10.370946,11.3669195,11.774363,11.548005,10.578441,8.718536,7.9413757,7.8017883,8.284684,9.1976595,10.182315,11.080199,10.223814,9.190115,8.83926,9.34102,9.857869,10.314357,11.042474,11.868678,12.098808,11.627231,11.038701,10.095545,8.650629,6.651138,4.395108,2.897376,2.323937,2.969056,5.2665844,7.748972,8.2507305,7.884786,7.284939,6.609639,6.3455553,6.2135134,6.156924,6.25124,6.700182,6.549277,5.674028,4.708236,4.014073,3.6783094,3.9763467,4.0593443,3.7990334,3.4255435,3.531177,4.055572,4.8742313,5.975838,7.250985,8.499724,7.956466,7.032173,5.772116,4.508287,3.8480775,3.3425457,3.108643,2.886058,2.7200627,2.9464202,4.323428,5.194905,5.643847,5.560849,4.6252384,3.591539,2.6332922,2.2258487,2.4031622,2.7728794,3.029418,2.7691069,2.3088465,1.8674494,1.5618668,1.7127718,2.1881225,2.5125682,2.4559789,2.0296721,1.3996439,1.5769572,2.1805773,2.8521044,3.259548,3.1237335,2.9728284,3.0105548,3.199186,3.2444575,3.1237335,3.108643,3.0407357,2.867195,2.637065,2.282438,1.8749946,2.003264,2.6898816,3.410453,4.0895257,4.3422914,4.1612053,3.5575855,2.595566,1.8334957,1.2298758,0.95447415,1.0035182,1.2223305,1.4637785,1.1317875,0.6828451,0.38103512,0.33576363,0.362172,0.3772625,0.43007925,0.5998474,0.97333723,1.539231,1.3619176,0.97710985,0.6752999,0.513077,0.3961256,0.27917424,0.21881226,0.21503963,0.21503963,0.17731337,0.1358145,0.1056335,0.094315626,0.10186087,0.15845025,0.18485862,0.16976812,0.19240387,0.40367088,0.59230214,0.38858038,0.1659955,0.08299775,0.10940613,0.20749438,0.44516975,0.845068,1.237421,1.237421,1.0110635,0.724344,0.4640329,0.29803738,0.24899325,0.7922512,1.0789708,1.0336993,0.7205714,0.35085413,0.16976812,0.16976812,0.241448,0.3169005,0.392353,0.27540162,0.181086,0.120724,0.120724,0.18485862,0.33953625,0.58475685,0.7469798,0.7696155,0.70170826,0.52439487,0.5583485,0.7922512,1.2298758,1.9089483,2.8106055,3.5500402,3.682082,3.2482302,2.7728794,2.252257,2.3805263,2.9615107,3.5839937,3.6443558,2.6144292,1.1506506,0.27917424,0.19240387,0.2263575,2.1956677,2.4522061,2.7200627,2.927557,2.9803739,2.746471,2.9313297,3.361409,3.8103511,3.942393,3.2972744,3.0746894,3.953711,4.285702,3.6066296,2.655928,3.2029586,3.6443558,3.9197574,4.1574326,4.67051,4.9987283,5.0439997,5.142088,5.4288073,5.8437963,6.379509,6.9189944,7.4169807,7.6584287,7.232122,7.4282985,8.054554,7.9489207,6.9189944,5.723072,6.013564,6.8661776,8.152642,9.352338,9.522105,9.81637,10.336992,11.32542,12.664702,13.8870325,13.041965,12.400619,12.083718,12.0233555,11.962994,11.59705,11.065109,10.729345,10.646348,10.574668,10.612394,10.914205,11.363147,11.559323,10.804798,10.925522,11.872451,12.653384,12.894833,12.849561,11.970539,11.18206,10.435081,9.97482,10.329447,10.868933,11.321648,11.004747,10.020092,9.261794,9.529651,9.276885,8.7600355,8.337502,8.484633,8.397863,8.296002,8.307321,8.382772,8.284684,7.809334,7.7829256,8.050782,8.567632,9.4013815,9.876732,10.167224,10.125726,9.880505,9.842778,10.257768,11.872451,14.237886,17.123945,20.492899,21.700138,21.647322,20.975796,19.828917,17.852062,14.396337,10.853842,7.635793,5.2779026,4.4101987,3.4934506,2.7426984,2.3465726,2.335255,2.5804756,3.2972744,3.3425457,3.187868,3.218049,3.7084904,3.9650288,4.08198,4.0593443,3.904667,3.6481283,3.1237335,2.3880715,1.720317,1.3543724,1.4637785,2.0372176,2.595566,2.7087448,2.41448,2.1805773,1.9994912,1.6335466,1.237421,0.9242931,0.77716076,0.694163,0.6526641,0.7809334,0.95447415,0.80734175,0.4074435,0.24899325,0.18485862,0.124496624,0.0754525,0.041498873,0.011317875,0.0,0.011317875,0.060362,0.120724,0.090543,0.041498873,0.02263575,0.0452715,0.033953626,0.041498873,0.071679875,0.14335975,0.29049212,0.44894236,0.35839936,0.20749438,0.094315626,0.0452715,0.0452715,0.03772625,0.02263575,0.011317875,0.0,0.0,0.018863125,0.03772625,0.0452715,0.0452715,0.02263575,0.0150905,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.0150905,0.02263575,0.033953626,0.0452715,0.1056335,0.17731337,0.15845025,0.060362,0.0,0.011317875,0.033953626,0.071679875,0.12826926,0.21503963,0.21503963,0.1659955,0.094315626,0.030181,0.030181,0.1056335,0.1056335,0.08677038,0.0754525,0.0754525,0.06413463,0.02263575,0.0,0.0,0.0,0.02263575,0.06790725,0.09808825,0.08677038,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.041498873,0.0754525,0.05281675,0.026408374,0.0150905,0.02263575,0.060362,0.1358145,0.14335975,0.13204187,0.120724,0.1056335,0.056589376,0.0452715,0.0754525,0.120724,0.120724,0.09808825,0.08299775,0.0754525,0.07922512,0.090543,0.07922512,0.0754525,0.06413463,0.071679875,0.1659955,0.32821837,0.62248313,0.84884065,0.9280658,0.91674787,0.80734175,0.6488915,0.5998474,0.67152727,0.73188925,1.6109109,3.8556228,5.4288073,5.692891,5.3873086,3.8593953,2.5917933,1.6561824,1.388326,2.3654358,2.9011486,2.2220762,1.7316349,2.022127,2.837014,4.5460134,5.715527,6.5643673,6.670001,4.9723196,3.6443558,3.5575855,4.002755,4.644101,5.523123,6.7944975,6.643593,5.80607,4.8138695,3.983892,3.6896272,4.0480266,4.285702,4.1800685,4.0593443,4.1310244,4.7648253,5.3609,6.0814714,7.828197,8.182823,6.2097406,3.9989824,2.686109,2.4408884,3.772625,5.1760416,6.379509,7.3792543,8.4544525,8.296002,7.6320205,7.5829763,8.537451,10.163452,11.589504,12.808062,13.822898,13.856852,11.351829,9.718282,9.0807085,8.571404,8.20546,8.850578,11.989402,12.936331,12.510024,11.834724,12.359119,12.691111,12.864652,12.879742,13.000465,13.732355,15.47908,15.226315,14.2077055,13.472044,13.902123,14.426518,14.70192,14.268067,13.223051,12.223305,12.4307995,13.35132,14.347293,14.758509,13.917213,12.061082,9.967276,8.526133,8.20546,9.046755,10.220041,10.340765,10.344538,10.86516,12.208215,12.193124,11.378237,10.106862,8.480861,6.3342376,3.8405323,2.4031622,2.0258996,2.9841464,5.828706,8.428044,9.903141,9.827688,8.416726,6.5002327,4.5460134,4.1612053,4.9459114,6.349328,7.6282477,7.3113475,6.590776,5.2288585,3.6292653,2.8219235,3.0558262,4.0291634,4.9421387,5.3382645,5.081726,5.119452,5.311856,5.4401255,5.6061206,6.2399216,7.0963078,7.5301595,7.484888,6.9869013,6.119198,5.1534057,4.1536603,3.187868,2.546522,2.71629,4.1197066,5.349582,5.9230213,5.515578,3.953711,2.6597006,2.0145817,2.1843498,3.0407357,4.164978,4.568649,3.663219,2.5087957,1.6976813,1.3430545,1.6976813,2.323937,2.6597006,2.444661,1.7240896,1.1129243,1.0978339,1.478869,2.0258996,2.5012503,2.4182527,2.1654868,1.8184053,1.4373702,1.0827434,0.97333723,0.94692886,0.87147635,0.73188925,0.6111652,0.5017591,0.5281675,0.694163,1.0299267,1.6184561,2.263575,2.8936033,3.1010978,2.897376,2.71629,2.093807,1.478869,0.965792,0.68661773,0.80734175,0.88279426,1.0751982,1.0601076,0.7884786,0.45648763,0.44516975,0.44139713,0.47157812,0.5470306,0.65643674,0.7432071,0.7997965,0.77338815,0.67152727,0.55080324,0.452715,0.42630664,0.48666862,0.5583485,0.47157812,0.32821837,0.23390275,0.181086,0.16222288,0.19994913,0.18485862,0.17354076,0.23390275,0.34330887,0.36594462,0.32821837,0.24899325,0.150905,0.060362,0.0,0.09808825,0.1961765,0.29803738,0.41876137,0.56589377,0.6149379,0.56212115,0.4376245,0.29803738,0.21503963,0.33576363,0.5017591,0.6451189,0.6451189,0.35085413,0.181086,0.18485862,0.26408374,0.35839936,0.44139713,0.29426476,0.17731337,0.08677038,0.06413463,0.19994913,0.331991,0.4376245,0.47535074,0.44516975,0.3961256,0.5319401,1.2600567,2.425798,3.6443558,4.304565,4.98741,4.515832,3.3764994,2.1164427,1.358145,1.4939595,1.5354583,1.5882751,1.6524098,1.6184561,1.116697,0.62625575,0.27917424,0.116951376,0.090543,0.8903395,1.1581959,1.3732355,1.6976813,2.0673985,2.1956677,2.3616633,2.6106565,2.7728794,2.6295197,1.9051756,2.0560806,2.6672459,3.138824,3.3350005,3.5953116,4.2894745,4.466788,4.3800178,4.244203,4.2291126,4.1008434,3.9725742,4.183841,4.708236,5.172269,5.7117543,6.3945994,6.937857,7.118943,6.779407,7.4169807,8.043237,8.367682,8.329956,8.103599,7.937603,7.699928,7.635793,7.8923316,8.533678,9.831461,11.140562,12.283667,13.075918,13.313594,12.81938,12.713746,12.864652,13.140053,13.392818,13.200415,12.875969,12.596795,12.510024,12.709973,12.551523,12.313848,12.351574,12.615658,12.657157,12.381755,12.668475,13.27964,13.687083,13.079691,11.92904,11.027383,10.242677,9.593785,9.242931,9.273112,9.21275,8.66572,7.7904706,7.2962565,7.145352,6.881268,6.677546,6.647365,6.8737226,6.79827,6.820906,6.7643166,6.6322746,6.6134114,6.741681,6.903904,7.2358947,7.8131065,8.643084,9.295748,9.918231,10.355856,10.612394,10.831206,11.038701,12.294985,14.030393,15.98084,18.199142,19.229069,19.681786,19.527107,18.674494,16.961721,14.618922,12.15917,10.355856,9.7069645,10.401127,8.45068,6.6020937,5.2967653,4.5988297,4.1762958,4.164978,4.266839,4.425289,4.606375,4.7836885,4.9421387,5.0854983,4.9949555,4.568649,3.8556228,3.1727777,2.7879698,2.516341,2.282438,2.1013522,2.4484336,2.795515,3.0030096,2.9841464,2.6823363,2.1088974,1.5580941,1.0827434,0.7130261,0.46026024,0.422534,0.47912338,0.6526641,0.7997965,0.5772116,0.271629,0.29426476,0.33576363,0.24899325,0.05281675,0.033953626,0.011317875,0.0,0.00754525,0.03772625,0.049044125,0.026408374,0.00754525,0.003772625,0.00754525,0.0150905,0.026408374,0.05281675,0.1056335,0.19240387,0.271629,0.22258487,0.13958712,0.071679875,0.033953626,0.033953626,0.030181,0.018863125,0.00754525,0.02263575,0.0452715,0.03772625,0.026408374,0.018863125,0.00754525,0.003772625,0.003772625,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0150905,0.026408374,0.018863125,0.0150905,0.018863125,0.02263575,0.05281675,0.116951376,0.13204187,0.090543,0.049044125,0.02263575,0.011317875,0.0150905,0.026408374,0.041498873,0.041498873,0.041498873,0.026408374,0.00754525,0.018863125,0.120724,0.14335975,0.13958712,0.13204187,0.11317875,0.08299775,0.030181,0.0,0.0,0.0,0.033953626,0.026408374,0.02263575,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.0150905,0.011317875,0.018863125,0.056589376,0.10940613,0.14713238,0.13204187,0.120724,0.1056335,0.090543,0.056589376,0.03772625,0.026408374,0.033953626,0.05281675,0.071679875,0.060362,0.060362,0.0754525,0.090543,0.090543,0.07922512,0.06790725,0.056589376,0.049044125,0.071679875,0.10186087,0.26408374,0.49044126,0.68661773,0.7432071,0.694163,0.55080324,0.44139713,0.40367088,0.41498876,0.6790725,1.9202662,3.2633207,4.142342,4.2894745,4.032936,3.561358,2.897376,2.2069857,1.8146327,2.2560298,2.2183034,2.052308,2.1051247,2.71629,3.7914882,5.3194013,6.7680893,7.5716586,7.1340337,5.3458095,4.7421894,4.640329,4.768598,5.2552667,5.802297,6.0739264,6.039973,5.775889,5.4212623,5.402399,5.6023483,5.8513412,6.1342883,6.598321,6.6624556,6.1116524,5.511805,5.304311,5.7909794,5.5382137,5.0553174,4.776143,4.5724216,3.772625,3.893349,4.991183,6.771862,8.511042,9.076936,6.7114997,5.855114,5.975838,6.620957,7.405663,8.492179,9.439108,9.842778,9.442881,8.130007,6.688864,5.8437963,5.723072,6.6850915,9.314611,11.23865,11.3820095,11.306557,11.668729,12.2119875,12.189351,12.1101265,11.498961,10.7218,10.985884,12.528888,13.7700815,14.2077055,13.856852,13.27964,12.857106,13.015556,13.226823,13.419228,13.981348,14.977322,15.181043,14.400109,12.713746,10.487898,9.137298,8.197914,7.8508325,8.311093,9.81637,11.185833,12.276122,13.12119,13.694629,13.902123,13.102326,11.717773,9.955957,8.035691,6.2097406,4.13857,2.727608,2.4672968,3.5877664,6.0626082,8.59404,9.265567,8.582722,6.907676,4.4743333,3.059599,3.2444575,4.38379,5.696664,6.2851934,5.9682927,5.3646727,4.5460134,3.5802212,2.5314314,2.5276587,2.9652832,3.429316,3.6858547,3.7009451,3.6028569,3.6858547,3.863168,4.1197066,4.5196047,5.093044,5.8400235,6.488915,6.8774953,6.9869013,6.851087,6.0739264,4.9760923,4.123479,4.304565,5.7570257,6.617184,6.228604,4.6818275,2.8181508,1.9240388,1.7240896,2.052308,2.7389257,3.6179473,3.5689032,2.9992368,2.2258487,1.6033657,1.5015048,1.7769064,1.8976303,1.8636768,1.7127718,1.4939595,1.4562333,1.5656394,1.7429527,1.9127209,1.9881734,1.8070874,1.6788181,1.6373192,1.6260014,1.4977322,1.448688,1.3694628,1.20724,0.9922004,0.8299775,0.72811663,0.70170826,0.72811663,0.79602385,0.8865669,0.94692886,0.9242931,0.8903395,0.9620194,1.2751472,1.4939595,1.20724,0.7582976,0.422534,0.41876137,0.55080324,0.6752999,0.6488915,0.482896,0.35839936,0.3772625,0.44894236,0.5470306,0.6413463,0.694163,0.7092535,0.7130261,0.6790725,0.6187105,0.573439,0.5357128,0.452715,0.362172,0.28294688,0.21503963,0.17731337,0.14335975,0.15467763,0.20372175,0.211267,0.17731337,0.17731337,0.211267,0.24899325,0.1961765,0.2263575,0.44139713,0.62248313,0.66020936,0.56212115,0.5017591,0.46026024,0.41121614,0.36594462,0.34330887,0.32444575,0.33576363,0.36971724,0.422534,0.482896,0.47912338,0.4678055,0.44516975,0.38858038,0.25276586,0.16976812,0.1659955,0.20749438,0.26408374,0.32067314,0.331991,0.3169005,0.26408374,0.1961765,0.17354076,0.32821837,0.40367088,0.38480774,0.3169005,0.2867195,0.43007925,1.0223814,2.1013522,3.3425457,4.0706625,2.7351532,1.7052265,1.1921495,1.1959221,1.5430037,1.5015048,1.3166461,1.1619685,1.0525624,0.8601585,0.47912338,0.271629,0.27540162,0.482896,0.84884065,0.52062225,0.73566186,0.91674787,1.1317875,1.3241913,1.3166461,1.358145,1.5015048,1.7580433,2.0296721,2.0975795,2.5238862,2.776652,2.8143783,2.704972,2.6295197,2.9539654,3.1840954,3.4330888,3.6971724,3.874486,3.561358,3.1840954,3.0105548,3.2105038,3.832987,4.4818783,5.240176,5.7909794,6.0739264,6.2851934,7.1604424,7.7301087,8.088508,8.341274,8.624221,8.620448,8.375228,8.152642,8.141325,8.424272,9.050528,10.121953,11.317875,12.325166,12.800517,13.490907,14.6151495,15.049001,14.66042,14.317112,14.535924,14.532151,14.4114275,14.132254,13.528633,12.985375,12.58925,12.717519,13.313594,13.8719425,13.604086,13.332457,13.162688,13.04951,12.826925,11.9064045,10.665211,9.495697,8.601585,7.964011,7.7414265,7.4282985,6.9265394,6.25124,5.523123,5.100589,4.938366,4.847823,4.772371,4.8025517,5.0515447,5.1156793,4.927048,4.6327834,4.6026025,4.7233267,4.8440504,5.2326307,5.9117036,6.670001,6.8963585,7.2962565,7.7678347,8.22055,8.586494,9.242931,10.623712,12.189351,13.72481,15.316857,16.365646,17.093763,17.482344,17.712475,18.157644,18.467,18.89708,19.074392,19.036665,19.24416,17.886015,16.74291,16.022339,15.264041,13.373956,12.170488,11.763044,11.227332,10.246449,9.114662,8.303548,7.2057137,5.885295,4.6252384,3.904667,3.3764994,3.0822346,2.8143783,2.493705,2.1466236,2.142851,2.1503963,2.1503963,2.0900342,1.8749946,1.50905,1.1959221,0.8865669,0.5696664,0.29049212,0.2867195,0.36971724,0.5281675,0.633801,0.42630664,0.241448,0.29426476,0.32067314,0.21503963,0.026408374,0.0150905,0.003772625,0.0,0.003772625,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.003772625,0.06413463,0.18863125,0.31312788,0.3055826,0.26408374,0.17731337,0.10186087,0.060362,0.041498873,0.026408374,0.02263575,0.018863125,0.02263575,0.041498873,0.049044125,0.026408374,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.018863125,0.018863125,0.0150905,0.018863125,0.02263575,0.041498873,0.071679875,0.090543,0.08299775,0.05281675,0.02263575,0.00754525,0.0,0.0,0.00754525,0.00754525,0.011317875,0.011317875,0.011317875,0.02263575,0.06790725,0.0754525,0.09808825,0.14335975,0.150905,0.08299775,0.026408374,0.0,0.0,0.0,0.0452715,0.02263575,0.00754525,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.026408374,0.060362,0.094315626,0.08677038,0.07922512,0.08299775,0.09808825,0.1056335,0.090543,0.071679875,0.05281675,0.03772625,0.03772625,0.071679875,0.071679875,0.0754525,0.08677038,0.1056335,0.120724,0.1056335,0.1056335,0.10186087,0.090543,0.08299775,0.06790725,0.1056335,0.30181,0.62248313,0.8865669,0.94315624,0.7432071,0.46026024,0.24899325,0.2263575,0.32067314,0.7997965,1.3770081,1.9051756,2.3654358,3.4066803,3.9725742,4.1574326,3.9914372,3.4255435,3.3651814,3.2972744,2.848332,2.2107582,2.1277604,3.138824,4.7421894,6.439871,7.6207023,7.5565677,6.7077274,6.2097406,5.783434,5.3571277,5.0968165,4.878004,4.983638,5.2062225,5.3194013,5.0854983,5.6476197,6.741681,7.6282477,8.024373,8.130007,6.5266414,5.062863,4.025391,3.7235808,4.5120597,4.9949555,5.4665337,5.6325293,5.27413,4.2706113,3.2520027,3.62172,4.9232755,6.3229194,6.6322746,5.3986263,4.5799665,4.3121104,4.5460134,5.0741806,6.149379,7.24344,8.062099,8.141325,6.8133607,5.4363527,4.8742313,5.3986263,6.960493,9.22784,10.257768,10.084227,9.631512,9.522105,10.035183,11.038701,12.536433,12.728837,11.604594,10.9594755,11.461235,11.351829,10.661438,9.914458,10.137043,9.8239155,9.488152,10.121953,11.853588,13.962485,15.362129,15.516807,14.381247,12.272349,9.865415,8.469543,7.6886096,7.4999785,7.9036493,8.937348,10.831206,12.396846,13.513543,13.9888935,13.577678,12.728837,12.038446,10.691619,8.5563135,6.1531515,4.459243,3.3764994,3.0407357,3.361409,4.0216184,5.0854983,5.7796617,5.7004366,4.776143,3.2520027,2.3088465,2.3390274,3.1161883,4.104616,4.432834,4.485651,4.4139714,3.9989824,3.218049,2.2560298,2.4069347,2.5276587,2.5012503,2.474842,2.8898308,2.9992368,2.9841464,3.0520537,3.2746384,3.5839937,4.0782075,4.798779,5.594803,6.25124,6.477597,6.19465,5.270357,4.2102494,3.482133,3.519859,5.100589,5.926794,5.772116,4.708236,3.108643,2.1390784,1.8938577,2.0447628,2.3654358,2.6898816,2.4522061,2.1088974,1.7429527,1.4600059,1.3845534,1.4750963,1.4109617,1.2864652,1.1695137,1.1317875,1.3241913,1.418507,1.4637785,1.5203679,1.6863633,1.6033657,1.3128735,1.1431054,1.1883769,1.2902378,1.3355093,1.327964,1.2600567,1.1280149,0.95824677,0.814887,0.7582976,0.76207024,0.80356914,0.83752275,0.6790725,0.482896,0.33576363,0.3169005,0.49421388,0.6790725,0.6111652,0.4376245,0.28294688,0.24899325,0.28294688,0.331991,0.33576363,0.29049212,0.26408374,0.2867195,0.35839936,0.452715,0.5470306,0.6187105,0.6187105,0.5998474,0.55080324,0.49044126,0.44139713,0.38858038,0.32067314,0.241448,0.15845025,0.08677038,0.0754525,0.060362,0.06790725,0.094315626,0.08677038,0.07922512,0.07922512,0.094315626,0.120724,0.1358145,0.271629,0.5093044,0.724344,0.845068,0.83752275,0.784706,0.67152727,0.5357128,0.392353,0.24522063,0.26031113,0.29426476,0.3169005,0.32821837,0.36594462,0.35839936,0.29426476,0.23767537,0.211267,0.19994913,0.16976812,0.17731337,0.21503963,0.2678564,0.30935526,0.3055826,0.24522063,0.181086,0.14335975,0.13958712,0.2263575,0.27540162,0.28294688,0.2678564,0.24899325,0.30935526,0.59230214,1.0827434,1.6146835,1.8976303,1.0525624,0.5696664,0.543258,0.94315624,1.5882751,1.8749946,1.841041,1.6448646,1.3317367,0.83752275,0.41498876,0.3055826,0.5319401,1.0412445,1.6976813,0.633801,0.8186596,0.9507015,1.0223814,1.0186088,0.9016574,0.86770374,0.9808825,1.3053282,1.750498,2.0862615,2.4974778,2.7426984,2.8143783,2.7502437,2.6106565,2.5691576,2.6634734,2.8785129,3.0935526,3.1048703,2.7540162,2.4220252,2.191895,2.2296214,2.776652,3.712263,4.515832,5.0213637,5.3344917,5.8437963,6.7831798,7.77538,8.443134,8.744945,8.990166,9.484379,9.469289,9.046755,8.544995,8.503497,8.529905,8.888305,9.544742,10.33322,10.948157,12.151625,13.494679,13.88326,13.340002,13.004238,13.468271,13.728582,13.905896,13.928532,13.536179,12.721292,12.189351,12.178034,12.51757,12.615658,12.117672,11.7555,11.4838705,11.41219,11.781908,11.027383,9.650374,8.024373,6.670001,6.273875,6.48137,5.9682927,5.311856,4.7308717,4.0895257,3.7914882,3.7499893,3.6707642,3.4783602,3.31991,3.500996,3.519859,3.3878171,3.2444575,3.350091,3.2784111,3.2331395,3.470815,4.006528,4.606375,4.8063245,5.1571784,5.624984,6.145606,6.617184,6.903904,7.5188417,8.66572,10.201178,11.631002,12.808062,13.81158,14.966003,16.7995,20.036411,23.43932,26.849771,28.464457,28.173964,27.600525,26.766775,25.8123,25.231316,25.103046,25.12191,24.8201,24.786146,24.016531,22.469755,21.058792,20.398582,18.331184,15.452672,12.170488,8.6732645,6.009792,3.7688525,2.505023,2.0900342,1.7278622,1.5580941,1.4449154,1.3468271,1.20724,0.9393836,0.7507524,0.6451189,0.51684964,0.33953625,0.16222288,0.15845025,0.20372175,0.29426476,0.3961256,0.42630664,0.35839936,0.271629,0.18863125,0.1056335,0.00754525,0.0,0.003772625,0.00754525,0.011317875,0.02263575,0.02263575,0.0150905,0.003772625,0.0,0.00754525,0.030181,0.12826926,0.3055826,0.44894236,0.32821837,0.211267,0.120724,0.071679875,0.05281675,0.0452715,0.02263575,0.011317875,0.0150905,0.026408374,0.026408374,0.026408374,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.02263575,0.02263575,0.02263575,0.02263575,0.041498873,0.05281675,0.05281675,0.0452715,0.026408374,0.011317875,0.003772625,0.003772625,0.00754525,0.00754525,0.0150905,0.0150905,0.011317875,0.011317875,0.02263575,0.02263575,0.041498873,0.08299775,0.1358145,0.15467763,0.090543,0.0452715,0.0150905,0.0,0.0,0.030181,0.0150905,0.003772625,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.018863125,0.03772625,0.0452715,0.018863125,0.030181,0.049044125,0.071679875,0.090543,0.090543,0.08677038,0.07922512,0.060362,0.049044125,0.071679875,0.090543,0.090543,0.08677038,0.094315626,0.11317875,0.10186087,0.094315626,0.090543,0.08299775,0.08299775,0.07922512,0.056589376,0.17354076,0.46026024,0.84129536,1.0186088,0.94692886,0.69039035,0.38480774,0.2565385,0.2263575,0.3169005,0.42630664,0.58475685,0.97333723,2.8181508,4.715781,5.772116,5.7570257,5.1345425,4.195159,3.712263,3.1048703,2.3088465,1.750498,2.425798,3.6028569,5.2628117,6.8925858,7.4811153,7.2283497,6.7643166,6.1305156,5.4778514,5.0553174,4.425289,3.9084394,3.8782585,4.187614,4.195159,4.5497856,5.828706,7.1679873,8.307321,9.590013,8.043237,5.704209,3.802806,2.9728284,3.2369123,4.006528,4.8327327,5.3571277,5.3759904,4.82896,3.7009451,3.1614597,3.470815,4.304565,4.7572803,4.678055,4.0103,3.2859564,2.9841464,3.519859,4.5460134,5.73439,6.688864,6.907676,5.7796617,4.8553686,4.640329,5.240176,6.507778,8.009283,8.873214,9.114662,8.926031,8.714764,9.0957985,10.702937,12.73261,13.588995,12.879742,11.415963,10.487898,9.258021,8.001738,7.2660756,7.8432875,7.8206515,7.6282477,8.533678,10.710483,13.223051,14.792462,14.894323,13.675766,11.45369,8.726082,8.269594,8.314865,8.786444,9.250477,8.918486,9.205205,10.242677,11.121698,11.310329,10.642575,10.499215,10.789707,10.627484,9.522105,7.3905725,5.643847,4.496969,3.832987,3.482133,3.2331395,3.1425967,3.5462675,3.9084394,3.99521,3.8556228,3.8141239,2.9728284,2.372981,2.3578906,2.5502944,3.6481283,4.7421894,5.0553174,4.534695,3.8593953,3.7914882,3.6292653,3.2444575,2.757789,2.5238862,2.5012503,2.4220252,2.6068838,3.059599,3.500996,3.953711,4.2781568,4.5761943,4.7610526,4.561104,4.08198,3.338773,2.7087448,2.3767538,2.3163917,3.2105038,3.7084904,3.8141239,3.4783602,2.6106565,2.161714,2.2711203,2.6068838,2.9351022,3.138824,3.0143273,2.5389767,1.9655377,1.5128226,1.3619176,1.3091009,1.2298758,1.2147852,1.2638294,1.3091009,1.3241913,1.3543724,1.3958713,1.4562333,1.5467763,1.3996439,0.94692886,0.6187105,0.5696664,0.66775465,0.73566186,0.77338815,0.784706,0.754525,0.6413463,0.5394854,0.5017591,0.5093044,0.5319401,0.56589377,0.43385187,0.30935526,0.19994913,0.12826926,0.1358145,0.14335975,0.15845025,0.16222288,0.15467763,0.14335975,0.124496624,0.13204187,0.14713238,0.15467763,0.1659955,0.19240387,0.24522063,0.31312788,0.38858038,0.4678055,0.482896,0.543258,0.6375736,0.70170826,0.5998474,0.47535074,0.36594462,0.26408374,0.16222288,0.071679875,0.06413463,0.049044125,0.033953626,0.018863125,0.011317875,0.0150905,0.018863125,0.030181,0.056589376,0.10940613,0.21881226,0.33576363,0.44516975,0.5281675,0.5583485,0.543258,0.4640329,0.362172,0.26031113,0.13958712,0.16976812,0.20749438,0.241448,0.26031113,0.24899325,0.23390275,0.1659955,0.120724,0.120724,0.16976812,0.15467763,0.15845025,0.181086,0.211267,0.23390275,0.211267,0.14335975,0.094315626,0.09808825,0.12826926,0.18485862,0.23013012,0.24899325,0.24899325,0.26408374,0.31312788,0.3734899,0.42630664,0.452715,0.4376245,0.33953625,0.362172,0.5885295,1.0072908,1.5128226,1.9127209,1.9730829,1.7957695,1.4260522,0.83752275,0.46026024,0.34330887,0.52439487,0.9808825,1.629774,0.7054809,0.87902164,0.965792,0.9808825,0.9620194,0.97710985,1.0035182,1.1355602,1.3543724,1.5505489,1.4939595,1.6637276,2.1202152,2.6823363,3.2067313,3.591539,3.4745877,3.3236825,3.1727777,2.969056,2.5804756,2.4182527,2.4069347,2.3692086,2.305074,2.3805263,3.2746384,3.953711,4.3649273,4.644101,5.1043615,6.1644692,7.8319697,9.031664,9.454198,9.548513,10.412445,10.303039,9.378746,8.303548,8.231868,8.314865,8.130007,7.9753294,8.00551,8.2507305,8.975075,9.507015,9.740918,9.854096,10.310584,10.767072,11.114153,11.563096,12.166716,12.849561,12.208215,11.631002,11.272603,10.967021,10.238904,9.329701,9.065618,9.133525,9.363655,9.740918,8.854351,7.798016,6.273875,4.7912335,4.6629643,5.323174,4.67051,3.85185,3.399135,3.259548,3.229367,3.180323,3.048281,2.8445592,2.6785638,2.505023,2.4672968,2.5314314,2.6898816,2.969056,2.848332,2.6974268,2.6823363,2.8822856,3.289729,3.8556228,4.3611546,4.8327327,5.27413,5.7004366,5.13077,4.6026025,5.1269975,6.677546,8.20546,9.507015,10.604849,12.253486,15.116908,19.753464,24.465473,28.875671,30.78462,30.343224,30.02255,29.675468,28.660633,28.05324,29.037895,32.889744,35.16841,36.545418,36.63596,35.836166,35.315544,35.60226,33.764996,30.271544,25.042685,17.47857,11.555551,6.462507,3.5877664,2.6785638,1.8448136,1.1846043,1.0450171,1.0412445,0.9016574,0.4678055,0.2565385,0.17731337,0.1358145,0.090543,0.060362,0.041498873,0.030181,0.049044125,0.15845025,0.45648763,0.4678055,0.23390275,0.05281675,0.0150905,0.00754525,0.011317875,0.02263575,0.033953626,0.0452715,0.071679875,0.06790725,0.03772625,0.0150905,0.00754525,0.0150905,0.06790725,0.150905,0.27917424,0.35839936,0.19994913,0.090543,0.05281675,0.041498873,0.041498873,0.041498873,0.02263575,0.011317875,0.011317875,0.011317875,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.003772625,0.0,0.0,0.003772625,0.0150905,0.026408374,0.026408374,0.02263575,0.02263575,0.011317875,0.033953626,0.041498873,0.030181,0.011317875,0.003772625,0.003772625,0.003772625,0.00754525,0.011317875,0.0,0.011317875,0.0150905,0.011317875,0.00754525,0.018863125,0.0150905,0.06413463,0.11317875,0.1358145,0.13958712,0.1056335,0.090543,0.06413463,0.018863125,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.02263575,0.0452715,0.056589376,0.056589376,0.056589376,0.06790725,0.090543,0.094315626,0.0754525,0.060362,0.08677038,0.07922512,0.06790725,0.071679875,0.08677038,0.0754525,0.05281675,0.03772625,0.03772625,0.049044125,0.06413463,0.05281675,0.0754525,0.20749438,0.55080324,0.814887,1.026154,1.0110635,0.7582976,0.43385187,0.23013012,0.23767537,0.3470815,0.48666862,0.5998474,2.3692086,4.983638,6.360646,6.1342883,5.6476197,4.266839,3.4217708,2.9351022,2.5578396,1.9579924,1.7731338,2.2598023,3.682082,5.6551647,7.152897,7.1038527,6.907676,6.379509,5.7419353,5.621211,5.2288585,3.9650288,3.187868,3.2972744,3.7273536,3.3840446,3.821669,4.961002,6.900131,9.944639,10.148361,7.575431,4.927048,3.2784111,2.0862615,2.1466236,2.7653341,3.802806,4.859141,5.2628117,4.847823,3.8065786,3.3651814,3.8103511,4.4705606,4.3686996,3.7499893,2.8898308,2.3692086,3.0897799,3.92353,4.889322,5.323174,5.0854983,4.561104,4.255521,4.2102494,4.3611546,4.776143,5.6476197,6.507778,7.424526,8.379,9.186342,9.465516,10.608622,11.6875925,12.528888,12.58925,10.974566,9.009028,7.77538,7.1302614,6.881268,6.79827,6.7077274,7.115171,8.103599,9.635284,11.555551,12.996693,12.951422,11.695138,9.522105,6.749226,7.756517,9.1825695,10.714255,11.389555,9.590013,7.1378064,6.832224,7.0472636,6.9454026,6.470052,7.326438,8.224322,9.167479,9.733373,9.046755,7.3151197,5.8966126,4.776143,4.0706625,4.0178456,3.9197574,3.832987,4.06689,4.6252384,5.198677,5.9192486,4.4215164,2.516341,1.3317367,1.3166461,3.4745877,5.624984,6.752999,6.7643166,6.507778,5.8437963,5.1345425,4.395108,3.4972234,2.1956677,1.8334957,1.7542707,2.1051247,2.7691069,3.380272,3.7575345,3.5877664,3.1765501,2.6785638,2.11267,1.7957695,1.5807298,1.539231,1.599593,1.5505489,1.358145,1.3468271,1.3920987,1.388326,1.2751472,1.6863633,2.3692086,3.1199608,3.802806,4.376245,4.587512,3.9310753,2.8936033,1.9579924,1.5958204,1.4713237,1.4298248,1.5505489,1.7655885,1.8749946,1.6071383,1.5203679,1.5430037,1.5467763,1.3430545,1.0336993,0.6149379,0.3055826,0.16976812,0.10186087,0.13958712,0.14713238,0.14335975,0.1358145,0.09808825,0.1056335,0.1358145,0.13204187,0.090543,0.0452715,0.0452715,0.03772625,0.026408374,0.0150905,0.018863125,0.00754525,0.00754525,0.0150905,0.03772625,0.060362,0.07922512,0.08299775,0.07922512,0.0754525,0.09808825,0.13204187,0.1659955,0.20749438,0.26031113,0.3055826,0.3470815,0.51684964,0.77338815,0.9620194,0.8111144,0.6488915,0.4979865,0.35462674,0.23013012,0.14713238,0.12826926,0.1056335,0.071679875,0.049044125,0.07922512,0.08677038,0.0754525,0.06790725,0.07922512,0.094315626,0.071679875,0.060362,0.0452715,0.030181,0.018863125,0.0150905,0.00754525,0.011317875,0.026408374,0.041498873,0.056589376,0.10186087,0.1961765,0.29426476,0.271629,0.19994913,0.14335975,0.116951376,0.13204187,0.19240387,0.16222288,0.13958712,0.124496624,0.11317875,0.1056335,0.1056335,0.1056335,0.116951376,0.14713238,0.18863125,0.27540162,0.32821837,0.32067314,0.2867195,0.32067314,0.41876137,0.41121614,0.3734899,0.35085413,0.3470815,0.4074435,0.5357128,0.7809334,1.1016065,1.3505998,1.5430037,1.5165952,1.3430545,1.0487897,0.63002837,0.41498876,0.29803738,0.3772625,0.6790725,1.1544232,0.1056335,0.241448,0.3470815,0.422534,0.52439487,0.7922512,1.0751982,1.1808317,1.237421,1.3015556,1.3732355,1.3845534,1.5618668,1.9768555,2.505023,2.8219235,2.969056,3.1350515,3.4217708,3.802806,4.1197066,4.67051,4.8063245,4.255521,3.2331395,2.4408884,1.8938577,1.9278114,2.2296214,2.6521554,3.2520027,4.9345937,6.537959,7.7037,8.473316,9.291975,9.74469,8.933576,7.960239,7.3905725,7.232122,7.4396167,7.6093845,7.515069,7.224577,7.1264887,7.1868505,7.5792036,8.13378,8.809079,9.688101,10.103089,10.325675,10.601076,10.9594755,11.216014,11.506506,11.491416,11.385782,11.314102,11.276376,10.533169,9.65792,8.699674,7.677292,6.590776,5.383536,5.1534057,5.3269467,5.27413,4.3347464,3.7235808,3.2331395,3.108643,3.2972744,3.4179983,3.0143273,2.686109,2.4031622,2.2409391,2.3503454,2.4484336,2.5087957,2.5314314,2.5427492,2.5804756,2.7615614,2.8634224,2.9049213,2.9841464,3.2670932,3.5462675,3.772625,3.893349,3.9197574,3.904667,4.1272516,4.45547,4.9760923,5.8626595,7.4018903,8.631766,9.061845,9.763554,11.159425,13.015556,13.920986,14.879233,15.8676605,17.086218,18.953669,20.783392,22.337713,24.046711,26.136745,28.64177,31.79191,34.489338,36.334152,37.13395,36.926453,36.30397,36.21343,34.75342,30.822346,24.107073,18.700903,13.860624,10.155907,7.352846,4.4101987,1.5430037,0.91674787,0.94692886,0.80734175,0.44139713,0.32067314,0.26408374,0.1961765,0.10940613,0.060362,0.060362,0.060362,0.07922512,0.12826926,0.21503963,0.21503963,0.1659955,0.11317875,0.06790725,0.030181,0.056589376,0.07922512,0.1056335,0.120724,0.120724,0.09808825,0.056589376,0.030181,0.026408374,0.0150905,0.026408374,0.02263575,0.02263575,0.041498873,0.0754525,0.0754525,0.049044125,0.030181,0.030181,0.030181,0.030181,0.030181,0.02263575,0.011317875,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.0,0.0,0.011317875,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.0150905,0.011317875,0.0,0.0,0.00754525,0.02263575,0.030181,0.030181,0.018863125,0.041498873,0.10940613,0.17731337,0.150905,0.116951376,0.16222288,0.1659955,0.09808825,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.071679875,0.12826926,0.1358145,0.1056335,0.090543,0.06790725,0.116951376,0.150905,0.1358145,0.060362,0.049044125,0.0452715,0.06413463,0.10186087,0.1358145,0.124496624,0.094315626,0.06413463,0.049044125,0.060362,0.049044125,0.03772625,0.041498873,0.120724,0.36594462,0.66020936,0.9620194,1.1506506,1.0676528,0.52062225,0.33576363,0.27917424,0.3734899,0.58475685,0.8526133,1.4637785,2.2598023,2.8445592,3.350091,4.425289,4.6554193,4.1197066,3.6028569,3.2972744,2.8219235,1.5656394,1.8297231,2.927557,4.357382,5.798525,7.213259,8.850578,9.208978,8.329956,7.7829256,8.465771,6.858632,4.82896,3.7273536,4.4101987,4.606375,4.304565,4.4215164,5.194905,6.19465,6.3908267,5.670255,4.6327834,3.4896781,2.0749438,1.1091517,1.1280149,1.8938577,3.0897799,4.274384,4.063117,3.8556228,3.8820312,4.093298,4.164978,3.7990334,2.837014,2.3880715,2.8936033,4.1498876,4.8100967,5.138315,4.961002,4.3875628,3.8141239,3.3123648,3.270866,3.3274553,3.2029586,2.71629,2.191895,2.8106055,4.9345937,7.4999785,8.024373,8.111144,8.820397,9.431562,9.544742,9.0957985,7.61693,6.2135134,5.3948536,5.0553174,4.45547,3.6971724,3.802806,4.515832,5.73439,7.492433,8.235641,8.424272,7.884786,6.990674,6.6360474,7.149124,8.631766,9.971047,10.114408,8.088508,6.2323766,4.7044635,3.904667,3.893349,4.395108,5.6513925,6.379509,6.828451,7.3000293,8.118689,7.8734684,7.043491,5.66271,4.191386,3.4934506,4.508287,5.070408,5.168496,4.817642,4.074435,3.7801702,3.6971724,3.059599,1.9994912,1.5731846,3.2331395,4.606375,5.670255,6.3719635,6.651138,5.7872066,3.874486,2.3126192,1.5731846,1.2223305,1.2562841,1.2562841,1.0978339,0.97710985,1.4034165,1.6712729,1.4449154,1.0940613,0.86770374,0.91674787,0.98842776,1.0336993,1.0223814,0.97710985,0.97710985,1.0374719,1.1732863,1.2864652,1.3241913,1.2525115,1.2525115,1.4524606,1.9240388,2.6446102,3.5085413,4.032936,4.0178456,3.62172,2.9501927,2.0598533,1.8297231,1.7882242,1.7769064,1.7655885,1.8599042,1.8485862,1.5241405,1.146878,0.8563859,0.67152727,0.5998474,0.51684964,0.41121614,0.32067314,0.32067314,0.41876137,0.38858038,0.30181,0.20749438,0.120724,0.15845025,0.23013012,0.24899325,0.20372175,0.1659955,0.21503963,0.19240387,0.13204187,0.06790725,0.030181,0.030181,0.030181,0.030181,0.03772625,0.060362,0.09808825,0.116951376,0.116951376,0.10940613,0.120724,0.14713238,0.16222288,0.181086,0.20749438,0.24522063,0.3055826,0.38480774,0.3734899,0.26408374,0.150905,0.17731337,0.211267,0.22258487,0.23013012,0.3055826,0.20749438,0.1659955,0.120724,0.116951376,0.27540162,0.35839936,0.27917424,0.17731337,0.120724,0.1056335,0.094315626,0.090543,0.09808825,0.1056335,0.090543,0.06790725,0.041498873,0.03772625,0.056589376,0.090543,0.1659955,0.23767537,0.29803738,0.331991,0.32067314,0.211267,0.1659955,0.18485862,0.25276586,0.35085413,0.30181,0.25276586,0.19994913,0.13958712,0.090543,0.090543,0.12826926,0.18863125,0.27540162,0.3961256,0.482896,0.513077,0.5017591,0.4678055,0.44139713,0.44139713,0.3961256,0.33576363,0.2867195,0.27540162,0.47157812,0.7205714,0.9016574,1.0110635,1.1431054,1.3166461,1.2487389,1.0110635,0.70170826,0.45648763,0.35839936,0.35462674,0.84884065,1.7165444,2.2899833,0.02263575,0.049044125,0.06790725,0.08299775,0.1056335,0.15845025,0.271629,0.41876137,0.6451189,0.9205205,1.1280149,1.2110126,1.4562333,1.7693611,1.9429018,1.6750455,1.5279131,1.6146835,1.8334957,2.1315331,2.4974778,2.938875,3.1954134,3.3350005,3.3538637,3.1727777,2.8106055,2.5767028,2.3314822,2.1692593,2.4559789,3.663219,4.447925,4.859141,5.1873593,5.9984736,6.5455046,6.5341864,6.571913,6.7831798,6.828451,6.72659,6.7379084,6.7077274,6.5530496,6.258785,6.2625575,6.6813188,7.17176,7.6282477,8.16396,9.310839,9.993684,10.303039,10.423763,10.642575,10.710483,10.438853,10.299266,10.514306,11.042474,10.378491,9.544742,8.692128,7.91874,7.3113475,6.571913,5.8173876,5.1458607,4.5497856,3.8820312,3.712263,3.6368105,3.7499893,3.9348478,3.8707132,3.4859054,3.2935016,3.1840954,3.1161883,3.1199608,3.1199608,3.1048703,3.1199608,3.1765501,3.2633207,3.3463185,3.4972234,3.6858547,3.9310753,4.2781568,4.29702,4.244203,4.3309736,4.5535583,4.6856003,4.644101,4.3800178,4.172523,4.266839,4.8855495,5.270357,5.383536,5.2590394,5.168496,5.617439,7.1264887,8.45068,9.688101,10.876478,11.981857,13.196642,14.569878,16.078928,17.663431,19.217752,20.06282,21.990631,24.695602,27.260988,28.136238,28.65686,29.181253,28.166418,25.182272,20.900343,18.372684,15.943113,13.687083,11.351829,8.341274,5.062863,2.8596497,1.5203679,0.8224323,0.56589377,0.47157812,0.4074435,0.35839936,0.34330887,0.392353,0.4678055,0.35085413,0.19994913,0.120724,0.12826926,0.14713238,0.1358145,0.1056335,0.08299775,0.1056335,0.17731337,0.24899325,0.3169005,0.3734899,0.40367088,0.33953625,0.241448,0.15845025,0.11317875,0.10186087,0.16222288,0.124496624,0.060362,0.02263575,0.041498873,0.049044125,0.0452715,0.041498873,0.041498873,0.041498873,0.02263575,0.011317875,0.003772625,0.003772625,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.003772625,0.0150905,0.003772625,0.00754525,0.011317875,0.011317875,0.011317875,0.003772625,0.003772625,0.003772625,0.003772625,0.003772625,0.02263575,0.033953626,0.030181,0.011317875,0.0,0.060362,0.0452715,0.033953626,0.041498873,0.041498873,0.041498873,0.1056335,0.16222288,0.181086,0.17731337,0.120724,0.10186087,0.071679875,0.030181,0.049044125,0.011317875,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.03772625,0.10940613,0.14335975,0.13958712,0.11317875,0.090543,0.08677038,0.1056335,0.120724,0.116951376,0.071679875,0.060362,0.06413463,0.08299775,0.1056335,0.11317875,0.10186087,0.090543,0.094315626,0.1056335,0.09808825,0.056589376,0.0452715,0.060362,0.11317875,0.23013012,0.60362,0.9695646,1.1883769,1.1695137,0.87147635,0.55457586,0.44894236,0.45648763,0.49421388,0.5017591,0.84884065,1.2449663,1.5958204,2.1353056,3.4255435,5.142088,5.20245,4.644101,4.123479,3.9197574,3.308592,2.9124665,2.6182017,2.5993385,3.2972744,4.606375,6.3229194,8.00551,9.046755,8.6732645,8.058327,6.809588,5.8588867,5.5457587,5.6061206,5.8890676,5.9117036,5.9984736,6.432326,7.4509344,7.364164,5.8173876,4.22534,3.1652324,2.3918443,1.4750963,1.146878,1.4071891,2.1503963,3.138824,3.350091,3.006782,3.0633714,3.8178966,4.8855495,4.617693,3.9159849,3.1124156,2.8181508,3.9310753,5.27413,6.017337,6.0776987,5.481624,4.353609,5.247721,6.5266414,7.1604424,6.677546,5.1798143,3.3576362,2.8822856,3.5689032,4.9685473,6.3908267,6.643593,6.4549613,5.9909286,5.4212623,4.919503,4.398881,4.0480266,3.9876647,4.0706625,3.893349,3.6066296,3.519859,3.6368105,3.953711,4.4403796,5.138315,7.111398,9.288202,10.63503,10.163452,10.27663,10.182315,10.242677,10.272858,9.514561,8.167733,6.477597,5.323174,5.2099953,6.2361493,7.0963078,7.575431,7.541477,7.149124,6.8246784,6.6662283,6.224831,5.670255,5.040227,4.22534,4.6742826,6.0701537,6.5832305,5.5797124,3.6330378,2.41448,2.3503454,3.0030096,3.5085413,2.5729303,1.7731338,1.7919968,2.0560806,2.293756,2.5767028,2.2183034,1.7731338,1.6335466,1.6712729,1.2713746,1.0148361,0.7997965,0.62625575,0.5394854,0.633801,0.7469798,0.80356914,0.90543,1.0676528,1.2449663,1.1808317,1.1695137,1.1431054,1.0714256,0.965792,0.94692886,1.0186088,1.177059,1.3241913,1.2525115,1.3204187,1.3468271,1.2562841,1.1280149,1.2034674,1.3845534,1.4901869,1.539231,1.539231,1.4864142,1.5580941,1.5845025,1.569412,1.5958204,1.8485862,1.9655377,1.9429018,1.8787673,1.7919968,1.6486372,1.3392819,1.1204696,0.9318384,0.77716076,0.69793564,0.6790725,0.6413463,0.5772116,0.49421388,0.42630664,0.38480774,0.36594462,0.3470815,0.30935526,0.25276586,0.22258487,0.22258487,0.23013012,0.23013012,0.21503963,0.21503963,0.2565385,0.23767537,0.15467763,0.10940613,0.1358145,0.10940613,0.090543,0.07922512,0.02263575,0.049044125,0.041498873,0.041498873,0.05281675,0.049044125,0.07922512,0.13958712,0.15845025,0.13958712,0.116951376,0.13204187,0.13204187,0.116951376,0.10186087,0.14713238,0.12826926,0.13204187,0.16976812,0.21503963,0.23767537,0.29426476,0.38480774,0.422534,0.38103512,0.29049212,0.27917424,0.27540162,0.27917424,0.27540162,0.21503963,0.18863125,0.19240387,0.19240387,0.16976812,0.12826926,0.124496624,0.13204187,0.14713238,0.15467763,0.16222288,0.16976812,0.241448,0.34330887,0.4376245,0.48666862,0.44516975,0.36971724,0.36971724,0.41876137,0.35839936,0.18485862,0.13204187,0.15467763,0.2263575,0.3470815,0.3961256,0.44516975,0.55080324,0.67152727,0.68661773,0.6073926,0.6073926,0.56212115,0.43007925,0.26408374,0.35839936,0.4979865,0.7696155,1.20724,1.7919968,1.961765,1.6222287,1.0601076,0.5696664,0.482896,0.69793564,1.0412445,1.6260014,2.335255,2.8030603,0.0,0.0,0.0,0.0,0.0,0.0,0.03772625,0.10186087,0.211267,0.36971724,0.5470306,0.7092535,0.95447415,1.1732863,1.2336484,0.98465514,0.633801,0.56212115,0.633801,0.784706,0.9997456,1.358145,1.7882242,2.2258487,2.6031113,2.8634224,2.3390274,1.9089483,1.5467763,1.3091009,1.2864652,1.7089992,2.04099,2.3314822,2.674791,3.2331395,3.9650288,4.82896,6.013564,7.0963078,7.039718,6.6586833,6.3644185,6.0211096,5.5985756,5.1534057,5.251494,5.5306683,5.775889,6.0248823,6.5568223,7.7301087,8.624221,9.22784,9.6051035,9.895596,10.03141,10.023865,10.144588,10.438853,10.729345,10.272858,10.137043,10.016319,9.623966,8.6732645,7.888559,7.213259,6.4738245,5.6853456,5.05909,5.247721,5.13077,4.851596,4.587512,4.561104,4.4215164,4.395108,4.436607,4.504514,4.5761943,4.644101,4.617693,4.5460134,4.4894238,4.5233774,4.538468,4.5761943,4.7346444,5.0439997,5.4476705,5.7192993,5.832478,5.8928404,5.87775,5.624984,5.089271,4.4139714,3.9122121,3.7877154,4.1197066,5.4476705,6.4134626,6.198423,5.1345425,4.7120085,5.3609,6.3417826,7.4811153,8.635539,9.699419,10.314357,10.929295,11.502733,12.095036,12.887287,13.626721,15.184815,17.327667,19.383747,20.255224,20.75321,21.03993,20.028866,17.723793,15.207452,14.264296,13.192869,12.027128,10.657665,8.846806,6.4474163,3.8443048,2.0145817,1.1959221,0.90543,0.8865669,0.8186596,0.7130261,0.6413463,0.7205714,0.7809334,0.62248313,0.43385187,0.30935526,0.24522063,0.35085413,0.39989826,0.35462674,0.2565385,0.24899325,0.31312788,0.39989826,0.47912338,0.5319401,0.5470306,0.39989826,0.2565385,0.1659955,0.14713238,0.17731337,0.24899325,0.19240387,0.10186087,0.041498873,0.030181,0.026408374,0.02263575,0.018863125,0.018863125,0.018863125,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.02263575,0.026408374,0.0150905,0.011317875,0.0150905,0.00754525,0.0,0.0,0.0,0.0,0.00754525,0.026408374,0.030181,0.02263575,0.0150905,0.00754525,0.06790725,0.06790725,0.0452715,0.033953626,0.056589376,0.026408374,0.049044125,0.06790725,0.094315626,0.18485862,0.150905,0.124496624,0.0754525,0.018863125,0.02263575,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0452715,0.08299775,0.090543,0.08677038,0.08299775,0.08299775,0.09808825,0.120724,0.120724,0.09808825,0.06790725,0.06413463,0.060362,0.056589376,0.05281675,0.05281675,0.0452715,0.05281675,0.071679875,0.09808825,0.116951376,0.09808825,0.08677038,0.090543,0.116951376,0.181086,0.40367088,0.6828451,0.8526133,0.8526133,0.7130261,0.5357128,0.47912338,0.5357128,0.6111652,0.5583485,0.5772116,0.7432071,1.056335,1.6260014,2.6521554,4.1612053,5.040227,5.221313,4.8855495,4.4441524,3.8820312,3.6443558,3.5047686,3.519859,4.025391,4.134797,4.429062,5.5683947,7.201941,7.960239,7.8508325,6.8359966,5.8702044,5.560849,6.187105,6.466279,6.911449,7.7942433,8.831716,9.205205,8.43559,6.63982,4.5837393,2.9124665,2.142851,1.478869,1.2713746,1.4939595,2.003264,2.5427492,2.6182017,2.938875,3.9310753,5.462761,6.832224,6.7944975,5.794752,4.9723196,5.0553174,6.356873,7.0812173,7.2396674,6.8397694,6.1078796,5.485397,6.436098,7.9526935,8.873214,8.578949,6.9793563,4.678055,3.3651814,2.9426475,3.2029586,3.8103511,3.99521,3.6330378,3.1350515,2.8181508,2.9049213,3.5236318,4.2592936,5.032682,5.572167,5.409944,4.3686996,3.9461658,3.85185,3.874486,3.8593953,4.610148,6.379509,8.503497,10.220041,10.661438,10.733118,10.020092,8.967529,7.9753294,7.4207535,6.628502,5.406172,4.395108,4.06689,4.7120085,6.405917,7.3453007,7.092535,5.904158,4.7233267,4.3121104,4.2706113,4.4101987,4.515832,4.353609,4.112161,4.357382,4.22534,3.4217708,2.252257,1.5015048,1.4260522,1.7769064,2.0560806,1.5128226,0.9620194,0.94315624,1.2336484,1.6184561,1.8749946,1.599593,1.2487389,1.0978339,1.1431054,1.1091517,1.056335,1.0525624,1.1016065,1.1996948,1.3317367,1.3656902,1.3166461,1.2713746,1.2902378,1.3656902,1.2751472,1.2034674,1.1431054,1.0714256,0.9507015,0.8639311,0.8563859,0.94692886,1.0789708,1.1129243,1.1921495,1.3166461,1.3468271,1.2826926,1.2940104,1.1996948,1.0751982,1.0299267,1.0789708,1.1053791,1.146878,1.1431054,1.1317875,1.177059,1.3619176,1.4864142,1.5015048,1.4449154,1.3543724,1.2864652,1.1921495,1.2449663,1.327964,1.388326,1.4449154,1.3656902,1.297783,1.2185578,1.1317875,1.0601076,0.97333723,0.7507524,0.5281675,0.362172,0.2565385,0.120724,0.094315626,0.124496624,0.16222288,0.150905,0.11317875,0.16976812,0.1961765,0.1659955,0.13958712,0.1659955,0.15845025,0.1358145,0.10940613,0.06413463,0.02263575,0.003772625,0.003772625,0.00754525,0.00754525,0.018863125,0.041498873,0.05281675,0.060362,0.08677038,0.15845025,0.23767537,0.362172,0.4979865,0.56589377,0.42630664,0.30935526,0.271629,0.3055826,0.36594462,0.43007925,0.52062225,0.60362,0.66775465,0.7092535,0.7432071,0.724344,0.6413463,0.52439487,0.4376245,0.45648763,0.47535074,0.44894236,0.36594462,0.23767537,0.271629,0.392353,0.47912338,0.47157812,0.35085413,0.27917424,0.31312788,0.3961256,0.46026024,0.45648763,0.35839936,0.2678564,0.23767537,0.24899325,0.2263575,0.13204187,0.09808825,0.10940613,0.14335975,0.20749438,0.24522063,0.2867195,0.36594462,0.4678055,0.5357128,0.543258,0.6111652,0.6149379,0.4979865,0.3055826,0.2678564,0.32444575,0.51684964,0.9016574,1.5241405,1.7316349,1.4034165,0.95447415,0.6526641,0.633801,0.8262049,1.5656394,2.6483827,3.3689542,2.516341,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.011317875,0.03772625,0.120724,0.24899325,0.41498876,0.573439,0.6488915,0.5583485,0.33953625,0.392353,0.5394854,0.6828451,0.83752275,1.056335,1.358145,1.5580941,1.6335466,1.7354075,1.2562841,0.9922004,0.8337501,0.68661773,0.48666862,0.4376245,0.5357128,0.77716076,1.1242423,1.5052774,2.233394,3.1954134,4.4177437,5.4967146,5.587258,5.300538,4.9421387,4.61392,4.349837,4.115934,4.2328854,4.3611546,4.436607,4.5912848,5.138315,6.0512905,6.9567204,7.865923,8.733627,9.446653,9.8239155,10.054046,10.20495,10.382264,10.759526,10.876478,11.151879,11.449917,11.521597,11.00852,10.1294985,9.431562,8.646856,7.6622014,6.537959,5.9418845,5.3194013,4.7233267,4.3649273,4.6214657,5.089271,5.564622,5.926794,6.1720147,6.417235,6.6850915,6.6850915,6.511551,6.25124,6.006019,5.96452,5.994701,6.2135134,6.6322746,7.1566696,7.828197,8.209232,8.333729,8.050782,7.009537,5.873977,4.7836885,4.22534,4.3007927,4.7120085,6.0286546,7.2585306,7.6282477,7.2170315,6.952948,6.911449,7.5603404,8.654402,10.001229,11.472552,10.736891,10.287949,10.291721,10.79348,11.691365,12.883514,13.283413,13.521088,13.751218,13.656902,13.604086,13.407909,12.513797,11.080199,9.982366,9.9257765,9.333474,8.605357,7.9753294,7.541477,6.0701537,3.832987,2.2258487,1.6146835,1.3317367,1.3543724,1.2525115,1.0714256,0.9318384,1.0374719,1.0299267,0.84129536,0.62248313,0.44894236,0.3169005,0.38858038,0.41876137,0.36971724,0.28294688,0.27917424,0.33576363,0.42630664,0.4979865,0.52062225,0.4979865,0.33953625,0.21503963,0.1659955,0.17731337,0.1961765,0.211267,0.15467763,0.08299775,0.033953626,0.018863125,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.011317875,0.02263575,0.026408374,0.011317875,0.003772625,0.00754525,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.0150905,0.02263575,0.0150905,0.00754525,0.00754525,0.00754525,0.041498873,0.056589376,0.041498873,0.02263575,0.049044125,0.030181,0.018863125,0.011317875,0.05281675,0.21881226,0.211267,0.13204187,0.056589376,0.0150905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.033953626,0.056589376,0.056589376,0.041498873,0.041498873,0.05281675,0.06413463,0.07922512,0.09808825,0.09808825,0.0754525,0.06790725,0.06790725,0.05281675,0.03772625,0.02263575,0.02263575,0.026408374,0.033953626,0.0452715,0.06790725,0.10940613,0.120724,0.10940613,0.1056335,0.124496624,0.16222288,0.23767537,0.35839936,0.42630664,0.43007925,0.4376245,0.47535074,0.56212115,0.69793564,0.814887,0.7922512,0.5394854,0.48666862,0.6752999,1.1506506,1.9391292,3.0369632,4.45547,5.4212623,5.6287565,5.198677,4.4630156,4.1197066,4.1272516,4.436607,4.9760923,4.930821,5.028909,5.794752,6.9567204,7.454707,7.5829763,7.0472636,6.2851934,5.8664317,6.470052,6.5832305,7.232122,8.416726,9.325929,8.337502,7.164215,6.119198,4.7006907,3.0709167,2.0447628,1.6939086,1.7089992,1.9844007,2.3880715,2.7691069,2.9464202,3.6896272,5.2967653,7.5603404,9.774872,9.280658,8.039464,7.277394,7.443389,8.20546,8.22055,7.756517,6.8737226,5.828706,5.0515447,5.670255,6.7454534,7.3490734,7.145352,6.387054,5.330719,4.2781568,3.5575855,3.2746384,3.3161373,3.199186,2.565385,1.9655377,1.7693611,2.1466236,3.561358,4.9534564,6.168242,6.7869525,6.1606965,4.825187,4.3083377,4.244203,4.3309736,4.3309736,4.7346444,5.5268955,6.579458,7.828197,9.246704,9.820143,8.971302,7.462252,5.9984736,5.221313,4.429062,3.5085413,2.727608,2.3880715,2.795515,4.564876,5.485397,5.304311,4.2819295,3.199186,2.8822856,3.059599,3.5085413,3.9763467,4.172523,3.5839937,3.0520537,2.565385,2.1088974,1.6524098,1.3619176,1.2411937,1.1506506,1.056335,1.0072908,1.3392819,1.5052774,1.6448646,1.7655885,1.7429527,1.5920477,1.50905,1.3694628,1.1883769,1.1204696,1.3770081,1.6222287,1.8485862,2.0372176,2.1466236,2.071171,1.7769064,1.4939595,1.3392819,1.3355093,1.2336484,1.116697,1.0035182,0.90543,0.7997965,0.7130261,0.7205714,0.8526133,1.1242423,1.5165952,1.4675511,1.4977322,1.6637276,1.8938577,1.9844007,1.6863633,1.3732355,1.1657411,1.0751982,0.995973,0.9620194,0.935611,0.91674787,0.90920264,0.9205205,0.94692886,0.9318384,0.87902164,0.814887,0.7922512,0.8337501,0.98842776,1.1280149,1.1996948,1.2411937,1.1883769,1.1242423,1.0525624,0.9808825,0.9393836,0.875249,0.6526641,0.42630664,0.27540162,0.21881226,0.08677038,0.05281675,0.06413463,0.08299775,0.0754525,0.05281675,0.07922512,0.09808825,0.09808825,0.090543,0.10940613,0.1358145,0.12826926,0.090543,0.08299775,0.0452715,0.049044125,0.05281675,0.05281675,0.06413463,0.049044125,0.030181,0.030181,0.049044125,0.094315626,0.16976812,0.33576363,0.59607476,0.8865669,1.0902886,0.965792,0.72811663,0.573439,0.5696664,0.66020936,0.73566186,0.8111144,0.91297525,1.0676528,1.2789198,1.4034165,1.3807807,1.2449663,1.0525624,0.9016574,1.0223814,1.0978339,1.0714256,0.935611,0.7130261,0.65643674,0.90920264,1.1431054,1.177059,0.95447415,0.60362,0.35462674,0.2678564,0.2867195,0.26031113,0.17731337,0.116951376,0.07922512,0.06790725,0.071679875,0.060362,0.05281675,0.056589376,0.06413463,0.07922512,0.1056335,0.14335975,0.1961765,0.26031113,0.32444575,0.35839936,0.41121614,0.43385187,0.39989826,0.31312788,0.24522063,0.24899325,0.3169005,0.5017591,0.8941121,1.1204696,1.1053791,1.0186088,0.9507015,0.91674787,1.056335,1.8938577,3.2821836,4.172523,2.6219745,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.06413463,0.17354076,0.27917424,0.26408374,0.5055317,0.91297525,1.1996948,1.3204187,1.4901869,1.6033657,1.5807298,1.3807807,1.0751982,0.8526133,0.6375736,0.6526641,0.6790725,0.5885295,0.33576363,0.20372175,0.20372175,0.331991,0.59607476,1.0148361,1.4939595,1.8033148,2.1051247,2.4823873,2.9049213,2.9652832,2.886058,3.006782,3.338773,3.5575855,3.6179473,3.6179473,3.640583,3.7952607,4.2404304,4.8553686,5.59103,6.5341864,7.635793,8.726082,9.295748,9.661693,9.759781,9.876732,10.646348,11.476325,11.872451,12.174261,12.566614,13.045737,12.30253,11.423509,10.465261,9.34102,7.7829256,6.066381,4.9685473,4.4101987,4.3800178,4.8930945,5.9117036,6.9152217,7.643338,8.13378,8.722309,9.390063,9.786189,9.918231,9.808825,9.484379,8.967529,8.688355,8.661947,8.888305,9.371201,10.11818,10.378491,10.33322,9.786189,8.126234,6.628502,5.300538,4.8327327,5.2250857,5.7909794,6.0324273,6.809588,7.9715567,9.144843,9.7069645,9.857869,10.536942,11.759273,13.392818,15.192361,13.355092,12.321393,12.404391,13.404137,14.57365,15.520579,14.305794,12.51757,10.963248,9.676784,9.088254,8.541223,7.914967,7.2962565,6.983129,7.0887623,6.379509,5.5495315,5.0968165,5.311856,4.38379,2.9728284,2.0258996,1.7316349,1.5505489,1.5656394,1.5015048,1.3694628,1.237421,1.2487389,1.1393328,0.9205205,0.67152727,0.4376245,0.26408374,0.24899325,0.24522063,0.25276586,0.26031113,0.2263575,0.23767537,0.3055826,0.35085413,0.33953625,0.29049212,0.22258487,0.20372175,0.2565385,0.3169005,0.22258487,0.10940613,0.05281675,0.018863125,0.0,0.0,0.011317875,0.011317875,0.00754525,0.0,0.0,0.0,0.018863125,0.03772625,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.011317875,0.011317875,0.011317875,0.011317875,0.0150905,0.0150905,0.00754525,0.0,0.0,0.003772625,0.018863125,0.02263575,0.018863125,0.0150905,0.02263575,0.0452715,0.041498873,0.030181,0.06413463,0.21881226,0.21881226,0.08677038,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.030181,0.0452715,0.06790725,0.049044125,0.033953626,0.033953626,0.041498873,0.049044125,0.0452715,0.0452715,0.049044125,0.060362,0.06790725,0.06413463,0.056589376,0.0452715,0.0452715,0.05281675,0.06790725,0.0754525,0.06413463,0.0452715,0.0754525,0.09808825,0.090543,0.08677038,0.1056335,0.13204187,0.15467763,0.14713238,0.124496624,0.13958712,0.26408374,0.452715,0.6828451,0.87147635,0.9808825,1.0148361,0.7092535,0.4678055,0.41498876,0.65643674,1.2600567,2.2786655,3.7499893,5.168496,6.0550632,5.9909286,5.1232247,4.432834,4.304565,4.817642,5.745708,6.436098,7.24344,8.039464,8.428044,7.7376537,7.594294,7.598067,7.375482,6.952948,6.7567716,6.5341864,6.851087,7.405663,7.375482,5.4288073,4.3196554,4.5196047,4.7044635,4.2102494,3.0143273,2.7841973,2.9803739,3.2557755,3.500996,3.8254418,4.5535583,5.3873086,6.911449,9.2844305,12.223305,11.242422,9.884277,8.83926,8.307321,7.9828744,7.665974,6.9793563,6.058836,4.9685473,3.7009451,4.0895257,4.425289,4.29702,3.953711,4.293247,5.0175915,4.8365054,4.4139714,4.187614,4.406426,4.236658,3.3764994,2.4823873,2.0070364,2.191895,3.6934,5.2364035,6.40969,6.741681,5.66271,4.772371,4.395108,4.4403796,4.7044635,4.8930945,4.7610526,4.5837393,4.561104,5.062863,6.6322746,7.9489207,7.5301595,6.387054,5.1798143,4.22534,3.2029586,2.354118,1.7580433,1.5656394,2.0070364,2.6898816,2.8785129,2.8898308,2.8558772,2.6974268,2.8256962,2.9803739,3.2859564,3.6292653,3.6669915,3.180323,2.8256962,2.584248,2.372981,2.0447628,1.7240896,1.5430037,1.4373702,1.4034165,1.4977322,2.0975795,2.191895,1.9202662,1.4750963,1.1280149,1.2223305,1.7391801,1.9957186,1.7769064,1.3392819,1.6146835,1.9127209,2.1692593,2.3201644,2.3013012,2.11267,1.6939086,1.3694628,1.2600567,1.2638294,1.1280149,0.98842776,0.84129536,0.70170826,0.6111652,0.5772116,0.6488915,0.8903395,1.3468271,2.052308,1.9353566,1.7995421,1.9730829,2.3578906,2.4522061,2.0862615,1.6637276,1.3166461,1.0978339,0.97710985,0.9280658,0.9280658,0.90543,0.83752275,0.7394345,0.6752999,0.66020936,0.6790725,0.7092535,0.7167987,0.7205714,0.7394345,0.6752999,0.5281675,0.3734899,0.33576363,0.2867195,0.2263575,0.17731337,0.19240387,0.1961765,0.16222288,0.1358145,0.14335975,0.1961765,0.17354076,0.16222288,0.13958712,0.120724,0.120724,0.1358145,0.10186087,0.056589376,0.030181,0.02263575,0.030181,0.06413463,0.060362,0.026408374,0.03772625,0.120724,0.1961765,0.23390275,0.23390275,0.21881226,0.19240387,0.1659955,0.16976812,0.19994913,0.21503963,0.211267,0.3961256,0.6828451,0.9997456,1.2789198,1.3317367,1.1657411,1.0148361,0.97333723,1.0035182,1.0148361,1.0374719,1.1016065,1.2751472,1.6561824,1.9730829,2.0787163,1.9844007,1.7391801,1.3920987,1.5467763,1.6675003,1.690136,1.5920477,1.3732355,1.177059,1.4939595,1.8448136,1.9466745,1.720317,1.056335,0.4376245,0.124496624,0.09808825,0.07922512,0.06790725,0.049044125,0.033953626,0.033953626,0.041498873,0.030181,0.02263575,0.018863125,0.0150905,0.011317875,0.026408374,0.06413463,0.124496624,0.18863125,0.21503963,0.19994913,0.16976812,0.19240387,0.2678564,0.34330887,0.3169005,0.27917424,0.24522063,0.26031113,0.38103512,0.5885295,0.9016574,1.1242423,1.1883769,1.1393328,1.3770081,2.052308,3.3350005,4.3649273,3.240685,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.02263575,0.0452715,0.80356914,1.3128735,1.2261031,0.7696155,0.73188925,1.0148361,1.0450171,1.1695137,1.5354583,2.1202152,1.8749946,1.4675511,1.1393328,0.9205205,0.6413463,0.32444575,0.362172,0.6149379,1.0299267,1.6637276,1.81086,1.6184561,1.599593,1.8674494,2.1353056,2.233394,2.5616124,3.0746894,3.6330378,3.9989824,4.146115,3.9612563,3.85185,3.9688015,4.22534,4.617693,4.9987283,5.3646727,5.723072,6.089017,6.4926877,7.277394,8.096053,8.703445,8.971302,9.997457,11.125471,11.793225,11.921495,11.887542,11.642321,10.997202,10.197406,9.480607,9.061845,8.552541,7.9941926,7.7037,7.748972,7.91874,8.480861,9.0957985,9.782416,10.650121,11.932813,13.422999,15.256495,16.90136,18.089737,18.859352,16.614641,14.6151495,12.985375,11.910177,11.642321,11.570641,10.661438,9.495697,8.360137,7.2472124,6.2097406,5.3571277,5.1345425,5.523123,6.013564,6.6360474,7.7602897,9.035437,10.197406,11.0613365,12.049765,13.102326,14.471789,16.022339,17.240896,17.338985,17.520071,17.77661,17.882242,17.395575,16.516552,15.067864,13.494679,12.0082655,10.604849,9.955957,9.337247,8.6732645,7.8621507,6.7756343,5.6891184,4.6290107,3.6896272,2.916239,2.3201644,1.9429018,1.6260014,1.3694628,1.1846043,1.0978339,1.1242423,1.4222796,1.6863633,1.6637276,1.1732863,0.91674787,0.754525,0.5470306,0.30181,0.1659955,0.33953625,0.52062225,0.6828451,0.70170826,0.33576363,0.150905,0.09808825,0.07922512,0.056589376,0.0452715,0.094315626,0.25276586,0.52062225,0.7092535,0.44139713,0.17354076,0.060362,0.018863125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10186087,0.18485862,0.181086,0.0452715,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.0150905,0.00754525,0.0,0.003772625,0.0150905,0.05281675,0.02263575,0.0,0.0,0.0,0.0,0.026408374,0.026408374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.030181,0.030181,0.056589376,0.0754525,0.071679875,0.060362,0.049044125,0.03772625,0.03772625,0.041498873,0.030181,0.018863125,0.041498873,0.071679875,0.10186087,0.1358145,0.16222288,0.1961765,0.15845025,0.06413463,0.0150905,0.026408374,0.030181,0.02263575,0.02263575,0.0452715,0.056589376,0.071679875,0.094315626,0.14335975,0.23013012,0.4376245,0.633801,0.8186596,0.97710985,1.0978339,1.1355602,0.94315624,0.7582976,0.69793564,0.7469798,1.5882751,2.7238352,4.214022,5.5382137,5.5985756,4.817642,4.678055,5.111907,6.270103,8.529905,8.420499,7.4207535,7.0812173,7.665974,8.179051,8.812852,8.695901,8.22055,7.696155,7.352846,6.6360474,5.794752,5.2137675,4.9534564,4.745962,3.8895764,4.3649273,5.855114,7.152897,6.1644692,5.492942,5.9003854,6.2361493,6.0248823,5.462761,6.8058157,8.231868,9.461743,10.465261,11.427281,12.049765,10.220041,7.9753294,6.458734,5.9192486,5.3609,4.7874613,4.5309224,4.640329,4.8968673,5.1798143,4.82896,4.2592936,3.904667,4.195159,3.953711,3.451952,3.029418,2.8822856,3.0520537,4.06689,4.1083884,3.5651307,2.9728284,3.0218725,3.7537618,5.2175403,6.187105,6.25124,5.798525,4.957229,4.561104,4.606375,4.8930945,5.0515447,5.1345425,4.315883,3.4594972,3.0445085,3.127506,4.6290107,5.885295,5.7381625,4.432834,3.6179473,3.4330888,3.0935526,2.7238352,2.4484336,2.4107075,2.0673985,1.4713237,1.4411428,2.0749438,2.746471,2.9539654,2.916239,2.7238352,2.5314314,2.516341,2.2862108,1.9089483,1.7542707,1.8976303,2.1051247,1.7278622,1.5241405,1.478869,1.4750963,1.267602,1.0827434,0.9922004,0.8865669,0.77338815,0.76207024,0.8865669,1.116697,1.4222796,1.6335466,1.448688,1.0601076,1.1280149,1.3392819,1.50905,1.5580941,1.4449154,1.2713746,1.2223305,1.3015556,1.3128735,1.1280149,0.9922004,0.88279426,0.7922512,0.73188925,0.7092535,0.7092535,0.79602385,0.9808825,1.237421,1.5769572,1.9391292,2.3277097,2.686109,2.867195,2.686109,1.9164935,1.1846043,0.7696155,0.6111652,0.56212115,0.56589377,0.6111652,0.663982,0.70170826,0.77338815,0.7922512,0.8111144,0.8639311,0.9620194,1.0714256,1.1883769,1.146878,0.935611,0.7167987,0.47157812,0.32067314,0.211267,0.14335975,0.1659955,0.19240387,0.20749438,0.21881226,0.23013012,0.24522063,0.27917424,0.29049212,0.29049212,0.29426476,0.3055826,0.23013012,0.15845025,0.10940613,0.094315626,0.1056335,0.1056335,0.1056335,0.06413463,0.0,0.0,0.2678564,0.5017591,0.6451189,0.67152727,0.55080324,0.56212115,0.6111652,0.6526641,0.65643674,0.59607476,0.47157812,0.56212115,0.73188925,0.83752275,0.7167987,0.83752275,1.1431054,1.3166461,1.2713746,1.1732863,0.8941121,0.6488915,0.48666862,0.58475685,1.267602,1.9730829,2.5276587,2.6068838,2.1466236,1.3430545,1.1846043,1.1544232,1.2826926,1.4826416,1.5580941,1.5920477,1.8674494,2.1353056,2.233394,2.0749438,1.3920987,0.7167987,0.35839936,0.31312788,0.27540162,0.21503963,0.150905,0.090543,0.041498873,0.030181,0.018863125,0.02263575,0.02263575,0.011317875,0.0,0.02263575,0.056589376,0.094315626,0.13958712,0.21503963,0.23767537,0.23390275,0.29426476,0.44139713,0.62625575,0.49044126,0.36594462,0.27917424,0.271629,0.38103512,0.5394854,0.6451189,0.73566186,0.8337501,0.9318384,1.4449154,2.11267,3.0331905,3.7914882,3.4481792,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.16222288,0.26408374,0.24899325,0.16222288,0.14713238,0.211267,0.23767537,0.3734899,0.63002837,0.875249,0.77716076,0.7507524,0.91674787,1.1695137,1.1544232,0.83752275,0.76584285,0.7432071,0.7167987,0.784706,0.784706,0.754525,0.90920264,1.327964,1.9278114,2.474842,2.9652832,3.5123138,4.123479,4.6931453,4.4403796,4.112161,4.0517993,4.2592936,4.398881,4.504514,4.6327834,4.7950063,5.149633,6.013564,6.9567204,7.809334,8.231868,8.231868,8.167733,8.341274,8.831716,9.473062,10.208723,11.068882,11.751727,12.106354,12.5326605,13.200415,14.045483,14.437836,14.735873,14.943368,15.339493,16.486372,18.12369,18.670721,18.821627,18.983849,19.266796,19.429018,19.711966,20.88148,22.93756,25.133228,26.04243,24.156118,21.005976,17.829426,15.596032,13.79649,12.434572,11.121698,9.650374,7.9941926,6.458734,5.455216,5.0439997,5.191132,5.7570257,6.620957,7.7301087,8.741172,9.484379,9.940866,11.212241,12.936331,15.520579,18.459454,20.353312,21.115381,20.730574,19.859098,18.742401,17.199398,16.214743,15.347038,14.441608,13.370183,12.034674,10.401127,9.363655,8.612903,8.009283,7.61693,6.530414,4.61392,2.916239,1.8259505,1.0638802,0.91674787,0.9393836,1.177059,1.4637785,1.4298248,1.2864652,1.4939595,1.629774,1.478869,1.0412445,0.8337501,0.67152727,0.49421388,0.3169005,0.241448,0.32444575,0.28294688,0.21503963,0.1659955,0.13958712,0.094315626,0.05281675,0.033953626,0.03772625,0.0452715,0.08299775,0.13204187,0.18485862,0.24899325,0.32067314,0.27540162,0.15467763,0.05281675,0.011317875,0.0,0.011317875,0.018863125,0.030181,0.033953626,0.02263575,0.003772625,0.018863125,0.03772625,0.03772625,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.003772625,0.011317875,0.011317875,0.02263575,0.030181,0.0,0.0,0.011317875,0.018863125,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.0150905,0.02263575,0.03772625,0.05281675,0.049044125,0.056589376,0.07922512,0.094315626,0.090543,0.06790725,0.033953626,0.033953626,0.0452715,0.071679875,0.1358145,0.181086,0.211267,0.21881226,0.19240387,0.124496624,0.08677038,0.049044125,0.030181,0.026408374,0.02263575,0.02263575,0.041498873,0.0754525,0.11317875,0.13204187,0.241448,0.43007925,0.6526641,0.875249,1.086516,1.056335,0.91674787,0.7469798,0.5998474,0.55080324,0.7997965,1.5505489,2.5314314,3.440634,3.953711,5.455216,6.7152724,7.069899,6.752999,6.8925858,6.647365,5.987156,5.617439,6.224831,8.495952,8.98262,8.326183,7.17176,5.9984736,5.119452,5.093044,5.1534057,5.3684454,5.798525,6.4926877,6.2625575,6.3417826,6.8133607,7.3905725,7.3981175,8.024373,8.201687,7.77538,6.934085,6.19465,5.342037,5.828706,7.0812173,8.75249,10.7218,11.627231,11.5857315,10.967021,10.095545,9.265567,8.518587,7.8508325,7.0057645,6.217286,6.1908774,6.5002327,6.94163,6.8397694,6.1606965,5.5268955,4.4705606,4.1272516,4.5988297,5.330719,5.100589,4.719554,4.772371,4.4441524,3.5839937,2.704972,5.0854983,7.220804,8.616675,8.892077,7.77538,4.776143,3.3236825,2.8143783,2.9539654,3.7575345,4.52715,4.5497856,3.5575855,2.123988,1.6637276,2.8898308,4.357382,5.3458095,5.485397,4.715781,4.4931965,4.2102494,3.8178966,3.3727267,3.0331905,3.3651814,3.1765501,2.686109,2.3465726,2.8332415,3.3538637,3.1840954,2.9539654,2.9916916,3.361409,2.8822856,2.252257,1.6863633,1.3204187,1.2261031,1.2298758,1.1129243,0.97333723,0.875249,0.8639311,0.8262049,0.8299775,0.95824677,1.1091517,1.0186088,0.87902164,0.8903395,0.8978847,0.8262049,0.6790725,0.8563859,1.3053282,1.8523588,2.372981,2.8030603,2.505023,2.5578396,2.7879698,2.9086938,2.5201135,1.8599042,1.4260522,1.1204696,0.9205205,0.87902164,0.9318384,1.0487897,1.3505998,1.8448136,2.444661,3.059599,3.4896781,3.7575345,3.783943,3.380272,2.6219745,1.7542707,1.1091517,0.784706,0.633801,0.5772116,0.58098423,0.6375736,0.7432071,0.8978847,1.086516,1.3543724,1.5015048,1.4562333,1.2789198,1.2336484,1.1355602,0.9997456,0.8563859,0.754525,0.65643674,0.52439487,0.41121614,0.34330887,0.33953625,0.31312788,0.27917424,0.28294688,0.32821837,0.3772625,0.49421388,0.66775465,0.845068,0.9318384,0.8186596,0.68661773,0.47535074,0.29426476,0.18863125,0.14335975,0.17354076,0.20749438,0.2263575,0.241448,0.32821837,0.5885295,0.8903395,1.1355602,1.2638294,1.267602,1.4373702,1.629774,1.659955,1.5015048,1.2525115,0.97710985,0.87147635,0.87147635,0.8639311,0.694163,0.63002837,0.69039035,0.77716076,0.814887,0.7469798,0.7507524,0.62248313,0.452715,0.47912338,1.0827434,2.0862615,2.9086938,2.9954643,2.2560298,1.0487897,1.1355602,1.4222796,1.7542707,2.0183544,2.1315331,2.1956677,2.2447119,2.2484846,2.1768045,1.9768555,1.448688,0.995973,0.7469798,0.663982,0.58098423,0.422534,0.28294688,0.18485862,0.13958712,0.17731337,0.18485862,0.1659955,0.13204187,0.08299775,0.011317875,0.018863125,0.0452715,0.09808825,0.15845025,0.19994913,0.21503963,0.20372175,0.19994913,0.23013012,0.29426476,0.3772625,0.60362,0.98465514,1.4147344,1.7014539,1.6637276,1.4600059,1.3468271,1.4222796,1.6373192,1.6448646,1.8485862,2.5729303,3.561358,3.9612563,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0150905,0.03772625,0.120724,0.241448,0.33576363,0.331991,0.331991,0.41876137,0.5470306,0.56589377,0.47157812,0.44894236,0.44139713,0.422534,0.39989826,0.32821837,0.32067314,0.43385187,0.724344,1.2449663,1.8599042,2.4295704,3.0256453,3.6594462,4.2894745,4.236658,4.183841,4.3007927,4.557331,4.7233267,4.8629136,5.0025005,5.1458607,5.3684454,5.8211603,6.670001,7.5037513,8.111144,8.431817,8.541223,8.635539,8.990166,9.537196,10.284176,11.314102,12.449662,13.404137,14.2077055,14.920732,15.618668,15.829934,16.207197,16.610868,17.342756,19.153618,20.756983,21.254969,21.21347,20.972023,20.673985,20.209951,19.666695,19.47429,19.753464,20.304268,20.643805,20.209951,19.202662,17.931286,16.807045,16.697638,16.90136,16.697638,15.629986,13.505998,10.280403,8.771353,8.167733,7.9941926,8.126234,8.013056,7.6848373,7.699928,8.14887,8.669493,10.005001,12.012038,14.818871,18.206688,21.609596,24.220253,25.186045,24.854053,23.511,21.379465,18.478317,16.003475,14.234114,13.102326,12.208215,11.427281,10.540714,9.639057,8.854351,8.348819,6.722818,4.3611546,2.4710693,1.4109617,0.694163,0.68661773,0.7092535,0.8111144,0.94692886,0.98842776,1.0412445,1.3091009,1.4071891,1.20724,0.8526133,0.70170826,0.6187105,0.6187105,0.633801,0.51684964,0.36594462,0.211267,0.090543,0.030181,0.056589376,0.041498873,0.018863125,0.011317875,0.02263575,0.03772625,0.060362,0.08299775,0.1056335,0.124496624,0.150905,0.181086,0.18863125,0.15467763,0.08299775,0.018863125,0.030181,0.03772625,0.041498873,0.041498873,0.030181,0.02263575,0.011317875,0.026408374,0.0754525,0.15467763,0.09808825,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.018863125,0.02263575,0.00754525,0.0,0.00754525,0.026408374,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.0150905,0.030181,0.03772625,0.049044125,0.06413463,0.071679875,0.06413463,0.049044125,0.033953626,0.026408374,0.026408374,0.05281675,0.10940613,0.12826926,0.14335975,0.14335975,0.12826926,0.1056335,0.07922512,0.049044125,0.026408374,0.02263575,0.02263575,0.018863125,0.02263575,0.0452715,0.0754525,0.08677038,0.150905,0.331991,0.5772116,0.8186596,0.9997456,0.98842776,0.9242931,0.814887,0.6828451,0.55080324,0.6187105,1.1280149,1.9240388,2.8030603,3.5123138,4.7610526,5.353355,5.3646727,5.149633,5.3571277,6.3153744,7.2057137,7.3000293,6.9491754,7.5792036,7.5603404,6.771862,5.704209,4.7421894,4.168751,4.4101987,4.779916,5.119452,5.462761,6.013564,6.5530496,7.654656,9.099571,9.948412,8.5563135,7.635793,7.043491,6.670001,6.5455046,6.85486,5.0025005,4.2064767,4.8553686,6.8359966,9.5183325,11.155652,10.853842,9.857869,8.846806,7.960239,7.635793,7.7338815,7.443389,6.802043,6.700182,7.3981175,7.575431,7.2924843,6.79827,6.5568223,5.715527,4.927048,4.8327327,5.240176,5.138315,4.236658,4.074435,4.4101987,4.7648253,4.447925,5.696664,6.6662283,6.888813,6.1531515,4.496969,2.7804246,1.9693103,1.7618159,2.123988,3.2859564,4.8402777,4.908185,3.9386206,2.5691576,1.599593,2.2598023,3.5538127,4.534695,4.8100967,4.561104,4.4441524,4.0895257,3.5387223,2.9728284,2.7125173,3.2218218,3.500996,3.1840954,2.4899325,2.203213,2.6332922,2.7841973,2.8332415,2.9916916,3.470815,3.5424948,3.3010468,2.8219235,2.1503963,1.3355093,1.2147852,1.1695137,1.0978339,1.0072908,1.0299267,1.5430037,2.003264,2.323937,2.41448,2.2107582,1.7089992,1.2864652,0.94315624,0.7092535,0.633801,0.7394345,0.9620194,1.2713746,1.6750455,2.2447119,2.6936543,3.4859054,4.2102494,4.4894238,3.983892,3.029418,2.1390784,1.4109617,0.9205205,0.724344,0.7507524,0.9205205,1.2562841,1.750498,2.3616633,3.0369632,3.5990841,3.8367596,3.6481283,3.0331905,2.1466236,1.4562333,1.0450171,0.875249,0.814887,0.79602385,0.8186596,0.86770374,0.95824677,1.1091517,1.2411937,1.3732355,1.4222796,1.358145,1.2034674,1.086516,0.98465514,0.91297525,0.8601585,0.80734175,0.76207024,0.68661773,0.60362,0.55080324,0.573439,0.633801,0.5885295,0.5093044,0.42630664,0.3470815,0.35839936,0.482896,0.66775465,0.8337501,0.9016574,0.965792,0.94692886,0.8299775,0.63002837,0.4074435,0.24899325,0.19994913,0.2565385,0.38103512,0.52062225,0.8941121,1.327964,1.6486372,1.81086,1.9089483,2.1579416,2.3390274,2.3013012,2.04099,1.7014539,1.3845534,1.2223305,1.1280149,1.0336993,0.8865669,0.7054809,0.58098423,0.56589377,0.62625575,0.66775465,0.814887,0.7582976,0.573439,0.43385187,0.62625575,1.3355093,1.9429018,2.1051247,1.7882242,1.2525115,1.448688,1.9051756,2.3956168,2.71629,2.686109,2.4597516,2.323937,2.2371666,2.1466236,1.9881734,1.6260014,1.267602,1.0035182,0.84884065,0.7205714,0.5281675,0.34330887,0.23013012,0.27917424,0.5998474,0.76584285,0.59607476,0.35462674,0.1659955,0.05281675,0.02263575,0.026408374,0.056589376,0.094315626,0.116951376,0.120724,0.11317875,0.10940613,0.116951376,0.13958712,0.23013012,0.48666862,0.88279426,1.3468271,1.7655885,1.9844007,1.8938577,1.8070874,1.8221779,1.8259505,1.3505998,1.177059,1.5015048,2.384299,3.7235808,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.033953626,0.08677038,0.17354076,0.3055826,0.30935526,0.23390275,0.17731337,0.1659955,0.16976812,0.1961765,0.26031113,0.36594462,0.49044126,0.5772116,0.49044126,0.34330887,0.271629,0.35462674,0.633801,1.0827434,1.5807298,2.1390784,2.7238352,3.240685,3.4217708,3.7952607,4.236658,4.6214657,4.8402777,5.0439997,5.2779026,5.4891696,5.6551647,5.798525,6.3342376,7.0057645,7.7112455,8.360137,8.884532,9.325929,9.857869,10.370946,10.876478,11.54046,12.5326605,13.411682,14.003984,14.32843,14.607604,14.626467,14.777372,15.011275,15.531898,16.803272,17.772837,18.240643,18.417955,18.414183,18.255732,17.89356,17.354074,16.686321,16.014793,15.531898,15.105591,15.264041,15.607349,15.901614,16.109108,17.40312,18.840488,19.945868,20.055275,18.316093,15.158407,13.475817,12.555296,11.974312,11.615912,10.714255,9.522105,8.710991,8.503497,8.661947,9.397609,10.933067,13.087236,15.905387,19.644058,23.22428,25.804754,26.974268,26.740366,25.4954,21.507734,17.984104,15.331948,13.70972,13.023102,12.672247,11.627231,10.54826,9.797507,9.416472,7.3679366,4.930821,2.8936033,1.5656394,0.7582976,0.70170826,0.6752999,0.6526641,0.6451189,0.7092535,0.87147635,1.1129243,1.1355602,0.9016574,0.63002837,0.543258,0.5772116,0.7469798,0.91674787,0.80734175,0.58098423,0.38858038,0.23390275,0.11317875,0.030181,0.018863125,0.0150905,0.0150905,0.0150905,0.018863125,0.026408374,0.049044125,0.0754525,0.090543,0.071679875,0.1056335,0.1659955,0.16976812,0.09808825,0.018863125,0.026408374,0.026408374,0.026408374,0.03772625,0.071679875,0.094315626,0.06413463,0.049044125,0.08299775,0.16222288,0.09808825,0.033953626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.00754525,0.00754525,0.003772625,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.00754525,0.0,0.003772625,0.018863125,0.030181,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.00754525,0.00754525,0.0,0.003772625,0.011317875,0.026408374,0.049044125,0.056589376,0.056589376,0.056589376,0.049044125,0.041498873,0.03772625,0.026408374,0.026408374,0.03772625,0.071679875,0.08299775,0.08299775,0.06790725,0.056589376,0.071679875,0.056589376,0.041498873,0.026408374,0.02263575,0.03772625,0.02263575,0.030181,0.041498873,0.060362,0.071679875,0.09808825,0.21503963,0.39989826,0.5998474,0.7432071,0.8299775,0.90543,0.94692886,0.91297525,0.72811663,0.69039035,0.95447415,1.5731846,2.4333432,3.2331395,3.7235808,3.6594462,3.399135,3.2633207,3.5236318,4.5422406,5.772116,6.187105,5.798525,5.6778007,5.7192993,5.330719,4.776143,4.323428,4.2404304,4.644101,5.0779533,5.342037,5.3646727,5.198677,5.7683434,7.3075747,8.948667,9.556059,7.7414265,6.4549613,5.9305663,5.8890676,6.0211096,5.9682927,3.9574835,3.289729,4.2064767,6.462507,9.2995205,9.918231,8.699674,7.4811153,6.8473144,6.126743,5.198677,5.523123,6.0362,6.258785,6.319147,6.749226,6.2927384,5.832478,5.783434,6.115425,5.832478,5.089271,4.5497856,4.38379,4.266839,3.5839937,3.9386206,4.9119577,5.794752,5.583485,5.5382137,5.251494,4.3611546,2.969056,1.6071383,1.4071891,1.418507,1.690136,2.3465726,3.5689032,4.9044123,4.8063245,4.08198,3.1840954,2.2107582,1.8523588,2.625747,3.8593953,4.776143,4.478106,4.0782075,3.5575855,2.987919,2.5012503,2.305074,2.7238352,3.3425457,3.5349495,3.1010978,2.252257,1.8184053,2.335255,3.127506,3.8480775,4.4516973,4.678055,4.4743333,3.8480775,2.867195,1.6410918,1.4864142,1.5618668,1.5543215,1.4298248,1.4449154,2.0485353,2.6710186,3.127506,3.3651814,3.4481792,2.7125173,1.9504471,1.3430545,0.9922004,0.91674787,0.8903395,0.8186596,0.8111144,0.9808825,1.4562333,2.2484846,3.180323,3.8367596,3.9688015,3.5160866,2.637065,1.8184053,1.1732863,0.7507524,0.5583485,0.543258,0.6413463,0.84129536,1.1317875,1.5128226,1.9881734,2.4295704,2.5993385,2.4333432,2.0258996,1.4939595,1.1619685,1.0035182,0.95447415,0.9318384,0.8941121,0.87902164,0.8941121,0.94315624,1.0374719,1.086516,1.0789708,1.0450171,0.995973,0.94692886,0.875249,0.845068,0.84884065,0.86770374,0.875249,0.8526133,0.8111144,0.7394345,0.66020936,0.633801,0.6790725,0.6451189,0.5583485,0.43007925,0.27540162,0.1961765,0.211267,0.31312788,0.4640329,0.5885295,0.72811663,0.9205205,1.0525624,1.0525624,0.87902164,0.6828451,0.5394854,0.513077,0.58475685,0.65643674,0.86770374,1.2261031,1.6146835,1.9579924,2.2296214,2.5767028,2.8294687,2.848332,2.6182017,2.2220762,1.9579924,1.7731338,1.5769572,1.3241913,1.0336993,0.76207024,0.65643674,0.68661773,0.8186596,1.0110635,1.20724,1.1996948,0.9997456,0.73566186,0.65643674,1.1204696,1.5128226,1.720317,1.7089992,1.539231,1.6675003,2.252257,2.7992878,2.9803739,2.6446102,2.2258487,2.0108092,1.9693103,2.0108092,1.9768555,1.7693611,1.4411428,1.1317875,0.90543,0.76207024,0.59230214,0.56589377,0.7092535,0.90920264,0.8903395,0.8563859,0.65643674,0.43385187,0.2565385,0.13204187,0.071679875,0.060362,0.06790725,0.0754525,0.071679875,0.07922512,0.090543,0.1056335,0.11317875,0.10940613,0.14335975,0.3169005,0.60362,0.9808825,1.4600059,2.04099,2.516341,3.127506,3.651901,3.399135,2.0372176,1.2638294,1.1129243,1.8070874,3.7537618,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0150905,0.08299775,0.23013012,0.45648763,0.42630664,0.331991,0.27917424,0.27917424,0.27917424,0.26408374,0.362172,0.543258,0.754525,0.95447415,0.87902164,0.59230214,0.36971724,0.3169005,0.3734899,0.573439,0.87902164,1.2826926,1.7089992,1.9957186,2.263575,2.927557,3.651901,4.2027044,4.466788,4.6290107,4.9044123,5.1835866,5.4212623,5.6589375,5.9418845,6.3342376,6.809588,7.3981175,8.194141,8.993938,9.748463,10.27663,10.559577,10.736891,11.208468,11.615912,11.864905,11.989402,12.151625,12.30253,12.272349,12.298758,12.46098,12.672247,12.96274,13.370183,13.86817,14.317112,14.441608,14.324657,14.143571,14.060574,14.166207,14.456699,14.667966,14.705692,14.747191,14.890551,15.165953,15.769572,17.184307,19.051756,20.432537,19.817598,18.651857,17.48989,16.418465,15.528125,14.909414,14.245432,13.321139,12.113899,10.895341,10.246449,10.012547,10.638803,11.649866,12.985375,14.999957,17.840744,20.930523,23.514772,25.163408,25.75571,22.639523,19.806282,17.282394,15.328176,14.426518,13.588995,12.23085,11.189606,10.782163,10.819888,8.903395,6.700182,4.4139714,2.41448,1.237421,0.80356914,0.7167987,0.7884786,0.91674787,1.0902886,1.2940104,1.4675511,1.2826926,0.7997965,0.45648763,0.43007925,0.543258,0.7582976,0.9620194,0.97333723,0.875249,0.70170826,0.48666862,0.2565385,0.030181,0.018863125,0.02263575,0.02263575,0.0150905,0.00754525,0.011317875,0.018863125,0.0452715,0.09808825,0.20372175,0.18863125,0.1358145,0.08299775,0.041498873,0.0,0.0,0.0,0.0,0.02263575,0.10940613,0.14713238,0.10186087,0.041498873,0.011317875,0.011317875,0.003772625,0.0,0.0,0.0,0.0,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0,0.011317875,0.011317875,0.003772625,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.011317875,0.0,0.0,0.00754525,0.018863125,0.033953626,0.06413463,0.06790725,0.0754525,0.07922512,0.0754525,0.071679875,0.05281675,0.03772625,0.026408374,0.030181,0.041498873,0.071679875,0.071679875,0.060362,0.049044125,0.056589376,0.041498873,0.033953626,0.030181,0.033953626,0.041498873,0.033953626,0.0452715,0.060362,0.06790725,0.056589376,0.056589376,0.08677038,0.15467763,0.26031113,0.3772625,0.56212115,0.7884786,0.965792,1.0035182,0.8111144,0.69793564,0.77338815,1.1808317,1.8900851,2.7087448,2.969056,2.9728284,2.6710186,2.191895,1.841041,1.7731338,2.0183544,2.305074,2.6974268,3.5764484,4.5196047,4.678055,4.466788,4.274384,4.466788,4.9723196,5.4288073,5.7004366,5.6287565,5.028909,5.1345425,6.436098,7.748972,8.096053,6.692637,5.832478,5.6778007,5.66271,5.2137675,3.7462165,2.4371157,3.0407357,4.666737,6.760544,9.152389,8.526133,7.0812173,6.255012,6.092789,5.2288585,3.4255435,3.7801702,4.9157305,5.8626595,6.0512905,5.6853456,4.7421894,4.1008434,4.0782075,4.406426,4.478106,4.436607,4.217795,3.8593953,3.5047686,3.187868,4.1272516,5.300538,5.938112,5.523123,5.311856,4.395108,2.957738,1.5656394,1.1431054,1.6675003,2.535204,3.3953626,4.1574326,4.991183,4.8930945,4.4403796,3.9084394,3.3651814,2.6597006,1.3317367,1.5845025,3.361409,5.3986263,5.2062225,4.587512,4.06689,3.4330888,2.7087448,2.1466236,2.2711203,2.9539654,3.640583,3.7914882,2.8822856,1.6561824,2.4408884,3.9159849,5.198677,5.855114,5.8211603,5.342037,4.4215164,3.2369123,2.11267,1.9693103,2.191895,2.2711203,2.082489,1.9240388,2.0296721,2.3201644,2.7540162,3.270866,3.8103511,3.2218218,2.4484336,1.7354075,1.2562841,1.0978339,1.056335,0.9016574,0.8111144,0.90920264,1.2487389,1.6939086,2.0598533,2.1088974,1.8485862,1.5241405,1.056335,0.8224323,0.7205714,0.6752999,0.63002837,0.56212115,0.49421388,0.482896,0.5357128,0.63002837,0.7922512,0.91674787,0.9695646,0.9695646,0.9620194,0.965792,0.9808825,1.0072908,1.026154,0.98465514,0.8639311,0.76584285,0.7205714,0.7205714,0.7432071,0.7507524,0.7394345,0.7092535,0.6790725,0.694163,0.7205714,0.7582976,0.8111144,0.875249,0.965792,0.9997456,0.98465514,0.91297525,0.784706,0.63002837,0.5281675,0.47535074,0.43007925,0.35462674,0.22258487,0.1659955,0.124496624,0.14335975,0.18863125,0.18485862,0.20749438,0.5281675,0.9997456,1.4449154,1.6486372,1.7731338,1.7844516,1.6033657,1.2713746,0.95447415,0.69039035,0.7167987,1.0336993,1.5316857,1.9730829,2.384299,2.7351532,2.938875,2.957738,2.776652,2.6408374,2.463524,2.1768045,1.7731338,1.3166461,1.056335,1.086516,1.2411937,1.4637785,1.8070874,1.9806281,1.9693103,1.7769064,1.5203679,1.4449154,1.7769064,1.9994912,2.0787163,1.9957186,1.7580433,1.8485862,2.5087957,2.9728284,2.8521044,2.1692593,1.780679,1.5618668,1.5845025,1.7542707,1.8184053,1.720317,1.4260522,1.1053791,0.8639311,0.7696155,0.6451189,0.7922512,1.1883769,1.4449154,0.80734175,0.452715,0.38103512,0.36971724,0.31312788,0.20749438,0.1358145,0.13204187,0.13958712,0.1358145,0.120724,0.14335975,0.181086,0.211267,0.21503963,0.18863125,0.15845025,0.24899325,0.452715,0.8526133,1.6260014,2.516341,3.5085413,4.7006907,5.587258,5.0477724,3.1161883,1.9278114,1.448688,1.9353566,3.9197574,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.071679875,0.21503963,0.33576363,0.3734899,0.362172,0.331991,0.29426476,0.24522063,0.20749438,0.24522063,0.35462674,0.5281675,0.7469798,0.663982,0.58475685,0.52062225,0.47157812,0.45648763,0.49421388,0.6413463,0.80734175,0.935611,1.0072908,1.4109617,1.9504471,2.516341,3.0256453,3.4179983,3.440634,3.6028569,3.8669407,4.191386,4.5460134,4.8025517,4.859141,4.979865,5.2779026,5.692891,6.375736,7.0057645,7.4735703,7.7716074,7.964011,8.088508,8.458225,8.922258,9.367428,9.737145,9.906913,9.97482,10.495442,11.465008,12.344029,12.528888,12.728837,12.955194,12.902377,11.962994,11.034928,10.518079,10.676529,11.6008215,13.200415,15.128226,16.7995,17.659658,17.497435,16.448645,14.373701,15.01882,16.659912,18.025602,18.278368,18.414183,18.485863,18.131235,17.425755,16.874952,17.753973,17.369165,15.7657995,13.702174,12.664702,12.113899,12.408164,12.438345,11.668729,10.11818,10.948157,12.355347,14.826416,17.674747,19.04421,18.346275,17.569115,16.720274,15.720529,14.388792,13.422999,12.789199,12.46098,12.306303,12.098808,11.0613365,9.367428,6.94163,4.304565,2.5314314,1.2261031,0.87147635,1.0186088,1.4562333,2.2107582,2.848332,3.2520027,2.6483827,1.2864652,0.44139713,0.4678055,0.52062225,0.59230214,0.7054809,0.9016574,0.935611,0.8262049,0.6073926,0.32444575,0.030181,0.018863125,0.0150905,0.0150905,0.018863125,0.030181,0.056589376,0.060362,0.1358145,0.32821837,0.65643674,0.48666862,0.1961765,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.011317875,0.00754525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.0150905,0.0150905,0.003772625,0.0,0.0,0.0,0.0,0.0,0.0,0.00754525,0.011317875,0.0,0.011317875,0.02263575,0.02263575,0.011317875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.003772625,0.0150905,0.041498873,0.071679875,0.10940613,0.1358145,0.120724,0.071679875,0.033953626,0.0150905,0.018863125,0.030181,0.07922512,0.090543,0.07922512,0.056589376,0.0452715,0.02263575,0.0150905,0.02263575,0.030181,0.030181,0.041498873,0.03772625,0.03772625,0.0452715,0.0452715,0.0452715,0.071679875,0.1056335,0.120724,0.120724,0.2678564,0.5055317,0.55457586,0.3961256,0.27540162,0.3470815,0.58475685,0.9507015,1.4600059,2.1805773,2.7691069,2.9313297,2.7615614,2.3163917,1.6335466,1.7919968,1.8863125,1.6675003,1.539231,2.565385,4.881777,4.859141,3.9725742,3.270866,3.3576362,3.6858547,4.172523,4.6554193,5.089271,5.553304,6.126743,8.322411,12.038446,14.6151495,10.819888,6.326692,4.406426,3.4557245,2.6710186,2.0598533,2.7426984,3.482133,3.8556228,4.2328854,5.783434,8.89585,9.242931,8.201687,6.458734,4.044254,4.2630663,6.5530496,8.175279,8.296002,7.9791017,7.564113,6.647365,5.1835866,3.6368105,2.9916916,2.806833,3.3840446,3.9461658,4.093298,3.7990334,2.9464202,2.2447119,2.8143783,4.4743333,5.7683434,6.477597,5.251494,3.169005,1.4750963,1.5731846,3.1576872,6.145606,8.231868,8.699674,8.409182,6.356873,4.772371,3.7763977,3.0860074,1.9994912,0.935611,1.3204187,2.5427492,4.353609,6.8661776,7.586749,7.6923823,6.307829,3.8556228,2.0749438,1.5731846,1.9164935,2.686109,3.199186,2.5012503,2.625747,3.6896272,4.617693,5.0138187,5.172269,5.587258,5.6363015,5.172269,4.3196554,3.4783602,2.7087448,3.0218725,3.4066803,3.2670932,2.4107075,2.0183544,1.7769064,1.8146327,2.0787163,2.335255,2.565385,2.2673476,1.6373192,0.98842776,0.73188925,0.56212115,0.5357128,0.73188925,1.1393328,1.6637276,1.8448136,1.8448136,1.5769572,1.1808317,1.0223814,1.0336993,1.146878,1.2525115,1.267602,1.1431054,0.9507015,0.7167987,0.5998474,0.6187105,0.65643674,0.72811663,0.7582976,0.76207024,0.77716076,0.83752275,0.91297525,1.0035182,1.0902886,1.1581959,1.20724,1.0336993,0.88279426,0.76584285,0.694163,0.65643674,0.65643674,0.65643674,0.6488915,0.63002837,0.59607476,0.63002837,0.694163,0.80734175,0.9507015,1.0978339,1.2713746,1.3505998,1.3505998,1.2525115,1.0223814,0.80356914,0.6111652,0.452715,0.32067314,0.19994913,0.24899325,0.2867195,0.29803738,0.27917424,0.24522063,0.21881226,0.7167987,1.418507,2.161714,2.9313297,3.7462165,4.5912848,4.3913355,3.1161883,1.7844516,1.0525624,0.62248313,0.452715,0.52062225,0.83752275,1.1317875,1.2713746,1.569412,2.1654868,3.0218725,3.0709167,2.9916916,2.7691069,2.4974778,2.3654358,2.3880715,2.3956168,2.4371157,2.6106565,3.0520537,3.138824,2.9954643,2.8596497,2.8106055,2.7615614,2.565385,2.2786655,1.8900851,1.6373192,2.0145817,2.5616124,3.1124156,3.31991,3.0105548,2.1805773,1.841041,1.599593,1.4939595,1.478869,1.4034165,1.3053282,1.1091517,0.88279426,0.73188925,0.7922512,0.7092535,0.48666862,0.31312788,0.26031113,0.26031113,0.43007925,0.482896,0.4074435,0.2678564,0.18485862,0.10940613,0.12826926,0.17731337,0.21881226,0.24522063,0.3055826,0.36594462,0.41498876,0.43385187,0.3961256,0.2867195,0.27917424,0.41876137,1.1016065,3.0671442,4.2517486,4.6554193,4.29702,3.361409,2.2296214,1.9466745,1.6373192,1.3015556,1.418507,2.9464202;
 } 
