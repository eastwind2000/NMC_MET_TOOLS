netcdf QPE_CPC_CMORPH.2018062900{
dimensions: 
 lat = 180; 
 lon = 281; 
variables:  
float lat(lat) ; 
   lat:long_name = "latitude" ;
   lat:units = "degrees_north" ;
   lat:standard_name = "latitude" ;
float lon(lon) ;
   lon:long_name = "longitude" ;
   lon:units = "degrees_east" ;
   lon:standard_name = "longitude" ;
float APCP_24(lat, lon) ;
   APCP_24:name = "APCP_24" ;
   APCP_24:long_name = "Total Precipitation" ;
   APCP_24:level = "A24" ;
   APCP_24:units = "kg/m^2" ;
   APCP_24:_FillValue = -9999.f ;
   APCP_24:init_time = "20180628_000000" ;
   APCP_24:init_time_ut = "1530144000.0" ;
   APCP_24:valid_time = "20180629_000000" ;
   APCP_24:valid_time_ut = "1530230400.0" ;
   APCP_24:accum_time = "240000" ;
   APCP_24:_FillValue = -9.99e8 ;
   APCP_24:accum_time_sec = 86400 ;
 // global attributes: 
 :_NCProperties = "version=1|netcdflibversion=4.4.1.1|hdf5libversion=1.8.12" ;
	:FileOrigins = "CPC_CMORPH_DAILY_PRCP" ; 
	:MET_version = "V7.0" ;
	:Projection = "LatLon" ;
	:lat_ll = "15.125 degrees_north" ; 
	:lon_ll = "70.125 degrees_east" ; 
	:delta_lat = "0.250000 degrees" ;
	:delta_lon = "0.250000 degrees" ;
	:Nlat = "180 grid_points" ; 
	:Nlon = "281 grid_points" ; 
data:
lat = 15.125,15.375,15.625,15.875,16.125,16.375,16.625,16.875,17.125,17.375,17.625,17.875,18.125,18.375,18.625,18.875,19.125,19.375,19.625,19.875,20.125,20.375,20.625,20.875,21.125,21.375,21.625,21.875,22.125,22.375,22.625,22.875,23.125,23.375,23.625,23.875,24.125,24.375,24.625,24.875,25.125,25.375,25.625,25.875,26.125,26.375,26.625,26.875,27.125,27.375,27.625,27.875,28.125,28.375,28.625,28.875,29.125,29.375,29.625,29.875,30.125,30.375,30.625,30.875,31.125,31.375,31.625,31.875,32.125,32.375,32.625,32.875,33.125,33.375,33.625,33.875,34.125,34.375,34.625,34.875,35.125,35.375,35.625,35.875,36.125,36.375,36.625,36.875,37.125,37.375,37.625,37.875,38.125,38.375,38.625,38.875,39.125,39.375,39.625,39.875,40.125,40.375,40.625,40.875,41.125,41.375,41.625,41.875,42.125,42.375,42.625,42.875,43.125,43.375,43.625,43.875,44.125,44.375,44.625,44.875,45.125,45.375,45.625,45.875,46.125,46.375,46.625,46.875,47.125,47.375,47.625,47.875,48.125,48.375,48.625,48.875,49.125,49.375,49.625,49.875,50.125,50.375,50.625,50.875,51.125,51.375,51.625,51.875,52.125,52.375,52.625,52.875,53.125,53.375,53.625,53.875,54.125,54.375,54.625,54.875,55.125,55.375,55.625,55.875,56.125,56.375,56.625,56.875,57.125,57.375,57.625,57.875,58.125,58.375,58.625,58.875,59.125,59.375,59.625,59.875;
lon = 70.125,70.375,70.625,70.875,71.125,71.375,71.625,71.875,72.125,72.375,72.625,72.875,73.125,73.375,73.625,73.875,74.125,74.375,74.625,74.875,75.125,75.375,75.625,75.875,76.125,76.375,76.625,76.875,77.125,77.375,77.625,77.875,78.125,78.375,78.625,78.875,79.125,79.375,79.625,79.875,80.125,80.375,80.625,80.875,81.125,81.375,81.625,81.875,82.125,82.375,82.625,82.875,83.125,83.375,83.625,83.875,84.125,84.375,84.625,84.875,85.125,85.375,85.625,85.875,86.125,86.375,86.625,86.875,87.125,87.375,87.625,87.875,88.125,88.375,88.625,88.875,89.125,89.375,89.625,89.875,90.125,90.375,90.625,90.875,91.125,91.375,91.625,91.875,92.125,92.375,92.625,92.875,93.125,93.375,93.625,93.875,94.125,94.375,94.625,94.875,95.125,95.375,95.625,95.875,96.125,96.375,96.625,96.875,97.125,97.375,97.625,97.875,98.125,98.375,98.625,98.875,99.125,99.375,99.625,99.875,100.125,100.375,100.625,100.875,101.125,101.375,101.625,101.875,102.125,102.375,102.625,102.875,103.125,103.375,103.625,103.875,104.125,104.375,104.625,104.875,105.125,105.375,105.625,105.875,106.125,106.375,106.625,106.875,107.125,107.375,107.625,107.875,108.125,108.375,108.625,108.875,109.125,109.375,109.625,109.875,110.125,110.375,110.625,110.875,111.125,111.375,111.625,111.875,112.125,112.375,112.625,112.875,113.125,113.375,113.625,113.875,114.125,114.375,114.625,114.875,115.125,115.375,115.625,115.875,116.125,116.375,116.625,116.875,117.125,117.375,117.625,117.875,118.125,118.375,118.625,118.875,119.125,119.375,119.625,119.875,120.125,120.375,120.625,120.875,121.125,121.375,121.625,121.875,122.125,122.375,122.625,122.875,123.125,123.375,123.625,123.875,124.125,124.375,124.625,124.875,125.125,125.375,125.625,125.875,126.125,126.375,126.625,126.875,127.125,127.375,127.625,127.875,128.125,128.375,128.625,128.875,129.125,129.375,129.625,129.875,130.125,130.375,130.625,130.875,131.125,131.375,131.625,131.875,132.125,132.375,132.625,132.875,133.125,133.375,133.625,133.875,134.125,134.375,134.625,134.875,135.125,135.375,135.625,135.875,136.125,136.375,136.625,136.875,137.125,137.375,137.625,137.875,138.125,138.375,138.625,138.875,139.125,139.375,139.625,139.875,140.125;
APCP_24 = 0.425,0.42222226,0.3,0.13333334,0.18888889,0.15833333,0.16666667,0.3,0.37777776,0.6333333,1.2333333,2.1222222,2.966667,2.977778,4.433334,5.511111,11.750001,13.611112,9.966666,4.658334,3.0222223,2.1916666,1.9222221,1.2083334,0.73333335,0.4888889,0.058333337,0.022222223,0.19166666,0.08888889,0.14166667,0.25555557,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.56666666,2.3333335,5.775,9.2,12.07778,15.866667,22.855553,20.091665,17.577778,14.141667,9.344444,7.35,8.833334,8.900001,8.700001,6.7999997,5.233333,3.8111115,2.6583333,2.0222223,1.1666666,1.6166668,8.488889,16.941668,21.333332,16.975,13.422222,15.666667,20.811113,20.744444,22.916666,25.255556,23.083332,17.08889,11.4,5.211111,2.2,0.34166667,0.6888889,0.80833334,0.65555555,2.1416667,5.055556,8.211111,12.049999,14.355555,14.75,14.400001,15.433332,17.188889,21.541668,27.622223,30.422224,28.941666,27.555555,26.366667,20.111113,15.625,14.144445,10.277779,8.533334,8.344444,11.375,17.6,22.375,16.4,8.025001,6.7666674,7.711111,2.7416666,2.0111113,7.6250005,8.555556,16.199999,37.044445,60.300003,58.091667,24.855558,4.2083335,5.8333335,5.475,15.188888,23.311111,22.858334,16.98889,11.125,7.7888894,7.3083334,13.633334,5.6916666,2.688889,0.0,0.0,0.13333334,1.3000001,0.0,0.0,0.0,0.0,0.0,0.0,0.20833333,0.5777778,0.44166666,0.9555557,2.4916668,13.655556,14.166666,12.316668,8.288889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333334,0.20000002,0.20000003,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38888887,0.6083333,0.39999998,0.29999998,0.6555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.14444445,0.1888889,0.37500003,0.36666667,0.18333334,0.033333335,1.1833334,4.5444446,7.9888887,11.416667,16.166668,22.2,30.611113,34.758335,33.622227,34.675003,32.766666,25.844446,21.441666,22.288889,24.575,26.366667,33.800003,28.444445,29.88889,38.683334,41.9,28.858334,32.41111,32.608334,28.88889,18.591667,7.9444447,2.4333334,1.2083334,0.26666668,0.49166673,0.31111112,0.008333334,0.37777779,0.5,0.05,0.044444446,0.175,0.41111112,0.39166668,0.17777778,0.0,0.0,0.0,0.0,0.0,0.0,0.9166667,0.67777777,0.72222227,0.35833332,0.2888889,0.3416667,0.43333334,0.85833335,1.4888887,2.4222221,3.5833335,4.711111,6.5666666,8.177778,10.849999,13.555557,17.275,13.755555,8.311111,2.05,1.0222223,0.6333333,0.5,0.3,0.18888888,0.33333334,0.20833334,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.2,0.14166668,0.24444443,2.5583332,5.588889,7.491667,9.822222,11.122223,14.525002,27.21111,28.283335,27.233332,23.075,15.944447,11.508333,11.877779,12.1,10.25,7.7555556,5.75,4.4,3.6,2.8666666,1.4000002,0.9166667,2.988889,9.55,16.544445,21.15,19.2,23.883335,27.933334,29.544445,31.383335,28.944447,26.80833,19.088888,11.8,5.9777775,2.5444446,0.6583333,2.0666666,2.0583334,1.7111111,2.025,3.3666666,5.0666666,8.341667,11.455555,14.408333,16.766668,22.858334,28.555557,33.433334,40.5,45.31111,39.649998,36.066666,31.108334,32.444447,27.058334,28.02222,22.68889,11.566667,8.244445,9.075,14.377779,23.90833,20.33333,7.233333,6.7222223,8.966667,3.75,2.8111112,6.3750005,12.433332,8.541666,9.388888,15.933334,37.141666,19.833334,0.7666667,6.266667,7.825001,4.588889,10.644445,16.0,14.688889,8.116667,4.288889,1.3083334,2.9666667,1.1,0.6111111,0.0,0.0,0.0,0.0,0.0,2.7,4.0111113,3.911111,1.0500001,0.06666667,0.13333334,0.51111114,1.2666667,2.0333333,2.6333337,8.255555,11.055555,8.408334,2.1888888,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.20000002,0.116666675,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.55,4.4666667,4.533334,3.825,2.8333335,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0333333,0.0,0.0,0.0,0.75000006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.53333336,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.18888889,0.23333335,1.1500001,2.5,1.55,0.48888892,0.9000001,4.3777776,8.766666,14.933332,11.555555,13.600001,24.6,33.7,29.98889,30.158333,25.722223,22.633333,21.6,23.577778,28.591667,26.711111,25.908333,24.344444,35.777782,39.416664,61.100006,43.65,29.466667,30.283333,31.488892,26.941666,13.588888,7.1111116,4.491667,2.4222221,1.1583334,0.24444446,0.075,0.5,0.31111112,0.0,0.24444444,0.4166667,0.6888889,0.18333334,0.05555556,0.055555556,0.0,0.0,0.0,0.0,0.0,0.38750002,0.43333334,0.65,0.625,0.64166665,0.7625,1.075,1.7375,3.0083334,3.8583333,5.4000006,6.708333,8.500001,12.233334,16.31875,17.041668,14.600001,8.700002,4.0083337,1.1999999,0.5666667,0.325,0.225,0.20000002,0.13333333,0.09166667,0.06250001,0.008333334,0.0,0.016666668,0.1625,0.15,0.0125,0.008333334,0.16666667,0.28750002,0.2916667,0.25,0.35833335,0.6125001,1.3083334,2.0249999,1.7000002,1.1333333,3.9875,8.866667,13.05625,13.833334,15.125001,14.818749,20.675003,24.856249,29.675001,35.425,30.133331,21.756252,20.558336,18.775,13.337501,11.341667,8.675,6.958333,4.8375,3.341667,2.4916668,1.8,2.475,4.50625,9.008333,14.375,17.666666,20.981253,29.483335,36.166668,32.36875,30.283333,25.599998,21.183332,11.3875,4.6,1.8999999,0.37500003,1.1083335,2.4250002,3.5,2.9499998,2.1083336,2.4166667,3.3937502,6.9000006,11.66875,18.383335,26.537502,36.16667,44.8375,53.741673,58.524998,66.11875,66.09167,67.524994,69.325005,33.43125,30.683332,35.05,18.7625,8.783334,7.6875005,7.7749996,13.156252,24.391668,10.8875,8.400001,12.891666,8.44375,2.9,3.8249998,8.108334,13.243751,9.433333,5.1666665,1.3750001,0.36666667,0.99375,3.2,4.88125,3.441667,3.1583335,7.5,9.291668,5.3000007,2.8083334,0.75625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30624998,2.2083335,2.658333,0.96874994,0.20833333,0.31875002,0.008333334,0.65625,1.7416668,5.1187496,8.575,2.108333,0.10625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,2.86875,9.924999,10.674999,8.79375,4.6000004,0.52500004,0.2916667,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.16875,0.0,0.0,0.75000006,2.53125,0.0,0.0,0.0,0.0,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.18750001,0.6,0.23750001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.056250006,0.075,0.23333335,0.975,2.775,4.81875,2.8833334,1.7624999,3.8333333,9.3,11.0625,11.2,13.700001,21.008333,26.825,28.2,24.206251,25.958336,21.3,18.262503,19.341667,25.312502,32.24167,38.949997,41.883335,58.241665,74.80001,63.183334,53.0625,36.75,29.34375,38.791668,42.9125,22.85,18.275,8.95625,4.0833335,2.1125002,0.625,1.30625,1.6416668,1.4416667,1.09375,1.0416666,1.6625,1.8166667,0.26875,0.15000002,0.13333334,0.0,0.0,0.0,0.0,0.0,1.4000001,1.8888888,2.2666667,2.391667,2.2666667,1.9333334,1.488889,1.3750001,1.6333334,1.8555557,2.3249998,2.8111112,3.5166664,5.066667,7.233334,9.188889,7.9166665,3.8999999,2.888889,2.4333336,1.6777778,0.49999997,0.3222222,0.16666667,0.17777778,0.08888889,0.05,0.022222223,0.0,0.14444445,0.21666667,0.08888889,0.033333335,0.08888889,0.44444448,0.16666669,0.033333335,0.08333334,0.1,0.25833336,0.9777778,2.8777778,5.15,4.233333,5.075,9.466667,7.708333,8.122223,10.722223,13.033335,17.222223,23.591667,31.499998,42.375,51.011112,51.56667,36.511112,32.944447,26.633333,21.922222,15.408334,9.433334,6.4249997,4.3777776,3.3,3.225,2.7444446,3.6916661,5.0333333,8.741667,13.222223,17.308334,25.61111,28.966665,28.975,22.533333,16.108334,13.166666,10.349999,5.7111115,3.8111112,2.1083333,0.9888889,2.0916667,3.6555557,3.825,2.411111,3.1555555,3.6333332,5.1777773,6.575001,10.9,19.741667,31.833334,48.733337,67.68889,79.77778,91.12501,88.26666,84.6,64.63334,30.891665,30.855553,28.877775,18.758333,8.222222,6.2583337,5.1222224,4.908334,9.166667,5.416667,10.377778,21.07778,23.525002,13.0,6.1666665,7.511111,11.575002,11.244446,5.5,0.475,0.011111111,0.09166667,1.3222222,1.0916667,0.95555556,1.9,2.7333333,4.2,0.9166666,1.4444444,2.366667,1.4666667,1.0416666,0.0,0.0,0.99999994,0.22222222,0.24166667,0.13333334,0.25,0.50000006,0.0,0.0,0.5777778,0.9416667,0.42222223,1.375,2.6666667,10.608334,15.866667,1.3333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.70000005,2.1222224,10.583334,21.455557,18.377779,9.966667,1.7222223,0.5666667,0.40000004,0.15000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7166667,4.9,0.0,0.0,0.0,0.0,0.26666668,0.4666667,0.044444446,0.075,0.1,0.044444446,0.06666667,0.055555556,0.025,0.022222223,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.033333335,0.075,0.18888889,0.35555553,0.8000001,1.6333334,4.5833335,4.7,4.3,7.377778,11.722222,19.133333,18.244444,18.766666,24.333334,27.491669,32.86667,32.408333,25.755556,28.166666,21.125,19.322224,21.283335,28.577778,36.625,35.211113,40.65556,39.11667,51.144447,47.508335,32.88889,23.95,35.477776,49.766666,30.300001,25.411112,15.108334,6.3111115,2.141667,0.9333333,3.0916667,6.8,7.9,4.3333335,2.7555556,3.225,3.0777779,0.94166666,0.48888886,0.5,0.016666668,0.0,0.0,0.033333335,0.1,1.3625,1.5416667,1.7,1.7625,1.8916667,1.6000001,1.1916668,1.0875,0.90833336,0.9833334,1.125,1.3166667,1.7562499,3.175,4.3562503,4.0833335,3.0812502,0.8083333,0.3666667,0.41874996,0.3916667,0.0375,0.0,0.0,0.10833333,0.14166667,0.0375,0.0,0.0,0.23333335,0.55625004,0.2,0.59999996,0.5666667,0.35000002,0.29375002,0.19166666,0.20625001,0.058333337,0.0375,0.3916667,1.2583334,3.28125,5.25,7.56875,11.733334,12.425,12.058332,11.841667,12.625001,14.441668,13.862499,15.966667,25.175001,32.016666,34.668747,35.408333,36.325,35.850002,32.325,22.85,13.466666,8.1625,4.408334,3.275,3.4,3.0333333,2.7625,2.3000002,5.4187503,11.050001,16.224998,26.458334,32.6,28.39375,19.833332,11.543749,7.208334,6.0937505,5.1333337,4.991667,5.29375,5.3083334,5.6062503,8.558333,9.418751,7.025,5.8083334,5.33125,8.308333,12.418751,17.141666,27.412502,41.566666,52.80625,58.875,75.23334,94.85625,88.89166,66.793755,42.575,23.78125,9.958333,8.058333,5.1375,3.5833335,4.9375,4.8500004,3.8625,1.0999999,0.6812501,4.3,15.766667,34.4125,38.841667,27.925001,14.508334,11.618752,8.641666,5.7083335,2.4812498,0.1,0.0,0.40833336,0.075,0.21666667,0.15,0.9437499,1.9166666,0.49375004,0.3166667,0.63125,0.083333336,0.0,0.0,0.0,0.25,0.1,0.61249995,0.27499998,1.31875,0.0,0.0,0.0,1.0833333,2.79375,5.7166667,13.025,17.316668,12.031251,5.6583333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.76875,3.8333333,16.35625,24.033335,14.9833355,7.61875,2.7583334,1.84375,4.475,1.0875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8000001,0.8000001,0.52500004,0.46666673,0.21666667,0.10000001,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,0.09166667,0.081250004,0.13333334,0.26666668,0.7375001,1.7249999,3.2562501,4.9416666,7.25625,14.791667,24.058332,28.887505,29.8,35.15625,41.475,42.799995,45.733337,47.768753,45.89167,47.38333,34.231255,22.083334,23.45,29.708334,29.743752,28.45,22.658335,18.525,26.258333,33.46875,29.475,32.143753,34.216667,47.4625,36.233334,31.266668,19.575,10.491667,2.2,0.93333334,0.725,6.541667,7.5250006,2.8875,5.0833335,4.6,2.3916664,1.675,1.075,0.76666677,0.0125,0.0,0.00625,0.20833333,1.13125,0.10000001,0.044444446,0.033333335,0.25833336,0.8888889,1.1416665,1.0333333,0.85833347,0.56666666,0.36666667,0.27500004,0.18888889,0.16666667,0.4,0.81666666,0.47777778,0.041666668,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36666667,0.60833335,0.06666667,0.46666667,0.2,0.0,0.016666668,0.022222223,0.016666668,0.011111111,0.0,0.15555556,1.3666667,2.9750004,5.177778,6.916666,8.311112,11.108334,14.466667,17.966667,17.233334,11.88889,12.066668,14.9,16.541666,23.200003,27.816668,27.733334,26.822224,26.508335,26.822222,23.875,19.133333,14.916666,6.933334,4.0444446,2.9750004,3.1666665,3.2833335,2.5666666,2.8166666,5.8333335,12.258333,23.47778,28.944447,24.600002,19.311111,12.825001,6.844445,4.491667,3.7000005,4.077778,5.6166663,8.0222225,10.133333,16.333332,18.641666,15.533335,13.444445,11.025001,12.044443,16.233334,22.733334,35.783333,46.98889,44.025,35.11111,35.18889,41.933334,42.011112,34.791668,27.322222,18.175001,9.711111,5.8111115,1.25,0.24444446,1.5500001,4.1777773,3.5416667,0.13333334,0.8166666,7.644444,17.233335,21.775,41.044445,51.533337,36.61111,20.766668,7.611111,4.4888887,1.2833332,0.51111114,0.0,0.0,0.0,0.19999999,0.26666665,0.075,0.32222223,1.0916667,0.3111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.56666666,1.1555555,4.4583335,3.488889,0.0,0.0,0.17777778,0.8333333,5.644445,16.833332,21.255556,13.058333,1.8222221,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,1.2555557,9.416666,22.5,25.877779,10.791667,16.177778,8.941667,14.044445,1.7666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,0.82222223,0.6,0.36666667,0.31111112,0.16666667,0.06666667,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.31111112,0.36666667,0.23333335,0.36666667,0.9666667,2.0555556,4.075,6.6000004,10.408335,19.1,33.555553,45.108334,42.666668,47.716667,55.9,61.091667,61.666668,59.775,56.644447,56.933334,45.533333,29.355556,21.658333,30.688889,40.691666,33.333332,30.422222,16.425,16.966665,27.166668,32.655556,56.233337,74.03334,67.78333,55.57778,55.211113,31.875004,20.077778,5.2833333,1.7444446,0.90000004,3.3111112,2.288889,0.26666665,3.5222223,4.825,3.0333333,3.6833334,2.522222,0.88888896,0.016666668,0.0,0.008333334,0.4222222,2.0083334,0.2875,0.48333335,0.52500004,0.5375,0.95,1.08125,1.3416667,1.39375,1.1999999,1.2750001,0.78125006,0.9250001,1.1125,1.925,2.875,3.0416667,2.1625001,1.6166666,0.9500001,0.6375,0.39999998,0.49375,0.375,0.25000003,0.24166669,0.64166665,0.64374995,0.05,0.0,0.0,0.0,0.083333336,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.375,1.0833334,1.9666666,4.1625,6.108333,7.8750005,9.433332,9.84375,10.833334,13.041666,15.468749,15.225001,13.7375,15.416667,17.425001,19.516668,22.3125,23.041666,22.875,23.225,25.35,24.712502,20.574999,17.85625,9.725,5.9333334,3.5687501,2.266667,2.3750002,2.4166665,2.7125003,4.441667,8.5,16.908333,21.733334,20.59375,16.5,10.6875,5.2750006,2.4312499,1.5749999,1.2666668,0.73125005,2.3,6.1500006,12.175001,17.312502,16.933334,15.425001,13.84375,12.741667,15.756249,22.983334,27.5375,29.516666,27.23125,21.166668,16.866667,14.8125,12.650001,9.975,11.766666,5.5,2.8166666,1.375,0.5187501,0.008333334,0.40625003,1.55,1.8874999,0.15,0.09375,2.1166668,11.883334,20.150002,19.241667,31.20625,43.466667,33.031254,13.183333,5.4583335,1.1187501,0.52500004,0.01875,0.16666667,0.12500001,0.26666668,0.6666666,0.0,0.0,0.10625,0.28333333,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.5375004,2.0416667,0.056250002,0.125,0.7875,0.26666665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.375,3.8875003,21.608334,24.666668,35.575,23.533333,11.387501,8.433334,1.65625,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108333334,0.45833334,0.10625,0.0,0.0,0.0,0.0,0.48333332,0.0,0.0,0.0,16.0875,0.9250001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.1875,0.275,0.46666667,1.0937502,2.7166667,5.0312495,8.283334,13.912499,22.775,37.233334,51.443756,60.008335,60.45,60.583336,62.449997,57.166664,59.9625,56.824997,51.274998,41.837498,40.85,31.056252,29.216667,38.6,42.350002,48.63333,25.125,16.15,34.09375,51.75,69.625,87.94167,67.193756,61.025,55.466667,34.44375,21.858334,6.8875,5.0166664,3.1062498,4.05,2.6166666,2.28125,3.1666665,3.7875,4.7833333,6.4937496,3.141667,0.5916667,0.0,0.0,0.0625,0.54166675,2.4750001,0.016666668,0.033333335,0.055555556,0.3333333,1.0444444,1.4083334,1.6111112,2.3500001,3.166667,3.5333335,3.8000004,4.933334,5.5916667,6.8444443,5.283334,2.3666668,1.2916667,0.67777777,0.3111111,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.45000002,0.28888887,0.15555556,0.033333335,0.08888889,0.5833334,0.96666664,1.9499999,3.3444445,5.333334,5.8500004,5.9555554,8.941668,12.577778,10.475,9.133333,12.088889,14.633335,14.944444,13.758332,13.911112,12.791667,16.033333,17.9,17.077778,15.622223,17.25,20.666668,18.941668,13.811111,13.283333,8.844445,6.666667,4.325,3.1555557,2.7250001,2.4555557,2.491667,2.9333334,5.183334,10.400001,15.766666,17.316668,15.533333,10.349999,5.8888893,2.6166668,1.2444444,0.51111114,0.22500002,0.73333335,2.441667,3.766667,6.283334,11.088889,11.944445,13.425,13.277778,19.349998,23.644447,27.858334,31.944447,33.458336,26.222221,14.422222,6.4333334,1.977778,0.6333334,0.14444445,0.033333335,0.35555553,0.3888889,0.0,0.0,0.016666668,0.5,0.33333334,0.0,0.0,0.033333335,1.3777778,12.416665,17.555557,13.333334,19.244448,28.283333,22.322224,18.133333,1.0,0.7777778,0.108333334,0.11111111,0.6,0.34444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.6166666,4.0111113,26.47778,52.099995,34.98889,7.9333334,11.111112,5.666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6111111,1.1111112,0.23333333,0.0,0.0,0.0,0.0,3.0,23.341667,5.3555555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.07777778,0.075,0.022222223,0.0,0.0,0.0,0.033333335,0.20000002,1.0416666,2.6111112,5.3500004,9.155557,17.025,28.91111,42.17778,59.425003,67.72222,72.84167,72.08889,61.93334,49.07778,45.183334,49.344448,46.955555,38.76667,40.81111,40.375,35.133335,31.741667,52.533337,64.14444,59.425,25.544445,27.191668,41.255554,59.775,61.56667,73.28334,64.48889,63.28889,46.933334,24.11111,11.641667,5.6000004,2.65,3.1,3.1444445,4.408334,5.2111115,5.508333,7.4666667,9.458334,2.3333335,0.22222222,0.0,0.0,0.033333335,0.8111111,3.0,0.0,0.033333335,0.17500001,0.7125,1.5916667,1.9437499,2.3166668,2.9125001,3.3083336,4.2999997,5.6875014,7.8083334,9.675001,10.741666,7.6000004,3.408333,1.48125,0.7083333,0.36666667,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8187501,2.4750001,2.7500002,4.1875,6.8,9.3,18.158335,18.631252,16.125002,13.083333,14.262501,16.983334,16.9375,22.733335,22.71875,16.358334,15.075001,15.025001,11.258333,9.26875,10.733335,11.606251,12.583334,12.031251,11.591667,10.783334,11.593752,14.091667,15.143751,11.95,9.8,8.7,7.1083336,5.33125,4.975,5.15625,3.3249998,1.84375,2.0916667,3.025,5.9583335,10.683334,10.975,9.916667,7.7625003,4.983333,3.0812502,2.0833335,1.4916668,0.7375001,0.26666668,0.23750001,0.425,3.1437502,7.0500007,9.291667,10.46875,11.025001,15.343751,22.566668,26.41875,31.833334,32.80625,23.408333,13.383333,6.3187504,2.6333332,0.84375006,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.86875004,0.84999996,0.025,0.0,0.016666668,1.2249999,6.3166666,14.031251,15.391666,9.912499,15.55,7.691667,0.45625004,1.5,1.3375,0.0,0.1,0.35000002,0.73333335,0.15625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108333334,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,2.2083335,11.466667,21.443748,27.2,12.762501,5.6666665,0.61875,0.0,0.025,1.3416667,1.0166668,0.09375,0.0,0.0,0.008333334,0.11875,0.775,1.0833334,0.46250004,0.0,0.15625,0.9916667,2.5750003,4.7,20.600002,2.8583336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.041666668,0.0,0.058333337,0.23125002,0.44166666,0.63750005,0.7333333,0.68125004,0.325,0.13333334,0.46250004,1.925,4.5875,9.225,18.649998,36.633335,55.48333,74.0875,85.66667,85.05,79.35,67.450005,51.025,37.293747,30.058334,31.583334,35.425003,34.958332,39.5,44.73333,53.725006,70.21666,70.65,59.437496,47.266666,32.8375,37.85,46.5625,45.61667,53.343754,70.51666,73.86667,51.55625,24.550001,12.95,4.3250003,0.92499995,1.0833333,2.2416666,4.0625,4.925,6.6499996,8.733334,6.875,1.4916668,0.008333334,0.0,0.28333333,0.825,1.3833333,2.625,0.38333333,0.2,0.2888889,0.45833337,1.0555556,1.1666667,1.0777777,0.9916668,0.78888893,0.9333334,1.0583333,1.1777779,2.1166666,2.6999998,1.5166669,0.73333335,0.33333337,0.24444446,0.11111112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05555556,0.65000004,2.5222223,3.0416665,1.9111111,2.5444448,5.9249997,7.822222,11.85,20.966665,21.041668,17.822222,18.7,20.0,21.1,19.316668,18.344444,19.4,19.044443,14.622223,10.516666,7.455556,4.4416666,5.9999995,7.9583335,11.222223,10.908334,7.5666666,8.488889,12.733335,14.822223,14.4416685,11.800001,10.391667,9.877778,9.088889,7.883333,7.3111115,8.141666,5.3,3.4,2.0555556,1.9250002,2.411111,6.0,8.6,6.111111,4.85,3.9222224,3.2250004,2.688889,2.766667,2.3000002,1.2777779,0.7166667,0.23333333,1.0,2.8444445,3.0555556,4.716666,5.777778,7.991667,14.300001,16.283333,15.611112,15.083334,15.577778,11.51111,6.6916666,3.0555556,2.6333332,2.188889,0.93333346,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.21666667,0.28888887,0.3,0.04166667,0.83333343,13.408333,25.755556,14.525001,5.033334,1.2444444,0.6333334,0.7222222,0.075,0.0,0.0,0.11111111,0.45555556,1.3666667,1.1444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,5.9333334,17.011112,15.808333,2.9,1.275,0.0,0.93333334,5.9222226,7.3222227,2.675,0.0,0.008333334,0.10000001,0.8583333,3.2999997,3.6888888,0.6,0.2777778,0.90833336,4.922222,2.55,3.2444446,5.366667,0.41111112,0.0,0.0,0.0,0.016666668,0.15555556,0.17500001,0.1,0.1,0.016666668,0.0,0.0,0.0,0.0,0.07777777,0.21111113,0.3333333,0.4888889,0.55833334,0.5888889,0.7416666,0.84444445,0.82500005,0.6666667,0.5222222,0.4166667,0.9555556,2.9916666,7.844445,22.875,47.044445,70.24445,86.51668,99.17778,99.48333,96.622215,81.433334,58.84444,42.58333,27.666666,23.966667,26.941668,31.455557,36.408333,41.066666,56.1,69.72222,70.51111,59.308334,47.366665,32.158333,26.300001,31.983334,36.822224,48.341667,83.288895,86.13333,59.466667,28.955555,15.5,4.8111115,2.6833334,4.022222,2.3444443,3.475,5.6555552,9.025,8.044445,3.9333334,0.8111111,0.0,0.0,0.32222223,1.5666666,3.0333333,5.2250004,0.0,0.0,0.011111111,0.26666665,0.8000001,1.1916667,1.3333333,1.1500001,0.9111112,0.9444445,0.93333334,1.1,0.6166667,0.43333334,0.24166669,0.17777778,0.083333336,0.044444446,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.6222222,1.6416667,5.0444446,11.3,13.877778,13.755555,18.791666,25.877777,20.016668,11.166668,10.275,11.255555,12.644445,13.408333,14.200001,14.55,15.644446,21.608332,20.911112,16.18889,12.908333,9.277778,7.0833335,7.5222225,6.825,5.3666673,5.8083334,6.4555554,8.133333,11.0,13.044446,15.5,14.933333,13.974999,11.755555,10.944445,11.508333,14.355555,17.341667,11.322223,7.066667,5.0222225,4.1000004,3.6111112,5.8444443,7.4,5.0,6.0,7.911111,8.416667,8.177778,7.822222,5.491667,3.8555558,1.9583333,0.9222222,0.9833334,1.4333334,2.3666668,4.55,7.5555553,7.7666664,10.255556,9.700001,8.066667,6.616667,7.0111113,5.6000004,3.575,2.3666666,5.05,5.388889,1.5583335,2.8444448,6.5888886,5.6583333,3.3555555,1.2083333,0.1,0.32500002,0.033333335,0.66666675,3.1777778,3.1333332,2.675,1.7333333,5.2083335,20.96667,17.675,9.933333,3.4333334,0.33333334,1.1666667,0.35,0.78888893,0.0,0.8444445,1.3000001,3.4583333,2.2222223,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2777778,2.2000003,13.099999,16.066668,16.433334,5.5,1.6999999,2.1583333,11.244445,7.2666674,6.9416666,1.1444445,1.2583333,1.1333333,2.0666668,7.655556,8.944445,0.7416667,0.0,0.16666667,2.288889,0.0,1.6888889,7.2666664,1.7555555,0.0,0.0,0.0,0.08333334,0.1888889,0.075,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.2888889,0.56666666,0.9666667,0.81666666,0.6111111,0.50000006,0.32222223,0.14166668,0.13333334,0.21111111,0.16666669,0.41111112,2.2416666,7.1222224,27.75,62.57778,92.700005,115.225006,116.8,109.9,99.166664,88.5,68.888885,54.800003,44.01111,38.52222,31.375002,33.155556,37.850002,39.744442,45.141666,55.477776,60.93334,57.65001,51.444443,33.975002,27.844444,32.175,44.08889,61.425003,81.688896,97.12222,67.78333,37.82222,18.258333,8.755556,6.7250004,7.2777777,3.7444446,4.408334,5.0666666,8.333333,5.6888895,2.7250001,0.4,0.0,0.008333334,0.4111111,1.7416667,3.677778,5.1083336,0.125,0.21666668,0.34166667,0.5625,0.85,1.1687499,1.5916668,1.5500001,2.2166667,2.4750004,3.5625,1.7916665,1.50625,0.9416666,0.64374995,0.041666668,0.0125,0.016666668,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.32500002,0.8625001,0.45833337,1.15625,2.7416668,3.7125003,7.1416664,9.6125,14.975,15.933332,14.425,10.683333,6.3812504,5.041666,5.875001,6.5249996,7.4250007,6.95625,6.7,6.7937503,12.525001,19.41875,19.433334,15.841665,12.612501,8.891667,5.83125,4.1666675,2.49375,1.5916667,3.7999997,6.95,8.983334,11.08125,13.116667,17.931248,20.0,20.40625,23.208336,25.333334,27.99375,29.683334,34.100002,37.708332,22.10625,15.258334,15.268749,11.858335,12.775,14.906251,12.0,11.793751,12.725,12.393749,12.900002,13.158335,11.575,8.408333,4.6187496,2.6416667,1.8812501,1.791667,2.375,4.8187504,8.266667,8.88125,8.991668,7.5875006,5.758333,5.20625,6.291667,6.416667,4.1875005,2.7083335,1.7125,0.85,1.9999999,2.0,3.9416668,4.46875,9.491667,6.4687495,2.6833336,0.91249996,0.36666667,0.68125004,3.3833337,9.791666,20.206251,35.141666,31.025002,13.391668,10.881249,5.7,0.7916667,0.0,0.0,0.0,0.42500004,0.06250001,1.1583334,1.4750001,2.6749997,2.4916666,0.99375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.3750002,7.29375,7.4,6.4,5.0333333,4.8125,2.175,1.7625,6.1750007,4.766667,8.98125,3.7249997,2.3000002,1.75,1.8562502,2.7416666,2.8916667,0.04375,0.0,0.0625,0.65000004,0.0,0.34166667,1.325,4.7,0.0,0.0,0.0,0.09375001,0.15833333,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.35000002,1.1250001,1.6666667,1.6187501,1.5166667,1.125,0.71666676,0.45625,0.20000002,0.1,0.0125,0.60833335,3.5625005,10.158333,33.63125,74.38334,107.25,138.43124,139.01666,129.45625,111.549995,93.25625,74.39167,61.49375,55.683334,56.958336,51.6375,48.21667,49.0125,46.425,41.3625,37.1,36.899998,35.51875,43.13333,36.743748,33.125,38.162502,53.25833,70.2125,82.816666,87.84167,82.987495,42.933334,18.4375,13.708334,10.918751,6.541667,3.9500003,3.2750003,4.475,7.9625,5.7083335,2.225,0.033333335,0.008333334,0.28125,1.1833334,2.8312497,4.2000003,4.50625,0.033333335,0.07777778,0.36666667,1.05,1.5444443,1.8000001,2.2333333,2.9583335,2.711111,2.8999999,5.2916665,7.3222218,6.9000006,2.988889,1.0083333,0.15555556,0.008333334,0.0,0.0,0.0,0.0,0.05,0.0,0.24166667,0.37777779,1.3555557,7.8,10.666666,10.208334,1.9333333,4.366667,5.8222218,7.816666,12.388888,11.733332,7.758333,7.0888896,5.2416663,2.3222222,3.0916667,4.3444443,3.6777775,3.4500003,3.222222,3.0666668,3.3444448,3.9333334,3.9444444,3.0666666,1.7916669,0.8999999,1.5416667,1.8222224,1.4666667,1.7111111,3.816667,6.277778,8.155556,10.608335,15.755556,24.058332,31.288889,36.899998,45.655552,52.877785,65.799995,64.27778,66.916664,40.277775,35.350002,30.466667,31.550005,29.033335,29.122225,27.1,24.2,24.766668,21.377779,14.116666,10.8555565,10.622223,9.375001,6.5888886,3.6333334,2.5555556,2.9083335,2.9,4.2222223,7.416667,9.588889,9.558333,8.744444,4.475,2.6333334,3.9916668,5.3222227,5.955556,3.8833332,2.4333332,1.7,0.66666675,0.5583334,0.42222226,0.8,0.4666667,0.25555557,0.041666668,0.0,0.0,0.08888889,0.53333336,0.64444447,4.5,22.29167,40.71111,43.541668,30.444447,13.425001,3.8555555,0.5777778,0.0,0.0,0.0,0.0,0.0,0.26666668,0.85555553,1.275,0.9444445,1.6666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,5.2222223,8.433334,1.9666666,1.1333333,0.35555556,2.7,4.233333,1.1833334,5.377778,2.5777779,2.308333,3.166667,1.3499998,0.2111111,0.1,0.0,0.0,0.0,0.0,0.083333336,0.0,0.0,0.45555556,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.23333333,0.68888885,0.40833336,0.36666664,0.21666668,0.11111111,0.06666667,0.0,0.0,0.016666668,0.9222222,5.4333334,14.611112,39.291668,81.922226,119.53334,143.36667,146.96667,141.25835,125.92222,108.725006,85.91111,66.03333,69.555565,87.47779,83.59167,75.94445,64.091675,53.933334,49.11667,30.966665,23.31111,22.575,44.63333,49.333332,35.766663,42.833336,61.344444,62.65,69.344444,90.94444,97.933334,45.31111,22.1,14.922222,12.758333,6.2111115,3.5555558,3.725,7.044444,10.616667,5.1444445,2.3416667,0.011111111,0.25555554,1.2166667,3.088889,4.7000003,4.611111,3.1833339,0.0375,0.108333334,0.47500002,1.14375,1.875,2.56875,3.3999999,4.5437503,4.925,5.183334,7.3624997,10.75,8.037498,3.6666667,0.75625,0.14166668,0.075,0.033333335,0.008333334,0.0,0.0,0.40624994,1.6750001,3.2749996,4.0833335,4.8749995,6.937501,12.083332,9.03125,3.6499999,4.39375,4.4,5.11875,5.058334,3.25,2.59375,3.766667,4.56875,4.0249996,3.3624997,4.175,4.7,3.0625,1.8333334,1.2624998,2.0083334,1.4437499,1.1583333,1.05,0.55,0.55833334,0.68125004,1.075,1.1812501,2.0,3.525,5.366667,6.9833336,10.075001,18.025,30.199999,37.56667,43.36875,57.64167,66.04167,77.5125,72.61667,71.137505,51.208332,47.031254,39.225002,36.287502,38.325,38.075,27.98125,22.81667,23.3125,18.741669,13.3,12.375001,11.958335,10.08125,8.166666,6.700001,5.8416667,4.9875,5.875,9.133334,11.400001,10.724999,8.0375,6.7666683,3.3249998,1.75,2.2937503,2.8333335,3.266667,4.2937503,6.583333,8.200001,6.9750004,4.0312505,0.43333334,0.3916667,1.1437501,0.9333334,0.43125004,0.033333335,0.0,0.0,0.0,0.083333336,0.34166667,5.3500004,18.858334,26.2875,26.583334,23.56875,10.425,1.45,0.0,0.0,0.0,0.0,0.21875,0.18333334,0.6833333,4.9312496,2.7333333,0.66249996,0.0,0.0,0.0,0.0,0.0,0.20833333,0.10625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7833334,0.0625,0.0,0.0,0.0,4.5125003,11.575,3.4250002,1.2500001,1.9333334,1.33125,0.6083333,0.45000008,0.45,0.34375,0.008333334,0.0,0.0,0.0,0.1,0.13333334,0.3,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.32500002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,1.4583334,6.4624996,17.666666,44.95625,98.28334,164.57501,218.4875,223.13333,208.85626,164.34167,131.34375,111.825005,101.96875,98.625,99.25832,98.23126,98.68333,83.76875,71.51667,60.356255,36.074997,24.2,20.1,24.474998,31.83125,24.483334,38.756252,58.783337,64.674995,82.21667,97.05,96.549995,53.833336,26.4375,16.633335,12.712501,6.449999,2.7500002,3.6749997,6.7250004,9.15625,3.4499998,0.94375,0.10833333,0.85833335,2.7,4.8583336,4.6000004,1.9916668,0.56874996,0.0,0.0,0.0,0.0,0.033333335,0.24166667,0.70000005,1.1500001,1.1444445,0.98888886,1.0666667,0.9444445,1.0999999,0.7888889,0.24166667,0.12222222,0.083333336,0.044444446,0.011111111,0.033333335,0.12222223,0.20000002,0.21111111,0.37499997,1.7555556,3.2111113,3.391667,3.8111107,3.9,3.1555557,5.4249997,5.8777785,5.9666667,6.133333,4.9111114,5.483334,7.422222,10.733334,15.355555,15.466667,10.777779,5.544444,4.125,2.3222222,2.2333333,2.6555557,1.5833335,0.85555565,0.75555557,0.52500004,0.62222224,1.4333333,2.3666668,2.4333334,3.0333338,3.125,3.4444444,5.9111114,9.866666,19.122223,32.208336,37.255558,38.800003,47.555557,56.322227,56.725002,50.233334,46.283337,39.855556,31.500002,25.622221,27.858334,30.855555,32.622223,24.808332,18.844444,14.691666,10.144444,7.7083335,7.0666666,6.833333,5.991667,5.011111,4.841667,5.4444447,6.3500004,10.655556,16.01111,19.366667,17.844444,13.249999,10.422222,5.733333,1.7444444,0.7666667,0.37777779,0.7222223,2.825,5.766667,6.658334,5.9444447,4.0166664,1.8666667,1.3555557,0.4166667,0.32222223,0.175,0.6666667,1.2416667,0.5444445,0.8333334,0.85555553,0.34444442,1.8416668,6.022222,13.333334,16.900003,4.383333,3.1666665,0.21111111,0.0,0.0,0.0,0.16666667,0.125,0.2777778,1.3555555,6.1833334,2.4666667,0.6583333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4666669,18.324999,9.577778,1.4583334,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,0.0,0.0,0.0,0.0,0.13333336,0.5333334,0.13333336,0.0,0.06666667,0.33333328,0.29999998,0.1,0.055555556,0.2,0.011111111,0.0,0.0,0.0,0.074999996,0.37777776,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,0.14166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,1.3444445,5.2583337,14.433332,36.274998,91.11112,167.11111,239.6,263.84445,299.4167,283.40002,174.96666,117.18889,93.54167,89.2,96.63335,100.841675,96.88889,63.025,63.7,69.375,46.911114,26.944445,23.133333,21.177778,17.491667,20.18889,34.575,52.255554,77.75833,81.36667,69.63333,64.98334,45.055557,29.341667,20.655556,9.616668,4.311111,2.0222223,2.4333339,7.166667,9.625,2.5,0.4166667,0.13333334,1.0333334,3.125,5.311111,4.5416665,1.5,0.36666667,0.0,0.0,0.016666668,0.075,0.10000001,0.45625004,1.4416667,2.4812503,2.625,3.4166663,3.6812499,2.9833333,3.0500002,2.358333,1.4562501,0.975,0.6812501,0.3416667,0.11666667,0.01875,0.058333337,0.17500003,0.34166667,0.65,1.15,2.875,4.8375,5.5166664,3.7125,1.925,0.83124995,1.0416667,2.125,3.1333337,3.3833332,3.1125,2.6583333,6.9,10.650001,10.8375,7.4333334,2.975,2.125,0.8333334,0.9125,1.2166667,0.9312499,0.83333325,0.8833333,0.65,1.7583333,2.1875,1.85,2.13125,1.7583333,2.1750002,3.2833335,5.4249997,10.456251,19.866667,32.712498,32.500004,31.206251,35.01667,36.30833,30.056253,24.383333,23.53125,19.85,14.856252,13.183333,16.56875,19.525002,19.783335,15.41875,10.291666,7.0062504,5.708333,6.4,7.2166667,7.166667,6.393749,5.7000003,6.0875,8.125,12.4,18.516666,21.816666,24.393751,23.325,21.1125,19.566668,11.762501,3.3916664,1.05,1.0250001,1.8416668,3.025,5.3500004,8.099999,5.916667,2.125,1.4416668,1.7583334,0.45000002,0.14999999,0.09375,0.9916667,2.8249996,3.916667,2.3937502,1.7166667,0.3166667,0.33125,0.9500001,3.6374998,4.0499997,1.475,0.0,0.0,0.03125,1.1999999,1.3062501,2.5083332,0.48125,1.175,0.94166666,4.0,4.5333333,0.99375004,0.05,0.0,0.0,0.25,0.20833334,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.4416666,12.512499,16.35,4.95625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.51666665,0.0,0.0,0.0,0.14999999,0.05,0.1,0.13333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43333334,0.01875,0.07500001,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31875,1.7416668,6.46875,20.508333,42.875004,84.0,138.29167,194.88126,215.32501,250.28749,241.10834,192.63126,119.93334,78.81875,63.38334,81.25833,95.893745,87.433334,71.60625,72.63334,74.987495,55.550003,31.475,17.9625,14.141666,12.062499,22.775003,44.68125,64.98333,73.11875,54.733334,54.483337,52.693752,37.333332,29.61875,17.041668,8.15625,8.541666,3.4583335,1.9375001,8.408333,8.731251,1.7166667,0.3625,0.016666668,0.375,1.18125,2.2,2.1125,0.5,0.79375,0.0,0.022222223,0.17777778,0.34166667,0.47777778,1.1333334,2.4111114,3.4916666,3.7777777,4.1,3.8083332,2.3222225,0.9750001,0.51111114,0.22500001,0.15555555,0.22500002,0.23333335,0.14444445,0.041666668,0.011111111,0.108333334,0.17777777,0.39166665,0.58888894,0.53333336,1.0333333,1.8888888,1.9416666,1.0444446,0.7583333,0.5,0.47500005,1.1666667,2.7111113,2.9833333,1.8777778,2.1916668,3.0111108,3.4083335,3.5000002,5.955555,4.9250007,1.6222222,1.85,2.411111,1.5916668,1.9777777,1.688889,1.3,0.9111112,1.0583333,1.3555558,0.5166667,0.9222222,2.1750002,2.6222224,3.7222223,7.283334,13.955555,25.766666,24.044445,19.633333,15.288888,12.455555,11.166667,10.9,9.983334,9.8,7.358333,7.377777,8.641666,7.7444444,5.577778,4.0833335,2.7777777,3.5083332,4.3111115,6.05,7.0666666,7.855555,7.8250003,7.2999997,9.741667,14.944446,22.558332,24.988888,23.955555,23.558334,25.133335,25.891668,24.0,19.766666,9.277779,2.1333332,0.53333336,0.92222226,1.4333334,1.9111111,2.9583335,4.2666664,6.758334,3.8333333,1.6888889,0.40833333,0.011111111,0.5,1.1,0.9583334,1.0888889,4.0666666,1.7666665,0.7666667,0.9583334,1.7666667,1.0166667,0.988889,0.0,0.0,0.0,0.083333336,9.8,3.925,4.3555555,7.975,5.5111113,2.977778,1.0333334,3.2222223,1.3666668,0.23333332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,10.277778,10.066668,1.1777778,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8333334,0.44444445,0.4166667,0.8,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4000001,0.008333334,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.49166673,1.7777779,5.1249995,17.300001,33.0,56.288887,86.35556,129.075,161.64445,223.29166,259.84442,185.44168,110.700005,73.52501,64.31111,75.03334,88.68334,81.33334,70.341675,89.37778,98.20001,79.144455,51.75556,27.658335,18.155556,18.766668,28.444443,36.375004,56.344448,47.51667,40.18889,31.822222,39.041668,55.36667,30.3,14.633334,12.391666,1.8666667,0.1,1.4833333,10.444445,7.8833337,1.3,0.09166667,0.0,0.0,0.0,0.0,0.0,0.055555556,1.3666668,0.0,0.022222223,0.16666669,0.35,0.6444445,1.0916667,1.9666666,2.7999997,3.6,4.188889,4.008333,4.0666666,3.1000001,2.2333333,0.9666667,0.21111113,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.8083334,1.5555556,2.475,1.9555556,2.4777777,2.916667,2.1333334,1.0083334,0.2777778,0.9,1.9666667,2.8111115,3.5500002,4.755555,10.358334,14.333333,7.8916664,3.9444447,2.988889,2.8833332,2.3666668,1.6000003,0.9888889,0.6499999,0.9,2.6333334,3.6555557,3.6777778,5.0333333,7.3222218,10.924999,18.62222,17.283333,12.799999,9.866667,10.241667,9.455556,11.691666,11.066668,7.5083337,5.088889,4.6749997,2.6333332,1.7555555,1.2166667,1.3222222,2.95,4.911111,6.7083335,8.944445,9.7,9.583333,8.711111,10.016666,15.166669,21.516666,22.166668,18.2,21.275,22.811111,26.333334,26.333336,20.841667,8.98889,1.7666665,0.51111114,0.56666666,1.3166666,2.4888887,2.5083334,2.3555558,2.3583336,3.0,1.9111112,0.41666666,0.033333335,0.0,0.033333335,0.108333334,0.28888893,2.7833333,2.4666667,0.42222223,1.7916667,3.0555556,3.25,1.5666667,0.0,0.0,0.0,0.0,0.0,1.9000001,0.06666667,0.7083334,0.0,0.2888889,0.21666668,0.13333334,0.0,0.0,0.175,0.044444446,0.0,0.0,0.13333334,0.175,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,51.391663,3.9333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.0,0.48333332,1.6,0.61666673,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,0.34444442,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,1.2222222,3.1333334,12.266666,25.475,44.355553,67.566666,108.83333,143.1,193.04169,234.82225,150.05,89.32223,72.38334,73.933334,74.5,78.79167,63.166664,61.83334,74.100006,81.03334,55.87778,43.866673,25.133333,14.966667,15.133333,20.266668,24.566666,39.877777,35.875004,28.844444,23.622221,34.15,65.46667,33.38333,21.033333,15.141667,6.5111113,1.1111112,4.325,9.866667,5.4666667,0.74444443,0.008333334,0.0,0.0,0.0,0.0,0.0,0.16666667,2.0333333,0.03125,0.11666666,0.20833334,0.28750002,0.49166667,0.53125006,0.9666667,1.75625,2.8166666,3.5750003,2.0,0.71666676,0.54375005,0.5,0.19375002,0.36666667,0.35625002,0.18333334,0.15,0.30625,0.19166666,0.025,0.14166668,0.44375002,0.6,0.77500004,1.3625001,1.475,2.4625,3.2000003,4.9437504,6.3750005,6.14375,3.6666667,2.1333334,2.30625,1.5666667,0.40625003,0.5833334,3.1250002,7.9666667,13.6,17.3375,18.150002,19.05,18.516668,11.1875,6.2833333,3.75,1.725,0.7166666,0.38125002,0.48333335,0.43750003,0.6833333,1.1812501,1.6,2.0083334,3.1124997,3.7083333,3.5187497,8.458333,16.256252,10.966668,10.025001,8.99375,5.55,9.06875,15.091668,11.112499,6.5083337,3.6625004,1.5583333,0.94166666,1.40625,2.3500004,4.9000006,5.783334,7.325,9.241668,10.133334,8.612499,7.408334,8.49375,11.375,10.700001,10.208334,9.525,10.76875,12.558333,12.543751,10.316667,5.2000003,2.2500002,0.50625,0.041666668,0.18333334,1.5937502,3.2,3.4437504,3.5,2.3999999,1.1416667,0.72499996,0.0625,0.0,0.0,0.058333337,0.24375,0.45,0.93125004,0.475,0.775,1.16875,3.3333335,2.625,1.0416667,0.0625,0.0,0.0,0.0,0.0,0.1125,0.05,0.0,0.0,0.0,0.01875,0.125,0.075,0.025,0.24374999,0.15833332,0.09375,0.0,0.025,0.09375,0.20833331,0.18749999,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18750001,0.85,0.47500002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,0.36666664,0.21875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.043750003,0.07500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.48333335,1.6875,4.775,15.725,26.058334,38.975,63.025,80.66667,101.850006,96.53333,78.51875,56.175003,53.13125,70.075,91.066666,74.14375,36.183334,39.6125,49.591667,55.581253,34.208332,24.758333,19.26875,10.666668,11.756251,13.641666,15.275002,29.691666,31.806252,19.775002,18.383335,41.09375,33.458332,26.025,20.333334,14.906251,16.949999,2.6833334,7.3125005,6.791667,2.5000002,0.11666667,0.0,0.0,0.0,0.0,0.0,0.05,0.44166666,1.66875,0.38333333,0.8666667,1.4222223,2.225,2.9555557,3.2416668,4.377778,5.4666667,8.966667,12.077777,10.766666,5.8333335,2.5833333,1.6444443,0.53333336,0.43333334,0.43333337,0.44444445,0.9777778,2.075,2.5555558,1.7333336,2.1444445,2.65,3.7222226,3.8000002,3.5666666,5.3444443,5.341667,4.9,6.266667,7.8222227,4.6333337,2.6555557,2.7888887,2.5416667,2.177778,2.0083334,1.6111112,1.4333333,4.022222,8.177777,15.25,17.711113,16.55,12.077778,6.7999997,3.622222,1.6333334,0.55833334,0.011111111,0.025,0.18888889,0.11666667,0.26666668,0.47500002,0.51111114,0.6333334,1.7166667,3.7444446,6.8166666,9.777779,8.075001,6.7,6.188889,7.5083323,4.4555554,6.425,7.866667,8.725,5.7222223,2.675,1.9666667,1.777778,1.9583334,3.0111113,5.6666675,6.9777775,9.325001,11.155556,11.777777,9.416667,7.577778,10.691668,13.455555,11.308334,5.4777784,3.9,7.991667,13.066668,12.891666,6.3111115,2.6333334,1.6777778,0.39166668,0.0,0.044444446,0.11666667,0.17777778,0.30833334,0.68888897,1.475,1.7777778,1.1222223,0.84166676,0.5,0.7083334,0.47777778,0.075,0.51111114,2.275,3.488889,3.5333333,5.9750004,3.6000001,3.9083333,3.5333333,1.2249999,0.36666667,0.14444445,0.0,0.0,0.0,0.13333334,0.06666667,0.0,0.4,0.15,0.19999999,0.29999998,0.0,0.05,0.06666667,0.175,0.033333335,0.0,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24444447,0.9666667,1.0555556,5.808333,15.111112,30.744442,44.283333,62.54444,64.90834,52.53333,36.158337,31.922224,40.325005,60.755554,97.288895,79.00833,31.022223,28.475002,39.78889,46.116665,23.255558,14.5222225,11.008334,8.333333,12.266666,10.833334,15.141668,27.155556,29.474998,19.733334,13.411112,23.033333,29.222223,25.216667,11.744445,5.2666664,3.3666668,1.4222223,1.925,2.1,1.8083333,0.4,0.0,0.0,0.0,0.0,0.0,0.36666667,1.2111111,2.9333334,0.35625,0.9,1.4666667,2.36875,3.7416668,4.3375,5.5000005,7.1187496,9.283334,12.058334,12.825,9.033333,4.38125,2.6583335,2.3000002,1.9916668,1.11875,0.55833334,1.2833334,3.34375,4.766667,6.5999994,7.5500007,7.9875,8.633334,7.0083337,6.7000003,7.0249996,4.81875,3.8000002,3.26875,2.641667,2.50625,2.8333335,3.5916665,4.63125,6.6666665,6.65625,4.1333337,2.1937501,2.225,2.6166668,2.5875,2.1833334,1.29375,0.40833336,0.087500006,0.016666668,0.033333335,0.20000002,0.625,0.95625,1.2333333,1.2500001,1.1333333,1.1874999,1.3666667,1.9416668,3.58125,6.025,7.4125004,6.7666664,6.4750004,7.541667,9.999999,9.75,5.6250005,3.75625,4.4000006,5.3937507,4.2749996,2.475,1.1583334,0.5416666,0.45625004,0.8416667,1.6875001,3.5000005,4.2625003,6.9916663,5.25,6.025,8.458333,11.887501,14.224999,16.125,11.5,8.3,7.3375006,7.6583333,5.3937497,2.15,1.6312503,1.7166666,0.65000004,0.06666667,0.0,0.0,0.0,0.0,0.09166667,0.75,1.6999999,0.85,0.5,1.1083333,1.475,1.2083334,1.1312501,1.1500001,2.76875,5.2250004,11.258333,13.375,14.083334,14.68125,15.275,13.3375,6.95,2.8583333,0.4875,0.4166667,0.22500001,0.075,0.0375,0.0,0.60833335,0.61875004,0.05,0.4125,0.69166666,0.28125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15833333,2.8999999,8.008333,30.541668,49.968754,58.641674,49.3375,28.35,27.400002,30.416664,41.61875,70.23334,114.45836,85.262505,40.31667,31.281248,36.36667,41.0625,24.425,16.275,19.718748,22.766666,28.94375,17.108334,29.181248,29.733335,28.112501,31.758335,30.358334,45.16875,45.833336,24.718752,10.316668,2.6375,0.55,0.125,0.28125,0.51666665,1.8624998,1.475,0.29375,0.0,0.0,0.0,0.041666668,0.5875001,1.3583335,4.68125,0.016666668,0.044444446,0.044444446,0.14166667,0.5555556,1.225,2.7,3.1916668,4.3000007,4.9222226,5.5833335,3.7111108,3.4083333,2.6666667,2.6166668,1.6777778,1.5416666,1.8444445,2.0777779,3.1666665,3.6,4.45,4.788889,3.925,3.688889,4.266667,5.125,3.9888885,2.6666667,2.5444446,2.2666671,2.2444446,2.1916668,3.5777779,5.4444447,7.216666,7.5888886,6.166667,5.611111,7.7666674,12.166666,12.9777775,9.616667,6.5333333,3.6750002,1.6555557,0.97499996,1.5,2.3555555,2.4916663,4.2,2.8166666,1.8000001,1.8666667,2.188889,2.4083333,3.2555556,4.2333336,5.616667,5.666667,6.158333,6.6333337,7.766666,8.966667,13.844443,11.783334,7.9000006,5.8166666,5.3888884,5.0499997,4.388889,3.2416666,2.3777778,2.9555557,2.1000001,1.5222223,1.5083334,1.4000001,1.8166666,1.9888889,2.6888885,2.6000001,3.3444448,4.8583336,8.200001,12.566668,8.088889,4.822222,4.675,2.8,0.9916667,0.37777776,0.19166666,0.73333335,0.57500005,0.10000001,0.044444446,0.10000001,0.26666668,0.175,0.011111111,0.0,0.0,0.044444446,0.016666668,0.055555556,0.6333333,1.3333333,1.6,1.9444444,3.0416663,2.5444446,5.7222223,14.266666,20.91111,19.44167,15.777778,17.791668,14.133333,10.9777775,4.65,8.911111,2.4166667,1.7444444,0.40000004,0.0,0.0,0.0,0.022222223,0.083333336,0.6333333,0.69166666,0.11111111,0.0,0.0,0.1,0.05,0.0,0.025,0.11111111,0.0,0.0,0.0,0.75,1.6666666,0.75,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39166668,1.0222224,14.411112,40.516666,36.6,31.583334,19.055557,19.841665,17.8,21.425001,18.877777,22.68889,29.158333,31.944443,32.983334,34.744446,34.483337,23.08889,26.955557,35.49167,30.577776,26.233332,23.233334,30.066664,30.599997,21.883335,26.944447,42.888893,46.74167,40.422222,32.616665,12.844445,2.8833337,1.1000001,1.2666667,1.3416667,1.5777779,1.2083334,0.73333335,0.4333333,0.0,0.0,0.0,0.06666667,0.66666675,1.3222222,4.15,0.0,0.008333334,0.008333334,0.04375,0.35833335,0.88750005,1.9166667,2.225,2.85,2.8,2.9375002,2.3000002,1.80625,1.4083333,1.15,1.1250001,1.8625,3.5333338,4.891667,7.0375004,8.166666,6.2875,4.5083327,1.8937501,0.5083333,0.6,1.5875,2.7833333,5.9500003,8.683334,6.637501,5.941667,4.85625,5.2916665,6.7333336,8.06875,6.666667,8.9625,10.816667,13.0875,16.466667,16.533333,12.8875,8.05,5.3812504,3.733333,3.9875,4.966667,5.341666,4.575,5.9500003,6.206249,4.4500003,1.5625,0.6166667,0.675,0.9916667,1.5666666,2.4125,3.3,4.2687497,5.758333,7.737499,9.35,7.5166674,5.0249996,3.1916668,1.76875,1.6500001,2.60625,3.4083333,3.3562498,3.6583335,3.65,2.9687498,2.4916668,2.1625001,1.7083334,1.4562501,1.2500001,1.1833334,0.89375,0.9416667,1.5937499,3.6833334,5.3625,4.1500006,3.25,2.6625001,1.25,0.54375005,0.083333336,0.075,0.06666667,0.0125,0.0,0.0,0.13125001,0.625,0.35625005,0.05,0.15,0.13333334,0.15833335,0.05,0.0,0.0375,0.22500001,1.2874999,1.8416666,3.4562502,2.75,2.5333333,5.6312504,12.2,16.43125,13.4,8.587501,6.825001,7.2666664,8.481251,3.1000001,0.6625,0.51666677,0.3625,0.075,0.0,0.056250002,0.30833334,0.0,0.0,0.70625,1.1166668,0.81249994,0.1,0.125,0.63124996,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16250001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,8.558333,25.79375,24.408333,23.193752,13.0,11.237501,10.808333,11.318749,4.0750003,2.1083333,2.76875,3.2833335,15.687499,24.558334,20.01875,15.583333,31.391666,42.475,26.208336,18.23125,32.75,27.45,14.425,14.299999,20.641666,24.291668,32.25,29.258335,23.662502,13.366668,4.4875,3.291667,3.025,3.64375,2.0083334,1.05625,0.0,0.0,0.0,0.0,0.0,0.016666668,0.20625001,0.52500004,1.61875,0.0,0.0,0.0,0.033333335,0.12222223,0.21666667,0.39999995,0.65833336,1.0222223,3.7333333,6.591667,6.122223,5.0916667,4.7222223,4.325,3.5444446,3.1500003,2.9666667,4.011111,2.8166668,1.6000001,0.70000005,0.26666668,0.3,0.23333333,0.6666667,1.625,3.1444445,4.775,5.233333,4.258333,4.1555557,4.5333333,4.5,4.7555556,4.1000004,4.133333,5.5333333,8.888889,10.266667,14.144444,15.477777,13.516667,10.922222,8.341667,7.3555555,8.358335,10.599999,11.788889,14.341666,11.211111,5.5249996,1.3666668,0.17500001,0.2,0.3416667,0.6,0.8888889,1.2083333,1.4666667,1.6416667,1.9666667,1.4,1.7222223,1.0666667,0.6333333,0.3,0.28333333,1.0666666,1.75,1.7222223,1.45,1.0111111,1.2333333,1.2416668,1.3555555,2.025,2.2222223,2.6,2.9666667,3.1555557,3.158333,3.4222224,4.4916673,5.4333334,6.375,5.588889,4.5111113,2.4083333,0.8333334,0.14166668,0.0,0.016666668,0.18888889,0.20833334,0.044444446,0.0,0.074999996,0.011111111,0.13333334,0.3,0.116666675,0.0,0.0,0.0,0.0,0.016666668,0.044444446,0.3,0.46666667,0.91666675,1.2555556,0.9444444,2.5500002,5.855556,9.466667,10.422222,6.833334,2.1444445,1.4222221,1.1083335,0.16666667,0.19999999,0.26666665,0.39999998,0.16666667,0.0,0.0,0.0,0.0,0.0,0.33333337,0.73333335,0.575,0.06666667,0.1,0.35833335,0.14444445,0.0,0.0,0.0,0.0,0.17777778,0.53333336,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7,10.183332,15.733334,11.791668,4.4000006,6.9833336,8.466665,10.258334,2.0666668,2.0222223,2.075,8.433334,17.65,24.955559,18.375002,21.300001,30.233334,29.416668,23.488888,34.308334,50.86667,33.31667,14.211111,8.741667,14.044444,28.377779,35.86667,30.144447,17.025002,14.611113,6.4333334,8.8555565,9.822222,6.4833336,2.3222222,0.825,0.0,0.0,0.0,0.0,0.0,0.055555556,0.25,0.2777778,0.33333334,0.0,0.0,0.05,0.25625,3.1249998,5.225,5.3583326,5.1125,5.4416666,5.6333327,8.6125,6.791667,5.59375,4.891667,4.9875,5.283334,6.0875006,6.766667,6.6333337,7.1125,8.658332,7.9625006,7.116667,6.1125,4.05,3.166667,2.5375,3.0333333,6.23125,11.15,11.093751,10.533334,11.88125,13.791668,15.700001,14.868751,13.45,13.275,12.391666,10.7375,9.366667,9.383333,7.2437496,4.3666673,2.9125,2.9750001,2.8312504,3.4083338,4.216667,4.20625,2.0500002,0.2875,0.06666667,0.118750006,0.18333332,0.2125,0.21666667,0.26666668,0.3125,0.35833332,0.3625,0.25,0.025,0.083333336,0.13333334,0.125,0.0,0.08125001,0.375,0.43125004,0.33333337,0.1875,0.24166667,0.275,0.5500001,1.0333334,1.46875,1.475,2.33125,3.3166668,4.008333,4.3312497,4.433334,5.16875,5.4333324,5.1124997,4.4083333,2.8833332,1.5062501,0.5583334,0.10625001,0.0,0.0125,0.20833334,0.25,0.041666668,0.0,0.056250002,0.008333334,0.0,0.0,0.01875,0.0,0.033333335,0.19375,0.625,1.03125,1.3333333,1.7875,2.3916667,1.53125,0.36666667,0.22500001,0.9250001,1.6166668,2.2437499,1.975,2.0125,0.8166666,0.39166665,0.05,0.05,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0875001,0.5083334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.17500001,2.7083333,10.768749,12.991667,6.21875,2.8333335,3.5125,4.5916667,6.38125,1.4083334,5.3333335,3.2875001,6.475,8.925,12.175,14.08125,20.216667,27.966667,25.38125,30.333332,17.206251,21.133333,20.81875,33.0,19.21875,21.016666,32.88333,42.3375,26.758333,12.1125,10.808333,5.9125004,2.9416666,1.925,1.44375,1.3666667,0.51875,0.0,0.0,0.0,0.0,0.375,0.75,1.4375,0.5083333,0.48125,0.0,0.0,0.0,0.0,0.099999994,0.26666668,0.2888889,0.275,0.3,0.16666666,0.225,0.17777778,0.16666667,0.21111113,0.35000002,0.7555556,1.6750002,2.9777777,4.588889,7.125,10.6,13.858334,14.366667,13.775,14.088888,12.933334,8.016667,3.7666667,2.125,1.9000001,2.7666667,4.822222,8.2,11.544443,12.422222,10.233335,7.9777784,6.4,4.3333335,3.7166667,4.5333333,4.3,1.9416667,0.41111112,0.14166667,0.022222223,0.016666668,0.022222223,0.022222223,0.016666668,0.0,0.0,0.0,0.0,0.13333334,0.15833333,0.3111111,0.7777778,0.8583334,1.6333332,1.1416667,1.288889,0.8583333,0.32222223,0.15555555,0.016666668,0.0,0.07500001,0.35555556,1.95,4.3555555,5.4083333,5.4,5.5555553,6.458333,5.4777784,2.591667,1.3222224,1.15,1.0666668,1.5777779,1.9083332,1.7,1.7416667,1.8333334,1.9000001,1.4444445,1.0111111,0.55,0.24444446,0.058333337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.06666667,0.011111111,0.3,0.97777784,3.3916664,7.233333,10.316668,11.844444,9.766666,4.2666664,1.3111111,0.6916667,0.51111114,0.9666667,0.022222223,0.0,0.0,0.0,0.14166667,0.18888888,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.40833336,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32222223,1.2166667,5.2888894,1.7833335,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14444445,0.09166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.033333335,0.18888889,9.091666,15.622221,6.5166664,2.766667,4.2999997,5.3111115,1.3916667,2.4333336,4.944444,5.1249995,4.288889,4.05,6.0,15.775001,30.344446,28.433334,19.383333,20.099998,11.299999,7.988889,18.974998,29.322224,25.408333,34.444447,45.233337,25.633333,6.3555555,6.966666,9.466666,3.1166666,0.53333336,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29166666,0.3888889,0.33333334,0.16666667,0.2,0.0,0.0,0.1,0.48333335,1.0333334,1.5416667,1.0555556,0.43333334,0.0,0.044444446,0.18333334,0.45555556,0.7833333,1.3777778,2.3166666,2.9,2.8333333,4.0111113,5.922222,8.541667,10.222222,10.691668,10.866667,11.758333,10.3111105,8.855555,6.566666,5.411111,5.491667,5.2333336,6.291667,9.055556,13.566667,17.077776,18.522224,16.866669,14.288888,8.05,3.5222223,1.9250001,2.588889,2.5666666,0.6166667,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.011111111,0.16666667,0.85555553,0.7416667,0.5111112,0.9444444,1.4166666,0.5888889,0.17500001,0.11111112,0.08333334,0.0,0.0,0.0,0.2,0.28333333,1.0333333,1.7166667,2.5444446,2.725,2.5222225,3.277778,3.4166667,2.8666668,2.3333335,1.7555556,0.85833335,0.3,0.3888889,0.38333333,0.3,0.30833334,0.25555557,0.25833333,0.16666667,0.07777778,0.12500001,0.21111113,0.52500004,0.48888892,0.38333333,0.2666667,0.125,0.14444445,0.16666669,0.025000002,0.1,0.058333337,0.08888889,0.15833335,0.15555556,0.0,0.19166669,0.5,1.4,1.6999999,1.275,1.2555555,4.1499996,6.6777782,6.788889,6.575,1.4666667,0.875,0.43333334,0.0,0.0,0.0,0.033333335,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05555556,1.3083334,2.0222223,0.7916667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,0.28888887,0.16666667,0.13333334,0.65555555,7.3,15.044445,11.741667,7.5000005,4.8583336,6.111111,2.1083333,1.888889,4.011111,5.758333,4.744445,4.1333337,9.266667,16.533337,17.844444,18.766668,16.2,8.555555,4.508333,6.855556,14.783334,16.58889,16.841665,19.977777,31.733334,14.358334,2.288889,1.3666666,2.7333336,2.0166664,0.4666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10000001,0.2916667,0.625,1.60625,2.7333336,3.5749998,3.0,1.6125,0.48333338,0.45000002,1.5125,2.9499998,4.1625,4.4333334,4.89375,4.816667,5.19375,4.9500003,4.5916667,4.7250004,6.5916667,7.4062495,8.141666,7.3312507,6.65,7.0833335,6.25,8.166667,8.3125,7.9750004,8.131249,9.916667,11.743752,13.541668,15.833333,16.706251,14.099999,7.7750006,2.8833332,0.94375,0.9583333,0.97499996,0.34375,0.22500001,0.118750006,0.06666667,0.075,0.033333335,0.7666667,0.95624995,0.80833334,0.79375,0.7583334,0.6250001,0.6,0.26250002,0.033333335,0.0,0.0375,0.033333335,0.025,0.0,0.0,0.0,0.0,0.0,0.075,0.88124996,1.6916666,1.1500001,0.50000006,0.5812501,0.55833334,0.53333336,0.59374994,0.70000005,0.93125,0.9166666,0.8937499,0.45000002,0.20833333,0.0,0.0,0.0,0.65000004,1.05,0.975,1.6583334,1.7999998,1.6666667,0.79999995,0.35000002,0.3125,0.20833334,0.2875,0.2,0.13333334,0.0375,0.125,0.050000004,0.016666668,0.0125,0.0,0.0,0.06875,0.20833334,0.75,1.3749999,0.35000002,0.008333334,0.18750001,1.4083334,3.3000002,3.7250001,3.8083332,2.4375,1.7083334,0.09375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.16666667,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4875,1.0833334,0.725,0.13333336,0.33333337,7.6499996,18.016666,17.925,9.766666,3.85,3.2083335,1.8625002,3.0833335,3.525,5.1750007,5.008333,5.2875004,5.7333336,6.9374995,15.008333,17.766666,9.2125,2.1833334,2.475,7.9833336,15.33125,18.5,14.543751,21.766666,15.916666,7.15625,1.575,0.0,0.65,0.875,0.55833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.08888889,0.14444444,0.26666668,0.4666667,0.73333335,1.2333333,0.8416667,0.39999998,0.0,0.1,0.2111111,0.5333333,0.7222222,1.1416667,2.0555556,1.7583333,0.8000001,0.7555556,0.9916668,1.2444445,1.3166666,1.2111111,0.875,0.41111112,0.36666667,0.95000005,1.511111,3.4916668,7.444444,9.866667,10.355556,12.800001,14.666666,16.422222,13.933333,12.755556,8.458333,3.1888893,0.9416667,0.8333334,2.8000002,2.9583337,4.2666664,4.5833335,3.6111112,4.5583334,5.7666664,5.255556,3.5083334,2.5888891,1.9583334,1.5444444,0.875,0.5111111,0.15,0.0,0.0,0.0,0.0,0.0,0.08888889,0.19999999,0.32222223,0.42222223,0.98333335,1.6333333,1.6916666,0.6777778,0.1,0.23333333,0.60833335,0.6222222,0.8777778,0.6,0.36666667,0.116666675,0.1,0.07500001,0.022222223,0.0,0.033333335,0.05555556,0.075,0.044444446,0.008333334,0.24444444,1.0111111,1.6500001,3.7000005,2.9666667,2.0444443,1.4166666,0.51111114,0.45833337,0.48888892,0.4,0.033333335,0.0,0.0,0.0,0.0,0.0,0.011111111,0.116666675,0.033333335,0.016666668,0.15555556,0.35000002,0.8777779,0.19166669,0.39999995,0.76666665,0.06666667,0.14444445,0.41666672,0.54444444,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39999998,1.3555555,1.575,0.36666667,0.13333334,3.9333334,8.288889,6.9333334,3.9666665,2.2000003,0.86666673,1.6583334,3.1555557,2.4111109,2.2583334,4.9444447,4.266667,1.888889,2.6416667,9.977778,9.655555,1.0666667,6.6444445,10.266666,15.611111,17.991667,24.1,17.4,12.8555565,6.255556,3.0583334,0.44444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.008333334,0.0,0.0,0.0,0.0,0.033333335,0.05,0.10833334,0.10625,0.19166668,0.11666667,0.30625,0.5833333,0.65625006,0.6083334,0.8375,1.6999999,1.625,0.8416667,0.8666667,0.9687501,1.275,1.625,1.8083332,1.4687501,1.6416667,2.325,3.6125004,4.6166663,5.8125,6.791667,7.8687496,7.9083333,5.6062503,6.625,6.3,6.04375,4.8,3.4812503,1.9083333,1.125,1.825,5.766666,7.5624995,7.875,6.5125,5.1166663,4.9125004,6.241667,5.925,3.0125,1.3916667,0.91875,0.5,0.23750001,0.108333334,0.01875,0.0,0.0,0.0375,0.14166668,0.38750002,0.45,0.6437501,0.90833336,0.7916667,0.70625,0.625,0.43124998,0.11666667,0.01875,0.06666667,0.081250004,0.108333334,0.06666667,0.1625,0.1,0.1625,0.20833334,0.118750006,0.033333335,0.0,0.05,0.15,0.6,1.625,1.975,2.4166667,2.3083334,1.15,0.69166666,0.91249996,0.9166667,0.95624995,0.7833334,0.58750004,0.6166667,0.7416667,0.36875,0.13333334,0.0,0.0,0.0,0.0,0.008333334,0.075,0.083333336,0.05,0.10000001,0.5812501,0.8,0.6375,0.058333337,0.025,0.0625,0.025,0.00625,0.016666668,0.0125,0.074999996,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28333336,1.3583333,0.36875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.34374997,0.06666667,0.0,0.0,0.0,0.0,0.0,0.00625,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,1.04375,2.016667,1.08125,0.13333334,0.0,2.1812503,3.2666667,2.6562502,1.75,0.32500002,0.06666667,0.5875,1.8083334,2.8083334,5.025,6.675,3.71875,0.8666667,0.5625,3.1833334,4.6916666,7.6937504,12.449999,11.900002,8.958334,9.88125,11.908334,14.49375,8.041667,2.591667,0.3,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19166668,0.38125002,0.0,0.0,0.0,0.0,0.17777778,0.65833336,1.477778,2.425,2.8555555,1.5444444,0.53333336,0.2777778,0.73333335,1.4111111,2.5,4.6111116,6.4500003,6.2777777,5.5000005,5.016667,2.7000003,1.3833333,0.42222223,0.1,0.7,1.7666667,3.141667,2.022222,0.42500004,0.5,0.6333333,0.40000004,0.22500001,0.20000002,0.6555556,1.4166666,2.2666667,2.9583335,3.4444447,3.6000001,3.7222223,3.888889,3.85,2.788889,1.4083333,0.7777778,1.6166668,3.6555557,5.144444,3.3333333,1.588889,0.5833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,0.09166667,0.07777777,0.016666668,0.0,0.0,0.0,0.3,0.31666666,0.46666664,0.5333333,0.46666664,0.35000002,0.26666665,0.1777778,0.15833335,0.055555556,0.0,0.0,0.075,0.099999994,0.31111112,0.0,0.0,0.0,0.31111112,2.3333335,5.1222224,8.222222,8.675,6.911112,2.2583334,0.90000004,1.5666668,1.3222222,1.3583333,1.3555557,0.8666667,0.5,0.5666667,0.20833334,0.06666667,0.008333334,0.0,0.0,0.0,0.022222223,0.23333336,0.35555556,0.8333334,0.8444444,0.32500002,0.033333335,0.011111111,0.033333335,0.16666669,0.20833336,0.2888889,0.108333334,0.08888888,0.25555554,0.25,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6666667,0.40000004,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.44444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,1.0916667,2.288889,1.35,0.43333337,0.15555556,0.016666668,0.0,0.15,0.0,0.3,1.3333334,4.5,4.688889,5.788889,7.983333,6.6777782,3.2833333,5.0555553,6.6333337,6.0666666,3.8222225,17.43333,19.088892,10.283333,6.4888887,6.6000004,16.444443,19.133333,9.744444,1.7333333,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.54444444,0.175,0.09375,0.31666666,0.25833333,0.6375,1.15,2.1,3.6833334,4.20625,3.991667,2.3666668,2.0,3.9166667,4.5750003,4.725,6.54375,7.291666,9.225,9.8166685,9.966667,11.406251,10.633334,5.2250004,2.1833334,1.1062499,1.4,1.7666668,1.8999999,1.5333334,0.76874995,0.475,0.75624996,0.7166667,0.91249996,1.6916667,3.516667,6.0937505,8.458334,8.725,9.116667,8.206249,7.1249995,5.825,3.8874998,2.4583333,1.2750001,1.05,1.9812502,3.4750006,3.9833336,3.475,1.3916667,0.23750001,0.0,0.0,0.0,0.0,0.0,0.13333334,0.76875,1.4666667,2.1,2.7583334,2.1125002,0.76666665,0.058333337,0.118750006,0.375,0.29375,0.11666667,0.1875,1.075,2.5875,2.7333333,1.8500001,2.175,2.0500002,1.9937501,1.8249999,1.55,1.2416667,1.0666666,0.50625,0.275,0.225,0.09166667,0.1,0.64166665,2.425,5.0312495,7.2,8.006249,5.5499997,1.8625,1.2083334,0.98125,1.1750001,1.3,1.3125001,0.8833334,0.4375,0.16666669,0.06250001,0.0,0.05,0.375,0.16666667,0.081250004,0.116666675,0.91875005,2.1083336,2.0625,1.3,0.575,0.40625,0.56666666,0.9187501,1.125,0.41875,0.125,0.050000004,0.4625,1.175,1.825,1.3666667,0.975,0.13333334,0.0,0.0,0.0,0.0,0.175,0.112500004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.75,0.5166667,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.175,0.21875,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3875,1.5916667,2.09375,1.4583334,0.6666666,0.15625,0.13333333,0.7875,1.1166667,0.39999998,0.6666667,4.3999996,3.8000002,5.6,7.1625004,5.5416665,4.21875,14.033333,18.475,12.166667,10.016666,12.4375,13.400001,16.58125,16.125,11.437501,18.841667,17.83125,11.766667,0.9583334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.0,1.6416668,3.4,4.9333334,6.641667,10.111111,9.808333,10.3111105,10.141667,8.566667,7.644444,8.325001,11.733333,14.691667,13.022223,9.908334,8.444445,9.133333,12.877779,18.455555,22.250002,16.522223,5.8749995,1.8222221,1.2333332,1.9222221,2.7222223,3.4916663,2.9888887,0.75,0.0,0.083333336,0.5222223,1.7666667,4.5333333,8.422221,10.808334,12.599999,11.724998,8.700001,6.366667,5.2999997,4.5777783,2.983333,1.2222223,1.025,1.1333333,1.3416667,1.2111111,0.98888886,0.64166665,0.24444443,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,1.2444445,2.7416666,1.5222223,0.14444445,0.19166668,0.16666667,0.15,0.13333334,0.10000001,0.1,0.0888889,0.033333335,0.0,0.0,0.0,0.008333334,0.0,0.022222223,0.15,0.6,2.6333337,5.488889,5.283334,2.8222222,1.2583333,0.5444445,0.39999998,0.71666676,1.2444445,1.025,0.7,0.36666667,0.17777778,0.18888889,1.325,2.8111112,2.0083332,0.81111115,0.76666665,0.28888887,1.7583333,2.1555555,1.8222221,0.775,0.5888889,0.85,0.19999999,0.06666667,0.15555556,0.17777778,0.50000006,2.2333333,4.766667,4.4444447,6.983333,0.9666667,0.23333335,0.016666668,0.0,0.0,0.0,0.1,0.12222223,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.51111114,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.08888889,0.25833336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28333333,1.3111111,1.9083333,1.1222223,0.53333336,0.18333335,0.15555556,2.25,3.166667,1.7,0.26666668,0.8333334,1.8555557,3.8888888,3.125,2.3555555,2.7833333,8.5,10.525,13.044445,20.733335,18.708336,18.355553,25.033333,24.144447,20.025002,16.866667,12.125,4.6666665,2.022222,1.4666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0833334,2.122222,2.9,4.1,6.577778,6.0249996,7.166667,12.391666,15.766666,17.800001,21.866665,27.7,34.925003,29.488892,15.308333,13.777778,17.366669,24.82222,25.57778,21.316668,11.722222,2.325,0.8111111,0.96666664,2.4555557,3.3333335,3.0249999,1.1333334,0.7416667,0.8111111,4.7,9.766666,12.708334,11.455555,9.888889,7.8166666,7.033334,5.091667,4.288889,2.475,1.5777779,1.7777778,1.4250001,1.3777779,1.625,1.5888889,0.55,0.44444442,0.17777778,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15555556,0.2888889,0.108333334,0.2,0.2916667,0.5555556,1.9666667,4.1333337,3.3333335,1.3333334,0.54444444,0.25833333,0.21111111,0.15833333,0.33333334,0.40833336,0.5,0.24444446,0.48333335,1.5000001,4.1333337,4.4111114,2.0083334,0.32222223,0.05,0.42222223,0.9777777,1.0166667,0.8666667,0.6166667,0.6666666,0.32500002,0.11111111,0.06666667,0.36666667,1.7888889,3.8916667,4.4444447,13.05,3.0999997,0.022222223,0.0,0.0,0.0,0.0,0.0,0.055555556,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.85555553,1.0666667,1.0111111,0.62500006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.425,1.2444445,1.2416668,0.44444448,0.14444445,0.041666668,0.0,0.7,0.6888889,0.5833333,0.0,0.43333334,2.3,4.377778,3.1666665,3.711111,3.5250003,11.866667,15.35,19.766666,24.500002,20.566668,12.844444,10.85,10.188889,9.974999,11.011112,5.716666,0.76666665,4.2777777,8.700001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10833334,0.7,0.10000001,0.0,0.0,6.3124995,6.0999994,6.1499996,4.78125,3.3333337,2.3187501,1.8416668,3.09375,5.3916664,7.6,11.599999,13.933332,12.3375,9.675,9.375,16.05,26.25,31.416668,28.849998,14.825,7.116667,2.6,2.541667,5.4875,11.941667,13.975,14.98125,18.008333,19.150002,23.449999,24.631248,24.95,19.8875,12.933333,9.608334,6.575,6.958334,7.33125,5.941667,1.95,1.4666667,0.76666665,0.52500004,0.52500004,0.52500004,0.38333338,0.35,0.24166667,0.47500002,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.083333336,0.118750006,0.225,0.75,1.3333334,1.4375,0.28333333,0.28333336,0.10625,0.14166668,0.11875,0.083333336,0.050000004,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.075,0.058333334,0.0375,0.13333336,0.29375,0.9916667,2.4499998,2.1333334,0.9166666,0.58750004,1.1833334,2.11875,0.8,0.53125006,0.425,0.5500001,0.21875,0.108333334,1.1437498,2.4166667,4.2000003,3.075,1.9874998,0.9416667,0.425,0.98125,0.56666666,0.35625,0.175,0.69374996,0.55,0.225,0.125,0.42500004,2.2062502,2.8833337,5.98125,8.916667,2.9583335,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.1,0.0,0.0,0.0375,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.033333335,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.20625001,0.13333334,0.18125002,0.0,0.033333335,0.06875,0.20833336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,0.525,0.20000002,0.008333334,0.0,0.0,0.0,0.0,0.23333333,2.5624998,4.0666666,3.3875,6.1,3.3333335,8.83125,14.941666,9.7625,10.799999,11.425001,12.608334,10.366668,9.225,5.2333336,6.3375,7.333334,7.55,3.2833335,1.3437502,0.76666665,2.2583332,3.8187504,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0,0.46875006,0.49166673,0.0,0.0,0.0,3.7333333,3.5222223,4.4888887,4.2166667,3.8111115,4.9833336,7.288889,12.166668,14.933334,18.011112,14.966666,12.433334,11.225001,9.711111,12.233334,19.58889,25.266665,24.666668,14.755556,5.75,1.7444444,1.375,3.6111112,9.091667,21.17778,28.266668,34.825,33.211113,33.658337,31.88889,24.266668,16.655554,8.183333,3.8333335,2.3222222,1.3250002,0.9888889,1.325,2.3,2.0416667,1.7888889,1.6,1.2416667,0.9444445,0.52500004,0.35555553,0.15,0.15555556,0.13333334,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2888889,0.41666666,0.9888889,1.575,1.8333333,2.641667,3.2888892,2.8833332,0.94444454,0.70000005,0.45833337,0.29999998,0.18333335,0.0888889,0.025,0.011111111,0.0,0.075,0.18888889,0.20833333,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.15555556,0.38333336,1.0777777,0.8,0.4166667,1.6888888,4.333333,3.4888887,1.3333334,0.1,0.13333334,0.31666666,0.1777778,0.008333334,0.44444445,0.8083333,1.7777777,2.8833334,2.8222222,2.1444445,1.0250001,0.35555556,0.15,0.06666667,0.28333333,1.0111111,1.3666668,0.55833334,0.07777778,0.70833325,1.8,0.9666667,5.6111107,7.133333,0.44166666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.06666667,0.033333335,1.2111112,0.23333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.17500001,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.34444448,0.5083333,0.3,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.6666667,2.8750002,2.3000002,1.7916667,0.18888889,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.1000001,4.844445,6.666666,8.4,5.588889,4.216666,2.1000001,4.425,9.599999,16.358334,17.744444,19.044443,14.283333,9.422223,5.45,4.1333337,8.983334,1.8666667,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21111111,0.2,0.0,0.0,0.0,0.0,0.0,0.92499995,2.2833333,3.3416667,4.5874996,4.991667,5.24375,5.116667,4.7500005,3.2416668,2.875,2.2187502,3.3083334,3.65625,3.6833334,5.0625,7.866667,8.2375,7.016667,3.2500002,2.15,2.9333334,8.925001,15.216667,19.53125,24.933334,29.483335,26.168747,22.508333,17.1375,10.391667,7.4624996,5.05,4.58125,5.433333,9.958334,12.756248,9.724999,8.46875,4.325,2.9625,1.8083334,1.7416667,0.9250001,0.43333334,0.15000002,0.0,0.06875001,0.083333336,0.075,0.043750003,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.9875,3.566667,5.2,6.4375,7.225001,7.1812496,7.2,6.6624994,5.6833334,4.3375,2.8499997,1.7083333,0.78125006,0.3416667,0.10625,0.050000004,0.03125,0.083333336,0.025,0.15000002,0.3166667,0.70625,0.6583334,0.88125,0.9083333,0.71666664,0.28125,0.0,0.13749999,0.775,1.2812501,1.2166666,0.9,0.3416667,0.21666667,0.63750005,2.025,4.6125,6.2250004,5.225,3.4166665,1.975,1.1,0.325,0.70000005,0.6333333,0.01875,0.33333334,0.55,1.4583333,1.7583334,1.4687501,0.93333334,0.3125,0.75833327,0.45000002,0.25833333,0.51666665,1.0625001,0.76666665,0.20000002,0.325,0.13125001,0.9416667,1.675,0.78125006,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.05,1.2,0.99375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.20625001,1.7666668,2.6312501,1.4916667,0.0,0.0,0.0,0.0,0.108333334,0.70624995,1.025,0.74375,1.2,1.1083333,0.11875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.7375,1.2083333,1.09375,0.083333336,0.0,0.0125,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.425,4.291667,1.7375001,1.3083332,2.9687505,4.2083335,5.0333333,7.3,6.3416667,4.3375,13.0,17.74375,16.25,12.583334,10.6625,10.766666,5.3875003,7.1666675,3.35,0.26666668,0.1875,8.366666,10.391667,6.9375,4.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,14.474999,12.555555,11.911112,8.85,3.8666668,1.2583333,0.3888889,0.43333334,0.81111115,1.1555555,1.5749999,1.4222221,1.1416667,1.2111112,0.85,0.34444445,0.22500001,0.88888896,1.5555556,2.6333332,5.2333336,11.341666,24.700003,26.366667,21.711111,17.3,11.058332,5.3777776,1.4250002,0.33333334,0.9333334,1.3888888,3.3083334,5.6555557,7.7333326,10.908333,14.48889,8.991667,5.322222,3.4666667,3.477778,2.5777779,1.4999999,1.3555558,0.9333333,0.022222223,0.041666668,0.06666667,0.1,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,1.0166667,4.533334,7.7555566,8.533334,11.822223,10.0,9.28889,7.075,6.088889,6.5250006,6.377778,5.5555553,4.666667,3.1888888,2.3166666,1.6111112,1.1999999,1.0333333,0.6222222,0.2916667,0.055555556,0.033333335,0.24444446,0.91666675,1.6444445,2.4,1.9666665,0.6333334,0.2916667,0.6111111,0.65833336,0.37777776,0.33333334,1.2444444,0.8888889,0.82500005,0.8,1.3249999,2.0444446,3.75,3.6888888,2.8333335,2.5666666,1.9333333,1.3416667,0.9777778,0.8833334,0.1777778,0.1,0.56666666,1.2,1.05,0.18888888,0.59999996,0.48888892,0.4833333,0.22222224,0.1,0.19166668,0.72222227,0.825,0.24444443,0.041666668,0.0,0.0,0.5833333,0.4222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22222224,0.57500005,0.34444445,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.39166668,0.2,0.65555555,0.15833333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7333333,3.0083332,0.7888888,1.7833333,5.366667,1.188889,2.9333336,3.9333334,12.35,3.7111113,2.675,2.0888891,0.6,0.0,3.466667,2.1333332,1.3555557,0.116666675,0.11111111,2.9833336,11.266666,14.566667,10.358334,6.2333336,0.050000004,0.0,0.06666667,0.36666664,0.36666667,0.0,0.0,0.0,0.0,0.12500001,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,22.987503,18.516666,15.875002,10.474998,5.091666,2.36875,1.4499999,2.1000001,3.4333334,4.0416665,4.9125,5.366667,6.9375005,5.6416664,4.46875,4.508333,6.875,8.591666,11.475,12.975,18.208332,23.1625,21.875,14.975,10.191668,7.058334,4.3625,2.4583333,1.7812499,2.6333334,4.15625,6.05,10.349998,16.375,20.833332,22.81875,18.866667,13.26875,11.6,11.1125,6.474999,2.9833336,0.90624994,0.60833335,0.34375,0.25833336,0.18125002,0.06666667,0.025,0.00625,0.058333337,0.10000001,0.25833333,0.31875002,0.30000004,0.2625,0.12500001,0.0,0.0,0.0,0.0,0.0,0.1125,0.77500004,1.6083332,1.4125001,2.8583336,3.0312502,1.3166667,1.025,0.65000004,0.4,0.3,0.3833333,0.45,0.6666667,0.47500002,0.38333333,0.2125,0.08333333,0.05,0.0375,0.041666668,0.0,0.016666668,0.13125001,0.108333334,0.48333332,1.0000001,1.4166667,0.59999996,0.35833335,0.7,0.9833333,1.33125,2.3416667,2.816667,3.1937501,4.25,5.7375,6.1916666,4.7375,4.266667,4.466667,4.3750005,3.15,4.5875,4.2666664,1.325,1.5416667,1.3312501,0.91666675,0.4583334,0.5875,1.2833334,1.16875,0.85833335,0.65,0.125,0.05,0.08125001,0.13333334,0.40625,0.6999999,0.33749998,0.075,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.36875,0.35000002,0.025,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17500001,0.08125,0.0,1.2625,2.6999998,1.5625,2.425,1.1500001,1.075,5.3166676,10.19375,6.558333,0.59999996,0.45,0.15,0.0,0.0,0.0,0.033333335,0.21249999,1.0,3.25,3.6750002,5.875001,4.3437505,1.2750001,2.5375001,10.016667,0.056250002,0.6666667,3.0333333,0.2625,0.041666668,0.043750003,0.21666667,0.425,0.23333335,0.041666668,0.0,0.0,0.0,0.0,0.0,37.15,25.800001,14.777778,7.533334,3.8666666,2.591667,4.8,9.091667,11.48889,11.044445,9.225001,6.477778,8.183333,7.866667,8.799999,8.933334,9.791666,14.222222,18.766666,23.008333,18.1,11.733333,7.8888893,6.7666674,5.7888894,6.5111113,10.533333,16.488888,17.583334,17.6,20.508335,19.800001,19.508333,21.433334,27.322222,28.583334,26.300003,16.891666,4.533334,2.3666668,2.6555557,4.5444446,4.775,1.0333333,1.5083334,1.2111111,0.89166665,0.25555557,0.84444445,1.0666667,1.0888889,1.0583334,0.7111111,0.42499998,0.16666669,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108333334,0.2777778,0.4333333,0.25555554,0.425,0.39999998,0.16666669,0.0,0.17777778,0.041666668,0.0,0.12500001,0.39999998,0.59166664,0.5111111,0.44444448,0.6750001,0.67777777,0.325,0.13333334,0.016666668,0.044444446,0.12222223,0.14166667,0.07777778,0.016666668,0.055555556,0.116666675,0.33333334,1.275,2.3888888,4.2444444,8.033334,11.200001,12.283333,13.144444,15.075001,15.511111,13.933332,13.400001,9.966667,5.8583336,5.9888887,5.925,3.088889,2.6,1.9666667,0.61111116,0.18333334,0.055555556,0.6333333,1.9111111,1.2666667,0.6777778,0.34444445,0.36666667,0.26666665,0.108333334,0.3222222,0.4583333,0.34444442,0.16666667,0.0,0.0,0.0,0.0,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19166666,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.1,0.23333332,1.425,2.155556,0.9333334,0.15,0.06666667,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14444444,0.108333334,0.0,1.2166667,4.177778,4.9166665,3.6666667,0.88888896,2.2833335,7.088889,6.6,3.2666667,0.40000004,0.044444446,0.06666667,1.6166668,4.933334,3.5750003,0.0,0.53333336,3.577778,7.275,3.3666668,1.0111111,0.29166666,0.033333335,0.0,2.277778,0.0,0.47777778,1.7444444,1.5749999,0.5666666,0.34166664,0.36666667,0.73333335,0.45555556,0.0,0.0,0.0,0.0,0.0,0.0,17.758333,7.211111,3.9888892,1.5416667,0.76666665,1.2583333,2.9555557,4.883333,5.5555553,4.266667,3.0583332,2.3444448,2.9166667,3.4333336,3.55,6.166667,12.475,28.866667,31.97778,21.525,12.244445,7.4,7.2555556,8.733334,10.888887,16.122223,23.841667,28.133335,26.59167,25.233335,24.925001,23.866667,24.175,22.744446,24.955555,22.825,16.844444,2.15,1.5666667,1.9666667,6.111111,7.055556,6.491667,8.144445,7.0333333,4.288889,1.9749999,4.611111,2.1666665,1.6,0.46666664,0.15,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.06666667,0.116666675,0.14444444,0.14166667,0.06666667,0.025,0.0,0.022222223,0.025,0.011111111,0.0,0.05555556,0.4666667,0.8333333,1.0333334,1.45,1.4222223,0.7083334,0.05555556,0.0,0.0,0.0,0.008333334,0.08888889,0.033333335,0.0,0.0,0.0,0.37499997,1.5222223,3.488889,7.1250005,10.133333,14.9,18.288889,20.075,24.522224,31.022224,34.541668,32.733334,14.825001,7.1555557,6.8499994,5.5777783,4.125,2.5111113,1.2888889,0.5416667,0.13333333,0.34166664,0.5666667,1.35,2.0555556,1.6555555,0.975,0.9333334,0.275,0.7777778,1.1166667,0.6888889,0.42222223,0.175,0.033333335,0.0,0.0,0.0,0.26666665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7583333,1.5555555,0.18333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.011111111,0.0,0.3555556,2.177778,0.18333335,0.07777778,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,1.3416667,2.6777778,4.883334,6.477778,3.7111115,1.4916667,3.322222,2.8083334,1.7444446,0.70000005,0.26666668,0.0,7.6499996,25.033333,5.833334,2.4666667,4.3166666,2.4,3.0,9.922222,3.4222221,1.8916667,0.13333334,0.0,0.0,0.30833334,0.7555555,2.733333,1.5416666,0.26666668,0.57500005,0.84444445,0.8166667,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,3.7624998,1.3833333,0.64166665,0.47500002,0.9583333,1.35,2.4333334,2.7000003,1.9250001,1.2916666,1.10625,1.3666668,1.4937501,2.4583335,4.1625004,11.175,20.28125,19.191666,15.033334,11.9,12.875,12.912499,13.216668,18.43125,27.800001,32.683334,37.893753,36.85,34.056248,34.0,28.268751,23.758335,16.1625,7.741667,5.583334,2.8562503,2.6166668,5.6375003,8.95,12.625,11.391666,10.166666,7.2812495,4.0,1.6187501,0.8166667,2.4625,3.4250004,1.5416667,0.3375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.112500004,0.42499998,0.425,0.3,0.14999999,0.043750003,0.0,0.0375,0.30833334,0.6625,0.6833334,0.25000003,0.20833334,0.17500001,0.15625001,0.125,0.00625,0.0,0.00625,0.30833334,1.1333333,1.75625,1.375,0.66875005,0.29166666,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108333334,0.30625,0.68333334,2.5416667,7.825001,12.933333,19.599998,22.816666,25.0375,22.483335,22.041668,27.275,29.116667,24.006252,18.225,7.5,7.075,7.66875,4.3916664,2.3500001,0.51250005,0.225,0.50625,0.43333337,0.9187501,1.25,1.5583334,2.6437502,1.8333334,1.3062501,1.0666667,1.7750001,2.6833334,2.3583333,0.63750005,0.05,0.0,0.075,0.03125,0.116666675,0.06875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,2.3,1.79375,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2916667,0.0,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.112500004,0.29999998,0.0,0.0,1.45625,3.8500004,7.8812494,3.4333334,1.8166671,2.21875,2.9666667,0.5375,0.45833337,0.6125001,0.88333344,0.5,0.05,1.8166668,3.18125,4.8333335,2.2,0.53333336,0.05,0.975,0.20000002,0.0,0.0,0.06875,0.8166667,2.1000004,3.6750002,5.6916666,5.375,0.3333333,0.575,0.4666667,0.13749999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.45555556,1.5555556,1.8416667,3.1777775,4.783334,4.811111,3.85,2.9444444,1.4333333,2.7166667,5.0111113,5.3083334,9.333334,16.141666,19.955553,14.925,12.622223,10.788889,10.966666,15.58889,24.166666,37.17778,50.725,48.81111,41.73333,34.441666,24.944445,20.95,16.233335,9.641667,4.5222225,3.7833333,3.5333333,2.9777777,2.6833334,3.2111113,5.2749996,8.822222,8.791667,5.633333,2.5,0.89166665,0.17777778,0.016666668,0.0,3.1583333,6.0000005,6.3777776,0.9250001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.022222223,0.033333335,0.055555556,0.09166667,0.022222223,0.008333334,0.86666673,0.72222227,0.6333333,0.5888889,0.29166666,0.11111112,0.24166667,0.51111114,0.26666668,0.25833333,0.26666668,0.15833335,0.011111111,0.050000004,0.0,0.011111111,0.30833334,0.5,0.43333334,0.11111111,0.06666667,0.13333334,0.26666668,0.45555556,0.7222223,1.7166668,3.5111113,11.050001,21.166668,27.441666,29.766666,25.855556,22.766666,21.38889,20.275,12.677778,5.133333,3.8555555,7.9166675,8.566667,5.133333,1.7916666,0.46666667,0.40833336,0.13333334,0.5,1.0777779,1.8444445,1.9083333,2.8111112,2.266667,1.2,1.5833333,2.5666664,5.2888894,5.7583337,3.0,0.27499998,0.12222222,0.26666668,0.07777778,0.09166667,0.08888889,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12222222,2.7916667,1.2888889,0.13333334,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.39999998,0.0,0.0,0.0,0.0,1.6000001,0.93333334,1.2333333,2.916667,6.188889,0.6666667,0.42222223,0.36666667,0.9333334,0.97777784,3.1,3.2444444,5.2333336,0.0,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.32500002,2.8000002,2.9250002,5.7,8.5,4.4083333,0.45555556,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.25833336,0.0,0.06666667,0.6333333,2.45,5.425,5.6812496,4.2250004,2.05,2.9583333,4.45,5.4687505,8.808334,16.206251,23.800001,23.80625,16.250002,10.39375,7.8166666,8.233334,12.381249,19.416668,24.443748,26.85,24.4125,19.008333,18.033335,18.78125,13.816667,7.6,5.108333,5.3999996,5.15,4.8125005,6.625,6.941667,6.54375,1.7833334,1.2375,2.1583333,2.0625,1.1166666,0.60833335,0.22500001,0.275,2.1000001,4.9333334,7.98125,9.049999,2.0916667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.043750003,0.16666667,0.34375003,0.5333333,0.6374999,0.44166666,0.2,0.05,0.016666668,0.056250002,0.13333334,0.19375001,0.108333334,0.11250001,0.15833333,0.21666668,0.19375001,0.16666669,0.125,0.5750001,0.4125,0.30000004,0.3083333,0.60625,0.82500005,0.8,1.0416667,1.3625,1.9083334,1.3875,1.5416666,2.1333332,2.3750002,1.1166667,2.1875,7.175,11.16875,16.458334,17.808334,13.36875,9.683332,11.69375,13.641666,11.51875,6.4416666,4.1687503,5.25,9.833333,8.212501,3.3666668,1.10625,0.425,0.29375002,0.56666666,0.85833335,1.2687502,1.8333333,2.15625,2.3333333,1.49375,1.1499999,1.5583334,4.675,8.750001,7.35,2.0,0.51250005,0.6,0.42499998,0.09166667,0.10000001,0.056250002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06250001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.375,3.7833333,2.5125,2.4083333,0.675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28333336,0.9437501,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.075,2.78125,1.9000001,4.6749997,1.3333334,0.16250001,0.43333334,0.7666667,4.4,11.033333,5.725,0.0,0.0,0.0,1.1,0.0,0.0,0.0,0.0,0.0,0.15,0.9625,1.6583333,2.6750002,1.0687499,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.44166666,2.63125,0.0,0.0,0.14444445,0.825,1.5555556,1.025,0.4666667,0.81666666,1.7111111,3.3888888,6.4750004,11.366667,12.291667,11.077778,12.2,12.133334,13.425,13.344445,15.655556,16.458334,16.722223,17.108334,16.588888,16.966667,17.47778,15.211111,9.683333,4.9555554,5.1,6.7666674,6.1833334,5.3555555,7.758333,8.466667,7.9555564,5.1916666,3.7111113,3.2166672,2.9,3.3999996,2.7222223,1.4555557,0.40833327,0.2888889,0.60833335,1.4222223,0.6916667,0.15555555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.055555556,0.14166667,0.11111112,0.16666669,0.11111111,0.22500002,0.27777776,0.6222222,0.55833334,0.22222222,0.1,0.3666667,0.6583333,1.0888889,1.1444445,1.025,1.5666666,1.8749999,3.4222221,5.4083333,7.6444445,7.125,5.7888894,3.9000003,2.5000002,1.3777778,0.51666665,0.51111114,0.87500006,2.5,4.5444446,3.7416668,4.7777777,5.091666,5.1,6.108334,6.2666664,3.85,2.4444447,2.011111,6.8250003,9.844446,5.5833335,2.2333333,0.84166676,0.32222223,0.54444444,0.8833334,1.1111112,2.0083332,1.577778,2.2166665,1.5222222,1.3555555,1.9166669,4.2777777,6.725,8.277778,2.9750004,1.7777779,3.1000001,2.488889,0.9555556,0.475,0.31111112,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14166668,0.12222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0500001,10.977778,3.7333333,5.6555557,3.6222224,0.5833333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2166667,0.11111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39999998,1.9916667,1.7111111,1.7,0.9111111,0.008333334,0.0,0.0,0.0,0.0,0.15,0.13333334,0.0,0.0,1.7833333,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15833335,1.2555555,1.5416666,0.0,0.0,0.0,0.0,0.083333336,0.225,1.0583334,3.3062499,6.4583335,7.741667,11.262501,14.341667,17.975,20.841665,22.006248,26.95,23.293749,18.0,17.466667,20.81875,22.46667,19.637499,22.25,20.693748,12.216667,6.2416663,6.0687504,8.941667,13.831251,17.025,9.418751,8.174999,8.21875,6.2916665,4.041667,6.231251,9.016666,10.91875,7.366667,3.7500002,0.76666677,0.083333336,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.6750001,0.7166666,0.0375,0.083333336,0.225,0.20000002,0.06666667,0.025,0.15833335,0.35625008,0.59166676,1.125,2.01875,4.1333337,6.41875,6.55,6.0875,6.8583336,8.668751,8.808333,6.616667,3.4375002,1.2416667,0.64375,0.80833334,0.84375006,0.6333334,0.9249999,1.06875,1.3583332,1.21875,1.2916667,1.2062501,2.1083333,2.0812502,2.575,2.2,1.68125,3.616667,6.1937494,6.083334,3.3249998,1.0333333,0.35833338,0.3,0.6666667,0.9312501,1.3333334,1.2937502,1.8333334,1.9833332,1.29375,1.4583333,3.0,6.708333,7.3,4.066667,4.90625,6.875,6.816667,4.59375,1.9333335,0.70000005,0.116666675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11250001,0.3,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0666666,1.9624999,1.3083334,3.4083333,1.5125,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.71250004,0.79999995,1.56875,0.6,0.95,0.9,1.4833333,0.75,0.71666664,1.05,0.48333335,0.0,0.0,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.6875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.15555556,0.5333333,1.5777779,2.7166667,3.077778,3.8833332,6.077778,11.08889,19.675001,30.888891,36.91667,43.455555,49.89167,48.188892,35.499996,27.611113,25.977777,22.166668,25.055557,25.233337,21.522224,16.233335,9.244445,7.0888886,8.241666,11.0222225,15.091666,5.2666664,3.6583333,6.411111,9.941667,12.155556,17.011112,21.158333,16.2,6.225,0.7222222,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.25555557,0.0,0.14444444,0.45555556,1.5666666,3.1333334,1.0583334,2.4444444,2.8666666,3.2222223,4.111111,4.1833334,1.0444446,0.025000002,0.0,0.29999998,1.7555555,2.5,1.8166666,1.5111113,3.4333334,5.0333333,5.216667,2.9444447,3.8833334,8.377778,11.911112,10.933334,8.522222,6.3500004,5.8444443,2.4166667,1.1222223,0.6888889,0.26666668,0.58888894,0.9833333,1.0666667,0.87500006,1.0777777,0.74166673,0.6888889,1.0222223,1.2833334,1.4222224,2.6833334,3.6000001,4.3666663,3.1111112,1.8222222,0.4666667,0.07777778,0.34166667,0.6111111,0.48333335,0.51111114,1.2888889,1.5083333,0.6111111,0.85833335,3.722222,6.908334,7.3888893,6.4833336,9.366668,8.188889,7.4416666,8.177777,3.3416667,0.37777779,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.044444446,0.0,0.0,0.016666668,0.21111113,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,0.2,0.2,0.36666667,0.1,0.0,0.05,0.033333335,0.0,0.11111112,1.1333334,1.6999998,0.2888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.022222223,0.5833334,3.0444446,3.125,10.8,13.866666,7.2666664,2.411111,1.7333333,0.68888885,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.31666666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.21666667,0.64166665,2.4312499,8.4,14.787499,25.041666,19.63125,22.249998,27.583336,34.675,42.108337,49.78125,59.008335,57.324997,51.691666,40.699997,34.725002,33.141666,30.631248,36.708336,25.65625,15.041668,9.8,5.8833337,5.3500004,5.06875,8.1,9.375,11.041667,10.9,11.341666,15.1375,19.2,22.891665,18.45,7.675,2.35625,0.95000005,1.05625,1.1833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18333334,0.8125,0.6166667,0.15,0.041666668,0.13750002,0.8666666,0.53749996,0.43333334,0.55833334,2.275,6.2833343,4.35,1.3166667,0.96250004,2.1750002,4.45,6.5000005,7.3250003,4.59375,2.3166666,1.0749999,1.45,1.3416666,1.0187501,0.90833336,2.525,6.933334,10.1625,9.375,7.0375004,5.0583334,7.875001,12.006251,14.641666,15.4875,15.475,9.943751,3.5333338,1.8499999,1.63125,1.3666666,0.41875,0.2166667,0.25,0.625,0.9187499,0.7166667,0.6583334,0.65625006,0.7083334,1.6875,3.483333,3.5375004,3.3083334,2.7749999,2.65625,1.1750001,0.43125,0.30833334,0.49374998,0.45833337,0.48333335,0.7187499,0.75,0.49375,0.50000006,3.11875,6.45,7.63125,8.533333,10.216667,8.88125,7.525001,8.75,2.85,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.27499998,0.39999998,0.0,0.0,0.025,0.32500002,0.17500001,0.00625,0.0,0.0,0.0,0.0,0.0,0.38125002,0.44166672,0.116666675,0.043750003,0.0,0.24375,0.058333334,0.0,0.058333337,0.55,1.31875,0.7916666,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20000002,1.1750001,2.0166667,2.6,3.2416666,4.9812503,15.525,17.233334,8.23125,2.375,0.875,1.0333333,0.625,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.112500004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.6,3.0888891,6.408334,7.9555554,14.508333,23.155556,33.408333,43.522224,51.799995,54.691666,55.65556,59.4,61.500004,57.675,62.622223,50.733337,39.77778,33.744442,28.916668,22.222223,14.291667,7.666667,4.6250005,7.744445,7.8888893,8.099999,9.411111,11.974999,10.5222225,11.083334,15.833334,19.741665,18.68889,15.28889,5.5833335,2.188889,1.5500002,0.92222226,1.35,0.8000001,0.4666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.016666668,0.0,0.0,0.0,0.0,0.05,0.3777778,0.44999993,0.32222223,0.32500002,0.17777778,0.083333336,0.15555558,0.0888889,0.14999999,1.3000001,2.65,2.177778,0.80833334,0.34444445,0.055555556,0.15,0.5777778,2.2500002,3.377778,1.8,1.3222222,1.2333333,0.525,0.6777778,1.8333334,4.822222,8.766667,12.6888895,12.874999,10.177778,5.1555557,4.2500005,8.655557,13.808334,15.788889,11.2,5.7555556,3.2444446,2.9166665,3.4,1.3083334,0.45555556,0.3416667,0.2888889,0.2916667,0.5555555,0.9666667,0.6416667,0.5666667,1.1666667,2.8555558,5.575,4.9777775,3.1777778,3.6750004,5.2000003,4.266667,1.3111112,0.38333336,0.42222223,0.6333334,0.4166667,0.3888889,0.8500001,0.92222226,0.47500002,1.8555557,5.3333335,10.222222,8.155556,9.791667,8.711111,6.108333,8.344444,1.4666668,0.20000002,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.025,0.17777777,0.2888889,0.48333332,0.37777776,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7166667,1.0888889,0.10000001,0.0,0.016666668,1.1,1.0555556,0.125,0.0,0.0,0.0,0.0,0.0,0.041666668,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44444445,0.9416666,0.9000001,0.15833335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,1.4666667,1.5111111,0.65,0.45555556,1.3500001,1.4666666,1.0888889,0.45000002,0.26666668,0.0,0.4888889,1.0333334,0.4222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.275,1.2444446,3.3444448,5.9083333,8.233334,16.308334,26.777775,41.84167,53.81111,62.31111,64.4,56.86667,49.06667,40.91111,39.516666,38.444443,29.016666,26.366669,24.733334,20.733334,11.777778,9.408334,9.444445,9.649999,9.533334,11.955556,15.166667,13.422223,13.258333,15.544445,19.366667,23.922224,23.533335,13.633333,2.6111112,0.90833336,0.5222222,1.3249999,2.7222223,1.9,1.3888888,0.76666665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.17777778,0.15,0.17777777,0.13333333,0.0,0.0,0.0,0.033333335,0.13333336,0.14444445,0.14166667,0.10000001,0.20833334,0.022222223,0.0,0.008333334,0.055555556,0.1,0.31111112,0.7333333,1.0666666,0.44444448,0.38333338,0.24444444,0.125,0.15555555,0.6583334,0.86666673,0.88888896,0.18333334,0.044444446,0.36666667,1.9555556,4.2500005,6.933334,10.525,12.655556,11.9,4.8416667,1.3333335,2.5,3.6000004,5.083333,6.533334,7.9222226,6.5583334,3.4333334,1.2083334,0.53333336,0.68333334,1.2777777,0.6166667,0.23333335,0.47777775,0.9083334,0.5555556,0.8833334,1.8222222,2.5083332,4.577778,4.5888886,3.5833335,5.6444445,9.758334,6.5888886,1.4250001,0.4666667,0.56666666,0.7,0.17777778,0.35833338,1.0111113,2.0916667,0.53333336,2.0416667,6.122223,9.977778,7.416667,8.444445,6.5,5.422222,4.1833334,1.0555556,0.47777778,0.0,0.0,0.0,0.0,0.008333334,0.044444446,0.0,0.11111111,0.79999995,1.4666666,1.522222,1.0333334,0.2888889,0.05,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0916666,1.5555557,0.24166667,0.0,0.0,0.3111111,1.2444444,0.46666667,0.21111111,0.375,0.0,0.0,0.0,0.0,0.0,0.05555556,0.041666668,0.011111111,0.0,0.0,0.0,0.0,0.044444446,0.3333333,0.25555554,0.041666668,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.0,0.0,0.26666668,0.13333334,0.0,0.33333334,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,0.0,0.0,1.2437501,1.825,3.4333334,4.90625,8.125,16.55,24.058332,30.112501,44.875,55.533337,58.8125,56.741673,52.381252,37.225,23.862503,21.35,20.018751,18.283333,13.983333,11.556251,9.408334,9.1625,15.525,15.393749,27.791668,28.575003,29.525,29.741669,26.625,19.824999,20.199999,16.241669,8.2,2.3833334,0.025,0.05,0.4166667,2.25625,3.3250003,3.04375,0.575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0125,0.0,0.041666668,0.025,0.050000004,0.3125,0.28333333,0.4375,0.57500005,0.625,0.1875,0.25000003,0.0,0.008333334,0.056250002,0.091666676,0.175,0.09166667,0.033333335,0.01875,0.008333334,0.03125,0.083333336,0.1625,0.5083333,0.68333334,0.57500005,0.108333334,0.33750004,0.26666668,0.33749998,0.05,0.0,0.03125,0.16666667,0.03125,0.06666667,0.43124998,0.89166677,1.7375,2.0666666,4.308334,5.5375004,2.1833334,0.70000005,0.41666666,0.59375,1.6666669,3.791667,4.1937504,2.033333,0.2875,0.14166668,0.69375,1.7750001,1.2250003,0.95000005,0.125,0.14375001,1.0583334,1.3937501,1.2083334,1.575,1.9666666,4.741667,6.94375,5.175,6.1812506,9.683334,6.7687507,2.6833334,1.0583334,0.36875004,0.68333334,0.3125,0.3,1.65,2.8833337,0.9125,1.5666666,4.8083334,7.45,5.25,6.6624994,3.5833335,2.3625,1.3249999,0.8249999,0.3375,0.008333334,0.0,0.0,0.0,0.0,0.0375,0.041666668,0.24999999,1.5875,3.0749998,3.1312501,2.2333333,1.0375,0.3166667,0.15,0.0375,0.05,0.0,0.0,0.0,0.116666675,0.25625002,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.55,2.3666668,0.51874995,0.0,0.0,0.0,0.0,0.0875,1.2833333,2.06875,1.7250001,0.0,0.0,0.0,0.73333335,0.9333334,0.8375,0.32500002,0.0,0.0,0.0,0.28333333,0.25833336,0.00625,0.0,0.0,0.0,0.075,0.1,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.0,0.1875,0.63333327,0.51666665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.1625,0.0,0.0,0.39166668,1.1888889,4.1777782,6.65,7.8,13.866668,23.533335,21.325,28.744446,47.76667,49.650005,48.144447,44.658337,28.644447,20.949999,19.333334,17.041666,13.066667,9.366667,6.0249996,6.1888885,15.016666,24.955555,30.466665,32.877777,28.82222,34.23333,32.022224,22.041668,13.244444,9.058332,1.1,0.008333334,0.022222223,0.2,0.033333335,0.41111112,1.3833334,2.8333333,1.2166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.044444446,0.15833335,0.06666667,0.011111111,0.11666667,0.25555557,0.45000002,0.56666666,0.9416667,0.6333333,0.41111112,0.86666673,0.31111112,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.058333334,0.13333334,0.05,0.0,0.108333334,0.16666666,0.37777779,0.8333334,0.41111112,0.2916667,0.14444445,0.6333333,0.9,0.6333334,0.27500004,0.011111111,0.041666668,0.0,0.10000001,0.22222222,0.16666667,0.47777778,0.53333336,0.6833334,0.82222223,0.275,0.055555556,0.0,0.0,0.0,0.0,0.022222223,0.041666668,0.111111104,0.09166667,0.15555556,0.45833334,0.8222222,0.17777778,0.025000002,0.53333336,2.15,2.1666667,0.8500001,1.0444444,1.5666667,4.9500003,7.2000003,5.708333,4.766667,7.058334,5.3333335,3.8222222,1.225,0.5444445,0.5416667,0.1888889,0.23333335,1.0888889,1.2,0.33333334,0.6444444,3.1166668,3.7333336,3.5833335,4.4666667,1.2583332,1.7222222,1.7666667,0.83333325,0.15555556,0.016666668,0.0,0.0,0.0,0.0,0.033333335,0.12222223,0.35,2.1333332,4.5,5.244445,3.3916667,1.8666667,0.58888894,0.44166672,0.5,0.0,0.0,0.0,0.35555553,0.49166667,0.25555554,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.0166667,3.2555556,0.76666665,0.0,0.0,0.0,0.0,0.34166667,2.822222,3.6083333,4.711111,0.0,0.0,0.0,3.1666665,1.5333334,1.6833333,0.24444446,0.0,0.12222222,0.025,0.66666675,0.6222223,0.0,0.0,0.0,0.0,2.0333333,0.7111111,0.12500001,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20000002,0.93333334,0.5333333,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.0,0.0,0.0,0.125,0.79166675,1.8333334,3.6125,5.366667,15.062499,13.325001,15.35,20.983334,34.266666,32.91875,28.633335,24.81875,20.083334,17.931252,14.216667,13.14375,8.9,6.2416663,9.45,17.358332,26.90625,28.133331,29.39375,32.633335,33.725,33.1125,24.291668,11.312501,4.7000003,0.9375,0.11666667,0.60625,0.6333333,0.25000003,0.025,0.21666665,1.075,0.625,0.056250002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09375001,0.22500001,0.1875,1.0166667,1.8500001,3.7,5.3583336,0.83124995,0.575,1.0187501,0.8166667,0.14166668,0.0125,0.008333334,0.056250002,0.075,0.0125,0.018181818,0.0,0.05,0.036363635,0.0,0.0,0.16875,0.475,0.66249996,1.1833334,0.55833334,0.5625,1.1500001,1.08125,0.6333333,0.21875001,1.0083333,1.7083335,1.95,1.0,0.0625,0.0,0.16250001,0.60833335,0.99375,0.2916667,0.25833333,0.10625,0.05,0.01875,0.0,0.0,0.0,0.0,0.0,0.1,0.275,0.29166666,0.28125,0.69166666,0.11875,0.075,0.016666668,0.0,0.083333336,0.88750005,1.8083333,2.0375,0.87500006,1.0999999,1.9625,4.7,6.7312503,6.1166663,5.5874996,5.291667,5.708334,4.25625,2.2749999,0.70000005,0.40000004,0.13125001,0.15833335,0.34375,0.058333334,0.033333335,0.4625,1.0833334,1.0062499,2.25,0.9312501,0.4416667,1.1583333,1.8500001,0.48333335,0.056250006,0.05,0.0125,0.0,0.0,0.016666668,0.13333334,0.33125,0.38333336,2.4437501,6.3999996,7.31875,5.0916667,2.9416664,1.05625,0.9166666,0.1875,0.0,0.0,0.21666668,0.75000006,0.28333333,0.27500004,0.025,0.0,0.0,0.0,0.0,0.0,0.0,2.41875,3.7916667,0.9250001,0.0,0.0,0.0,0.21666667,1.7125,2.1166668,3.7875,0.53333336,0.0,0.0,1.6125001,1.325,1.1083333,0.65000004,0.075,2.5875,1.5666667,0.0,1.1583333,0.8666666,0.0,0.0,0.05,2.8000002,3.125,0.0,0.112500004,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.375,1.15,0.7,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777778,0.24444446,0.6083334,4.4666667,9.908334,12.011111,14.758334,17.1,16.511112,13.8,13.700001,13.516667,15.300001,14.858335,11.666666,7.691667,4.2555556,5.8,12.808333,16.055557,23.916668,22.78889,22.816668,29.977781,29.288889,21.150002,9.566667,3.5333338,0.0,0.05,0.6,0.625,0.08888889,0.0,0.48333335,0.67777777,0.39166665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777778,0.25833336,0.72222227,2.6916666,2.3222225,1.5111113,2.1833336,0.14444444,0.6583333,0.0,0.016666668,0.011111111,0.044444446,0.0,0.29999998,0.43333334,0.5,0.53333336,0.65555555,0.8666667,2.2333333,1.4222223,0.44166666,0.08888889,0.0,0.06666667,0.71666664,1.2375001,2.1486113,2.5194445,2.427778,3.1,3.123611,1.6833334,0.73333335,1.0444446,2.6083333,2.1111114,1.0833334,0.0,0.025,0.011111111,0.23333332,0.62222224,0.5666667,0.23333335,0.21111111,0.06666667,0.0,0.0,0.0,0.0,0.0,0.18888889,0.5083333,0.6333334,1.6083333,1.3444445,1.0916667,0.22222222,0.0,0.0,0.0,0.06666667,0.6333334,2.425,3.5444443,1.5444444,0.85,1.8555555,4.5666666,6.244445,4.6500006,6.0444446,8.555555,11.808334,8.155557,3.3416667,0.56666666,0.25000003,0.16666667,0.108333334,0.2,0.0,0.016666668,0.34444445,0.24166669,0.5444445,0.4166667,0.10000001,0.35555556,0.8166667,1.0222223,0.058333337,0.055555556,0.14166668,0.011111111,0.0,0.0,0.011111111,0.2916667,0.5666667,0.475,2.5222225,8.575,9.877778,7.4555564,3.566667,1.1111113,0.93333334,0.0,0.0,0.044444446,0.7916667,0.75555557,0.33333334,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,2.8166668,4.5111113,1.2250001,0.0,0.0,0.15555555,1.0444444,1.2833334,2.988889,0.36666667,0.0,0.0,1.2,0.8333334,0.8333333,0.23333332,0.0,0.5333333,4.958334,0.47777778,0.0,1.2333335,0.7777778,0.0,0.0,0.05,1.9666667,0.0,0.0,0.083333336,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.075,2.2916667,4.3875,6.3,13.075001,16.416666,5.6083336,6.60625,8.416666,12.25,12.341667,10.4875,7.350001,2.76875,2.4666665,4.2333326,11.449999,11.758334,16.162498,16.858334,24.55,21.95,20.525002,7.7,3.466667,0.06875,0.116666675,0.61875,0.90833336,0.58125,0.083333336,0.23333333,1.03125,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10000001,0.8333334,0.825,0.26666668,0.225,1.8499999,0.76250005,0.81666666,1.4562502,0.20833334,0.008333334,0.0,0.0,0.006666667,0.016666668,0.725,0.083333336,0.05,0.3375,0.9166666,2.3125,2.65,2.34375,4.0916667,6.0250006,6.4249997,5.708333,3.9624999,2.6166668,1.4375,1.0833334,0.9,2.325,7.084091,9.7195835,12.058333,10.450001,9.438636,7.2625003,3.5583334,1.725,1.74375,1.1250001,1.7687501,1.6166668,0.26875,0.0,0.0,0.20000002,0.15833335,0.0125,0.008333334,0.0,0.0,0.0,0.0,0.0,0.00625,0.18333334,0.71875006,1.1750001,2.18125,2.3083334,2.9875,1.9583334,0.625,0.125,0.0,0.0,0.0,0.35625,1.4333334,2.175,1.26875,0.33333334,0.8000001,1.8999999,2.5000002,3.5666666,5.291667,8.64375,9.9,6.5312505,3.4916668,1.0999999,0.6333333,0.35625002,0.06666667,0.17500001,0.18125,0.033333335,0.00625,0.14166667,0.19375002,0.033333335,0.09166667,0.06875,0.20833334,0.13750002,0.06666667,0.05,0.12500001,0.1125,0.0,0.0,0.112500004,0.275,0.7687501,0.80833334,3.4312499,10.066667,12.741667,9.6,2.5083334,1.5312499,0.85,0.0,0.0,0.20000003,1.125,1.1750001,0.54375,0.0,0.0,0.0,0.0,0.0,0.0,2.13125,6.283334,1.8437501,0.0,0.0,0.116666675,0.39999998,1.13125,0.23333335,0.0,0.0,0.3125,0.3,0.25,0.1,0.0,0.0,0.083333336,0.94375,0.3416667,0.15625001,0.5916667,0.79166675,0.20625001,0.13333333,0.06875,0.4416667,0.0,0.0,0.0125,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17777778,0.22500002,0.3888889,0.7666667,1.9666668,3.0666668,2.8111112,3.8333335,4.9916663,6.6666665,9.216667,10.422222,7.7500005,3.2555556,2.4833336,2.9,4.133333,5.2999997,6.166667,10.541666,14.577779,17.658335,13.5222225,7.888889,5.766667,0.8444445,0.14166667,0.8,3.266667,1.388889,0.92499995,0.43333334,0.56666666,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.74444455,4.3,5.311111,3.9333334,1.9583335,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.23472221,0.48553032,2.6555557,5.533334,0.35555553,0.13333334,0.22500001,0.93333334,3.0249999,6.988889,8.5,7.338889,9.208334,13.844444,13.455555,11.591667,8.177778,5.533334,3.9777777,3.25,4.3444443,5.422222,9.458334,12.411111,11.400001,13.211112,13.6,10.044445,9.0847225,4.2499995,2.663889,0.975,1.8777779,0.73333335,0.011111111,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108333334,0.8555556,2.4416666,4.211111,5.158334,3.611111,0.96666664,0.9,0.18888889,0.25,0.0,0.0,0.11111112,0.54444444,1.3333334,1.1666666,0.06666667,0.4888889,0.59999996,0.97777784,3.3777776,5.5621214,6.8888893,5.366667,2.4111114,2.5666666,2.3111112,1.2083333,0.011111111,0.033333335,0.42499998,0.36666667,0.041666668,0.022222223,0.058333337,0.0,0.0,0.0,0.033333335,0.19166669,0.18888889,0.17500001,0.13333334,0.083333336,0.16666667,0.06666667,0.85,0.84444445,0.30833334,1.1000001,1.0916667,4.077778,14.033333,16.691668,9.222222,2.325,1.9777778,0.51666665,0.0,0.0,0.36666667,1.9222223,1.0999999,0.26666668,0.0,0.0,0.0,0.0,0.0,1.6833333,3.4777775,2.2333336,0.0,0.0,0.11111112,0.07777778,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0,0.0,0.075,1.4,1.9333333,1.4,1.4833333,1.7333335,2.022222,1.2416666,0.43333337,2.766667,2.9222224,0.875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,0.20833334,0.11111111,0.20000002,0.82222223,0.6416667,0.2,1.8444444,2.9250002,5.055556,5.558334,3.8222222,2.7583337,4.5,2.6166663,1.4,3.8888888,6.8999996,10.500001,12.041667,13.133333,17.150002,16.88889,6.0666666,0.8,0.1,0.4,1.988889,1.2833332,0.5,0.725,1.2222222,0.9111112,0.0,0.0,0.083333336,0.0,0.008333334,0.0,0.0,0.041666668,0.12222223,6.641667,14.4777775,12.766667,4.088889,0.62222224,0.0,0.0,0.0,0.0,0.05,0.06666667,1.3416667,2.2125,1.6222222,1.6371213,2.5,2.075,2.2555556,1.6833334,1.0222222,0.7111111,0.9166667,2.288889,4.0,8.044445,10.441667,14.1,12.75,12.333333,15.3,15.083333,11.500002,7.858333,4.211111,2.8833332,2.1111112,2.3305554,4.025,5.2111115,3.3999999,2.7222223,8.6,10.377778,8.299999,13.041668,7.8111115,5.8166666,2.6888888,1.2583333,0.6666666,0.041666668,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,1.4916667,4.7222223,6.8,5.711111,2.6333334,1.0166668,1.0333334,0.94166666,0.3111111,0.0,0.0,0.08888889,0.65,1.3666668,0.7416667,0.044444446,0.13333334,0.07777778,1.2888889,9.753031,13.766666,9.708334,4.3333335,2.0,2.7333333,2.5416667,1.0111111,0.11111112,0.30833334,1.2,0.325,0.0,0.06666667,0.0,0.0,0.0,0.0,0.033333335,0.22222224,0.23333333,0.2,0.19166666,0.1,0.37777779,0.9,1.1999998,1.2749999,1.4555557,2.4416666,3.1,9.666667,19.433334,17.911112,8.183333,2.688889,1.3833334,0.0,0.0,0.13333334,1.611111,1.7333333,0.17777778,0.0,0.62222224,0.19166668,0.0,0.06666667,5.4750004,6.488889,1.2,0.06666667,0.17500001,0.6111111,0.044444446,0.0,0.0,0.05,0.33333334,0.22500001,0.0,0.06666667,0.06666667,0.6,2.3416667,6.1000004,6.6,8.455556,9.791668,6.1777782,4.711111,4.2749996,3.0333333,17.916668,16.022224,3.225,0.2777778,0.36666667,0.32222223,0.3,0.7166667,2.211111,1.825,1.9222221,2.25,0.9111111,0.044444446,0.075,0.13333334,0.09166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.11666667,0.28750002,0.22500002,0.075,0.14166668,0.112500004,0.26666668,1.1750001,2.3874998,2.8166668,1.125,2.1333332,3.03125,3.3666668,2.71875,2.1166668,3.3416667,9.575001,14.666666,23.818748,27.158335,21.893751,9.233334,0.49166667,0.53749996,0.48333335,0.4,1.1249999,2.1687498,1.575,1.3874999,1.8166666,1.7833335,0.8874999,0.14999999,0.24375,0.20000002,1.6125,3.8500001,5.2000003,8.075,15.025,19.7625,15.625001,5.0625,0.98333335,0.725,0.725,0.050000004,0.03125,0.85,1.51875,2.1083333,1.5562501,2.8416667,4.3916664,7.30625,8.766667,9.40625,9.166666,8.606251,7.391667,4.9083333,2.8041668,1.7666667,3.30625,5.5583334,7.3937507,9.816668,11.506249,10.891666,11.875,16.3625,14.408335,11.431251,5.3416667,2.5562499,3.0083332,3.075,2.56875,2.6083333,1.15,0.30833334,1.6125,3.5749998,4.183333,5.55625,6.508333,5.5141025,5.425,1.9375001,0.45833337,0.4875,0.4083334,0.058333337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,0.97499996,5.2750006,9.343751,8.408334,6.416667,4.39375,2.4916668,2.2125,0.7083334,0.0,0.0,0.0,0.1375,0.3416667,0.41874996,0.25,0.10000001,0.23333333,0.9522728,7.166894,19.625,18.562498,10.566667,3.1875,2.7166667,3.54375,3.1083336,0.43333334,0.86875,1.1166666,1.7874999,0.45833334,0.087500006,0.0,0.0,0.0,0.0,0.0,0.0,0.18125,0.44166666,0.25625002,0.20833334,0.38333336,0.7875,0.5833334,1.1375,0.92499995,1.0687499,3.9666662,7.483334,15.775,25.050003,14.681251,4.9250007,3.5562503,0.6166667,1.175,3.5916667,8.208333,6.5375,2.175,1.05625,1.2583334,1.00625,0.73333335,1.7083333,5.74375,5.0083337,0.5375,0.7666667,1.2437501,0.98333347,0.7166667,0.81249994,0.0,0.1375,0.64166665,0.2875,0.108333334,0.25,1.4666667,19.025,21.287498,20.25,20.3375,30.883335,38.16875,18.075,12.716667,11.30625,5.4,3.71875,2.75,3.9250002,5.3583336,6.54375,7.7833333,8.608335,10.53125,11.25,13.45,15.475,14.19375,7.425,3.7416663,1.38125,0.40833333,0.21875,0.008333334,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.10833334,0.26666665,0.25,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.06666667,0.15,0.10000001,0.3,0.3666667,0.4416667,2.3333337,1.8111111,1.0416667,0.5888889,0.35,1.4777777,1.9666665,1.3444445,1.9750003,3.8222222,5.555556,11.733334,21.444447,24.458334,25.522223,11.75,4.188889,2.2444446,1.4833335,0.67777777,0.26666668,1.1888889,1.0416667,2.0777779,1.0583334,1.9666666,2.5444446,1.4499999,0.70000005,1.0416666,1.2222223,5.9,11.811111,14.0222225,16.066668,12.0222225,5.95,0.7444445,0.73333335,1.1333333,0.90000004,0.0,0.0,0.083333336,0.9111111,2.9250002,2.4555557,1.4916668,2.2111113,4.3444443,9.641666,14.911112,20.358334,27.144445,30.158333,25.533333,20.444445,13.366666,4.9,2.4333336,3.288889,6.2166667,9.088889,7.9500003,5.377778,6.588889,12.575001,16.9,11.658334,7.077778,5.8666673,6.2888885,7.966666,6.6601515,3.9708335,3.9916668,0.7777778,0.3,1.7111111,3.5666666,2.266667,0.43472221,0.9265151,1.9347222,1.2750001,1.6444445,0.0,0.08888889,0.044444446,0.033333335,0.0,0.0,0.0,0.016666668,0.0,0.0,0.016666668,0.033333335,0.10000001,0.07777778,1.1416667,4.377778,8.000001,7.955556,7.0333333,5.825,5.377778,2.55,1.7222223,0.33333334,0.055555556,0.011111111,0.36666667,1.011111,0.8416667,0.055555556,0.09166667,0.2,0.6333334,4.8833337,12.955555,21.658333,19.18889,6.816667,4.5,6.391667,5.5444446,1.8,1.3916668,2.6111112,2.9250002,4.1222224,0.725,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.49166667,0.5222222,0.75555557,2.6166668,1.7555556,1.3916668,1.4888889,0.88333344,2.5,6.288889,15.283335,23.022223,17.9,7.833333,7.0249996,3.7111113,3.725,3.2222223,10.08889,14.083334,8.922223,3.658333,3.9222224,5.016667,3.4222221,3.3000002,3.9750001,4.388889,2.2916665,3.211111,3.7416668,8.344444,7.1444445,4.858333,0.13333334,0.47499996,0.53333336,0.52500004,0.29999998,0.33333337,12.888889,63.155556,50.74167,31.566666,27.96667,42.11111,45.71667,24.28889,19.033333,15.208334,6.7999997,2.8416667,2.1777778,2.9499998,3.077778,2.9333334,3.9444447,7.166667,8.183333,5.244445,8.208334,15.333335,19.483334,26.4,31.022224,14.333333,4.555556,1.0500001,0.54444444,0.26666665,0.044444446,0.0,0.0,0.0,0.0,0.0,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,0.2777778,0.52500004,0.3111111,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18333334,2.1125,0.7083334,0.26875,0.21666668,0.38333336,0.59375,0.5666667,0.48125002,0.30833337,0.39999998,0.6833334,2.4125001,4.566667,7.291667,10.606251,15.491666,16.306252,12.666667,9.36875,4.708333,1.4999999,0.59374994,0.45833334,0.9749999,0.92499995,0.59375,1.7,3.3062503,2.8166664,2.4083333,1.68125,1.85,2.2375002,4.7916665,5.3937497,3.7333333,5.383333,3.8125,1.7666665,0.1375,0.15,0.0125,0.06666667,0.0,0.0,0.033333335,0.12500001,0.033333335,1.66875,7.0583334,10.924999,8.983333,7.633333,7.8095837,10.150001,12.7375,14.425756,13.512085,11.933333,12.916666,14.469167,11.325001,7.1749997,5.9416666,5.3500004,6.166667,9.550001,9.016666,6.241667,6.425,8.391666,8.900001,7.2250004,4.1000004,3.5966666,9.828031,16.413332,15.868938,7.8250003,4.7166667,1.5062501,0.8666667,0.85833335,3.3,4.635606,3.3218184,1.73,1.1255682,4.105303,1.11875,0.48333335,0.23333335,0.05,0.0,0.0,0.008333334,0.0375,0.0,0.0,0.0,0.025,0.21875,0.6083334,0.9437501,2.8000002,7.8562503,10.541667,7.4166665,4.25,4.05,4.14375,1.4666666,0.33125004,0.06666667,0.016666668,0.0125,0.68333334,1.71875,2.1499999,0.8625,0.29999998,0.275,0.8125,2.1750002,11.331249,20.849998,12.94375,9.133333,10.575001,8.558334,4.1083336,0.66875005,3.4166667,5.475,5.3000007,5.0312505,0.49166664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.575,1.0833335,5.35,7.808334,5.9187503,5.8500004,2.7749999,1.4166666,4.4416666,19.55,25.383335,19.518751,11.3,13.7625,12.966667,12.081251,3.6833334,8.066668,14.087502,7.016667,6.2875,11.266666,13.343751,15.058332,8.925,4.09375,5.908333,6.0,8.533333,8.8375,13.050001,9.049999,8.218751,0.86666673,1.23125,1.3166666,1.7625,1.7666668,7.8375,45.308334,62.16667,39.574997,28.616669,38.84375,51.825,36.675003,24.6,22.600002,21.10625,13.1,6.20625,3.0083332,1.98125,1.9583333,1.49375,2.35,10.216667,12.175001,7.233333,8.481251,15.275002,29.306252,41.800003,43.19167,34.28125,25.391665,19.706251,8.541666,2.9375,0.8083333,0.49166667,0.55,0.25000003,0.20000003,0.20000003,0.18750003,0.0,0.0,0.033333335,0.13333334,0.05,0.041666668,0.00625,0.0,0.0,0.016666668,0.1416667,0.46875003,0.60833335,0.56875,0.65,0.225,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.33333334,0.8500001,0.2,0.65833336,0.97777784,0.87777776,0.6416667,0.65555555,0.6166667,0.8666666,1.1750001,1.5222223,3.8666668,6.455556,11.388888,9.9,9.8,11.075,16.911114,20.991669,11.944445,3.7333333,1.5416666,1.0111111,0.65,0.31111112,1.15,6.4333334,4.9833336,3.1222224,3.3666666,3.0083334,2.822222,3.0583336,5.1555552,6.0833335,4.966667,4.8555555,2.2583332,0.31111112,0.0,0.0,0.0,0.0,0.0,0.0,0.67777777,0.9000001,0.022222223,1.1916667,2.2777777,6.308334,16.744444,14.48889,6.616667,7.0444446,4.416667,2.6666667,0.95,2.011111,5.7111115,10.258333,8.588889,6.8916674,2.4333334,1.0666666,1.4555556,1.0416666,3.4444447,7.7222223,7.608334,10.311111,11.474999,12.588889,12.725,6.6555557,0.5911111,8.001667,18.133333,12.358335,4.936111,3.2083335,1.2222222,0.82222223,0.34166667,3.3666663,5.125,6.866667,0.9333334,3.1222222,2.2666667,0.5,0.33333334,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.033333335,0.0,0.88888896,1.4416667,4.4111114,7.5333333,13.5,10.8111105,3.1583335,2.2,3.0333333,3.022222,0.97499996,0.033333335,0.0,0.116666675,1.1111112,2.6666665,3.6111112,2.575,1.2666667,0.2111111,0.60833335,0.5777778,1.6416667,8.944446,15.999998,17.811113,14.55,15.977778,11.333334,1.45,2.5,7.666667,8.677777,3.7999997,2.588889,0.18888889,0.0,0.0,0.0,0.0,0.0,0.0,0.31666666,0.57777774,1.0333333,6.3250003,13.700002,14.8166685,14.0,7.2666664,2.1888885,2.4444447,22.833332,30.233334,19.100002,14.888889,21.983334,28.0,21.216665,7.244445,8.5222225,12.65,3.6000004,10.675,24.188889,28.150002,35.655556,18.788889,7.55,9.8,13.283334,17.722223,17.241667,13.244445,10.288889,12.366667,1.8444445,2.0333335,2.7333336,4.691667,8.600001,28.691666,29.633333,21.744446,25.575,54.13333,71.86667,65.4,34.891666,18.922222,14.6,20.158333,23.08889,11.924999,6.6333337,6.2500005,7.144444,6.241667,7.666667,16.922222,40.95,31.611113,18.708332,25.344446,32.38333,38.833336,44.07778,52.583332,53.666668,48.15834,38.455563,23.625,11.9777775,6.355556,4.991667,2.1666665,1.1999999,0.26666668,0.15833335,0.06666667,0.10833334,0.15555556,0.15555558,0.25000003,0.12222223,0.06666667,0.0,0.0,0.0,0.022222223,0.2916667,0.8111111,1.5166668,0.8111111,0.008333334,0.32222223,0.13333334,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20000002,0.26875,0.0,0.10625,0.25,0.13333334,0.21875,0.47500002,0.70000005,0.57500005,2.01875,1.9666667,5.18125,7.9916673,11.500001,8.1125,4.225,6.95,12.075,16.03125,17.850002,17.133333,3.9687498,1.8583332,0.30625,0.75,1.64375,7.616667,5.2875004,3.8166668,4.366667,3.5687501,2.1,2.7375,4.6613636,2.435577,0.4965909,0.80833334,0.375,0.0,0.0,1.0083334,0.0,0.0,0.0,0.0,0.20000002,0.45,0.116666675,1.09375,5.5333333,8.543751,7.5666666,3.3666668,2.80625,2.1916668,2.5125,4.4666667,9.018751,15.008332,16.0,11.950002,9.408334,12.674999,20.883331,8.74375,3.916667,3.875,2.9666667,4.0333333,4.1499996,2.7583332,4.03125,5.1749997,4.075001,1.6416668,0.94166666,2.0986743,5.2749996,8.653265,6.1166673,2.9250002,2.6166668,2.0916667,1.84375,2.8166668,5.81875,2.5886362,1.3308333,0.0,0.18125,0.075,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.025000002,0.1125,0.20833334,2.2749999,4.525,9.843751,17.041666,15.075001,3.5375,0.55,1.5624999,2.3583333,1.4187499,0.47500002,0.058333334,0.25625002,0.30833334,4.74375,6.6416664,3.3249998,1.8416667,0.20833334,0.0375,0.058333334,0.53125,4.2916665,12.875,21.758333,20.856249,30.449999,23.349998,3.6812503,2.0500002,6.65,8.725,4.8,2.7250001,0.875,0.33124998,0.0,0.0,0.0,0.075,0.10000001,1.8937502,5.566666,3.3666663,5.7562504,15.016666,22.8375,21.35,14.175,5.766667,2.325,16.5375,32.108334,18.79375,17.766666,24.300001,37.25,24.44375,14.900001,17.05,13.34375,3.4666667,14.424999,41.141666,49.256252,51.23333,25.325,9.64375,14.033334,21.63125,29.000002,30.8125,21.475002,11.4,11.212502,2.8833334,2.45,3.375,11.4125,22.258331,17.012503,14.991667,21.125,29.243752,31.658333,34.63125,43.20834,31.20625,24.85,18.933332,12.68125,7.541667,6.5875,9.149999,14.150002,20.95,20.550001,30.525002,44.450005,72.19375,66.1,56.518753,50.641663,52.081253,57.008335,60.466667,64.06875,67.96666,70.168755,58.158337,51.6875,34.64167,23.25,12.74375,8.925,7.0875006,3.8083332,2.5687501,1.3416667,0.58750004,0.22500001,0.13333334,0.20000003,0.06666667,0.01875,0.0,0.0,0.0,0.008333334,0.14375001,0.69166666,1.2312502,1.2833334,0.0,0.0,0.0,0.025000002,0.15833333,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3,0.5333334,0.0,0.016666668,0.07777778,0.044444446,0.22500001,0.84444445,0.8416667,0.88888896,1.6333333,1.7777779,7.0333333,11.655555,13.877778,6.308334,1.5333335,3.6416667,7.922223,17.841667,18.333332,20.922224,6.575,1.2,0.525,4.266667,4.75,5.3222227,5.208333,2.5777776,3.6444447,5.141667,4.2000003,2.6500003,1.0708334,0.18333334,0.011111111,0.0,0.0,0.0,4.475,13.266665,2.641667,0.0,0.0,0.0,0.0,0.0,0.0,0.22500001,2.6555555,6.1833334,3.855556,3.3444445,8.825001,9.28889,11.000001,20.43333,26.141666,19.722223,13.799999,11.691667,9.2,21.75,34.144447,8.383333,6.077778,6.8416667,8.944445,8.977778,7.058334,4.8888893,3.7833335,2.1000001,1.0999999,1.3555555,2.722222,15.108335,16.911114,1.025,0.45555556,2.1750002,7.3555555,6.833333,7.4416666,6.5,5.2999997,2.7682538,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.20833334,0.14444445,0.25833336,0.73333335,0.9166667,2.9,5.7166667,13.355555,16.788887,6.225,0.35555556,0.28333333,0.9111111,0.97499996,0.8333334,0.25555557,0.24166669,0.24444446,4.4249997,6.0,3.3500001,1.5444444,0.22222222,0.041666668,0.0,0.14166667,1.5333333,10.433332,27.366669,26.291668,28.911112,27.966665,10.366669,2.0777779,4.516667,6.966666,6.4916663,4.5666666,4.466666,4.55,2.4777777,0.6666667,0.0,0.60833335,0.2777778,2.3666666,9.933332,6.722222,4.05,9.077778,16.724998,32.32222,18.849998,9.977778,5.3555555,7.266667,23.677776,17.75,15.033335,21.716667,34.333332,21.55,25.366669,26.3,14.241668,5.7222223,13.566668,51.32222,58.36667,52.255558,24.777779,8.766667,17.733332,28.891666,38.37778,40.750004,24.644444,13.055556,9.958334,3.5222225,2.7500002,6.0666666,16.116667,14.255555,14.475,14.677778,12.266666,12.800001,10.311111,17.208332,41.85556,45.291668,25.788887,12.888889,9.150001,16.222223,18.6,21.488892,20.841667,17.1,18.141666,21.855555,24.555555,44.79167,62.15556,79.433334,91.6,107.275,116.77778,122.8,113.100006,99.399994,101.75834,85.95555,74.75833,51.63333,38.111115,30.266666,20.2,17.483334,15.08889,11.083333,5.8222227,2.35,0.7777778,0.31111112,0.20000003,0.08888889,0.0,0.0,0.0,0.0,0.0,0.016666668,0.3,0.7416666,0.68888897,0.3,0.0,0.0,0.0,0.42222226,0.35000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33333337,0.05,0.0,0.044444446,0.35833335,0.7222222,1.3833333,0.82222235,1.0916667,2.9555557,9.741667,15.0,17.5,6.7833333,2.6111112,3.05,7.755556,17.516666,25.577778,20.28889,11.2,3.2333333,2.4916668,4.966666,3.9666667,5.4444447,6.0833335,4.7555556,3.9000003,2.2190475,1.6,0.28500003,0.08888889,0.008333334,0.022222223,0.0,0.32500002,1.1,1.2916666,2.4888887,0.33333334,0.0,1.2888889,0.8666667,0.0,0.0,0.0,0.19166668,2.0666666,1.1583333,0.6333334,1.7777778,8.541667,9.844443,4.7916665,12.5222225,11.183334,5.066667,1.8777779,8.808333,7.577778,14.325,7.611111,0.32500002,1.7666667,6.4500003,3.7666667,2.2555554,1.6742424,1.5333333,1.6333332,2.6888888,5.475,2.8222222,1.4555556,9.158334,11.78889,5.8666673,2.6777778,1.6916666,8.822223,12.4,10.15,10.733333,4.575,1.7444446,0.55833334,0.033333335,0.0,0.0,0.0,0.0,0.0,0.11666667,0.1,0.4098485,0.62222224,1.2333333,1.2,0.2777778,0.17500001,2.1625,5.1833334,2.588889,4.2333336,7.2222223,10.511111,5.2916665,0.8333334,0.3,0.56666666,0.3,0.3555556,0.3,0.2916667,0.18888889,2.791667,3.9222224,2.3166668,1.1666667,0.08888889,0.05,0.0,0.275,0.47777778,3.916667,11.555555,17.608334,17.144444,22.722221,11.450001,2.2555556,2.9750001,5.7,5.641667,4.8888893,7.222222,12.016666,12.855555,4.55,0.23333335,0.81666666,2.1555557,1.6166668,11.222221,9.811111,4.8583336,5.0111113,6.7000003,30.07778,22.883335,11.066668,8.6,3.9499998,17.177778,14.75,10.5222225,19.099998,28.522224,16.741667,29.144445,28.666668,15.116667,7.3444448,10.783334,52.688885,51.93334,42.46667,19.51111,7.791666,22.455559,36.15,45.33333,43.141666,28.599998,14.699999,10.408334,3.2222223,3.3083332,7.922222,12.816666,13.922222,14.041666,7.833334,6.7666664,7.541666,8.111112,19.058334,39.155556,33.9,23.233335,17.833332,18.583334,27.266665,35.658333,39.65556,24.325,20.755556,17.266666,16.766666,17.611113,28.908335,46.544445,48.958336,54.28889,75.70833,96.41112,110.18889,112.083336,102.01111,100.13334,94.45555,79.875,63.022224,53.9,49.483334,39.31111,25.883337,15.444445,14.783333,11.4,6.208333,2.3333335,0.88888896,0.4166667,0.34444445,0.13333334,0.11111112,0.016666668,0.0,0.0,0.008333334,0.16666667,0.6416667,1.4666667,0.975,0.0,0.0,0.37777776,1.0444444,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.2125,1.25,0.75,0.0,0.050000004,0.45000002,3.1166663,1.9687501,1.125,1.83125,5.416667,14.775002,20.841667,18.891666,7.7125006,3.6416667,7.6562505,14.033333,26.868753,36.31667,26.350002,13.0375,5.558334,4.3937497,3.8666666,5.99375,6.983334,5.09375,5.1833334,2.2183332,0.25,0.23333332,0.01875,0.0,0.00625,0.108333334,0.375,0.37500003,0.0,0.0,0.0,0.0,0.0,0.43333334,0.475,0.0,0.0,0.16666669,1.56875,0.40000004,6.225,8.133333,4.55,5.80625,3.233333,1.0812501,9.116667,6.7937503,1.6250002,0.025000002,2.50625,8.625,8.1,5.5833335,2.0,1.2166667,5.1000004,7.658333,14.375001,8.993751,4.25,1.48125,1.3166666,3.3812501,3.0583336,1.6083335,4.7374997,6.758334,4.80625,7.708333,13.197084,6.675,14.1,16.78125,8.433334,4.3937497,0.55833334,0.043750003,0.0,0.0125,0.025000002,0.875,1.09375,0.30833334,0.22625001,1.9833333,2.0500002,2.7483766,4.9227276,3.4610667,0.7083333,0.30625,1.8575758,9.28125,10.691666,10.337501,3.9916668,2.4916668,2.1374998,0.17500001,0.43125,0.9916667,0.118750006,0.075,0.28333336,0.38750005,0.20833336,1.6812501,1.8499999,1.0849999,0.47500002,0.050000004,0.0,0.0,0.44375002,0.125,0.24375,1.675,5.14375,7.183333,11.716666,11.25,5.1,2.875,3.0500002,4.24375,4.8250003,6.3333335,16.38125,27.258335,20.51875,3.2833335,1.73125,5.391667,2.75,4.7416673,8.075001,4.7125,6.833333,4.75,15.133334,28.075003,14.766667,9.075,2.875,10.983334,12.9125,7.2916665,15.231251,24.391666,13.862501,21.733334,27.700003,17.993752,7.916666,9.700001,48.4,41.1,30.916666,13.2,7.4187503,31.558332,46.106247,52.266666,45.218758,28.7,14.791667,9.60625,3.458333,3.5875003,8.016666,13.050001,14.050001,10.700001,6.283333,6.4583335,9.462501,8.941667,23.925,36.166668,31.1625,26.016665,23.283335,20.40625,26.925,28.781254,26.366665,31.599998,35.475,35.78125,27.675,22.258333,22.625,24.158333,24.7125,27.766666,42.212498,60.9,73.56667,89.20625,103.916664,113.3125,108.65833,93.525,80.325,77.025,73.11876,62.958332,43.481255,23.108332,14.525001,11.408334,6.46875,4.3750005,1.8916669,1.075,0.52500004,0.3125,0.7083333,0.85,0.7166667,0.21666668,0.0,0.041666668,0.18750001,0.075,0.0,0.0,0.043750003,0.16666669,0.8666667,0.83750004,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3,0.49166667,0.1,0.083333336,0.0,0.0,0.7083333,1.7555555,0.46666667,0.06666667,0.825,2.5333333,7.3416667,13.544445,9.311111,4.875,4.911111,13.341666,22.5,42.483334,46.666664,34.45555,17.866667,8.033333,7.3333335,8.122223,6.591666,5.8555555,2.496667,0.9263889,0.5444445,0.16363636,0.0,0.0,0.0,0.0,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.34444445,0.6166667,1.6111112,1.8333333,0.82222223,3.7749999,4.377778,0.14444445,0.425,3.688889,0.56666666,1.2555556,0.56666666,1.3333335,1.3222224,0.9333334,3.2888892,0.95833343,0.7555556,0.6583334,0.7111111,4.525,3.5,1.9888891,2.2083333,1.2555556,5.941667,0.7888889,2.4416666,6.1777782,8.333334,10.908335,12.98889,5.4083343,3.955556,9.841667,14.944443,5.9444447,7.8166666,3.2555556,1.9416666,0.3,0.016666668,0.13333334,0.0,0.34444445,4.1333337,6.9916673,1.8111113,0.65318185,3.1383333,8.464395,6.4624996,13.436111,12.641666,5.711111,1.5666666,1.9194446,9.85,16.833332,18.925001,9.777778,1.0666667,0.43333334,0.099999994,0.16666667,0.4666667,0.17500001,0.0,0.022222223,0.5500001,0.5555556,1.6666666,1.3555555,0.4666667,0.22222224,0.28888887,0.125,0.0,0.65,0.14444445,0.116666675,0.23333335,0.16666667,1.2444445,2.7555556,3.9083333,6.366667,3.516667,1.3666668,2.0916667,4.7222223,4.633333,11.799999,30.51111,35.191666,15.066667,2.5916667,7.4888887,6.4,2.9888887,3.9444442,4.008333,6.333334,5.591667,7.900001,26.675005,15.188889,7.3,2.7916667,7.744445,11.266666,5.9111114,11.225,17.177778,12.416667,15.044445,23.400002,18.158333,7.666667,9.316668,39.077774,30.966663,22.400002,9.3111105,11.341667,31.8,49.25,49.51111,43.800003,27.18889,13.555556,7.925,3.9222221,4.141667,10.511112,13.500001,15.266666,11.308334,7.5555553,7.4777775,10.083332,15.644445,27.05,37.622223,26.533335,26.933334,22.044445,15.158333,15.533335,13.833334,15.755556,10.691667,8.744445,8.833333,7.833334,6.3111115,6.4583335,6.477778,7.4666667,12.477778,14.608334,18.277779,28.566668,43.625004,61.566666,79.0,89.06667,95.06667,100.05556,102.0,96.683334,87.28889,68.899994,40.622223,22.816666,15.677779,9.591667,6.2333336,3.5666664,1.8083334,0.6666667,0.7,1.7,1.7666665,2.0333333,0.8111111,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.033333335,0.011111111,0.76666665,0.6333333,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.225,0.36874998,0.4,0.2625,0.05,0.075,0.63124996,0.225,0.90000004,0.9916666,0.1625,1.325,2.5375001,4.758334,7.925,4.10625,4.3583336,17.468748,35.200005,48.331253,56.875008,42.71667,20.706251,12.566668,9.768751,8.733334,4.358928,2.5,0.6,0.0,0.22500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.06666667,3.0187502,2.1083336,0.00625,0.083333336,0.1875,0.48333335,0.13333334,0.025,0.0,0.0,0.36666667,0.85625005,0.66666675,0.69166666,0.75625,2.5333333,1.76875,0.108333334,0.325,0.4166667,3.5312498,0.31666666,0.275,0.33125,4.1250005,23.51875,6.275,7.1375003,6.7749996,13.016667,17.31875,17.300001,8.356251,3.075,3.2937498,5.391667,7.2,6.125,2.5416665,2.3625,1.3583333,0.075,0.041666668,0.49374998,1.7749999,3.6962125,6.1125,5.108333,1.2687501,0.9568435,5.5206094,10.950758,7.6916666,12.891603,13.902122,7.2062497,3.7666667,4.5625,7.591666,12.05625,5.4249997,1.5916668,0.21875,0.5083333,0.55625004,0.16666667,0.25,0.09166667,0.074999996,0.61875004,1.2166667,1.5250001,1.8916669,0.77500004,0.38333336,1.3333333,0.90625,0.0,0.325,0.25833333,0.6125,1.1666667,1.0312501,0.23333333,0.17500001,1.25,3.516667,2.61875,2.125,1.5187502,3.65,4.3916664,6.0937505,21.608334,36.437496,26.575,6.4312496,7.0583344,8.693749,4.583334,4.116667,4.3,4.666667,5.2812505,5.8,21.4125,11.65,4.85,1.3499999,4.808334,7.612499,3.5833335,7.025,6.9000006,7.46875,14.525,18.766668,15.23125,4.783334,6.45625,28.666668,21.6,14.633332,7.1,11.85625,26.541668,40.875,38.674995,32.075,19.358334,11.133335,6.1562495,4.875,6.375,13.516666,14.968752,15.783333,12.087502,9.158332,13.183333,15.275,22.758335,35.63125,38.291668,27.824999,23.833332,18.091667,15.281251,14.633334,13.65625,17.916668,12.262501,7.866667,5.4125,7.3416667,5.6833334,6.575001,5.441667,7.2375,7.133333,7.1250005,7.608333,10.9,17.65625,30.316666,48.287502,59.158337,73.38125,101.90834,115.81667,110.99375,107.208336,95.69375,67.700005,50.13125,35.24167,21.30625,10.691667,5.891666,3.3812504,1.1916666,0.6249999,1.1,1.1812501,2.7833335,2.6166668,1.0125,0.016666668,0.0125,0.0,0.0,0.0,0.0,0.0,0.033333335,0.1,0.78333336,0.80625004,0.083333336,0.025,0.0,0.0,0.175,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.24444444,0.108333334,0.22222222,0.6555556,0.8083334,1.3555555,1.3166668,1.4000001,0.5083333,0.53333336,1.4000001,4.3111115,7.755555,3.7083335,5.1333337,22.508333,46.522224,52.3,58.833332,43.56667,23.65,16.433334,9.983333,4.9333334,0.39333332,0.0,0.15833335,0.0,0.0,0.058333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.23333333,0.24444444,0.05,0.0,0.8666667,0.5666667,0.44444445,0.0,0.0,0.016666668,0.16666667,4.366667,15.058333,3.8444448,0.70000005,0.76666677,6.0666666,5.0222225,2.1583333,2.266667,1.0,1.7083334,1.8111112,11.883334,1.3666668,3.475,3.9222224,6.9666667,11.6916685,17.666666,8.108333,3.2333333,4.1,0.98888886,1.4222223,3.3166666,7.044445,6.512121,8.1,2.125,0.022222223,0.40000004,3.661111,5.3597226,2.6083333,0.33888888,0.25833333,0.26666665,0.33333337,4.749207,7.122024,2.4602523,16.872223,21.733334,8.0222225,4.016667,5.0666666,4.0583334,1.911111,2.977778,0.86666673,0.4,1.0583333,0.5555555,0.13333334,0.5222222,0.76666665,1.4583333,2.5777779,2.216667,4.111111,2.0666668,0.90000004,3.2611113,2.3810606,0.0,0.25833333,0.6,1.1250001,2.688889,2.1333334,0.0,0.0,0.39166665,2.411111,2.6749997,3.3666666,1.9499999,1.9666667,4.9111114,4.991667,11.766666,27.733332,30.288887,13.033332,4.8888893,7.733334,5.533334,5.0555553,4.9583335,4.188889,3.5583334,4.2444444,22.258331,8.944445,2.3333333,0.375,2.1888888,4.1333337,0.9444445,1.425,1.3222222,3.7250001,8.2,11.01111,7.016667,1.7333333,4.275,18.733334,13.241667,7.7888894,4.0111113,6.8750005,17.833332,24.775002,13.544445,11.916666,8.9777775,5.533333,3.8333337,5.9111114,9.466666,13.688889,16.358334,15.833333,12.916667,13.633333,19.844444,24.400002,29.933334,38.5,36.100002,33.275,25.222223,19.97778,17.224998,16.97778,15.691667,20.055557,15.325001,9.566667,5.916667,4.8,4.1444445,3.3916664,8.644445,16.383333,15.700001,13.258334,13.200002,11.477777,12.625,23.133335,37.64167,49.97778,57.033333,64.46667,82.2,97.200005,98.288895,97.12501,99.94444,89.96666,67.95556,42.525,19.56667,10.733333,5.1499996,2.711111,1.1833334,1.4444444,1.7416667,3.8111112,4.4555554,4.3500004,1.1111112,0.30833337,0.0,0.0,0.0,0.0,0.0,0.011111111,0.116666675,1.1888888,0.98333335,0.62222224,0.89166665,0.08888889,0.0,0.23333333,0.39999998,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.025,0.025,0.19166666,0.5875,1.1999999,1.1812501,1.4583334,0.35000002,0.20833334,1.15625,3.775,9.441667,4.825,6.2833333,33.96875,48.133335,55.025,56.58333,44.225,27.437443,19.850002,7.0795836,2.165,0.112500004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333334,0.40625,1.0416667,0.83750004,0.0,0.36666667,4.1875,2.3583336,0.0,0.0,0.043750003,0.18333334,0.6166667,3.56875,8.533334,4.7875,1.5833334,1.2,0.3416667,0.1,0.15,1.075,2.7687502,4.666667,6.4624996,9.308333,10.28125,10.15,11.275002,8.2625,11.625,12.887501,11.900001,9.2625,1.1666666,0.36666664,2.1937501,7.05,12.050001,9.950002,3.4016669,2.2500002,0.35000002,1.2750002,4.541667,0.8375001,0.075,0.0,0.043333337,0.06363636,2.563889,6.841667,6.546667,7.067425,22.862501,22.508333,7.6875,6.883333,5.76875,4.208333,4.658334,3.6312501,0.05,0.83125,1.3750001,0.475,0.26666668,1.2750001,2.7999997,3.5416665,3.04375,4.666667,3.4083333,2.1250002,4.4992433,3.7124999,0.32500002,0.78392863,1.375,2.0258334,4.4249997,3.3624997,0.0,0.0,0.55625,2.6249998,2.85,2.25,4.1125,2.275,4.916667,6.05,8.425,18.081251,27.44167,15.88125,4.9000006,6.1874995,5.775,4.4083333,2.9625,1.9166667,2.45625,3.2583334,8.912499,3.483333,0.85,0.050000004,0.8333333,1.425,0.10000001,0.043750003,0.0,2.35,4.0916667,5.0833335,1.45,0.16666669,2.18125,9.749999,6.35625,3.3083334,1.1083332,2.9125,13.583333,10.587501,2.2666667,2.7250001,2.841667,2.8250003,3.6687498,5.616667,6.0375,8.458334,10.506251,9.55,10.26875,15.483335,17.391666,29.28125,35.025,46.0625,39.300003,33.6875,26.233334,23.633333,21.537502,19.375,20.281252,21.408333,18.050001,10.208334,7.3125,6.025,5.0916667,11.200001,23.308334,24.925,26.975,19.206251,16.616667,16.866667,18.106247,20.841665,27.881248,47.766666,56.000004,52.79167,57.75833,68.30625,79.2,90.4625,95.91667,93.26875,77.59167,61.225006,44.208336,30.533333,12.724999,7.0583334,3.0187502,2.3333333,2.4375,4.5249996,8.083334,14.6875,18.866665,11.3,1.3000001,0.0625,0.0,0.0,0.0,0.0,0.23750001,0.98333335,1.4125,1.55,1.325,0.66666675,0.033333335,0.025,0.19999999,0.19999999,0.0,0.15,0.29999998,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15555556,0.42499998,0.055555556,0.12222223,0.31666666,0.18888889,2.5333333,1.5555557,0.21666668,0.14444445,0.5916667,4.533334,13.555555,6.7916665,8.8,25.516666,40.744446,50.875004,44.93333,34.3875,19.664091,9.293333,2.891667,0.7955556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,1.6000001,2.6333334,1.6916666,0.11111111,0.0,0.0,0.0,0.0,0.011111111,0.20833334,0.9666667,2.788889,6.4249997,8.98889,6.008333,1.1222223,0.025757577,0.0,0.0,0.21111113,1.4777778,4.6250005,3.3777778,3.7,5.566667,9.583332,10.966666,5.688889,4.6916666,8.055555,9.150001,7.488889,10.025001,4.7000003,2.977778,4.6916666,2.0111113,2.656667,8.9317465,3.2257578,0.5444445,1.375,0.0,0.022222223,0.058333334,0.0,0.0,0.0,0.0,2.8333333,5.145833,5.6333337,7.0111113,10.624999,15.711111,9.108334,6.0444446,4.4416666,2.3777778,4.588889,5.4083333,0.87777776,0.78333336,1.5222223,0.9416667,0.26666668,0.65555555,3.8583336,4.744445,3.7833335,5.288889,4.166667,1.8444446,4.288889,4.7333336,1.4777777,2.5083332,3.0333333,3.2333333,6.2000003,4.6833334,0.0,0.0,1.4916668,2.1666667,2.075,1.4333335,4.8999996,3.177778,4.7,7.0916667,6.811111,12.000001,20.944447,13.925,5.5,5.2833333,5.4,2.8666666,1.3666667,0.6666667,1.0916666,1.5444446,2.275,0.2777778,0.0,0.0,0.06666667,0.13333334,0.0,0.0,0.0,2.0583336,2.4666667,0.4333334,0.075,0.0,0.7833333,3.2666667,1.6333334,0.7444445,0.22222222,2.6333334,12.622221,6.0416675,0.4777778,1.3166666,2.2333336,2.188889,3.6666667,6.588889,10.691668,13.644444,13.916666,9.244445,12.299999,16.022223,13.777779,26.133337,29.077778,43.21667,35.188892,28.1,27.1,26.533335,28.31667,23.4,22.55,20.433334,14.933333,10.777779,9.2,9.48889,12.788888,16.166666,25.711111,23.416666,23.355558,18.608334,16.222223,18.455557,20.791664,21.711111,31.183332,51.633335,65.39167,53.266666,46.03334,49.125004,59.844448,63.283333,63.388885,72.125,78.58889,83.35834,80.8,73.04445,50.683334,27.0,11.366666,6.477778,3.0416667,1.6555555,2.3888888,5.5166664,9.922223,15.250001,6.533333,0.95,0.044444446,0.0,0.0,0.0,0.06666667,1.1777779,0.975,1.9000001,1.4000001,1.1777778,0.48888892,0.6166667,0.88888896,1.6333333,0.40000004,0.26666668,0.24444446,0.06666667,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,0.63750005,0.06666667,1.7375,2.1083333,0.6625,0.25,0.36875,2.9416668,9.566667,11.8125,11.716667,18.28125,30.075,44.956253,34.533333,24.125,8.253395,3.8388891,2.5346842,0.9566667,0.0,0.0,0.28750002,0.116666675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,1.3083334,1.3062501,2.6833334,0.6166667,0.025,0.0,0.7,0.9666667,0.47500002,9.283334,4.175,1.8625001,2.0583334,2.66875,0.81666666,2.34375,0.38333333,0.0,0.0,0.13333334,4.0375004,2.9416666,1.2499999,0.06666667,0.58750004,1.0333334,0.575,0.7437501,3.208333,2.2625,1.5999999,5.375,4.4999995,5.658334,3.9250002,2.234091,0.00625,2.8516672,1.8037878,1.604762,3.832124,3.1611114,0.36212122,0.34375003,0.0,0.0,0.008333334,0.01875,1.2,4.2,1.8875,5.108333,12.575002,7.562728,5.852083,3.9780307,5.16875,4.4333334,6.208333,6.7249994,4.7666664,5.6500006,3.9083333,0.99375,0.6583333,0.825,5.2625,6.2166667,4.6875,5.525,3.8875,1.0666666,4.175,4.40625,4.1666665,6.0375004,5.8500004,6.3,9.674999,2.2437499,0.0,0.0,1.4437499,1.0750002,0.8625001,0.97499996,4.9125004,4.3166666,3.2333333,5.3500004,4.35,5.6312494,9.783334,7.1625004,3.825,3.71875,3.8083334,1.3833333,0.6,0.3,0.13125001,0.35,0.4125,0.0,0.0,0.0,0.0,0.00625,0.0,0.0,0.0,1.08125,1.5500002,0.6666667,0.0125,0.0,0.13125,0.55833334,0.18125,0.033333335,0.1,2.5812502,5.8166666,2.05625,0.275,0.65625006,0.8916666,0.9250001,6.3625,13.708333,30.400003,30.891666,29.087498,12.225001,13.124999,13.516667,7.1583333,10.89375,14.124999,21.6625,19.350002,22.2125,27.783333,34.908337,33.39375,19.999998,17.312502,13.133334,9.2875,11.091666,15.88125,17.208332,18.208334,20.425001,22.166668,21.893751,20.85,21.29375,23.541668,26.233334,29.706251,32.36667,32.524998,33.791668,37.775,44.191666,47.225002,48.13751,46.95,46.324997,44.158337,54.331245,66.36667,82.40625,99.716675,111.3,104.387505,91.75,62.687492,37.583332,20.406252,14.766666,7.8500004,4.4125004,3.2250001,4.9312506,5.1833334,1.7250001,0.40833333,0.03125,0.0,0.0,0.0125,0.033333335,0.6125001,1.25,0.25,0.10000001,0.15,1.0000001,1.7833333,5.5250006,4.433333,0.95000005,0.2,0.90000004,1.1333334,0.73333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24999999,0.11111111,0.0,0.0,0.0,1.1666666,2.5333333,2.9499998,1.2444445,0.65833336,2.6333332,11.388888,17.475,15.777779,15.775001,21.0,33.9,28.533333,16.851986,4.516558,2.2,1.4825002,0.0,0.05,0.0,0.98333335,1.2666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,1.1666666,0.41666666,0.0,0.11111111,0.21666667,0.26666668,2.0,0.88888896,0.0,5.277778,2.411111,5.541666,3.8555555,0.0,0.98888886,12.758333,11.433333,5.383333,3.666667,0.0,0.23333335,0.3888889,0.0,0.0,0.0,0.0,0.0,0.84999996,0.22222222,0.14166667,0.0,0.6833334,1.4777777,3.1986113,3.060606,0.099999994,0.008333334,0.28373018,1.4492425,12.5847225,18.283333,9.133333,3.8333333,1.1,0.033333335,0.0,0.22222222,0.625,1.0968254,2.7194443,3.1750002,4.866667,10.474999,4.9222226,6.7166667,4.9222226,7.5333343,6.4777775,6.3444448,7.433333,8.333333,9.808333,6.8222218,0.84166676,0.71111107,1.9666666,6.2416677,6.477778,4.041667,5.077778,2.7,0.56666666,3.6555555,3.641667,6.0222225,8.941668,7.8777776,10.983333,10.41111,0.31666666,0.0,0.0,0.6666667,0.15555556,0.16666667,0.5,2.5833335,1.4333334,0.5,1.0416666,0.6555556,0.5833334,0.5444445,0.71666664,0.9111111,1.3166667,1.1333332,0.33333337,0.15833335,0.06666667,0.0,0.022222223,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.9666667,2.3666668,1.3333334,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.9333334,0.0,0.05,0.055555556,0.20000002,0.36666667,0.4888889,9.708334,19.077778,42.816666,40.01111,35.875,12.777779,16.708332,16.766666,9.7,9.333334,12.366667,23.575,28.022223,26.125002,28.711113,38.088886,29.741667,14.6,9.383333,7.8222218,13.091666,15.533334,14.933333,19.433332,20.722221,19.68333,17.522223,13.666668,12.6888895,13.891668,17.022223,20.355556,29.125,34.944443,37.250004,38.43334,39.675,44.02222,46.244446,49.908333,49.477783,44.625,40.344448,44.708336,53.67778,66.35,81.17778,94.45556,108.075005,111.05556,112.85,110.87778,90.091675,70.01111,57.744446,34.216667,14.566667,8.608334,9.744445,8.633333,8.733334,2.8000002,0.07777777,0.0,0.0,0.0,0.0,0.011111111,0.0,0.0,0.044444446,0.38333333,2.2444444,2.7333333,1.6666667,0.8166666,0.79999995,0.8166667,1.2,0.8,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.11111111,0.0,0.0,0.37777776,1.625,2.9,0.78333336,0.9888889,0.7583333,0.97777784,10.944445,19.833334,19.788889,16.166668,15.155556,25.033337,21.17778,8.0125,5.593701,0.0,0.3118687,0.011111111,0.20833334,0.0,1.45,0.37777779,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17777778,0.0,0.0,1.2,1.375,0.0,0.06666667,0.08888889,0.39166668,1.4666667,1.9333335,6.5166674,1.311111,0.5666667,0.5777778,7.0083337,24.566666,15.933333,1.2888889,0.0,0.19166668,1.8111112,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.6888888,2.975,0.6555555,0.5333334,0.3888889,1.825,7.6555557,15.4,3.1333334,1.4222223,1.1861111,0.51111114,0.025,1.4527777,1.4401515,0.75555557,2.5194445,4.258333,2.2777777,3.2750003,3.1666667,4.2916665,4.8444443,10.425,7.422222,5.9111114,7.675,9.111112,11.875002,8.044444,0.75,0.92222226,2.711111,4.0333333,4.588889,1.5250001,2.5333333,0.9916667,1.2666667,4.133333,4.7833333,6.044444,8.825001,8.411112,13.725,10.611111,0.9333334,0.0,0.0,0.43333334,0.022222223,0.1,0.3,0.4416667,0.24444443,0.011111111,0.14166668,0.14444445,0.058333337,0.0,0.40000004,0.84444445,1.0500001,0.11111111,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.79999995,1.5333333,0.3666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.1,7.533334,15.355557,33.758335,28.822224,23.0,10.911112,24.766666,26.211113,18.644445,19.991667,22.222223,25.258333,38.15556,33.783333,23.388887,28.066666,23.216667,14.622222,9.633334,13.633333,13.375,14.233332,15.733333,13.177778,10.233334,10.791666,10.755557,12.0,14.922221,15.975,17.611113,18.811111,21.1,27.533337,34.441666,39.02222,43.54167,48.933334,54.433334,56.458336,52.344444,50.191666,44.144444,44.116665,47.62222,54.691666,67.03334,87.27779,96.658325,96.76667,102.075005,119.6,135.39166,135.24445,112.41112,88.54167,42.5,20.191666,16.466667,26.241667,20.58889,15.499999,1.7666667,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.53333336,0.35,0.51111114,2.4333334,0.08888889,0.51666665,0.44444442,1.0333333,1.0222223,0.40000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5083332,2.6875002,3.2083335,0.98125005,0.6,0.48125,1.3083334,9.266666,19.0875,20.383335,15.1625,11.225,12.393749,8.115909,3.5383842,0.96250004,0.22500002,0.16875002,0.16666669,0.00625,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.5916667,0.55625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14166668,0.4875,0.0,0.0,0.0,0.14375,1.1416667,0.5,0.0375,1.225,1.23125,0.05,1.7750001,4.808334,1.9375,0.13333334,0.0,0.0,0.38333336,0.28125,0.0,0.0,0.0,0.0,0.0125,0.32500002,0.00625,0.0,0.9717857,1.1924242,1.7916666,2.41,1.375,1.9624999,0.1,0.325,2.141667,13.362499,4.741667,0.5583334,2.825,2.3333333,0.45458335,1.9792424,0.7329167,0.32916668,3.9237375,4.8,0.25833336,1.15,1.4863636,5.14375,7.5916667,12.456249,9.233334,4.7166667,9.331249,9.675,11.54375,7.2166667,1.0250001,2.1,3.25,1.3625,1.4583335,0.9250001,0.9416668,0.6,1.9916667,4.525,5.30625,3.1000004,7.9437504,9.858334,9.918751,5.575,0.43750003,0.0,0.0,0.25625002,0.116666675,0.15,0.12500001,0.12500001,0.041666668,0.050000004,0.12500001,0.116666675,0.0125,0.0,0.14375001,0.5,0.82500005,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.3,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,2.54375,4.608333,11.8875,10.675,11.00625,7.7749996,28.85625,34.183334,26.666664,29.6625,22.558334,20.262499,27.883335,29.26875,16.708334,15.175,14.825001,16.216667,14.281251,12.566667,17.54375,17.125002,11.468749,8.083334,9.258333,10.818748,13.308333,14.24375,15.933335,18.331251,19.758333,22.283335,25.425001,28.741667,31.156248,34.63333,38.08125,40.816666,44.991665,50.775005,52.924995,56.375,57.73333,53.05,52.15,54.475002,58.224995,58.35,62.28125,69.78333,79.825,98.01667,123.137505,137.99167,146.05833,139.1875,103.61667,62.90625,34.816666,27.96875,31.916668,29.30625,13.483333,2.5083332,0.36875004,0.016666668,0.01875,0.016666668,0.0,0.11666667,1.3166667,5.2375,1.575,0.0,0.24999999,0.15,0.6,0.425,0.4166667,0.28333336,0.025,0.35000002,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1333333,4.0750003,4.1444445,1.6833334,2.0333333,3.425,4.3,8.800001,13.85,15.1,10.891666,6.744445,3.391667,0.0,0.6333334,2.3416667,0.7650794,0.20833333,0.36666667,0.325,0.0,0.033333335,0.0,1.0555556,0.48333335,0.0,0.0,0.7,1.5000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,2.488889,0.3,0.0,0.0,0.0,0.05555556,0.32500002,0.044444446,0.99166673,1.3555555,2.9083335,2.488889,0.0,0.0,0.0,1.0333333,0.0,0.0,0.033333335,0.16666667,0.5166667,0.54444444,0.09166667,0.0,3.591667,6.0111113,4.333334,4.3083334,0.35555556,0.15,0.011111111,0.5083333,2.1222222,10.875001,5.888889,0.32222223,9.533335,6.7222223,0.14833334,1.5916667,0.85277784,0.62222224,7.643056,5.9416666,0.0,0.58555555,1.6888889,8.133333,7.055556,12.725001,9.833333,4.666667,11.783333,9.788889,11.624998,6.8,1.6500001,3.7333333,4.6333337,1.2333332,1.5111113,1.7,1.7333333,1.2,1.5888889,3.3222222,3.7749999,1.9222223,6.2500005,6.4555554,2.2999997,0.35555556,0.0,0.0,0.0,0.075,0.8888889,0.7333334,0.0,0.016666668,0.011111111,0.15555556,0.20000002,0.11111111,0.0,0.0,0.0,0.9444444,0.5416667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.0,0.9166667,2.622222,5.816667,9.933333,26.408335,30.21111,22.6,19.783337,10.422222,12.783333,16.966667,12.733332,12.466667,10.944444,17.066666,15.722221,10.825001,11.222222,11.941668,7.133333,1.9916664,3.8777776,5.9666667,5.991667,7.822222,9.508333,9.744446,10.200002,10.966666,12.866667,15.491667,17.98889,20.091665,22.877779,26.658335,32.32222,40.01111,48.225,36.288895,35.433334,49.411114,66.025,77.100006,79.40001,73.65555,65.05556,57.09167,61.022217,70.48333,85.04446,99.375,110.755554,129.70001,160.33333,167.62222,137.55835,98.45556,55.300003,43.11111,45.875,37.922226,16.166668,2.875,0.11111112,0.033333335,0.0,0.0,0.0,0.0888889,0.45,0.33333337,0.041666668,0.5333333,0.14999999,0.0,1.7666668,6.4222226,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.60625005,1.0500001,1.7916667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.37500003,1.1083333,2.01875,0.84166664,0.80625,0.4666667,3.4833336,6.5125003,9.233334,5.150833,2.0916667,0.34374997,0.058333337,1.6316669,2.3491669,2.6575756,1.4937501,1.875,1.1437501,0.23333335,0.0,0.0,1.0916666,1.06875,0.0,0.0,0.05,0.0375,0.0,0.0,0.0,4.8833337,0.45,0.0,3.5812502,2.4166667,0.0,2.23125,1.4916667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.7333333,0.61249995,0.0,0.0,0.0,0.0,3.08125,0.0,0.33124998,0.82500005,7.075,10.058334,1.0,0.0,0.0,0.51686186,0.0,0.0,0.025,2.1750002,0.9625,0.4333334,0.22500001,0.10000001,2.4375,3.0500002,1.9250002,0.2,0.0,0.0,0.0,0.13125001,1.5083333,2.3937497,2.875,4.9416666,8.906251,2.7291665,3.2487411,7.252273,5.2510757,3.0000002,6.3803034,2.605682,0.0,0.19375,1.7204546,4.9437504,5.4333334,12.05625,8.383333,6.1333337,12.862499,6.8833337,6.3625,3.1833334,2.4624999,5.116667,5.5500007,1.45,2.0166667,2.7749999,2.0833333,1.3312501,0.6,1.5,1.4875001,0.83333325,1.5687501,1.5083332,0.275,0.0,0.0,0.0,0.0,0.3125,2.6916666,1.2062501,0.0,0.0,0.041666668,0.20000003,0.2,0.041666668,0.0,0.0,0.00625,0.9,0.1125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5000001,3.8166666,7.018751,15.941668,24.868748,18.358334,15.400001,6.58125,6.9916673,8.231249,11.766667,12.931252,17.291668,24.883333,20.04375,11.775002,8.18125,6.8166666,3.2375002,0.5583334,0.925,1.3166668,1.7583336,2.5375,4.125,5.6250005,6.6,8.125001,9.141666,10.366667,11.831248,14.116667,17.768751,22.05,25.062502,28.375002,32.025,34.281254,29.41667,23.512499,29.675,41.73125,52.816666,63.993748,74.71667,75.51667,67.69374,63.699997,67.3625,72.13332,81.84375,89.899994,109.808334,146.38126,172.325,184.54376,177.11665,118.23126,75.433334,73.24376,76.50833,48.225,20.912502,2.6333332,0.2125,0.0,0.0,0.0,0.0,0.46875003,1.1916668,0.46875,0.275,0.6375,0.4416667,0.35000002,1.5666667,0.0,0.21875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.32222223,1.825,1.7555556,0.8083334,0.24444443,0.82222223,1.6416667,2.1761906,1.1733334,0.47777778,0.4416667,0.8777778,1.5444446,1.1280303,3.5499997,4.2250004,3.9222221,3.8166666,0.92222226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5777778,0.0,0.0,4.308334,1.1555556,0.0,3.241667,0.18888889,0.3666667,2.0444446,0.0,1.5111113,4.4666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.0,0.0,0.6666667,2.2250001,3.611111,0.8666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.6444445,0.42499998,0.18888889,0.0,0.21111113,1.7222223,0.13333334,0.0,0.0,0.0,0.050000004,1.1999999,0.033333335,0.26666668,1.6,8.283334,7.666667,4.706061,8.911111,15.708335,6.422222,2.847619,0.083333336,0.0,0.058333334,0.5444445,1.3901515,5.0111113,9.391666,6.9555554,6.666667,14.558332,7.1000004,4.4666667,0.34444445,1.9083335,4.8555555,5.866667,1.3166666,2.2444444,2.8666668,2.0333335,1.1583333,0.25555557,0.43333334,0.11666667,0.08888889,0.058333337,0.011111111,0.0,0.0,0.0,0.0,0.0,0.6166667,2.3666668,0.275,0.0,0.0,0.033333335,0.13333334,0.13333336,0.022222223,0.0,0.0,0.025,0.64444447,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35555556,1.9166666,3.9222226,8.116667,19.433336,16.383333,11.088889,6.7000003,3.0083332,4.177778,9.808333,16.011112,23.075,34.244446,26.266666,13.158334,7.2000003,4.633333,1.7444445,0.98333335,0.9444445,0.9499999,1.0111111,1.1444445,1.5666667,1.8555555,1.6333332,1.5666667,2.5166667,3.977778,5.7666664,8.341667,10.755556,13.974999,17.944445,20.925003,22.155556,23.277777,22.675,21.055557,18.666666,17.6,19.475,25.377777,35.091667,41.922222,47.733334,53.033333,55.033337,57.333332,60.48889,67.025,73.666664,83.0,104.675,126.36667,156.26666,169.04446,150.80002,116.53333,88.316666,65.655556,51.466667,28.033335,6.2777777,1.1416667,0.08888889,0.0,0.0,0.0,0.17500001,0.06666667,0.07500001,0.16666667,0.35833335,0.16666669,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24444446,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.112500004,0.4,1.8625,2.625,1.925,1.0083334,0.3666667,0.8375,1.0333334,0.24375,0.44999996,0.90625006,0.6166667,1.6500001,1.5,1.1583334,1.60625,1.3499999,1.56875,2.1833334,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35833335,0.081250004,0.0,0.0,0.0,0.17500001,3.45,1.3499999,1.8562499,0.6,0.0,1.7333333,0.9125,5.3000007,6.2625003,0.48333332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17500001,0.1375,0.46666667,0.95000005,0.39999998,2.4312503,0.75,4.6875,3.275,0.0,0.0,0.65000004,0.725,0.65833336,1.3062501,3.8083332,0.75000006,0.0,0.20000002,0.4875,0.78333336,0.3125,0.16666667,0.32500002,0.0,0.033333335,0.9375,7.633333,2.1437497,6.675,1.8375,0.0,0.7719697,5.1687503,6.1833334,5.3949995,5.775,8.501667,4.183334,0.80833334,0.0,0.008333334,0.18124999,0.025000002,0.6,2.8833332,8.1875,6.65,10.75,19.7,9.566667,5.037501,0.058333337,1.8687501,4.1916666,4.9833336,2.0625,2.4333336,1.9187499,1.4250002,1.4375,0.45833337,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.23333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.15000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.575,2.0749998,2.8666668,8.925,12.458333,6.99375,3.6416667,0.6916667,1.2874999,10.408333,21.225,18.908333,25.699997,26.458334,16.616667,8.20625,4.6250005,2.3812504,1.3,0.6437499,0.39166665,0.45624992,0.49166667,0.30833337,0.10000001,0.16666667,0.35625005,0.52500004,0.40624994,0.6833333,1.2749999,2.425,3.075,5.6187496,8.466667,12.368751,15.916668,17.491667,17.46875,14.941667,13.44375,12.858334,12.981251,13.525,16.300001,18.541668,21.95,27.025,29.925001,35.83125,47.05,56.506252,62.833336,67.375,72.13125,86.76667,116.17501,114.03334,111.98126,103.13333,95.493744,71.433334,49.325,34.7125,15.441668,5.40625,0.8166666,0.043750003,0.0,0.0,0.0,0.0,0.0125,0.008333334,0.0625,0.8333333,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.0,0.10000001,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.8777778,0.92499995,0.74444443,2.3333335,0.9444445,0.33333337,0.5166667,0.7333334,0.25833333,0.2,0.82500005,0.70000005,1.0333333,0.9916667,0.07777778,0.15833333,0.7222222,1.0083334,0.21111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.3666668,1.4083334,0.0,0.0,0.0,0.0,3.6333334,0.2,0.32500002,2.4444444,0.0,0.0,0.0,0.27777776,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22222222,5.5111113,2.3083334,1.2444445,4.775,8.433334,6.633333,1.2333333,4.2583337,0.7444445,0.23333333,0.09166667,0.0,0.13333334,0.2888889,1.2666667,6.566667,2.0666668,0.0,0.17777778,1.5166667,2.7,1.5833333,0.67777777,0.0,0.0,0.37777779,15.9,44.22222,11.708332,16.31111,1.3166667,0.0,3.022222,5.516667,2.4333336,0.95000005,3.5555556,3.1583335,3.3666668,0.044444446,0.0,0.05555556,0.59999996,0.06666667,0.20000002,2.1666665,8.716667,8.044444,10.733334,14.583335,8.566667,4.008333,0.0,0.40833333,1.4888889,2.1999998,2.275,2.6555552,2.1666665,2.0111113,1.8166668,0.75555557,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.5888889,1.1833334,1.6666667,5.4583335,4.688889,2.8083334,0.07777778,0.18888889,1.0166667,5.811112,8.408334,10.244444,11.591668,10.655556,7.666666,4.45,2.6666665,1.1916667,0.51111114,0.108333334,0.033333335,0.05,0.022222223,0.13333334,0.42500004,0.9555556,1.8166668,2.0222223,1.7250001,1.3888888,1.1777778,1.45,2.5666666,5.2749996,8.933333,12.0,14.544444,16.211111,15.516667,14.233334,11.366667,9.844444,9.616668,10.133333,10.016665,9.922223,9.6888895,11.608334,13.177777,17.533335,27.4,38.933334,50.05556,55.966667,56.75,60.288887,72.95833,72.04445,72.71667,89.17778,94.058334,83.933334,72.51111,47.449997,24.58889,13.775001,4.8111115,0.77500004,0.2777778,0.011111111,0.0,0.0,0.0,0.14444444,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15833333,1.5666667,0.7916667,0.26666668,1.2666667,1.5777779,0.50000006,0.11666667,0.31111112,0.5916667,0.23333335,0.075,0.7555556,0.6333334,0.5083333,0.06666667,0.04166667,0.022222223,0.0,0.12222223,0.11666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,3.0833335,7.1555557,0.0,0.0,0.0,0.06666667,0.08888889,0.0,0.0,0.0,0.0,0.0,0.15,0.0,0.0,0.0,0.0,0.0,1.6222222,0.96666676,1.9444444,2.9583335,12.677778,6.558334,2.0111113,1.5416669,0.35555556,1.3333333,1.5916668,0.18888889,0.0,0.022222223,0.3628788,5.5666666,1.5444443,1.6416667,0.41111112,0.68333334,0.44444442,0.51666665,0.17777778,0.0,0.0,0.2888889,26.483334,34.066666,5.5333333,2.6111112,0.0,0.0,0.73333335,1.2666667,0.022222223,0.34166667,1.488889,1.4931818,1.9777777,0.06666667,0.016666668,0.044444446,0.7492424,0.87777776,2.3083334,6.922222,13.241666,6.188889,4.5333333,4.975,3.9999998,1.2666667,0.0,0.0,0.08888889,0.4666667,1.0833334,1.2666667,2.0083334,2.2,1.45,0.5,0.33333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.22222222,0.29999998,0.17777778,2.0666666,1.1999999,0.30833334,0.28888887,1.2111111,3.3416672,3.9222226,7.85,14.688889,4.966667,4.4111104,3.7444446,1.825,0.6555556,0.22500001,0.07777778,0.12500001,0.14444445,0.17500001,0.21111111,0.70000005,1.2416666,2.0444443,2.275,2.2555554,2.1583335,1.8666667,1.8333333,2.8666668,5.7333336,7.4333334,6.233333,5.916667,6.4,8.477779,11.324999,12.622222,9.891667,7.7222214,8.083333,7.9555554,8.5,8.98889,9.900002,8.975,9.766668,12.541666,17.911112,23.616669,31.411114,42.744446,54.45,66.333336,74.54167,72.833336,69.55,72.75556,76.01666,80.21111,86.8,83.50833,53.81111,27.808334,16.97778,6.0916667,1.3,0.35555556,0.016666668,0.022222223,0.025,0.055555556,0.16666669,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.73125,0.0,1.3583332,0.0,0.0,0.0,0.0,0.0,0.14999999,0.0,0.3,1.0999999,0.19999999,1.4666667,0.29375,0.025000002,0.51875,1.2166666,0.23333335,0.112500004,0.5500001,0.9562501,1.3916667,1.0125,0.89166677,0.7477273,0.24375,0.0,0.0,0.025,0.05,0.0,0.01875,0.0,0.0,0.0,0.0,0.0,1.0166668,2.53125,0.13333334,0.008333334,0.0,0.0,0.35,0.15,0.9375,0.775,0.40000004,0.25,0.075,0.925,3.725,0.33125,0.0,0.0,0.0,0.0,1.7375001,4.966667,1.5625,0.033333335,0.0,0.0,0.0,0.5,4.225,11.987501,8.516666,7.2750006,10.825001,9.10625,2.266667,1.5666667,4.5624995,3.3416667,1.39375,0.77500004,0.33125,0.8666667,0.38333333,2.1312501,0.72499996,1.1625,1.0166667,0.83125,0.15833333,0.0,0.0,0.0,1.5875,2.1166666,0.0,0.0,0.0,0.0,0.15833335,1.5250001,2.6166666,1.5500001,1.6181818,1.73125,1.0333333,0.36666667,0.25,1.8083334,3.0062501,2.1833334,2.94375,4.0,5.19375,0.91666675,0.70000005,0.8999999,0.9166666,0.425,0.0,0.0,0.0,0.09166667,0.1875,0.46666667,1.0,0.73333335,0.29375,0.13333334,0.15833336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.1875,0.18333335,0.00625,0.575,3.2750003,7.3125,7.083334,5.5312495,1.9666668,1.5500001,1.0749999,0.6750001,0.16250001,0.0,0.0,0.0,0.01875,0.125,0.42499998,0.8416667,1.2916666,1.79375,1.9916668,1.5250001,0.975,0.9375,0.8250001,1.1750001,2.6,6.0416665,7.3750005,8.258334,7.75625,6.0750003,5.2333336,5.425,7.2249994,6.9750004,6.125,6.0624995,7.05,7.99375,8.166667,8.166667,7.8249993,8.625,10.631249,13.483335,18.1375,22.975,29.733334,43.562504,58.333336,70.33125,71.90834,73.175,77.60834,78.8375,78.15,79.100006,81.53125,72.74167,52.825,37.291668,25.525,10.725,2.5500002,1.18125,0.16666667,0.28750002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7166667,0.0,0.0,0.0,1.488889,0.36666667,0.0,0.0,0.0,0.54444444,0.4166667,2.0222223,0.8083333,0.0,0.5333333,0.0,0.0,0.5333333,0.45555556,1.2333333,0.2777778,0.5,0.7777778,0.10000001,0.97777784,1.2138889,0.0,0.0,0.0,0.08888889,0.275,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2111111,2.5,0.51111114,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,1.2166668,0.92222226,0.2916667,3.322222,0.70000005,0.0,0.0,0.0,0.0,0.0,0.3111111,1.5916667,0.9777777,0.45833334,0.06666667,0.0,0.041666668,0.34444445,3.6333337,7.633333,10.3,5.922222,2.5,4.411111,3.8555555,6.5575757,4.2444444,2.5583334,2.5,0.3416667,0.3333333,0.7222222,0.9916667,1.2555556,1.5250001,0.0,0.0,0.0,0.1,0.21666668,0.10000001,0.09166667,0.0,0.0,0.0,0.0,0.0,2.5222225,4.8500004,1.9555556,1.7666668,1.4555556,1.0416667,0.8666667,1.6111112,2.3,3.3809524,1.8636364,0.8819445,0.43333334,0.975,0.36666667,0.07777777,0.8111111,2.0666668,2.7555559,0.22500001,0.0,0.0,0.022222223,0.0,0.15,0.12222223,0.125,0.011111111,0.016666668,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,2.5666666,6.8555555,5.675,3.6222222,1.4916668,1.7,1.0916667,0.6444444,0.33333334,0.11666667,0.0,0.0,0.0,0.0,0.20000002,0.45833337,0.4555556,0.36666667,0.33333337,0.38888893,0.35833332,0.3,0.13333334,0.0,0.08888889,0.6000001,2.5777776,5.5499997,10.622221,6.533334,5.622222,8.122222,10.058334,5.733333,4.1000004,4.1555557,5.383334,6.577778,7.1,7.1888885,7.188889,6.491667,5.7,8.066667,11.655557,14.266666,18.788889,22.100002,31.241665,45.77778,60.55,69.73334,73.958336,78.477776,80.925,81.55555,76.67778,72.7,71.13333,66.59167,56.488888,37.758335,22.333334,11.544445,4.4333334,1.7111113,1.0000001,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.11111111,0.0,0.2875,0.43333334,0.76666665,0.0,0.5833334,0.8625,0.90833336,0.0,0.8166667,1.6916667,0.19999999,0.15,0.8812501,0.083333336,0.0,0.0,0.2875,0.26666668,3.9916668,2.2250001,0.06666667,0.175,0.2,0.49999997,0.33939397,0.25227273,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4125,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32500002,0.18125002,0.0,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.11875,1.225,0.50625,1.425,0.5583333,0.14375001,1.4333334,2.2125,4.583333,5.793751,4.2749996,1.19375,0.7416667,3.35,14.206248,10.025002,0.78125,0.19166668,0.09107143,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.26875,0.26666668,0.06875,0.0,0.0,0.0,0.0,0.0,0.28333336,0.63125,0.675,0.8625,1.1500001,1.375,2.6,3.516667,2.4625,3.7166667,1.54375,0.625,0.20625,0.016666668,0.0,0.23333333,0.54166675,3.31875,2.05,0.13125,0.0,0.0,0.0,0.0,0.043750003,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.0,0.0,0.05,0.26666668,3.2749996,2.4750001,0.09166667,0.17500001,1.3833334,1.70625,0.79999995,0.39166668,0.05,0.0,0.0,0.0,0.00625,0.033333335,0.01875,0.0,0.0,0.0,0.0,0.07500001,0.08333334,0.03125,0.0,0.0,0.00625,0.033333335,0.23750001,0.8,1.9312501,5.9,10.508334,11.787499,8.683332,6.3375,5.3,4.36875,5.416667,6.6812496,6.7083325,6.6000004,7.3625,7.0916667,6.5812507,6.975,9.249999,12.283333,15.816668,24.41875,36.99167,51.8125,60.73334,70.087494,80.733345,86.3,84.49999,80.441666,73.45,67.200005,61.60625,59.34167,58.231255,51.81667,31.416666,11.050001,4.1500006,2.60625,0.975,0.5,0.30833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17500001,0.275,0.0,1.6333333,1.4222221,0.0,0.0,2.3888888,0.0,0.0,0.0,0.0,0.41111112,1.0666666,0.56666666,0.55,0.17777778,1.8333334,2.5666666,0.72499996,0.12222223,1.4666666,1.0340909,1.0,0.16666667,0.25555557,1.3431818,0.0,0.0,0.47651517,1.1777778,0.4666667,0.0,0.0,0.0,0.0,0.08888889,0.40000004,0.26666668,0.022222223,0.016666668,0.0,0.0,0.0,0.10000001,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.37777776,0.075,0.24444443,0.2916667,0.0,0.0,0.0,0.0,0.0,0.099999994,0.375,2.1888888,4.033334,1.7333333,1.1555556,3.625,3.466667,4.1,3.3777776,0.14166668,0.0,0.07777777,0.85833335,1.3999999,1.0833335,4.3111115,2.9666667,1.2,0.022222223,0.0,0.0,0.0,0.0,0.0,0.31111112,1.9444444,2.6333337,1.7888889,1.7916667,1.1888889,0.058333337,0.18888888,0.033333335,0.0,0.0,0.0,0.055555556,0.20833334,0.33333334,0.45833337,0.43333334,1.0,3.1583335,4.5,1.3249999,0.022222223,0.0,0.0,0.0,0.033333335,1.0888889,2.8833334,0.33333334,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777777,0.0,0.0,0.0,0.0,0.0,0.35833335,0.0,0.041666668,0.41111112,0.23333335,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.2888889,0.016666668,0.0,0.0,0.0,0.0,0.1,0.62222224,1.275,2.6111112,6.444444,10.200001,9.011112,8.8,8.98889,6.8,5.144445,6.7916665,7.9888897,7.9111114,9.641667,10.477778,10.566667,9.088889,7.3916664,7.6222224,9.733334,14.991667,26.855556,40.458336,51.844437,60.391666,69.26667,81.26668,87.22222,84.44444,76.45,71.55555,66.26667,60.000008,60.24167,60.622223,47.444443,33.0,17.355556,11.616667,7.055556,3.333333,2.688889,1.35,0.3888889,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.6666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28750002,1.6083333,2.8500001,0.89374995,0.98333335,0.69374996,0.49166667,0.0,0.0,1.0333333,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.675,0.76666665,0.35625002,0.73333335,0.2375,0.0,0.38125002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,0.7526785,0.34583333,0.11875,0.13333334,0.2125,0.0,0.075,0.1375,0.058333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.033333335,0.2125,0.35833335,2.01875,0.64166665,0.2,0.0,0.0,0.0,0.0,0.0,0.4166667,1.4333333,1.9187499,0.21666667,0.69375,3.0583334,6.1875005,10.375,0.4375,0.0,0.53333336,0.5875,0.24166666,0.73125005,0.98333323,0.6375,0.8666666,0.23000002,0.0,0.0,0.0,0.0,0.0,0.0,0.43333334,2.9,4.3,2.08125,0.825,0.58125,0.3166667,0.04375,0.0,0.0,0.0,0.0,0.0,0.033333335,0.081250004,0.0,0.38333336,1.9312501,1.0083334,0.15625001,0.0,0.0,0.0,0.0,0.26666668,0.85833335,0.925,0.0,0.0,0.0,0.0,0.0,0.0,0.056250002,0.050000004,0.1,0.36666667,0.0375,0.0,0.0,0.0,0.016666668,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.0375,0.0,0.0,0.0,0.0,0.043750003,0.79999995,0.275,0.0,0.0,0.0,0.0,0.0125,0.15833333,0.7687501,1.2083334,1.4250002,1.8625,2.391667,4.1,6.0916667,7.40625,7.508333,6.5999994,6.333333,7.066666,8.3375,16.258333,16.587502,14.758334,12.5625,9.650001,8.075,8.89375,13.858334,23.325,34.0,43.749996,54.366665,65.4875,73.65,79.89166,76.7625,69.55,61.843754,58.891663,58.750004,54.8,38.541668,35.71875,30.391666,24.962502,22.399998,12.325,4.7416663,3.4562497,2.475,2.5583334,1.3375001,0.30833337,0.0375,0.0,0.275,0.3,0.13333334,1.3937501,1.8833333,0.20625001,0.16666669,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9166667,0.56666666,1.7555556,0.35833335,0.36666667,0.43333334,2.8222222,0.5416667,1.4444444,0.25555557,0.0,0.7111111,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.65555555,0.15,0.0,0.0,0.0,0.0,0.0,0.34027776,0.72916675,3.1222222,0.93333334,0.31111112,0.14444445,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777778,0.025,0.0,0.0,0.044444446,0.05,0.11111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.15555556,0.06666667,0.0,1.409091,4.2555556,0.82500005,0.0,0.57777774,0.9583334,1.5222223,0.48712122,0.06666667,0.16060606,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5222222,0.65833336,0.65555555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3416667,0.5222223,0.116666675,0.0,0.0,0.0,0.0,0.24444446,0.23333332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.575,0.16666667,1.4833333,2.0555556,0.016666668,0.0,0.022222223,0.058333334,0.18888889,0.15,0.044444446,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.41111112,0.3222222,0.19166666,0.15555555,0.0,0.13333334,0.29166666,0.0,0.0,0.0,0.0,0.025,0.044444446,0.27500004,0.4666667,0.6444444,0.48333332,0.44444445,0.79166675,0.62222236,1.5916667,3.9111109,5.1916666,5.1777782,3.877778,3.3666668,7.233333,17.491665,21.833334,18.85,15.68889,13.044444,10.874999,11.144445,14.875001,20.777777,26.616667,34.666668,45.516666,57.644447,61.955555,63.091667,62.911114,58.475,54.61111,54.591667,54.100002,44.13333,35.258335,35.888885,35.600002,31.355556,19.366665,6.1666665,5.075,5.588889,5.766667,2.4083335,1.3000001,0.6583333,0.14444445,0.45833328,0.3111111,1.2555556,3.8083336,3.8,1.9416667,1.3222222,0.19166668,0.9111111,0.11111111,0.033333335,0.0,0.0,0.0,0.0,0.0,0.19166668,1.4000001,0.0,0.0,0.0,0.0,1.75,0.5416667,2.925,0.23750001,0.0,0.225,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16250001,0.06666667,0.0,0.3,0.0,0.0,0.0,0.0,0.0,0.0,0.21666667,0.55625004,0.59999996,4.3250003,2.0416667,1.0333334,0.40625003,0.008333334,0.0125,0.0,0.0,0.0,0.0,0.0,0.14166667,0.23125,0.26666668,0.0,0.06666667,0.14374998,0.19166666,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.5833334,1.41875,1.7083335,1.4660027,0.60833335,0.175,0.0,0.10000001,1.0374999,2.141667,1.4812502,0.39166668,0.05267857,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.14166667,0.3625,0.39166668,0.975,1.3062501,0.058333337,0.0125,0.0,0.0,0.0,0.01875,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4083334,1.4250001,1.1666666,6.9750004,1.0083333,0.0,0.48333335,0.7916667,1.1999999,1.2750001,1.5250001,0.8083333,0.10625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.32500002,2.24375,3.5250006,3.9333334,4.3,1.4749999,0.23124999,0.13333334,0.112500004,0.0,0.05,0.050000004,0.25000003,0.5375,0.875,0.77500004,0.7916666,0.9833334,0.69374996,0.5083333,0.425,0.22500001,0.11250001,0.13333334,1.4875,2.5916665,2.9833333,2.5499997,1.9583334,2.88125,7.6750007,11.399999,10.558332,10.775,11.093751,12.75,13.325,15.266666,21.03125,25.641666,31.06875,40.275,48.433334,56.437496,59.541664,59.18125,57.733334,52.2,42.850002,45.341667,41.85625,38.36667,37.66875,35.691666,24.575,18.2,9.55,9.341666,13.466667,14.04375,2.716667,1.9312501,0.6416667,0.17500001,0.033333335,1.1583333,2.05625,3.3583336,4.14,3.3833334,1.4250001,1.3333333,0.5833333,0.46875,0.77500004,0.24375002,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.40833333,0.0,1.4083333,0.7222222,0.65555555,0.46666664,0.2,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20000002,0.39999998,0.08888889,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7777778,2.9583335,2.2666667,2.3500001,1.5888889,0.53333336,0.108333334,0.11111112,0.19166668,0.17777778,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,1.3888888,3.8972223,6.8111115,6.125,5.1000004,2.0916667,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28333333,0.5555556,0.6,0.22222222,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5833334,2.3777776,1.25,0.64444447,0.70000005,0.0,0.0,0.0,0.2777778,0.35833335,0.033333335,0.041666668,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,1.4777778,2.4444444,0.8583334,4.3444448,4.175,0.11111111,0.7166667,2.7888892,3.6222222,3.216667,3.722222,4.8750005,0.9555556,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14166667,2.4222221,6.3749995,12.122223,10.78889,4.5,0.88888896,0.45833334,0.022222223,0.025,0.0,0.15555556,0.28333333,0.5888889,1.25,1.7555557,1.525,1.1888889,1.1333333,1.0583333,0.8333333,0.4666667,0.65555567,0.19166668,0.044444446,0.20000002,0.7111111,1.7111112,2.1000001,2.0555556,1.5583334,1.4777778,2.9583335,4.7666664,5.9000006,6.2666664,7.8888893,10.95,12.4777775,13.391666,16.58889,18.975002,22.266665,28.677778,39.283333,49.5,56.80834,58.08889,54.658333,52.666664,54.211113,56.0,50.855556,45.108334,38.966667,32.06667,28.966663,24.633333,29.188889,37.266663,32.274998,8.0,2.9833338,1.088889,0.875,0.5,0.6000001,0.925,1.6777779,3.7166665,3.5333333,2.6,1.3000001,0.70000005,0.16666667,0.0,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,1.7888889,0.36666667,0.36666667,0.0,0.7222222,0.73333335,0.5833334,0.0,0.45,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.08888889,0.0,0.22222224,1.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,3.4333334,5.8333335,4.533334,4.322222,1.9555557,1.3416667,1.6666667,0.9000001,0.33333337,0.18333335,0.0,0.0,0.0,0.0,0.016666668,0.14444444,0.8666667,1.0,0.68333334,0.46666673,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.85,5.033334,7.8999996,5.2222223,2.858333,0.35555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5111111,1.5250001,1.2222222,1.1583334,0.34444445,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44166672,1.1888888,0.09166667,0.41111112,0.0,0.0,0.0,0.0,2.2333333,0.43333334,0.055555556,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.52500004,1.988889,1.688889,1.0833334,3.7666667,1.0166667,0.41111112,5.1499996,6.311111,5.577778,3.7000003,7.5777783,4.591666,0.7444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32500002,2.6444445,4.6333337,7.533333,9.591666,6.1666675,2.3555555,0.6,0.11111111,0.033333335,0.033333335,0.1,0.1,0.41111112,0.9166667,1.2222222,1.3249999,1.8777779,2.1666667,1.8777779,1.4222224,1.3333334,1.3666667,1.0666666,0.5222222,0.9333334,0.022222223,0.016666668,0.10000001,0.42222223,1.2416667,1.7,3.3083334,3.9,1.7916667,1.2555556,1.7555557,3.233333,4.288889,5.475,6.888889,7.2416663,7.8888893,9.574999,11.555555,14.9,22.016665,27.611115,34.3,44.744446,51.166664,56.199997,67.72223,67.75,68.01111,58.441666,45.61111,31.933332,24.566666,26.691666,33.22222,39.32222,48.94167,29.466667,3.3416667,0.6555556,0.975,1.5222222,1.288889,1.025,1.3333334,1.0333334,1.888889,2.275,3.7555556,2.5666666,0.7583333,0.1888889,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.15,1.1187501,0.38333336,1.8874999,0.53333336,0.2,0.3625,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,2.6625001,4.383333,2.325,1.2416668,0.99999994,1.93125,3.8250003,6.0562496,2.875,0.59375,0.041666668,0.1,0.15,0.0,0.28750002,0.7166667,1.5749999,2.7583332,3.5562499,3.0583336,2.4416666,1.575,0.17500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40535718,1.125,0.6504487,0.21818182,0.10833334,0.14375,0.7916666,2.0125,0.84166664,2.58125,0.0,0.0,1.53125,4.2,4.5125,3.2749999,1.7624998,0.43333334,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.016666668,0.0,0.0,0.0,0.0,0.0,0.2625,0.3,0.0625,0.025,0.25,0.14166668,0.06666667,0.05,0.1,0.15,0.058333337,0.38125002,0.65,1.2416667,1.06875,1.5250001,1.4312501,6.1916666,9.856251,5.9083333,4.75,4.3125,7.0666676,2.5499997,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.10000002,0.008333334,0.01875,0.008333334,0.0,0.0,0.0,0.05,0.35625,0.47500002,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.15,0.008333334,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.80625,1.0833334,0.46875,0.575,0.14375,0.075,0.0,0.0,0.0,0.1125,0.38333333,0.056250002,0.6333334,0.75000006,1.75625,3.7083335,3.2812498,2.5416665,2.625,2.1083333,1.9083333,1.66875,1.4666668,1.2374998,0.7333333,0.31250003,0.17500001,0.3125,0.3666667,1.2166667,2.3999999,2.8166668,2.5687501,4.4,4.7125,1.9416667,1.3166666,1.3750001,1.55,2.1062498,2.9083333,2.5062501,2.4166667,3.7062502,4.4833336,5.6583333,8.337501,9.633333,12.143749,15.416667,24.125004,32.25,40.475002,45.875,50.566666,46.193752,37.000004,31.881248,26.900002,24.937502,25.791666,40.524998,59.481255,41.55833,15.450001,6.275,1.74375,1.4749999,2.1250002,2.3125,2.5500002,1.66875,2.1916668,2.4125001,3.4666667,2.8583336,1.49375,0.975,0.46250004,0.050000004,0.1875,0.0,0.0,1.0666667,0.40000004,0.22222224,1.175,0.25555557,0.19166668,0.44444445,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25555557,0.041666668,0.53333336,0.6111111,1.1166668,1.1222222,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20833334,0.6333334,2.1166668,1.8222222,1.011111,1.0916667,2.1111112,2.8666668,6.211111,3.4916668,1.2555556,0.29999998,0.39166668,0.22222224,0.09166667,0.4222222,1.5499998,3.122222,5.316667,5.7444444,4.6000004,3.0083334,1.6222222,0.90000004,0.18888888,0.20833334,0.044444446,0.0,0.0,0.0,0.075,0.033333335,0.108333334,0.28571427,0.033333335,0.0,0.0,0.275,1.3222222,5.133333,13.266667,12.433335,1.0333333,0.25555557,0.5083333,0.56666666,0.77500004,0.5111111,0.35000002,0.055555556,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40000004,0.13333334,0.033333335,0.0,0.7777778,0.7000001,0.6,0.74444443,1.1750001,1.5777777,0.95000005,1.0000001,2.391667,5.233333,2.6222224,4.5,4.7444444,6.416667,10.211111,5.3749995,3.3111112,2.3666668,4.2666664,1.8,0.3,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.14444445,0.31666666,0.21111113,0.14444445,0.15000002,0.055555556,0.0,0.0,0.0,0.22222222,0.5833334,0.3555556,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.05,0.06666667,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.18888889,0.5416667,0.62222224,1.2666667,3.241667,7.6222224,5.8416667,2.9111116,2.9333334,2.0111113,0.9444445,0.45000005,0.12222223,0.95,2.2555554,0.55,1.8888891,3.425,6.2444444,5.188889,6.616667,8.544444,6.8333335,5.288889,2.925,1.8888888,1.7444445,1.525,2.3222222,3.3166666,3.611111,2.5083334,1.5,0.73333335,0.67777777,1.4333333,2.4750001,3.9,3.9750004,4.033334,5.5166664,10.433333,18.144445,25.766666,31.877779,31.833336,28.666666,27.016668,26.28889,25.158333,27.644445,34.9,42.508335,39.82222,25.116669,11.400001,4.966667,2.3555558,1.8333334,2.6999998,3.277778,1.7833333,1.4888891,2.7083335,3.7444444,4.0444446,3.2333333,2.4444444,2.025,1.4222221,1.0250001,0.0,0.0,1.4916667,3.5125,1.325,0.63750005,0.0,0.2625,0.78333336,0.45,0.15,2.7333333,0.0,0.0,0.0,0.0,0.0,0.15,0.0,0.0,0.0,0.0,0.0,0.08125,0.95000005,1.2750001,0.75625,0.5083333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.2,0.275,0.29999998,0.25,0.59375,1.0833334,1.7562499,2.325,2.8500004,2.1,1.4000001,0.88750005,0.33333334,0.20625001,0.16666669,0.35,0.89166665,1.8999999,3.5249999,4.1749997,3.2812502,1.475,0.6125,0.59166664,1.075,0.62500006,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,0.72499996,0.9250001,0.13333334,0.06875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.23333335,0.15,0.0,0.0,0.0,0.2125,1.9083333,1.4812499,1.925,2.8250003,4.01875,4.275,3.5375001,7.258333,11.637501,9.625,9.258333,7.9125,6.2416663,6.9124994,4.3416667,2.38125,1.9,1.9666666,0.3625,0.0,0.075,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0375,0.025000002,0.23750001,0.7833333,0.86875,0.9333334,0.55,0.16250002,0.0,0.15625001,0.23333335,0.27499998,0.5,0.1875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,2.2250001,5.5499997,7.8750005,10.358333,10.868752,11.608335,13.062501,13.758333,9.599999,5.11875,1.5083333,0.3125,0.8833333,2.59375,8.95,17.012499,12.575001,15.033333,16.64375,16.316668,14.437501,11.991667,8.28125,6.7916665,7.625,7.55,8.241668,10.0875,9.233334,5.725,2.6833334,1.1312499,0.47500002,0.25,0.56875,1.6750001,2.4500003,2.4083333,2.6937501,3.2666664,6.3666663,11.743751,18.533333,24.575,27.591667,28.0,25.85,25.2375,24.866667,28.783333,31.037498,31.441668,33.525,29.191668,17.612501,7.9999995,4.6333337,3.40625,3.2916665,2.1000001,1.15,1.7812499,2.6583333,3.0416667,3.7687502,4.491667,4.7562504,4.175,2.8875003,0.0,2.4444444,1.3444445,1.5750002,1.4777777,0.38333336,0.8777778,0.49166667,0.22222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.9333333,4.777778,0.96666664,1.2444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.011111111,1.5583333,0.8555555,0.2,0.5249999,1.3000001,1.7000002,1.7777779,2.0750003,2.4444447,2.6999998,3.5249999,3.744445,2.1499999,0.18888889,0.1,0.16666667,0.8166666,1.5555556,1.8777778,2.4250002,2.5444446,3.1666665,2.5,2.6,1.7111113,0.50000006,0.38333336,0.26666668,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.36666667,0.425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.16666667,0.111111104,0.025000002,0.0,0.0,0.0,1.6174244,2.7319446,3.0666668,3.377778,4.0222216,3.8916664,3.1555557,5.175,9.0222225,9.191667,8.622223,6.2666664,4.6000004,3.9666667,3.2666667,1.6333334,0.8666667,0.5222222,0.06666667,0.17500001,0.07777778,0.11666666,0.0,0.0,0.0,0.0,0.06666667,0.22222221,0.35000002,0.34444445,0.9166667,1.2666667,1.5250001,0.8777778,0.37777779,0.058333337,0.11111112,0.16666667,0.14444445,0.175,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.06666667,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6666667,2.1333334,2.641667,7.1222224,14.241667,19.777777,16.133333,8.544444,6.088889,3.525,1.7111111,0.5500001,0.42222223,0.85833335,3.4888892,8.241667,12.255556,19.733334,26.016666,21.444445,13.283334,12.933333,14.075001,13.366668,13.444444,12.891667,10.211112,8.208334,7.5666666,9.349999,7.177778,3.0249999,1.0555556,0.37777779,0.13333334,0.11111111,1.4416666,1.8666667,1.7666667,1.9777778,2.6000001,4.8,8.244446,13.866667,18.611113,23.858335,26.100002,24.783335,23.455557,25.68889,28.341667,26.233332,26.216667,31.266666,30.141665,22.411112,14.3555565,6.4083343,3.3888888,1.6083333,0.92222226,0.65833336,0.5444445,1.3555557,2.6000001,2.5222223,3.458333,5.3555555,5.675,0.0,1.7166667,1.1083335,0.46875,0.9083334,1.75,0.4666667,0.0,0.5416667,0.0,0.0,0.0,0.0,0.0,0.0,0.275,1.66875,0.0,0.0,0.3875,0.6916666,0.0,0.19999999,0.875,0.98333335,0.16666669,0.0,0.0,0.0,0.016666668,0.087500006,0.14999999,0.20625001,0.28333336,0.30833334,0.09375,0.016666668,0.0,0.0,0.3875,1.2416667,1.3416667,0.125,0.57500005,2.03125,3.3999999,2.4750001,2.0333335,1.6833336,2.28125,5.383333,6.1250005,3.975,1.0625001,0.09166667,0.1125,0.45000002,0.7166667,1.4062499,0.8416666,0.7625,1.8749999,3.5375004,4.691666,4.7000003,3.53125,2.35,0.95000005,0.15,0.0,0.0,0.00625,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056250002,0.46666667,0.53125006,0.14166667,0.033333335,0.0,0.0,0.0,0.0,2.6062498,3.1,2.5187502,1.175,2.1666667,3.05625,3.2,5.83125,7.9500012,5.9375,3.7,2.6583335,2.3937502,2.3500004,1.4562502,0.68333334,1.6687499,0.7166667,0.25833336,1.225,0.1,0.0,0.0,0.0,0.025,0.30625,0.84999996,1.3249999,0.96875,0.9916667,1.5000001,1.7416668,1.1312499,0.6666666,0.375,0.25,0.16666669,0.075,0.0,0.0,0.0,0.0,0.0,0.05,0.0,0.0,0.0,0.0,0.0,0.033333335,0.13333333,0.06875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9583334,1.8500001,2.4583333,2.05625,2.6166668,3.2833335,2.5000002,1.325,0.37500003,0.31666666,0.71875,2.9583335,8.9875,16.883335,24.833334,26.862501,26.858332,23.58125,20.975002,24.13125,23.733334,20.525,13.993752,8.35,5.1625004,4.075,5.1,6.3833337,5.76875,3.8333337,1.5583334,0.5750001,0.15833333,0.10625,0.5416667,0.58750004,0.44166666,1.2833333,2.7124999,4.675,7.0437503,10.941667,14.906251,19.291668,23.46875,23.633333,22.55,24.5125,29.933334,30.100002,28.133335,28.15625,28.091667,27.4,21.806252,11.216666,4.1875,2.5000002,1.7125,1.2083333,1.2666667,1.075,0.53333336,1.0312501,2.95,4.76875,0.0,0.0,0.17777778,1.0666667,1.3555555,2.4750001,0.85555553,0.6,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.95,0.6222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.34444445,0.56666666,0.5666666,0.18888888,0.083333336,0.0,0.0,0.08888889,0.1777778,0.5083334,0.29999998,0.025,0.4,1.9416668,2.277778,1.0888888,1.2583333,1.5333333,3.2583332,6.1000004,5.233333,2.0555556,0.6333333,0.21111111,0.22222224,0.625,0.5,0.27500004,0.13333334,0.825,3.5444446,4.6888885,5.4166665,5.444445,3.3500001,0.7111111,0.0,0.1,0.09166667,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.26666668,0.20000002,0.0,0.0,0.016666668,0.11111111,0.13333333,2.6111112,1.7833334,2.0208335,1.5,4.244445,5.777778,4.6,8.322222,6.6666665,2.9,2.675,1.5,1.5333333,1.0916667,0.7444445,0.20833334,1.2,2.8500004,0.46666664,0.77777773,1.2500001,0.0,0.016666668,0.0,0.033333335,0.6888889,1.4416666,2.2666667,2.0111113,1.1,1.8666667,1.7500001,1.0,0.92499995,0.7222222,0.4555556,0.14166668,0.07777778,0.0,0.0,0.0,0.0,0.0,0.08888889,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,0.17777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,5.083334,10.211111,11.811111,7.241667,3.2,0.6833333,0.14444445,0.71666676,2.9333334,9.841667,19.466667,25.1,27.358335,29.800001,29.991667,28.62222,29.674997,26.377779,20.255556,14.25,9.311111,6.008333,3.7222223,3.5333333,3.1555557,2.9750001,3.6444445,3.7,1.9166666,0.58888894,0.15,0.011111111,0.0,0.0,0.044444446,0.7166667,2.0111113,3.6499999,5.1444445,6.9,10.6,14.500001,18.522223,19.044445,19.425001,21.98889,25.85,27.233334,24.008333,22.355555,24.56667,28.550001,25.81111,13.533335,6.2,4.883333,3.3888888,2.2555556,2.0833335,1.1333334,0.41666663,0.13333334,0.6916667,0.0,0.7111111,1.8444446,0.6166667,0.54444444,1.9083335,0.3111111,0.4,0.0,0.0,0.0,0.0,0.0,1.4444444,0.0,0.0,0.0,0.0,0.0,0.6,0.6777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.2888889,0.3,0.48888892,0.3416667,0.0,0.0,0.21111113,0.64444447,0.25,0.011111111,0.008333334,0.0,0.108333334,0.99999994,0.9555556,0.6916666,1.3111112,1.0166667,1.3111112,3.7666667,4.733333,3.041667,1.2222223,0.6333333,0.87499994,0.6666666,0.37500006,0.033333335,0.0,0.15555556,0.54444444,1.3833333,1.8000002,0.55,0.2,0.0,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5666667,0.44444445,1.8333334,4.3333335,5.3250003,7.633333,7.4083333,5.8333335,6.4750004,7.0111113,5.7,5.3583336,4.533334,3.1083336,2.6555555,0.9083333,0.8111111,0.24444444,0.39166668,0.14444445,0.20833334,1.2666667,0.6666666,0.12222222,0.6444444,0.475,0.14444445,0.05,0.011111111,0.65833336,1.2888889,1.9500002,1.977778,1.0444446,1.4750001,1.6111112,0.8666666,0.5555556,0.6083333,0.32222226,0.06666667,0.1,0.011111111,0.0,0.0,0.0,0.0,0.0,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1777778,0.6,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4416667,4.811111,8.58889,8.516667,7.166667,2.75,0.61111116,1.3083334,4.477778,13.716667,20.933334,23.11111,24.216667,26.633331,30.650002,33.522224,28.000002,17.833334,10.577778,8.900001,7.522222,4.7166667,4.2999997,4.1833334,2.5111113,2.15,1.9,2.0666666,2.2749999,1.3111112,0.45000005,0.011111111,0.0,0.0,0.0,0.083333336,0.4666667,1.1833334,2.011111,3.7166667,5.8111115,9.525001,12.844444,15.711112,16.966667,18.155556,19.666666,20.944447,21.71667,25.233334,23.211111,22.875,23.000002,23.425001,13.7,7.2166667,5.5444446,4.7333336,3.4166665,1.5,0.425,0.011111111,0.041666668,0.23125,0.60833335,0.0,0.1,0.0,0.74375,0.31666666,0.2625,0.9,0.0,0.0,0.46666664,0.0,4.8916664,0.8125,0.0,0.0,1.1583333,1.225,1.3125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.10625,0.033333335,0.05,0.0,0.0,0.18333335,0.32500005,0.41875005,0.15000002,0.0125,0.0,0.075,0.6999999,1.2916666,1.825,0.7833333,0.49375004,0.65000004,1.0937501,1.7666668,2.88125,2.5333335,1.3333334,0.58124995,1.5166667,1.93125,2.3999999,1.475,0.39166665,0.5583333,0.51875,0.22500001,0.0,0.0,0.0125,0.025,0.06875,0.041666668,0.041666668,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.91875,5.183333,8.400001,10.15,11.933334,10.200001,8.808333,6.7625,5.716667,4.1875,4.2250004,3.983333,2.5000002,2.091667,1.5812501,0.64166665,0.5500001,0.25833333,0.40833333,0.14999999,0.2916667,0.19375001,0.7166667,0.44999996,0.058333337,0.175,0.35000002,0.23333335,0.76875,0.52500004,0.675,0.54999995,0.6562501,0.45,0.5333333,0.6749999,0.3,0.13125002,0.15833335,0.06875,0.016666668,0.05,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5666666,0.91666675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.06666667,0.5833333,1.575,2.4333334,2.075,1.9250001,3.7125,7.791667,16.41875,19.991667,21.716667,21.08125,20.716667,23.16875,18.508333,11.6625,5.4333334,2.6750002,3.0374997,3.291667,3.15625,5.908334,7.3187494,4.816666,2.78125,1.4833335,1.2,1.0562502,1.0666667,0.75000006,0.20000003,0.043750003,0.0,0.0,0.0,0.041666668,0.056250002,0.46666667,1.5812501,3.241667,4.825001,7.158334,9.875,13.24375,16.941666,19.2,20.791666,20.4375,24.191668,22.933332,20.975,19.0,18.6625,19.891666,16.1125,10.025001,8.075,8.562501,6.758333,2.55,0.4166667,0.025,0.78333336,3.3777778,5.4,4.3,1.0666666,0.95000005,0.0,0.0,0.0,0.0,0.46666664,1.9333334,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4,0.73333335,0.21666667,0.055555556,0.28333336,0.15555556,0.008333334,0.0,0.3888889,1.7666667,2.0777779,1.3833334,1.0444444,0.53333336,1.1666667,1.525,1.6666666,1.0,1.1750001,0.4888889,0.85,1.2333333,1.8249999,1.6333334,1.3222224,1.0250001,0.9222222,1.8333334,2.5000002,1.1416667,0.87777776,0.52500004,0.22222225,0.14444445,0.12500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.58888894,2.711111,4.316667,5.555556,1.475,1.4111111,1.5166664,2.1333332,2.0916665,3.1666667,2.9777775,1.2166668,0.73333335,0.35000002,0.4888889,0.35,0.0,0.07777777,0.47500005,0.1,0.22500002,0.2,0.10833335,0.11111111,0.7444445,0.78333336,1.3555555,0.85,0.36666667,0.06666667,0.011111111,0.0,0.0,0.06666667,0.033333335,0.0,0.0,0.0,0.0,0.10000001,0.05555556,0.0,0.0,0.0,0.0,0.058333334,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.2916667,0.0,0.0,1.2888889,0.8111112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.23333335,1.6444446,1.5,0.9777778,2.9,8.177778,12.733334,10.744445,13.766666,15.766666,14.2,14.491667,11.477778,6.9333334,5.933334,4.4,2.0555556,1.011111,1.4333334,1.6777779,2.8583333,4.377778,6.783333,5.9888887,5.841667,3.6222224,1.5333334,0.73333335,0.63333344,0.37500003,0.36666667,0.15833333,0.0,0.0,0.0,0.06666667,0.125,0.10000001,0.14166668,0.66666675,2.1166668,3.8333335,5.7333336,7.766667,10.933333,14.591666,16.5,19.266666,20.08889,24.22222,24.108334,22.244444,18.3,15.422221,18.375,17.088888,14.855556,11.283333,14.48889,10.4,2.311111,0.45000002,0.61875004,1.3833334,0.9416667,2.14375,1.0166667,1.83125,1.0583334,0.44374996,0.23333332,0.46666664,0.68125,0.18333334,0.0,0.0,0.0,0.41666666,0.43125,0.0,0.0,0.0,0.33333334,0.43750006,1.4666666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.025,0.18333334,0.50625,0.425,0.1,0.033333335,0.15,0.13125001,0.7,2.5875,2.6333337,2.3249998,1.325,0.74375004,1.5166667,1.9083333,1.9687501,1.0,0.85625005,1.3000001,1.53125,1.5916667,1.7583333,1.9187499,2.525,3.0,3.275,2.35625,2.025,2.125,1.4083334,0.725,0.23125002,0.05,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10000001,0.0,0.0,0.13333334,0.975,2.7,1.8124999,1.2333333,1.0250001,0.66249996,0.2916667,0.45000008,0.2666667,0.09375001,0.06666667,0.11666667,0.1125,0.016666668,0.112500004,0.24166667,0.53125,1.6833332,1.4166665,1.1,1.2583333,0.48124996,0.041666668,0.0,0.0,0.10625001,0.13333334,0.016666668,0.0,0.0,0.0,0.0,0.01875,0.041666668,0.008333334,0.0,0.0,0.0375,0.25833336,0.31875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333333,1.1812501,0.32500002,0.0,1.1666666,0.6666667,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,1.0125,1.9583335,0.44374996,0.21666667,1.4062499,5.9249997,14.758334,22.79375,27.558336,19.462502,16.0,17.175,10.775,6.36875,6.725,7.016667,8.225001,8.333334,4.76875,2.4416666,1.675,1.5,1.4333333,0.9875,0.60833335,0.61875004,0.35,0.61875,2.8333335,4.1937504,3.8416667,2.8666666,1.4812499,0.5666668,0.2625,0.15000002,0.05625,0.0,0.0,0.0,0.041666668,0.081250004,0.13333334,0.13750002,0.19166668,0.30625,1.075,2.4833333,3.7812502,5.791667,7.6875005,9.841667,13.73125,18.491667,20.866667,23.475,22.216667,21.6125,20.858335,17.81875,19.633333,16.841667,14.23125,12.074999,9.0375,4.05,2.65,0.0,0.0,0.0,0.0,0.0,0.85,0.44444448,1.275,0.9444445,0.73333335,1.9000001,0.6,0.31666666,0.0,0.0,0.0,1.4083333,1.8888891,0.34444445,3.025,4.3444443,2.1333334,2.2888887,0.35,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.08333334,0.0,0.31666666,0.71111107,0.27500004,0.2888889,0.14444445,0.008333334,0.1888889,0.49999997,1.6444445,1.7916667,2.9333334,2.0166667,1.5888889,1.7666667,2.3083334,2.7777777,1.6416668,1.3111112,0.9250001,1.6666667,3.2555556,4.041667,5.6111116,5.416667,3.9333332,3.375,3.9444444,3.175,2.4,1.7666667,1.0,0.11111111,0.11666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.47777778,1.325,0.6333333,0.49166667,0.011111111,0.0,0.0,0.0,0.0,0.0,0.175,1.6888889,2.375,1.5000001,1.2,1.2888889,0.8222223,0.50000006,0.53333336,0.35833335,0.1777778,0.14166668,0.05555556,0.0,0.0,0.0,0.15833335,0.54444444,1.8833334,1.8,0.6444445,0.85,0.6777778,0.09166667,0.0,0.0,0.17777777,0.3166667,0.0888889,0.0,0.0,0.0,0.0,0.0,0.025,0.011111111,0.0,0.0,0.0,0.06666667,0.36666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.050000004,0.25555557,0.06666667,0.0,0.0,0.022222223,0.022222223,0.0,0.0,0.0,0.25555554,2.025,0.7111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,1.175,10.444445,5.6999993,1.0333334,7.4,40.17778,45.04445,34.508335,31.566668,21.05,15.8111105,17.625,6.3666673,3.8000002,2.288889,5.2222223,2.9833333,0.8222222,0.7166667,0.6777779,0.6,0.56666666,0.79999995,0.82500005,0.35555556,0.5833333,0.033333335,0.033333335,0.011111111,0.09166667,1.5666666,2.2222223,1.8166666,1.488889,0.36666664,0.10000001,0.016666668,0.0,0.0,0.0,0.0,0.0,0.022222223,0.075,0.033333335,0.16666669,0.24444446,0.37777779,1.2750001,2.4222221,3.5250003,5.488889,8.608333,12.511111,15.011112,19.175001,21.38889,22.991669,21.900002,19.033333,23.37778,21.166668,17.95,11.066667,5.3,4.8,4.6,4.24375,0.6,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21666667,0.22500001,0.0,0.0,0.0,0.475,0.7583334,1.46875,2.0,1.1333333,2.6812499,4.608333,4.325,4.7583337,5.5812497,2.6,0.175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.93333334,0.48125002,1.0666666,0.058333337,0.08125,0.30000004,0.35625002,0.35833335,2.0125,3.291667,2.70625,1.9416668,2.3166666,2.85625,2.075,1.5500001,1.1083333,0.78125,1.0416666,1.625,4.375,7.0,7.8249993,7.5916667,5.8624997,6.466667,5.25625,4.2166667,3.4499998,1.9999999,0.95000005,0.39375,0.125,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.15,0.22500002,0.28750002,0.23333335,0.16875002,0.17500001,0.083333336,0.19375,0.40833333,0.4,0.56666666,1.15625,1.9833333,1.4499999,0.85,0.675,0.55,0.4583333,0.33749998,0.28333333,0.14375001,0.05,0.0,0.0,0.05,0.31875002,0.925,1.1500001,0.5916667,0.60833335,0.4,0.041666668,0.0,0.016666668,0.19999999,0.51666665,0.25,0.0,0.0,0.0,0.0,0.0,0.05,0.03125,0.0,0.0,0.0,0.0,0.15625,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.10000001,0.15,0.1,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.125,0.17500001,0.3625,1.0583334,0.31875,0.033333335,0.025,0.18333334,0.116666675,0.0,0.0,0.0,0.52500004,3.2125006,1.2583334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.9375001,21.15,8.975,1.425,14.731251,47.666668,34.925,7.999999,15.350001,16.6,22.333334,11.200001,7.5499997,10.39375,6.575,0.0,0.15,0.15,0.0,0.16666667,0.26874998,0.041666668,0.0,0.0,0.0,0.43125,0.575,0.39375,0.008333334,0.0,0.0,0.3083333,1.1250001,1.5583334,0.85625005,0.19166668,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.118750006,0.13333336,0.21250004,0.21666667,0.2833333,0.38124996,0.9666667,1.9000001,2.8000002,4.25625,6.616667,8.341667,10.606251,13.700002,17.06875,17.95,16.05625,14.525002,14.391666,16.725002,13.775,9.875,4.441667,3.7875004,2.5,0.79999995,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777777,0.0,1.9555557,3.011111,0.6333333,0.122222215,0.99166673,1.4666667,4.2166667,4.6888895,4.7222223,2.1083333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.81666666,1.5333333,0.36666667,0.525,0.15555556,1.125,0.7555556,0.5416667,0.78888893,0.7416668,1.4111111,2.722222,3.816667,4.9555554,3.516667,2.4555554,1.5666667,1.7444444,1.3111112,1.9666667,3.0666666,3.1916666,4.9555554,5.2333336,6.088889,4.8166666,3.6000001,1.7888889,1.2416667,1.0111111,0.46666664,0.13333334,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.15555556,0.1,0.058333337,0.07777778,0.058333334,0.044444446,0.008333334,0.044444446,0.3333333,0.925,1.0666667,1.325,2.1555557,2.6166668,1.4666667,0.90833336,0.75555557,0.6333334,0.5,0.43333334,0.3833333,0.07777778,0.18333335,0.011111111,0.0,0.0,0.06666667,0.38333336,0.68888897,0.6666667,0.5222223,0.14444445,0.0,0.05555556,0.075,0.43333337,0.6,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18333334,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.21111111,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25833333,0.7222222,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666669,0.4666667,0.3,1.7833335,1.8666667,0.44166666,0.022222223,0.16666667,0.32222223,0.13333334,0.0,0.0,0.0,0.8333333,3.8500001,1.8222222,0.05,0.11111111,0.14444445,0.25,0.26666668,0.0,0.0,0.0,0.0,1.7333333,0.4666667,10.9,6.0916667,5.6444445,12.133333,13.055555,14.588888,10.641667,14.666668,6.2666674,4.3999996,5.808334,11.222223,25.85,15.088888,2.5111113,2.1166668,0.0,0.0,0.13333334,0.8583334,0.7666667,0.24444446,0.0,0.0,1.1166667,1.8111112,1.2333333,0.6666667,0.016666668,0.0,0.0,0.025,0.26666668,0.4416667,0.011111111,0.0,0.0,0.0,0.033333335,0.06666667,0.16666669,0.2,0.2916667,0.44444445,0.2166667,0.21111113,0.21111113,0.1,0.29999998,0.56666666,1.1888889,2.2833335,3.7777777,4.4888887,6.191667,7.922222,9.258333,10.744444,12.458333,12.055556,11.566667,10.733334,9.566667,12.450001,12.811111,8.291668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6222222,0.875,1.2111112,1.5694445,0.25833333,3.3666668,3.4833333,0.4666667,0.0,0.31111112,0.7,2.1750002,4.8111115,1.1583334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31111112,1.0166667,0.15555556,0.2916667,0.16666667,0.7111111,1.1,0.08888889,0.6666667,1.3111111,1.3916667,1.2777778,0.9583333,0.9111111,1.888889,3.0833333,2.5333333,1.8083334,1.8555555,2.0333333,1.9555557,1.5888889,1.1666667,1.4666667,1.5916667,2.2555556,4.133333,5.088889,3.9499998,2.288889,0.98888886,0.8916667,0.65555555,0.30833337,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.2888889,0.45,0.41111112,0.32222223,0.26666668,0.24444446,0.17500001,0.08888889,0.1,0.40000004,0.64444447,1.3083334,2.1555552,2.8249998,2.811111,2.15,1.888889,1.6250002,0.90000004,0.5777778,0.5166667,0.4555556,0.108333334,0.16666667,0.016666668,0.033333335,0.055555556,0.24999999,0.6333333,0.975,0.8333334,0.5166667,0.15555556,0.011111111,0.05,0.14444444,0.525,0.6222222,0.18333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24444444,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.60833335,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.37499997,0.5555556,0.94444454,3.6750002,2.0,0.26666668,0.055555556,0.5083333,0.37777779,0.022222223,0.0,0.0,0.008333334,0.33333334,2.666667,1.4888889,0.21666665,0.5222222,0.67777777,1.0416667,0.8777779,0.0,0.0,0.0,0.0,0.0,0.06666667,3.5444446,2.8999999,12.988888,15.991667,23.2,39.811108,7.6333337,16.744444,7.9666667,3.4111114,4.0333333,11.066668,17.833334,9.877778,6.788889,6.2666664,2.8777778,3.4416666,0.8333334,0.62500006,0.73333335,0.055555556,0.0,0.0,0.93333334,2.3444443,2.5499997,1.1444446,0.125,0.0,0.0,0.0,0.044444446,0.19166669,0.044444446,0.0,0.0,0.0,0.1,0.16666669,0.22500002,0.22222224,0.12500001,0.07777778,0.125,0.06666667,0.099999994,0.033333335,0.0,0.39999998,0.988889,1.3916669,2.3111115,3.3333335,4.3416667,5.566667,6.533334,7.9444447,9.099999,9.900001,10.48889,10.391666,11.5222225,10.4,9.955556,11.349999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.14166667,2.75,0.725,0.75000006,0.6625,0.05,0.025,0.0,0.087500006,0.18333334,0.5083334,0.6750001,0.8333333,1.98125,1.1333334,0.625,0.3416667,0.0375,0.025,0.041666668,0.05,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.31666666,1.2125001,1.5333333,0.39999998,0.32500002,0.48333332,0.725,1.6666665,1.41875,0.43333334,0.13125001,0.28333333,0.5250001,0.24166667,0.54166675,0.74999994,1.0083333,1.7062501,1.3916667,1.0375,0.9916667,0.74166673,0.8499999,0.8833334,1.0687501,2.0166667,6.7625003,6.05,4.95,3.7166667,3.141667,2.275,1.4749999,0.74375004,0.2166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.06666667,0.15,0.26666665,0.42499998,0.375,0.44375,0.5833333,0.5416667,0.35625,0.275,0.112500004,0.2,0.49375,0.83333343,1.1666667,1.41875,1.4250001,1.1312501,0.9250001,1.0562501,0.9166667,0.8875,0.6999999,0.4416666,0.21875003,0.19166668,0.15,0.008333334,0.09375001,0.35000002,0.8166667,1.1374999,1.4666666,1.06875,0.47500002,0.10625,0.016666668,0.10833335,0.4375,0.9166666,0.575,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.34166667,0.2625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,0.81250006,0.66666675,4.2333336,5.50625,1.3,0.17500001,0.24166667,0.68750006,0.25000003,0.058333337,0.0375,0.0,0.09375,0.375,2.0937502,1.2416667,0.45,1.1750001,1.35,1.9375,1.6166667,0.0,0.0,0.0,0.0,0.0,0.0,0.28333333,0.2,2.7583332,10.54375,23.566666,17.066668,3.71875,4.108333,3.1937501,0.33333334,7.7125,10.500002,7.1124997,8.408334,11.925,10.40625,7.025,7.425,7.6333337,8.075,1.6583334,0.008333334,0.0,0.0,1.1187499,2.8083334,2.29375,3.225,4.5375,4.4916663,1.7333333,0.23125,0.1,0.27500007,0.14166668,0.09375001,0.108333334,0.116666675,0.10000001,0.16666667,0.087500006,0.05,0.0125,0.0,0.0,0.0,0.025,0.075,0.025,0.0,0.23333335,0.48749998,1.0250001,1.3916668,2.43125,3.3333335,4.74375,6.558333,7.775,9.541667,10.041667,10.0375,11.758333,12.625002,12.041666,10.956251,0.0,0.0,0.86666673,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.475,1.0,1.3416667,0.033333335,0.12222222,0.05,0.0,0.0,0.0,0.0,0.025396826,0.3333333,0.625,0.9111111,0.79166657,0.06666667,0.0,0.122222215,0.6333333,0.1777778,0.4333333,0.65,0.21111113,0.116666675,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,1.1111112,0.25833336,0.0,0.22222222,0.1,0.2,1.1416667,1.5777779,0.55833334,0.6666666,0.73333335,0.61111116,0.4777778,0.325,0.45555553,0.43333334,0.5,0.31666666,0.4222222,0.8555555,0.69166666,0.7777778,0.43333337,0.24444446,0.3416667,0.2888889,0.90000004,1.0111111,1.1999998,1.3166667,1.1222222,0.4666667,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.18333335,0.32222223,0.48333335,0.7444445,1.075,1.0444446,1.3416667,1.4999999,1.5333334,1.1250002,0.8888889,0.4083333,0.23333335,0.28333333,0.34444445,0.41111112,0.625,0.8777779,0.89166665,0.7111111,0.39166665,0.23333335,0.4666667,0.3222222,0.2777778,0.18333334,0.022222223,0.0,0.14444445,0.65,1.4333334,1.8000002,1.8000002,1.1444445,0.49166667,0.011111111,0.083333336,0.18888889,0.8222222,1.2666665,0.4,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.28333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,0.26666668,0.6555556,0.6416666,0.122222215,0.05,0.022222223,0.0,0.0,0.0,0.0,0.0,0.058333337,0.1,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.7444444,1.0916666,2.4666667,9.288889,5.0583334,0.5111111,0.058333334,0.9111111,0.5333333,0.011111111,0.12222222,0.008333334,0.0,0.26666668,0.31111112,1.4,0.8444445,0.28333333,0.9888889,1.0444444,1.4499999,1.1777778,0.0,0.0,0.0,0.0,0.0,0.0,0.11111111,0.0,1.0888889,9.808334,6.9111114,5.5000005,1.1416667,1.1222222,7.2583337,5.7000003,4.85,12.300001,3.916667,4.1444445,19.111113,18.866669,16.055555,9.433333,4.9444447,5.283333,4.0111113,3.0777779,1.0166667,0.0,0.52500004,2.4888892,5.5416665,3.5777779,3.3000002,6.844444,4.6888885,0.5166667,0.3666667,0.3916667,0.36666667,0.32500002,0.47777778,0.4888889,0.39166668,0.37777779,0.17500001,0.07777778,0.0,0.0,0.0,0.011111111,0.0,0.0,0.011111111,0.0,0.0,0.0,0.11111111,0.055555556,0.24166669,0.9555555,2.4083335,4.5444446,6.516667,8.955556,9.366667,10.066668,10.466667,11.450001,14.511112,13.275001,0.17500001,2.0083334,0.24166666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.16666667,0.0375,0.86666673,0.62500006,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.0,0.016666668,0.20625001,0.375,0.51250005,0.15,0.075,0.13333334,0.225,0.2916667,0.6666667,0.45000002,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.48333335,0.925,0.3,0.15,0.0125,0.008333334,0.275,0.76666665,1.1187501,0.95,1.0,1.8166666,2.266667,1.8375,0.8166666,0.8312501,0.77500004,0.70625,0.39166665,0.22500001,0.19375001,0.275,0.38124996,0.7,0.60625005,0.4166667,0.3625,0.80833334,0.13333334,0.26250002,0.44166666,0.275,0.18333332,0.33125,0.21666668,0.30833334,0.27499998,0.29999998,0.25,0.033333335,0.0,0.0,0.016666668,0.112500004,0.26666668,0.38125002,0.6333334,0.88125,1.0333334,1.1937501,1.2416666,1.3416666,1.025,0.7333334,0.41875,0.19166668,0.0125,0.0,0.033333335,0.118750006,0.22500002,0.3125,0.25833333,0.275,0.2833333,0.26874998,0.23333335,0.075,0.081250004,0.14166667,0.79375005,1.8416667,2.23125,2.4416666,1.9500002,1.1,0.37500003,0.056250002,0.1,0.46874997,0.95833355,0.59999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.3125,0.675,0.84375,0.975,0.9749999,0.7374999,0.4166667,0.16250001,0.016666668,0.0,0.0,0.0,0.0,0.0,0.03125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3875,0.94166666,1.46875,7.0833335,12.1,3.875,0.31666666,0.10000001,1.1666667,0.53125,0.083333336,0.050000004,0.0,0.0,0.33749998,0.15833335,0.5625,0.4166667,0.0375,0.125,0.19166665,0.26249996,0.18333332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24375,4.3083334,6.33125,4.1750007,0.325,0.0,0.0,0.0,2.4750001,7.7874994,6.3583336,4.28125,3.1,14.241667,11.625,8.308334,7.8812504,2.1083333,1.9749999,4.25,6.491667,5.0937505,3.3666668,6.0250006,2.2416668,2.2375002,2.3416667,2.85,2.9416666,1.5500001,0.81875,1.05,0.9875001,1.1916666,1.0125,0.52500004,0.5666667,0.725,0.55833334,0.56874996,0.30833334,0.20000002,0.13333334,0.12500001,0.13333334,0.083333336,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.20625001,0.8833333,2.7999997,4.975,6.7916665,7.7687507,8.625,10.05625,11.291667,11.987499,0.0,0.0,0.0,0.0,0.32222223,0.8000001,1.8333335,3.0333333,0.0,0.0,0.0,0.0,0.0,0.37777776,0.70000005,0.27777776,0.0,0.0,0.34444445,0.18333334,1.2,0.6666666,0.46666664,0.2916667,0.4222222,0.13333334,0.016666668,0.0,0.041666668,0.14444445,0.14166667,0.24444446,0.36666667,0.50000006,0.31111112,0.75,0.23333335,0.033333335,0.17777778,0.21666668,0.0,0.0,0.0,0.0,0.0,0.055555556,0.23333333,0.08888889,0.44444445,0.5,0.36666667,0.2916667,0.24444446,0.69166666,1.6555556,1.0083334,0.9777778,1.5888889,1.4,0.98888886,1.25,1.1777778,0.53333336,0.48888886,0.31111112,0.4,0.3555556,0.5166667,1.5666668,1.9083333,0.9111112,1.8583333,3.477778,2.0555558,1.275,1.0444444,0.57500005,0.5222222,0.9916667,1.0666666,1.4444444,1.175,1.2333333,0.96666676,0.11111112,0.016666668,0.0,0.0,0.008333334,0.0,0.025,0.16666669,0.3,0.47777778,0.52500004,0.7888889,0.9888889,1.0166668,1.1222223,1.0583334,0.90000004,0.48333335,0.44444448,0.17777778,0.175,0.06666667,0.05,0.0,0.008333334,0.044444446,0.41666666,0.8777778,1.3777778,1.6833334,2.0222223,2.6833336,2.6888888,2.7833333,2.233333,1.3444445,0.375,0.15555556,0.1,0.06666667,0.0,0.0,0.17777778,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20833334,0.7,0.8333333,0.8111111,0.8249999,0.6666667,0.47777778,0.32500002,0.20000002,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.65,1.5222223,2.6499999,11.733335,13.977778,3.6916666,0.4,0.14999999,1.6666667,0.77500004,0.12222223,0.0,0.0,0.0,0.39999998,0.11111113,0.29999998,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,1.7666668,3.675,5.788889,11.444445,0.625,0.0,0.0,0.78888893,0.0,0.0,0.0,0.0,2.5111113,14.799999,4.855556,1.0333333,1.3111111,1.4833332,0.5222222,0.099999994,4.508333,11.811111,13.2,7.5888886,2.9416668,2.477778,2.7333336,3.1222224,2.3888888,1.5999999,1.4000001,1.725,1.5555556,1.375,0.8000001,0.6888889,0.8666668,0.96666664,0.90000004,0.6888889,0.7833334,0.78888893,0.40833336,0.3666667,0.1888889,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,0.23333335,0.5222222,0.6583334,1.5111111,3.0111113,5.425,7.1111116,6.858333,7.688889,7.783334,0.37500003,1.2333333,2.425,1.3812499,0.0,0.55625004,3.9267676,17.92125,14.843183,5.6166663,1.9625001,0.40000004,0.3125,0.21666667,0.425,1.1833334,2.2125,0.10000001,0.5833334,0.625,7.6416674,5.5,1.4416666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.90625006,0.45833334,0.05,0.11666667,0.4583333,0.9625,0.7583333,0.20625,0.49166667,0.83750004,0.5916667,0.5,0.13125001,0.16666667,0.05,0.083333336,0.225,0.4666667,0.575,0.30000004,0.275,0.13750002,0.19999999,0.41875002,0.69166666,0.725,0.8166666,1.6166666,1.8187499,1.4166667,1.11875,0.9916667,0.6,0.51666665,0.38333336,0.29375,1.7833335,6.5375004,3.6166668,1.075,0.58333325,1.4625,2.3333333,3.0750003,2.7875001,2.05,1.51875,1.3583335,1.2500001,1.3666667,1.4333334,0.95,0.6666667,0.49375,0.083333336,0.05,0.025000002,0.083333336,0.05625,0.18333334,0.35000002,0.7166667,1.2,1.9833333,2.9187503,3.6166666,4.6916666,4.9125,5.533334,5.3875,5.141667,4.80625,4.7250004,3.9583335,3.10625,2.7166667,1.0250001,0.34166667,0.31875,0.91666657,1.6249999,2.0583336,2.0416667,1.73125,1.4416667,1.2500001,1.2833333,0.9625,0.45833337,0.16666669,0.081250004,0.025,0.0,0.033333335,0.61875004,1.0666667,0.24166667,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.5083333,1.1749998,1.4333332,1.1875,0.9166667,0.6875,0.62500006,0.40000004,0.26250002,0.050000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056250002,0.19166668,1.33125,2.4166667,7.23125,16.933334,13.183334,3.2062497,0.35000002,0.44375,1.625,0.66249996,0.17500001,0.0,0.0,0.0,0.61875004,0.116666675,0.43750006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.65000004,1.6,0.5916667,0.0,0.0,0.0,0.6166667,0.425,0.0,0.0,0.0,0.06666667,10.643749,13.458334,2.8187501,2.825,2.56875,9.874999,16.783333,20.0375,15.891666,3.14375,6.3333335,8.568751,6.4666667,4.1625,3.4416666,2.4583335,1.6062499,1.3916667,1.7749999,1.375,1.4375001,0.8333334,0.5916667,0.70625,0.9083334,1.5812501,1.4166667,1.69375,2.8166666,1.21875,0.43333337,0.27500004,0.15625003,0.083333336,0.09375001,0.025000002,0.00625,0.0,0.0,0.0,0.0,0.056250006,0.25833336,0.70000005,1.0833335,1.5000001,2.0125003,3.5666666,4.9875,5.991667,6.5000005,0.0,1.988889,3.2555556,2.85,3.0777779,4.8916664,1.977778,1.85,4.81746,7.2763886,6.8944445,8.506945,3.315909,1.4444444,0.6166667,0.011111111,0.20833334,1.8111112,1.1666667,0.70833343,0.0,0.0,0.0,0.0,0.0,0.111111104,0.083333336,0.0,0.24166667,0.44444445,0.23333335,0.7,0.5083333,1.2555556,1.2666668,3.8083332,3.955556,1.0,0.15555556,0.075,0.0,0.1,0.52500004,0.2888889,0.56666666,0.8555556,0.6333333,0.0,0.0,0.0,0.0,0.075,0.7222222,0.9916667,0.9333334,2.6666667,2.9000006,1.688889,1.1833334,1.0666666,1.3666666,1.3111111,1.1750001,0.9333334,0.6333334,0.35000002,0.26666665,2.4666667,2.7,1.0833334,0.7777779,0.2916667,0.4555556,0.88888896,1.7166667,2.6444445,3.0583334,3.3777778,3.1583335,2.8333335,2.511111,1.6083333,0.8111111,0.9666666,1.1777779,1.6333336,1.6444446,1.5444444,1.1250001,0.9444445,1.2583333,1.3444445,1.2833333,2.111111,2.8,3.1222227,3.822222,3.8750002,4.644445,4.366667,4.533333,4.358334,4.3333335,3.4111114,2.25,1.3111112,0.45833328,0.5,0.73333335,0.71111107,0.425,0.3888889,0.13333334,0.05,0.0,0.033333335,0.0,0.0,0.022222223,0.044444446,0.025,0.0,0.083333336,0.58888894,1.1583333,0.14444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22222222,0.525,1.3444444,1.6888889,1.3083334,0.74444443,0.95,0.87777776,0.62500006,0.3888889,0.41111112,0.225,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.25833336,0.4555556,2.1499999,3.4555557,13.124999,20.811111,9.922223,1.6416668,0.31111112,1.0500001,0.8777777,0.18333334,0.2666667,0.0,0.041666668,0.0,0.83333343,0.12222222,0.60833335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7833335,0.8666667,0.0,0.0,0.0,0.0,0.0,0.0,2.3888888,5.541667,0.0,0.0,2.0416667,8.7,3.4083333,0.0,0.0,15.600001,37.67778,12.125,4.022222,1.3083336,1.7333333,3.6083333,10.811111,9.833334,9.58889,4.8444443,0.775,1.6,2.4166667,1.4111111,1.2583332,0.8333333,0.31111112,0.5833334,0.34444445,1.1666667,3.7666667,3.7083335,2.1777778,2.7000003,1.0111113,0.45555556,0.16666667,0.11111113,0.13333334,0.22222222,0.20833334,0.2888889,0.14444445,0.0,0.0,0.0,0.022222223,0.19166666,0.5222223,1.1777778,1.8916669,1.8888888,2.125,3.4444444,4.733333,0.0,0.0,0.99999994,1.7,0.72499996,0.275,0.15,0.00625,0.14166667,0.42878792,0.9660714,1.3066666,3.7169647,5.013788,2.7384067,1.5613637,2.1937501,2.2416668,2.4916666,0.6625,1.1750001,0.39999998,0.25833336,0.25,1.075,2.9083333,3.0625,10.508333,2.4437501,0.7833333,1.1812501,1.55,1.6624999,1.8333335,2.5083334,3.0562499,3.175,1.6500001,2.2083335,0.74375004,0.14166668,0.10833334,0.24375,0.0,0.16250001,0.25833333,0.70625,0.8916667,0.51666665,0.59375,1.0083333,0.79375005,0.6833333,1.46875,1.8666668,1.75,1.4666667,1.9166669,1.18125,0.79999995,0.34375006,1.3416667,2.0875,1.9833335,1.9333334,1.825,0.98333335,0.26250002,0.3,0.3,0.36666667,0.39375,0.4666667,0.45,0.34375,0.47500002,1.1687499,2.2,2.6562498,2.9833333,2.9083333,4.1375003,4.6416664,4.2,4.3000007,5.10625,4.858333,5.1583333,5.01875,3.6583335,2.9374998,2.0000002,1.8062501,1.4916667,1.3812499,1.0166667,1.1666667,1.1500001,1.1666667,1.1,0.8833332,0.7749999,0.76666665,0.7416667,0.53125,0.41666672,0.15625001,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.05,0.05,0.00625,0.016666668,0.13750002,0.31666666,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1375,1.1249999,2.1125,2.125,1.425,0.46250004,0.28333336,0.4375,0.57500005,0.45625007,0.38333336,0.09166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.14166667,0.19375001,0.73333335,4.2625,7.641667,16.81875,14.116668,4.4166665,1.39375,1.8250002,1.5875001,0.68333334,0.3125,0.1,0.06666667,0.17500001,0.10833334,1.04375,0.2,0.72499996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2,1.2166667,0.8833333,0.0,0.0,0.0,0.0,0.325,0.96666664,1.5000001,0.0,0.0,0.025,0.17500001,0.31875002,0.016666668,0.0,9.925001,8.200001,3.8125002,1.3416667,0.15,0.0,0.01875,0.5833334,6.1062503,9.066668,4.225,2.29375,2.1583333,1.61875,1.0583334,0.85625005,1.5916667,1.8416668,1.7187501,1.2666667,0.7937499,0.39166668,2.00625,1.975,1.9187499,1.0,0.4666667,0.1125,0.116666675,0.6625,0.9,1.0937499,1.1833333,1.2833333,0.6125,0.19166666,0.0125,0.0,0.0,0.11666667,0.45,0.83125,1.0666668,1.1687499,2.075,3.21875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,1.4555557,2.7222223,1.4083334,0.7666667,0.7083334,1.4222223,2.775,3.2444448,2.3333335,2.0666666,1.1666666,0.22500001,0.43333334,0.28333333,0.25555554,0.083333336,0.17777778,0.0,0.0,0.0,0.0,0.0,0.3,2.5666666,3.225,1.6555556,2.1555555,3.4916668,5.1,3.6250002,3.677778,3.075,1.5777779,1.8111112,1.3499999,1.4111112,0.7166667,0.11111111,0.125,0.10000001,0.13333334,0.19166668,0.64444447,0.6750001,0.88888896,1.475,1.8777778,2.375,2.1222222,1.2777778,0.95000005,0.76666665,0.225,0.22222224,1.05,0.33333334,0.78888893,0.7833334,1.0888889,0.9583333,0.44444445,0.95833343,0.6333333,1.0916667,2.5,1.5333333,2.2416668,0.67777777,0.125,0.43333334,3.3000002,6.6444445,2.988889,5.1333337,8.3555565,6.3666663,5.455556,5.375,8.155557,11.211112,10.616667,14.422223,11.499999,11.944446,8.991666,5.7000003,4.241667,3.988889,3.6333337,3.4250002,2.6333334,2.1833334,1.8666667,1.5166668,0.94444454,0.5555556,0.19166668,0.044444446,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.116666675,0.10000001,0.0,0.0,0.0,0.0,0.0,0.6,2.1888888,2.3833332,1.5444443,0.93333334,0.44166666,0.06666667,0.20833334,0.22222224,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666665,0.42222223,0.4583333,2.6666665,4.825,10.211111,12.916666,6.766667,1.6,1.6583333,3.0666666,2.5083334,1.5333335,0.8083332,0.0,0.2888889,0.19166666,0.05555556,1.0833334,0.22222224,0.6999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.07500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.8888893,4.1222224,0.0,0.0,0.0,0.0,0.0,0.0,0.825,1.7000002,4.577778,3.1833332,1.1555556,1.1833333,0.0,0.041666668,0.2777778,2.4666667,1.2166668,0.888889,0.45000002,0.07777778,1.0833334,2.0111113,4.116667,3.6666665,1.9222223,0.85833335,0.6666667,1.7166668,1.988889,1.9833333,2.2333333,2.4666667,1.9583335,1.4555557,0.8833333,0.24444444,0.008333334,0.022222223,0.08888889,0.2,0.22222224,0.083333336,0.47777775,1.45,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.48888892,1.1,0.925,0.5777778,1.2833333,1.6,0.6583333,0.73333335,0.3916667,0.33333334,0.26666668,0.21666667,0.28888893,0.51666665,0.7111111,0.625,0.6333334,1.0333334,0.43333334,0.11111111,0.19166666,0.5,0.0,0.0,0.42499998,0.8555556,0.8111111,2.4583333,4.0333333,5.116667,5.9333334,4.4,3.5777779,2.8000002,3.4416666,4.155555,5.2000003,3.0444443,0.73333335,0.18888889,1.2222222,2.25,0.62222224,0.21666667,0.0,0.016666668,0.24444446,1.3416666,1.3111111,0.9666667,0.6000001,0.50000006,0.4666667,0.4666667,0.6833334,1.2555554,1.7555556,0.6,0.07777778,0.058333337,0.044444446,0.65000004,1.1666667,2.6249998,4.122222,5.077778,5.325,3.2444444,1.5416667,1.0444444,0.4166667,1.0000001,1.4333334,4.3583336,5.955556,6.2166667,7.088889,7.533333,8.1888895,7.144444,6.8000007,5.1000004,6.175,5.888889,5.75,5.5,4.7666664,3.9111114,3.888889,3.05,2.3555555,1.6333333,1.3777778,1.45,1.0,0.47777775,0.275,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.14166667,0.2777778,0.20000002,0.06666667,0.0,0.0,0.0,0.0,0.7111112,1.9416666,2.0555556,1.5833333,1.4555556,1.2111112,0.47500002,0.07777778,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333333,0.95555556,1.8416668,3.5444448,3.7583337,5.8666673,6.9916663,2.7333336,2.8222222,2.9666667,2.7444444,2.3666666,1.3333334,0.21666667,0.13333333,0.46666667,0.24166667,0.099999994,1.0666667,0.21111113,0.7749999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.19999999,0.67777777,0.058333337,0.0,0.70000005,0.37777779,0.05,0.0,0.16666667,0.083333336,0.033333335,0.0,0.0,0.25000003,2.0444446,3.775,3.8666666,4.011111,2.8500001,2.4333334,2.9916663,3.0333333,2.4083333,3.1111112,3.6333332,3.4499998,2.1333334,1.8500001,1.3444445,0.87500006,0.36666667,0.06666667,0.0,0.37777779,0.3416667,0.0,0.33333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.22499998,0.0375,0.10833333,0.0,0.008333334,0.056250002,0.16666667,0.45833337,0.39999998,0.2916667,0.1875,0.35000002,0.55,0.45833334,0.85,1.23125,1.4499999,0.85625005,0.9083333,0.25625,1.075,2.5875,2.9416666,4.35,3.66875,2.6666665,3.225,4.6833334,11.04375,10.85,10.233334,7.88125,4.825,4.2062507,4.0000005,2.7874997,1.3416667,0.45000002,0.475,0.9666667,0.89375,0.8166667,0.5375,0.09166667,0.8625001,0.6333333,0.33333334,0.25000003,0.34166667,1.075,1.0666666,0.6875,0.5250001,0.24166667,0.23750001,0.29166672,0.056250002,0.0,0.1875,0.28333333,0.55625,0.8083334,1.475,2.2,3.0166664,2.71875,1.3916667,0.46250004,0.15833333,0.016666668,0.41875,1.5166667,2.4437501,3.666667,4.05,4.4500003,5.625,6.1499996,5.9750004,5.5562496,5.2,4.99375,4.8250003,4.4437504,4.025,3.4499998,3.5125003,2.5583334,2.66875,2.7250004,2.2312503,1.0083334,0.32500005,0.23125002,0.058333337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.125,0.081250004,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.125,0.31875002,0.51666665,0.5437501,0.33333337,0.081250004,0.0,0.0,0.0,0.15,1.1187499,1.8666667,1.6312501,1.4166669,1.4500002,1.075,0.6666667,0.11875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,1.3416667,4.2374997,4.4750004,3.1687498,3.0583334,3.825,1.8166666,2.7333336,2.9187498,3.2083333,2.0749998,0.36666667,0.025,0.5083333,0.40833336,0.28750002,0.20833333,0.22499998,0.15833332,0.14375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.225,0.3375,0.15833335,0.050000004,0.09166667,0.016666668,0.0,0.43333334,0.26875,0.025,0.09375001,0.016666668,0.0,0.0,0.0,0.25625,0.19999999,0.025,1.1583334,3.7749999,3.7416668,3.3000002,3.8,4.2,4.25625,3.9416668,3.2437499,3.0,4.7833333,4.95625,4.0166664,3.6750002,2.8333333,2.59375,2.05,1.6833334,1.04375,0.65,0.575,0.31666666,0.45625,0.033333335,0.0,0.07777778,0.19166668,0.15555556,0.14166668,0.022222223,0.0,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.022222223,0.19166669,0.51111114,0.7333334,1.0416666,1.1555555,1.1416667,0.9111111,0.6583333,0.5888889,0.0,0.0,0.24444446,0.8583334,0.73333335,0.33333337,0.51111114,2.575,3.4444444,3.4555557,3.5416667,1.9,0.56666666,0.24444446,3.75,6.922222,7.122223,5.025,3.4,2.8666666,0.88888896,1.025,1.5999999,1.8666667,1.4166667,0.8555556,0.24166667,0.011111111,0.20000002,0.26666668,0.075,0.2777778,0.44444442,0.7583333,0.7111111,0.98333335,0.988889,1.2416668,0.7888889,0.2888889,0.0,0.0,0.19999999,0.6888889,1.0833333,1.2444444,1.0250001,0.9111111,0.88888884,1.0833333,1.8555555,2.25,1.2888889,1.2666667,0.25555557,0.07777778,0.108333334,0.23333335,0.125,0.21111113,0.28333333,0.73333335,1.0000001,1.7750001,2.544444,2.8500004,3.3111115,3.275,3.8111115,3.75,3.8,3.9222221,3.4416668,3.222222,2.75,2.5333333,1.8166667,0.5222222,0.27777776,0.06666667,0.15555556,0.28333333,0.71111107,0.9000001,0.5777778,0.13333334,0.1,0.15555556,0.225,0.22222221,0.108333334,0.011111111,0.016666668,0.07777778,0.022222223,0.0,0.022222223,0.050000004,0.0,0.0,0.0,0.0,0.025,0.11111111,0.008333334,0.0,0.0,0.011111111,0.083333336,0.3,0.67777777,1.0166667,0.92222226,0.425,0.033333335,0.0,0.0,0.0,0.425,1.3111112,1.3583333,1.2666668,1.3249999,1.2555556,0.78333336,0.2888889,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40000004,1.9333335,4.266667,3.822222,2.4916666,1.8333334,1.8666666,1.3444444,2.0222223,4.366667,3.3111107,0.5666666,0.23333333,0.14166667,0.70000005,1.011111,0.75,0.5888889,0.48333335,0.47777775,0.23333333,0.06666667,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11111112,0.71666664,0.5,0.775,1.3777778,2.188889,2.7083333,0.18888888,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.13333334,0.016666668,0.0,0.84999996,2.2777777,2.3333335,2.4583337,3.988889,6.2750006,5.922222,4.025,3.2666667,2.6222224,4.591667,4.2222223,4.3500004,4.2555556,4.5166664,4.1333337,3.7555556,3.025,2.5777779,2.5249999,2.0,1.4166666,1.35,0.9083333,0.45,0.40624997,0.36666667,0.43124998,0.15,0.0125,0.025,0.083333336,0.21875003,0.13333334,0.10625,0.29166666,0.36875004,0.17500001,0.0125,0.125,0.26666668,0.53124994,0.9666667,2.3687499,2.4583333,0.63125,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0375,0.0,0.19375,0.56666666,0.6,0.44999996,0.95000005,0.76250005,0.0,0.01875,0.25,0.5916667,0.64375,0.40833336,0.325,0.35,0.056250002,0.16666667,0.26666668,0.60625005,1.0416667,0.59375,0.09166667,0.13125001,0.058333334,0.118750006,0.116666675,0.36666667,0.60625005,0.5666667,0.4125,0.6916667,0.8062499,0.38333333,0.75,0.84374994,0.725,0.33125,0.9916667,1.8375,1.4083333,1.4624999,1.2,1.0666667,1.29375,1.8166667,1.43125,1.0166668,0.65625,0.016666668,0.075,0.11875,0.12500001,0.16250001,0.18333335,0.19999999,0.125,0.116666675,0.25000003,0.5583334,1.28125,1.5083334,1.7187501,2.0,2.09375,2.4666667,3.0500002,3.2624998,3.275,2.8375,2.325,1.225,0.625,0.35000002,0.2125,0.075,0.10625,0.26666665,0.35625,0.24166667,0.06875,0.050000004,0.016666668,0.01875,0.0,0.0625,0.083333336,0.075,0.04166667,0.06666667,0.112500004,0.033333335,0.00625,0.0,0.0125,0.108333334,0.23333335,0.112500004,0.0,0.0,0.0,0.08125,0.28333333,0.68125004,1.2,1.4416667,1.0187501,0.43333334,0.10625001,0.0,0.0125,0.108333334,0.44166666,0.89375,0.925,0.99375004,1.1083333,0.9062501,0.4083334,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46249998,3.291667,2.6749995,2.4000003,1.1812499,0.9333334,0.57500005,1.6416668,2.8583336,8.00625,2.6,0.075,0.033333335,0.45,1.9750001,2.3666668,1.75625,0.70000005,0.41875002,1.4916667,1.7062503,0.325,0.075,0.0,0.0,0.0,0.0,0.00625,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.74375004,1.9166667,3.4,4.5125,2.2416666,0.26875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.5833334,0.90624994,2.1166666,4.4875,5.7250004,4.55,3.775,3.0333335,2.3625002,2.9666662,3.3875003,3.8250003,4.34375,4.558334,4.0916667,4.225,3.5333333,3.15625,3.0500002,2.8249998,1.3083334,1.5888889,1.8111112,3.1166668,3.6666665,3.3416667,1.6222223,0.60833335,0.4,0.47777778,0.21666665,0.16666667,0.10000001,0.18888889,0.9833333,0.65555555,0.3,0.022222223,0.0,0.0,0.0,1.0583333,4.7666674,4.0416665,4.3333335,7.244445,3.825,2.3777778,0.2,0.5666667,1.0583334,0.39999998,0.008333334,0.0,0.0,0.0,0.0,0.1,0.08888889,0.35,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.07777778,0.275,0.37777776,0.9166666,1.7777779,1.725,0.8555556,0.9888889,0.6166667,0.53333336,0.90833336,0.6,1.2583333,1.8555555,2.7111113,3.725,3.8,3.3500001,3.0222225,1.9166669,1.8222222,1.5916667,0.9111111,0.7777778,0.9666667,0.4111111,0.6416667,1.5999999,1.4583334,0.6666667,0.35555553,0.35833335,0.39999998,0.26666668,0.21111113,0.39166668,0.47777778,0.5,0.4166667,0.65555555,0.7750001,1.2555554,1.1750001,1.0444443,1.1083333,1.288889,1.4444445,2.0166667,2.0555553,2.3416667,1.4777778,0.7583333,0.45555556,0.21111113,0.09166667,0.011111111,0.0,0.0,0.0,0.0,0.0,0.022222223,0.033333335,0.15,0.23333333,0.058333337,0.42222226,0.675,0.72222227,0.3222222,0.10000001,0.0,0.0,0.06666667,0.64166665,0.7222222,0.17777778,0.025,0.0,0.008333334,0.25555554,0.64166665,1.3,1.9833335,1.9111111,1.0777779,0.48333335,0.22222221,0.36666667,0.19999999,0.25,0.53333336,0.5555556,0.61666673,0.77777785,0.86666673,0.6555556,0.25833336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1333334,0.3416667,1.9666667,0.80833334,0.6777778,0.6500001,0.6888889,1.1583332,1.7222222,3.4,4.25,1.011111,0.10833334,0.022222223,1.6416665,2.788889,2.511111,1.1166666,0.3666667,0.7583333,4.0111113,2.0,0.8111112,0.45,0.0,0.0,0.0,0.0,0.10000001,0.41111112,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.73333335,0.65833336,0.46666667,0.10000001,0.36666667,0.10000001,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.175,0.21111111,0.0,0.0,0.008333334,0.0888889,0.011111111,0.033333335,0.66666675,1.5083333,2.7555559,3.8083334,4.2666664,3.4555554,2.5333335,2.011111,1.8166666,1.9222225,2.6333334,3.2222223,3.4444444,3.6166668,3.522222,2.9750001,2.4444444,1.5249999,0.0,0.0,0.19166666,1.00625,2.25,3.4875,1.9333334,1.3437501,1.2416667,1.1166667,1.325,1.0166668,0.78125006,0.49166664,0.23750001,0.17500001,0.18750001,0.10833334,0.15000002,0.050000004,0.0,0.3375,4.7583337,10.88125,13.275,17.533333,16.212502,7.1916666,2.4812498,2.2083335,4.73125,5.799999,3.8624997,0.43333334,0.0,0.0,0.058333337,0.2875,0.125,0.425,0.73333335,0.4,0.2,0.0,0.0,0.0,0.0,0.13333334,0.06666667,0.0,0.0,0.14375001,0.64166665,1.075,1.8833334,0.775,0.30833337,0.116666675,0.0125,0.16666667,0.40625003,1.1416667,1.6062502,2.075,3.15,4.20625,5.4,4.5062504,3.7916667,2.325,1.6916668,1.48125,1.8916669,2.0416667,1.2437501,1.0166667,1.16875,1.5166668,1.3187501,1.1166667,0.90000004,0.98125,1.2166667,0.575,0.34166664,0.38750002,0.30833334,0.40000004,0.65000004,0.96666676,0.975,1.2333332,1.15,1.1333333,1.03125,0.5916667,0.35000002,0.8000001,0.9833333,0.6999999,0.2916667,0.1625,0.09166667,0.025,0.0125,0.11666667,0.05,0.016666668,0.075,0.21666667,0.7375001,1.3,1.15,0.8000001,1.0500001,1.0437499,0.9416666,0.38125002,0.17500001,0.041666668,0.4,0.45000002,0.4,1.2500001,0.8499999,0.125,0.0,0.0,0.116666675,0.5125001,1.1916668,2.075,2.5583332,2.0562499,1.15,1.1333332,1.0937501,0.8666667,0.8125,0.6916667,0.53125,0.3916667,0.47500002,0.57500005,0.5500001,0.43125004,0.19166666,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7166667,0.29375,1.2916666,1.26875,1.475,1.9312501,2.275,6.09375,4.1583333,4.466666,3.0499997,1.2416667,0.325,0.5,2.69375,3.1166668,4.0583334,0.38750002,0.0,1.05625,3.266667,2.2125,1.1583332,0.475,0.0,0.0,0.0,0.0,0.80625,0.8416667,0.48125,0.42499998,0.40000004,0.09375001,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7166667,1.3874999,2.6833334,0.225,0.0,0.275,0.5,1.1999999,1.8125,1.8833334,1.3874999,0.025,0.31250003,0.48333332,0.19375,0.5416667,0.71666664,0.9625,0.21666665,0.17500001,0.008333334,0.00625,0.041666668,0.08333334,0.056250006,0.075,0.2875,0.9583334,0.9875001,0.35833335,0.03125,0.0,0.0,0.0,0.0,0.18125,2.2166667,4.0750003,3.65,2.7666667,2.5375,1.9916666,2.0124998,1.7416667,1.3750001,1.5416667,1.825,2.5124998,2.7916667,2.8187501,2.2666667,1.43125,0.0,0.0,0.0,0.0,0.0,0.041666668,0.055555556,0.008333334,0.044444446,0.12222222,0.28333333,0.70000005,0.76666677,0.9888889,0.82500005,0.40000004,0.275,0.22222224,0.13333334,0.06666667,0.0,0.0,0.0,1.3166667,4.7666664,6.555556,5.616667,4.0444446,2.6083333,1.9555557,4.5416665,8.333333,8.408333,5.4333334,3.6666667,1.3666668,0.23333332,0.625,1.1444445,0.85833347,1.1666665,1.3555555,1.7,3.2444444,2.325,0.13333334,0.041666668,0.011111111,0.08888889,0.0,0.0,0.0,0.0,0.5916667,0.16666667,0.025,0.011111111,0.0,0.0,0.011111111,0.09166667,0.18888888,0.5083333,0.85555565,0.9666667,1.55,2.9666667,3.4249997,3.3333335,2.425,1.888889,1.2083334,1.1333333,1.5555556,1.6166668,1.9111114,2.3500001,2.1111114,2.1666665,1.8777777,1.4777777,1.0916667,0.67777777,0.35000002,0.12222223,0.016666668,0.033333335,0.011111111,0.050000004,0.033333335,0.7916666,1.2666667,1.9916667,1.9666667,2.9416668,2.8111115,2.3777778,2.5,2.711111,2.4416666,1.7888889,1.4666667,0.7111111,0.17777777,0.19166668,0.67777777,1.0083333,1.1111112,1.5500001,1.8222222,1.6333333,0.8888889,0.8555556,1.2500001,0.6333333,0.3166667,0.11111112,0.18333332,0.36666667,0.5777778,0.46666664,0.42222223,1.1916667,0.65555555,0.09166667,0.022222223,0.06666667,0.225,0.92222226,1.85,2.8,3.0666668,2.1444447,1.5083334,2.411111,1.7,1.5583332,1.6000001,0.9083334,0.2888889,0.19166668,0.54444444,0.5444445,0.3666667,0.34444445,0.116666675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41666672,1.6777776,1.9083332,1.3333333,1.9250001,3.6555557,11.266667,6.966667,5.3888893,2.8333328,1.3444445,0.23333335,1.2111111,6.6250005,5.877778,2.6222222,0.20833333,0.0,0.5999999,3.4222221,2.5916665,1.6888889,0.18333334,0.0,0.0,0.0,0.0,1.1500001,1.2555556,1.7083334,2.0444446,1.4666667,0.90000004,0.31111112,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0333334,3.125,5.8888893,0.0,0.0,0.0,0.0,0.35555553,1.225,0.6222222,0.31666666,2.288889,0.9666667,1.4,0.6833334,1.5222222,3.2222223,4.225,1.2444444,0.25833336,0.11111111,0.26666668,0.41111115,0.16666669,0.20833334,0.3888889,0.20833334,0.17777778,0.20833334,0.3,0.29166666,0.13333334,0.033333335,0.0,0.0,0.0,0.6888889,3.025,4.1222224,2.8888888,2.4333334,2.3333335,2.4666667,2.6222222,2.1833334,1.6111112,1.3666667,1.4583335,1.7888889,2.0083334,1.9333334,1.2666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.24444446,0.14166668,0.2777778,0.78333336,1.0888889,0.78333336,0.2111111,0.033333335,0.025000002,0.0,0.0,0.0,0.0,0.0,0.5111111,2.5083332,4.0333333,3.9916666,4.5000005,5.5666666,6.3888893,5.816666,5.3111115,6.5444446,6.591667,2.6222224,1.4,2.0222223,1.9,1.7444446,2.4,1.4583334,2.6111112,9.508334,6.055556,1.25,0.044444446,0.0,0.15833335,0.65555555,0.21666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.06666667,0.2,0.6333333,1.6777778,2.5583334,3.0444446,3.3500001,2.9666667,2.75,2.4111114,2.1222224,1.9166666,1.5666667,2.0333333,1.7,1.6416669,1.4666667,1.2111112,1.1083332,1.0777779,1.175,1.0222223,0.89166677,0.7,0.54444444,0.44166666,0.22222224,0.08333334,0.62222224,0.85833335,1.1777778,2.5333335,2.266667,2.6777778,3.283333,4.288889,4.991667,4.6444445,3.6166666,2.6333337,2.2666667,2.7333336,3.3,2.6833334,2.0666666,1.7166666,1.5222222,1.2833333,1.5777776,1.1888889,0.98333335,0.6222223,0.30000004,0.12222224,0.06666667,0.17777778,0.044444446,0.17500003,0.84444445,0.9,0.17777778,0.13333334,0.14444445,0.31111112,0.9416666,1.7555556,2.558333,3.1111112,2.6250002,1.5777779,2.6916666,1.8666667,1.8333334,1.6833334,0.73333335,0.26666668,0.2,0.36666667,0.28888887,0.10000001,0.28333336,0.33333334,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333332,1.0666666,1.2333335,0.85555553,1.3416666,2.522222,7.1166663,3.4777777,2.2000003,0.40000004,0.31111112,0.8333333,3.211111,7.425,5.6222224,2.6,0.8333333,0.15555556,1.0916667,5.6111107,3.1000004,0.4666667,0.0,0.0,0.0,0.0,0.0,1.4333334,2.466667,3.733333,3.5777779,3.0555553,1.4166665,0.3555556,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777778,1.7333333,2.7222223,0.0,0.0,0.26666668,0.0,0.0,0.13333334,0.0,0.14166668,1.3444445,1.125,1.7666667,0.325,0.6666666,2.4444444,1.9833333,0.78888893,0.5416666,0.34444442,1.3416667,4.0111113,2.1111112,1.0166667,1.0777777,0.65000004,1.1555556,1.6916667,1.4,0.108333334,0.15555556,0.26666668,0.1,0.0,0.0,0.0,1.2083334,4.5666666,4.688889,3.6500003,3.1444445,2.6750002,2.5444446,2.4416666,2.188889,1.4222224,1.0333333,1.1,2.0,2.0777779,1.0416667,0.1375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06875,0.23333335,0.55625,0.5583333,0.96875,1.0833334,1.30625,0.9166666,0.2,0.0875,0.0,0.0,0.0,0.0,0.0,0.48333338,2.4875,6.250001,10.775001,10.183333,7.3312497,5.075,3.5187497,3.7333333,6.683334,7.4,5.633333,2.0375001,1.3666667,1.30625,0.85833335,0.38333336,0.49999997,1.25,1.41875,1.0833334,0.45625004,0.083333336,0.17500001,1.275,2.266667,3.1375003,1.6416667,0.4875,0.25,0.0125,0.0,0.0,0.01875,0.41666666,0.35625,0.083333336,0.025,0.18333334,0.51666665,1.1312499,1.9250002,3.0625,3.7333333,5.2999997,6.3416667,6.0437503,6.216667,5.8999996,5.45,6.025,5.4625,3.1583335,1.16875,0.5416667,0.4333334,0.31250003,0.2666667,0.25000003,0.15000002,0.05625,0.041666668,0.016666668,0.09375001,0.21666668,0.32500002,0.42499998,0.54375,1.3833333,2.0187502,4.0083337,6.0083337,7.45625,9.025001,9.618751,8.45,6.9375,6.008333,5.1166673,4.6062503,4.025,3.9437497,3.7500002,3.06875,2.4499998,2.0375001,1.4666667,0.95000005,0.5812501,0.37500006,0.27500004,0.125,0.25625002,0.5083333,0.6833334,1.1812499,0.76666665,0.17500001,0.1,0.33125004,0.7666667,1.1583334,1.8375,2.3666668,2.5874999,2.3666668,2.08125,2.5583334,1.8125001,1.9416666,1.7083333,0.71250004,0.30833337,0.25625002,0.275,0.1,0.13333334,0.26666668,0.41250002,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.25833333,0.36874998,0.0,0.43125,1.0666665,3.5937502,0.7916667,0.083333336,0.0,0.075,0.78124994,4.9666667,6.15625,3.9500005,3.975,2.6875,2.7666667,5.01875,3.6499999,2.5562499,0.14166667,0.0,0.0,0.0,0.0,0.0,1.7375,3.341667,5.4,5.075,2.5916667,0.79375005,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45624998,0.775,2.15625,7.7666674,3.5187497,0.15833333,0.24166666,0.38125,0.0,0.70000005,0.85,0.20000002,0.12499999,0.1375,0.275,0.49166667,0.75,1.2166667,1.0625001,0.2,0.0375,0.7666667,2.4,3.0562499,3.6333334,2.7812502,2.425,2.3312497,1.75,1.0875,0.18333334,0.0,0.10625001,0.20000002,0.0375,0.0,0.0,1.0583333,2.2250001,4.05,3.8916667,3.6375,3.0,2.61875,2.275,1.8083334,1.1624999,1.2583334,1.4437501,1.4333334,0.6625,0.033333335,0.06666667,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.20000002,0.2888889,0.64166665,0.7111111,2.475,2.1777778,1.5888888,0.48333338,0.06666667,0.0,0.0,0.0,0.0,0.0,0.25833336,2.1000001,5.441666,6.2888885,6.75,7.9555554,6.7583337,6.377778,4.6555552,5.1333337,6.055556,6.541667,4.611111,4.075,3.5333333,2.6111112,1.0500001,0.6111111,2.2166667,3.3222225,1.5083333,0.44444445,0.055555556,0.44166666,0.7111111,0.40833333,0.62222224,0.55,0.3333333,0.05,0.0,0.0,0.0,0.08888889,0.0,0.0,0.45,0.99999994,1.3555557,1.7833335,1.9111111,2.3000002,4.1555552,7.3999996,9.733333,10.808334,7.5222225,5.455555,4.4166665,3.8555555,3.4750001,1.9555554,1.25,0.51111114,0.37777776,0.19166668,0.13333334,0.083333336,0.055555556,0.0,0.0,0.0,0.0,0.0,0.025,0.055555556,0.20833334,0.18888889,0.40000004,2.3333333,4.5222225,7.116667,8.055555,9.025,9.411112,8.791666,7.677778,7.3,6.125,4.833334,3.8333335,2.977778,2.3833332,1.577778,0.98333335,0.5888889,0.40000004,0.21666668,0.29999998,0.45833337,0.7777778,1.3166667,1.5555556,1.5333333,0.9416667,0.6111111,0.60833335,0.72222227,1.1666667,1.6777779,2.2444444,2.9416668,3.3555555,3.1416671,2.688889,2.2833335,1.8333333,1.9999999,1.2777778,0.7111111,0.4416667,0.43333334,0.21666667,0.033333335,0.19166668,0.33333334,0.3888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2416667,0.6666667,1.8083334,0.0,0.0,0.0,0.22222221,1.0999999,4.9444447,4.0166664,3.7111113,4.5111113,5.691667,7.866667,8.191668,5.3,5.891667,0.87777776,0.18333334,0.0,0.0,0.0,0.0,3.3166666,5.611111,6.783334,2.8333335,1.1666666,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.15,2.1333332,0.23333335,0.08888889,0.4888889,0.55,0.0,3.4,2.911111,0.39166668,0.17777777,0.016666668,0.17777777,0.5777778,2.2083335,0.8,0.15,0.0,0.0,0.0,1.3777778,3.2499998,4.2777777,4.4333334,2.8222222,2.0166667,1.2777778,1.3833334,1.6555556,0.022222223,0.0,0.0,0.05,0.011111111,0.0,0.0,0.044444446,1.8166667,3.0888891,2.5000002,2.1444445,1.2249999,0.7555556,1.0777779,0.6833334,1.2555556,1.2416668,1.1000001,0.29166666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.13125001,0.175,0.25,0.7416667,0.52500004,0.85,0.64166665,0.26250002,0.0,0.0,0.0,0.0,0.0,0.008333334,0.63125,1.5333333,2.6437497,5.375001,10.418751,13.258334,9.599999,5.8499994,3.6250005,2.99375,3.566667,4.9875,7.9083333,9.033333,6.6125,6.791667,4.163393,1.9825758,1.9616668,1.1250001,0.9833333,0.70624995,0.31666666,0.0,0.0,0.0375,0.025,0.0,0.0,0.0,0.0,0.0,0.125,0.175,0.20625001,0.29166666,0.46666667,0.70625,0.52500004,0.58750004,0.95000005,2.0125,4.425,6.40625,5.8833337,6.0916667,4.85625,3.891667,3.1625,2.0083334,1.5312501,0.4416666,0.36666667,0.21875,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.14166667,0.16874999,0.15000002,0.0375,0.6750001,1.1250001,2.3624997,4.0499997,7.66875,9.566667,9.793751,9.858334,9.616667,8.793751,7.025,5.8000007,4.6833334,3.49375,2.2333336,1.5312499,1.2333332,1.1333334,1.3812501,1.8583331,1.9625,2.6583335,2.375,2.0416667,1.9999999,2.11875,1.9083335,2.09375,2.1916666,2.40625,2.4,2.641667,2.7625003,2.6333332,2.54375,1.9583335,1.78125,1.4583335,1.0250001,0.75,0.5333333,0.18750001,0.050000004,0.09375,0.175,0.19375,0.1,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.10625,1.1500001,1.1750001,0.7916667,2.125,1.11875,1.0083333,2.3937502,3.958334,2.5874999,1.1416667,3.2,4.50625,7.3750005,7.975001,10.183332,10.374999,2.3999999,0.125,0.13333334,0.0,0.0,1.2,4.40625,5.958334,3.7375002,0.9749999,0.175,0.0,0.025,0.7937499,0.40833333,0.0,0.0,0.0,0.01875,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.5833333,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.66875005,1.425,0.28125,0.15,0.15,0.28125,0.0,0.0,0.0,0.0,0.0,0.06666667,0.8375,1.075,3.35625,1.775,0.8062499,0.39166668,3.7625,6.083334,3.7000003,0.16250001,0.025,0.043750003,0.0,0.0,0.0,0.008333334,0.2125,1.4666667,1.4,0.35000002,0.0375,0.0,0.041666668,0.35625005,1.0333334,1.1437502,1.2500002,1.1750001,1.1083333,0.15555556,0.055555556,0.23333333,0.25555557,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12222222,0.041666668,0.055555556,0.20833336,0.12222222,0.055555556,0.0,0.0,0.0,0.0,0.26666668,0.8666667,3.0083334,7.888889,13.422222,12.991667,5.255556,2.8666663,2.4666667,1.4916667,2.6555557,4.677778,5.9333334,3.2333336,2.3500001,3.088889,4.34697,2.5333333,0.6888889,0.6750001,0.9111111,1.1583332,0.17777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.2,0.33333334,0.40000004,0.775,1.2444445,1.2499999,1.5222222,1.9333334,2.5416665,2.211111,1.1500001,0.91111124,0.725,0.33333334,0.13333334,0.083333336,0.044444446,0.008333334,0.0,0.016666668,0.0,0.044444446,0.0,0.0,0.016666668,0.044444446,0.0,0.0,0.05,0.34444445,0.65555555,1.4583334,2.2333333,4.7333336,7.3444443,8.258333,8.155556,7.177778,5.9333334,4.733333,3.775,3.2555554,2.891667,2.411111,2.3083334,2.3777778,2.6888893,3.291667,3.477778,4.1,5.622222,2.1916668,2.0111113,2.3999999,3.0416665,3.2222223,2.591667,2.877778,2.016667,1.611111,1.2444446,1.0833334,1.4111112,1.8666666,1.8222222,1.475,1.111111,0.7416667,0.4555556,0.26666665,0.075,0.24444444,0.16666667,0.044444446,0.016666668,0.055555556,0.033333335,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.025,2.2888892,2.775,7.9000006,10.044445,7.3416667,4.388889,6.8083334,5.6,0.98333335,0.22222222,2.0444446,6.358333,4.7555556,1.7416667,3.7999997,6.6083336,2.1444442,1.3416665,0.8888889,0.0,0.1,2.3777778,4.3416667,5.0444446,1.5249999,0.6222222,0.14444445,0.4416667,0.2,0.16666667,0.0,0.0,0.6444444,1.6888889,2.0916667,1.1333333,0.25833336,0.75555557,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.14444445,0.0,0.0,0.5222222,0.625,0.0,0.16666667,0.26666665,0.3333333,1.0555556,1.525,0.7777778,0.4888889,1.0749999,2.1777778,0.0,0.0,0.0,0.0,0.0,0.033333335,0.2,0.13333334,0.011111111,0.7583334,0.9,2.875,3.6111112,3.0555558,1.0,0.48888886,0.7583333,1.1,1.4499999,0.24444443,0.0,0.0,0.0,0.3333333,1.0555556,0.55833334,0.06666667,0.10000001,0.3916667,0.8222223,1.3833332,1.7666668,1.35,0.3375,0.40000004,0.15833333,0.43125,0.69166666,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.18124999,0.29999998,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.375,1.2916666,1.675,5.0937505,8.149999,7.1687503,4.3583336,3.2312498,2.3333335,1.5250001,1.58125,1.2083334,2.23125,5.283334,8.5375,9.316667,4.766667,1.4562501,1.6000001,2.5249999,2.8,1.9125001,0.925,0.26875,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0625,0.108333334,0.0625,0.050000004,0.083333336,0.075,0.1,0.10625,0.033333335,0.025,0.041666668,0.116666675,0.14375001,0.2,0.24375,0.325,0.36875004,0.5,0.4916667,0.38125002,0.125,0.025,0.0,0.0,0.0,0.0,0.0,0.075,0.16875003,0.375,0.81875,1.6750001,2.03125,2.1166666,2.1166668,2.5437498,2.0583336,1.4625001,1.4833333,1.90625,2.3416667,2.3250003,2.325,2.2833333,1.8312501,1.5166667,1.8000001,1.5916666,1.1875,1.3083333,1.5749999,1.63125,1.1583333,0.69375,0.79166675,0.80625,0.8000001,0.85833335,1.2624999,1.9333333,2.0249999,1.75,1.3562499,1.1,1.1812501,0.78333336,0.3416667,0.16250001,0.05,0.043750003,0.075,0.11250001,0.108333334,0.10000001,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,0.275,0.0,0.008333334,0.050000004,0.0,0.77500004,1.225,4.9812503,8.516666,11.31875,14.625,12.291668,9.06875,9.150001,5.6062503,2.0833333,0.15,0.5916667,8.05,9.262501,2.8500004,0.95000005,2.4500003,1.4499998,0.65833336,1.0250001,1.1083333,0.975,1.16875,2.8166666,3.0187502,2.125,0.38125002,0.80833334,1.4833333,1.09375,0.083333336,0.0,0.0,0.43750003,1.7083333,2.0083334,2.33125,1.075,0.08125,1.3833333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5666667,0.8833333,0.0,0.0,0.85625005,1.5083333,2.7125,1.1,0.69375,0.45833334,1.1,3.3250003,2.1833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.98749995,3.7000003,0.475,0.325,2.8000002,5.041667,3.575,3.9625,1.8916667,0.63125,0.17500001,0.1875,0.0,0.0,0.0,0.0,0.03125,0.38333333,1.1374999,1.3416667,1.3666668,2.4125,3.1083336,3.2937503,2.6666665,0.47500005,0.0,0.13333334,0.31111112,0.6,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.5222222,0.48333335,0.16666667,0.14166667,0.055555556,0.033333335,0.4,0.67777777,3.141667,5.5222216,6.4333334,4.5555553,2.5555553,0.89166665,0.5,4.0416665,16.033333,26.258331,18.811111,7.088889,3.041667,1.2444445,2.3833334,3.4222221,2.9166667,3.8777778,3.5000002,2.2111113,0.53333336,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.22222221,0.2,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.033333335,0.07500001,0.055555556,0.058333337,0.1,0.075,0.22222222,0.51666665,0.21111111,0.34444442,0.0,0.0,0.0,0.033333335,0.15,1.1444445,1.5333334,2.4083333,1.9888889,2.358333,2.5333335,3.1166668,3.6888888,3.4666667,2.822222,2.0,1.3083334,0.6111111,0.20833334,0.16666667,0.17500001,0.07777777,0.055555556,0.05,0.16666667,0.65833336,0.7222222,0.79166675,1.5111111,2.1888888,2.4249997,2.0555556,1.8000002,1.8333333,2.0500002,2.0333333,1.075,0.36666667,0.13333334,0.083333336,0.15555556,0.29166666,0.26666668,0.15,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.13333334,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.083333336,0.0,0.0,0.008333334,0.26666668,4.5583334,6.911112,10.416666,11.922221,16.916666,13.622223,11.599999,11.958334,6.9111114,0.85833335,0.6777778,0.0,3.3333337,9.444445,4.0166664,1.3333335,1.05,6.444444,1.8666668,0.13333334,0.20833334,1.2,1.9666666,0.91666675,1.811111,1.4666667,0.45555556,1.0916667,2.6000001,2.4,0.09166667,0.0,0.083333336,0.08888889,0.68333334,0.2777778,0.26666668,0.0,0.15555556,1.15,1.4666668,0.16666667,0.28888887,0.0,0.0,0.0,0.0,0.0,0.55,2.988889,2.5583334,1.3111111,0.34444445,0.0,0.0,0.51666665,1.9000001,3.2416668,0.65555555,0.7583333,1.2555555,1.8111112,3.9166667,7.577778,4.9750004,0.0,0.0,0.0,0.0,0.0,0.0,0.23333332,1.0222223,2.8999999,2.0,5.025,11.244444,10.0,11.133333,10.855555,4.841667,2.6333334,0.0,0.033333335,0.06666667,0.0,0.0,0.008333334,0.044444446,0.56666666,1.7000003,1.8777778,2.3500001,2.588889,2.775,2.1777778,1.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.66666675,1.95,2.733333,2.9166665,3.811111,2.8833332,1.9777777,1.6888889,1.6166667,2.5444446,3.1000001,6.133333,8.716666,6.9888887,5.158333,6.677778,7.0222225,1.0166668,0.1,0.3,0.22222222,1.4749999,3.3222225,2.7,2.975,2.1444445,1.9500002,5.622222,17.875,17.47778,10.055555,3.7333333,1.2333333,2.075,1.9333334,3.1749997,3.2888892,4.025,4.233333,2.3888888,0.68333334,0.0,0.0,0.011111111,0.1,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.36666664,0.625,0.7111111,0.6333333,0.3555556,0.23333335,0.13333333,0.05555556,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12222222,0.055555556,0.0,0.0,0.0,0.0,0.0,0.033333335,0.0888889,0.16666669,0.32222223,0.65,1.1333333,1.5166667,1.8444445,2.0166667,2.4,2.4888887,2.2166665,1.9000001,1.4416667,1.0222223,0.40833336,0.1777778,0.06666667,0.2,0.8666667,1.025,0.6666667,1.5916667,2.6444445,2.4,2.1416664,2.5222223,2.516667,2.0555556,1.7500001,1.0111111,0.5833333,0.77777773,0.46666667,0.38333336,0.53333336,0.4583334,0.18888889,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.31111115,0.15555556,0.7833333,1.2555556,0.48333332,0.46666664,0.0,0.0,0.0,0.008333334,0.06666667,0.058333337,0.19999999,0.175,0.0,0.0,0.23333335,2.3222222,10.833334,10.666667,10.933333,9.611112,15.341665,14.555555,13.777778,5.8083334,1.0555556,0.28333336,0.83333343,0.6,5.755556,6.7666664,1.7416666,0.7,2.4666667,8.588889,1.0583334,0.22222222,0.3166667,1.0888889,1.2777778,3.1166668,2.111111,0.75000006,0.8000001,3.2083335,3.4888887,0.17777778,0.025,0.14444445,0.6833334,0.6,0.9333333,3.0333333,2.8777778,0.3,2.8222222,4.6583333,1.611111,0.6166666,0.9444444,0.34166667,0.0,0.0,0.0,0.0,0.25833333,1.7777778,1.3833334,0.6777778,0.15555556,0.0,0.0,0.0,0.011111111,0.5416666,0.14444445,0.55,0.8444444,0.6666667,0.475,1.2222223,2.1666667,1.5555556,0.55,0.0,0.0,0.0,0.0,0.0,0.0,1.4000001,1.6777779,1.575,4.577778,6.9,7.1833334,5.3222227,6.125,3.4666667,1.8333334,0.8,0.13333334,0.0,0.0,0.0,0.0,0.27500004,1.2111112,1.6888889,0.9250001,0.93333334,1.4250001,1.9000001,1.9583333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2625,2.4333334,5.3812504,8.566667,16.34375,15.091667,8.700001,4.3125,3.6833334,4.2312503,4.541667,7.3687496,8.133333,5.9874997,5.3083334,7.3500004,8.724999,5.4416666,1.5812501,0.20833333,0.03125,0.033333335,0.75833327,3.0749998,5.216666,6.36875,2.8,1.91875,3.7583332,5.116667,5.0375004,5.7250004,2.91875,0.73333335,0.41875,1.2583334,2.2937503,3.4916666,3.5833333,2.2375,0.8583333,0.175,0.95000005,1.3187501,0.97499996,0.041666668,0.0,0.025,0.1875,0.22500001,0.0,0.0,0.0,0.0,0.016666668,0.0875,0.16666667,0.3,0.375,0.41875002,0.35833338,0.25000003,0.16250001,0.083333336,0.025,0.016666668,0.00625,0.0,0.0,0.0,0.0,0.0,0.008333334,0.081250004,0.26666668,0.3875,0.4,0.43333334,0.47500002,0.45,0.2875,0.34166664,0.12500001,0.06666667,0.1,0.112500004,0.07500001,0.081250004,0.008333334,0.13125,0.13333334,0.17500001,0.13333333,0.18333334,0.21875,0.29999998,0.21875,0.25000003,0.4375,0.5583334,0.8833333,1.4562501,1.7583334,2.2875001,2.6,2.5249999,2.3,2.4416666,2.675,1.8916665,1.3937501,0.9166666,0.6125001,0.6083334,1.06875,1.3083334,0.9416667,0.96250004,0.8,0.4124999,0.11666668,0.03125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12500001,0.20833334,0.10833333,2.3937502,2.3416667,1.2124999,0.5166666,0.0125,0.075,0.116666675,0.47500002,0.81666666,1.2687501,1.125,0.89375,0.47500002,1.8916668,4.45625,9.458333,11.062501,12.258334,9.06875,7.0249996,10.293751,9.958334,4.4500003,1.15,0.4583333,0.26875,0.35833332,0.50625,3.9333334,4.483333,1.7937502,0.23333333,4.9249997,3.0083334,0.2125,0.9083333,0.75000006,2.266667,1.9666667,4.46875,1.7333336,0.81250006,3.8833332,3.4125004,0.22500001,0.083333336,0.43750006,0.7583334,2.6812499,2.091667,6.48125,12.058332,12.133333,8.66875,11.608334,15.037499,9.466667,2.48125,0.25833336,0.0375,0.0,0.0,0.0,0.0,0.0,1.5000001,0.6875,0.55,0.93333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1333333,1.9250001,1.6083333,1.78125,0.008333334,0.008333334,0.0,0.0,0.0,0.25833333,3.3000002,8.375,10.84375,7.316667,6.1083336,10.275,7.7833333,3.13125,1.2583333,0.55625004,0.17500001,0.15833335,0.51875,0.5416667,0.06875,0.0,0.10625001,0.52500004,1.75,1.6750002,2.4583335,2.55,3.0583334,3.0687501,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5222222,1.55,3.588889,3.6222224,2.4,1.1111112,0.25000003,0.23333332,0.48333338,0.34444445,0.7000001,0.7111112,0.5,0.425,0.62222224,1.4333333,0.90000004,0.09166667,0.0,0.0,0.0,0.1,0.25833333,0.5222223,0.45833337,0.05555556,0.3222222,2.9416666,6.211112,3.3416667,1.2222222,0.14166667,0.17777778,0.5333333,1.4000001,2.777778,5.741667,5.6000004,2.891667,1.977778,1.8833334,0.7666667,0.3333333,0.016666668,0.59999996,0.3,0.0,0.9333334,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15833332,0.39999998,0.55833334,0.57777774,0.5777778,0.80833334,0.5666667,0.42500007,0.54444444,0.19166669,0.14444447,0.10000001,0.075,0.044444446,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.10000001,0.26666668,0.32222223,0.93333334,1.8555555,3.1111114,3.1333334,3.266667,5.466666,6.4666667,6.0416665,5.2444444,3.1666667,2.108333,1.9777778,1.1916668,1.2666668,1.2166667,2.2555556,2.525,2.2,1.8444445,0.7250001,0.2888889,0.09166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.116666675,0.022222223,0.76666665,2.5083337,1.7222222,0.86666673,0.06666667,0.041666668,0.39999998,0.51111114,1.625,2.1444445,2.6833334,2.2666667,1.3083333,4.1444445,6.8,9.608335,10.122223,10.5666685,8.6,6.2500005,6.577778,10.408334,5.388889,1.4777777,0.33333337,0.2777778,0.35000002,0.14444445,0.425,2.8888888,3.2333336,1.2833334,0.31111112,4.391667,0.5777778,0.45833334,0.73333335,1.6416667,3.7888885,3.2000003,6.8,2.0333333,1.3333334,2.2555556,2.216667,0.122222215,0.3888889,0.93333346,1.9111114,3.95,9.833333,20.066666,27.611113,27.877777,26.391666,13.322223,5.7333336,3.1222224,0.65,0.23333335,0.008333334,0.0,0.0,0.0,0.0,0.15,1.5444446,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.37777779,0.8416667,0.4,0.0,0.0,7.4416666,12.955557,10.491667,5.133333,6.5222225,5.916667,4.6222224,2.7000003,2.1333332,3.766667,2.7888887,1.1666666,0.85,0.49999997,0.06666667,0.0,0.008333334,0.2888889,1.3222222,3.0500002,3.711111,3.866667,3.9222224,4.291667,0.0,0.25,0.59999996,0.58124995,1.1333332,1.01875,0.375,0.10000001,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.14375,0.14166667,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.39125,1.0583333,1.4687501,0.5833334,0.29375005,0.32500002,0.3375,0.5,0.6833334,1.925,3.3166666,5.5,4.866667,6.01875,7.3500004,6.0166664,1.8125,1.2583334,6.0125,5.4666667,4.7375,1.0333333,0.1875,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.083333336,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10625001,0.15,0.44375,1.025,3.4187503,5.2999997,8.258333,10.93125,12.008334,11.049999,7.366667,5.8312497,6.0666666,4.1250005,4.0,4.3083334,3.1750002,3.2,2.725,2.7916667,2.3062496,1.3000001,0.52500004,0.15625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.18333335,0.087500006,0.94166666,2.15,1.53125,0.7833333,0.25624996,0.025000002,0.54999995,1.4,2.4500003,2.99375,4.066667,3.4124997,1.4333333,3.18125,7.891667,9.408333,9.35625,9.691667,7.9437494,6.9833345,8.668751,15.375001,12.225,2.7583334,0.56666666,0.15625,0.19166668,0.25625,0.15,0.0625,0.09166667,0.041666668,0.325,0.20833333,2.9125004,0.22500001,0.5125,0.95000005,6.375,5.6333337,2.9499996,2.9,2.8583333,1.8562498,0.7833333,0.31874996,0.45833337,0.91666675,1.2312502,2.7916667,6.0562496,22.841667,36.993748,41.416668,37.025,24.631248,11.783333,2.9625,0.18333334,0.10625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.8333333,3.44375,2.3916667,0.30624998,0.42499998,3.1375,9.95,6.8562503,0.5,3.7166665,5.09375,5.775,6.7187505,7.9750004,5.0687504,4.1000004,3.166667,3.725,2.2749999,0.225,0.0,0.0,0.025000002,0.27500004,2.475,5.183334,6.51875,6.2833333,6.5687504,0.050000004,0.0,0.22222222,0.51666665,0.73333335,0.5083333,0.24444446,0.20000002,0.07777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.17777778,0.375,1.3888888,1.9749999,1.7111113,1.6777778,1.1333333,1.5777777,2.4333334,2.2222223,3.0500002,4.3222227,5.4,5.0,3.6777778,1.7083335,3.888889,7.8416667,3.5666666,1.1500001,0.17777778,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.30833334,0.6111111,1.5,3.7444446,8.958334,12.677778,13.511111,11.633334,8.677778,6.4,5.444445,5.383333,4.688889,3.5777779,2.8666663,3.0666666,2.4333334,2.777778,3.6416667,2.111111,0.92499995,0.3111111,0.06666667,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.10000001,0.33333334,2.2444444,1.7222222,0.9,0.27777776,0.075,0.5222223,1.8416667,3.7888892,4.233333,5.1,4.888889,2.0416667,1.5333333,5.8583336,7.7777786,7.911112,8.691667,7.6555557,6.7833333,9.577778,15.108335,12.300001,4.7166667,0.2888889,0.5666667,0.47500002,0.13333336,0.108333334,0.0,0.0,0.0,0.0,0.0,0.0,1.1833334,0.1,0.29166666,1.2666667,3.3500004,1.7333333,0.93333334,1.0,1.9,0.7916667,0.51111114,0.55833334,1.0777777,1.0333334,2.1583333,3.5666666,13.333335,36.488888,45.9,44.77778,35.344448,19.141666,5.688889,0.92499995,0.0,0.0,0.0,0.0,0.0,0.0,0.13333333,0.4222222,0.033333335,1.1111112,2.7833335,1.7333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.19999999,1.0333334,2.8416667,2.9222224,4.8833337,2.6777778,4.6000004,4.0333333,5.1555552,5.408334,6.122222,5.641667,2.3111112,1.4444444,1.625,0.13333334,0.0,0.0,0.0,0.0,0.0,0.47500002,3.0555558,5.7333336,7.4777784,8.783334,0.0,0.0,0.0,0.0,0.0,0.0125,0.05,0.05,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.1,0.175,0.18333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1125,0.8666667,2.9250002,5.166667,3.6,3.0249999,1.6666666,1.1500001,1.2500001,1.4812499,1.9583334,2.3083334,2.0625,1.75,0.425,0.0,0.00625,0.125,0.20000002,0.083333336,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.13333334,0.125,1.1687499,1.7,4.1000004,5.716667,7.6687503,8.666668,6.250001,4.48125,4.3583336,5.1000004,7.058333,6.0499997,3.6583338,5.333333,6.70625,4.4333334,3.5125005,2.8249998,1.7437501,0.7666667,0.39999998,0.175,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.087500006,0.025,0.83125,1.3000001,0.7333333,0.36875004,0.016666668,0.66875005,2.0833335,4.6625004,5.6916666,6.491667,5.906251,3.575,1.525,3.7833333,5.7,6.1416674,6.6916666,6.256251,5.4750004,9.05625,12.450001,9.631249,3.8333335,0.5875,0.083333336,0.85833335,1.9687501,1.4000001,0.49375004,0.033333335,0.0,0.0,0.0,0.0,0.0,0.06875,0.058333337,0.5500001,1.3083334,0.68125004,0.20833334,0.525,1.4750001,1.0916666,0.99375004,0.525,3.14375,7.333333,5.6416664,7.90625,9.799999,24.500002,34.71667,37.262497,36.633335,27.933334,15.54375,3.9,1.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.16250001,10.691666,2.3625,5.35,8.69375,3.991667,0.7583333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10000001,0.3,0.3416667,0.44375002,0.57500005,2.15625,5.1,5.6166673,4.875,4.075,2.3562498,1.2916667,2.8874998,4.1083336,4.825,2.39375,0.18333334,0.0,0.0,0.0,0.0,0.0,0.0125,0.8333334,3.5312502,6.7000003,9.35,0.0,0.0,0.0,0.016666668,0.08888889,0.15,0.06666667,0.016666668,0.0,0.022222223,0.075,0.011111111,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19166666,1.011111,1.3888888,0.8833333,0.39999998,0.0,0.0,0.0,0.022222223,0.11111112,0.275,0.24444444,0.23333335,0.7111111,2.3000002,5.6,12.941667,23.266666,8.055556,3.7000003,2.6666665,2.2916667,1.3333335,1.1,0.5777778,0.4888889,0.8416667,0.32222223,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.57777774,4.3111115,11.683332,3.5111113,0.51666665,0.0,0.0,0.31111112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7000001,0.7888888,0.53333336,0.5083333,1.0111111,1.8416667,2.655556,4.1083336,4.577778,3.3333335,3.275,4.6000004,7.033334,8.6,5.016667,7.9,10.033334,7.425,2.7,1.1083332,0.6333333,0.79999995,0.44444448,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.9,0.5555555,0.34444442,0.12500001,0.17777778,2.2833333,4.955555,7.016666,7.877778,7.4666667,6.4833336,1.3777777,3.0750003,3.5222225,3.7083335,4.6222224,4.822222,4.3333335,7.033334,9.825001,6.755556,2.741667,0.18888889,0.033333335,2.3222222,6.255555,5.333333,1.588889,0.29166666,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.10000001,0.20000002,0.18888889,0.1,0.32222223,1.1666666,2.4416666,2.688889,3.7083335,1.7555555,12.908334,18.444443,19.255556,20.300001,18.344444,25.016666,24.466667,21.616663,17.3,13.333334,9.883333,4.0777783,0.89166665,0.0,0.0,0.0,0.0,0.0,0.0,0.85833335,12.355556,5.2083335,5.077778,1.8000001,2.9888892,3.7111113,0.8833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.058333337,1.3666669,2.3999996,1.2583333,0.2,0.14166668,0.36666667,1.2666667,5.0555553,5.1222224,2.4833336,0.5888889,0.0,0.0,0.0,0.0,0.0,0.0,0.25555557,2.8166668,5.8111115,8.616667,2.14375,0.73333335,0.4166667,0.1,0.041666668,0.05625,0.025,0.03125,0.18333334,0.3166667,0.14375001,0.075,0.06250001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.20000002,0.7333334,1.7624999,1.7166666,1.0749999,0.49999997,0.125,0.0,0.0,0.32500002,1.2666667,1.84375,2.875,6.7375,14.333333,15.4125,7.95,3.633333,1.4750001,1.0083333,1.5375,1.7,1.1999999,1.4000001,1.1416667,0.69375,0.10000001,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.85,6.06875,10.225,3.1875,1.9083333,10.825001,9.191667,1.3124999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10000001,0.225,0.47500005,1.04375,2.4333332,3.59375,4.008333,4.2833333,7.4937506,9.658333,15.85,16.133333,12.54375,6.8583336,3.233333,2.63125,2.1083333,1.5250001,0.75,0.18125,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.22499998,0.116666675,0.033333335,0.0,1.7249999,4.1562505,8.658333,8.8,9.758334,9.3,4.375,2.3333335,2.71875,1.8083332,2.175,2.7333333,3.4166667,5.675,8.275,5.4875,2.3083334,0.33125,0.0,1.04375,2.6583335,2.1750002,0.4625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23750004,0.45000005,0.33125,0.31666666,0.31666666,0.96875006,1.9166666,6.0812497,4.1833334,15.875001,26.900002,35.216667,22.9125,20.391668,19.331251,10.008333,9.3375,5.8166666,3.5583334,3.46875,1.9833332,0.41250002,0.0,0.0,0.0,0.0,0.18333334,0.975,4.45625,17.858334,7.75,3.525,1.4625,1.8500001,3.9,1.6312501,0.175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44166666,2.9687498,7.1166673,6.1666665,2.3687503,1.3333334,3.675,3.0666668,4.0625,5.05,4.3,1.625,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.54375005,1.9000001,4.4937506,2.55,3.6555557,4.3555555,2.5666668,1.1666667,0.52500004,0.23333332,0.06666667,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.21111111,0.6,0.88888884,1.0583334,1.4666667,0.8500001,0.36666667,0.22222224,0.016666668,0.0,0.31666666,0.14444445,0.033333335,0.2777778,0.5583334,0.06666667,0.0,0.0,0.0,0.0,0.15555556,0.39999998,0.90000004,0.6777778,0.3416667,0.05555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1583333,1.5888889,0.55,0.0,0.0,0.2888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38333336,1.4111111,0.6166666,0.033333335,0.0,0.15555555,0.116666675,0.0,0.0,0.0,0.14444444,0.15833333,0.98888886,0.19166666,0.044444446,0.0,0.975,0.3,0.1,0.0,0.0,0.0,0.0,0.0,0.3111111,0.45000002,1.6777778,1.7333333,0.6666667,1.0666666,3.1444445,6.2333336,10.641667,15.211111,21.425,24.633335,17.708332,5.6000004,2.088889,0.94166666,0.39999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.5666667,4.4222217,6.975,8.633332,7.816667,6.788889,7.8777776,2.2083333,2.522222,1.4250001,1.1,1.4249998,1.8444445,4.4888887,6.341667,4.2666664,1.8166666,0.17777778,0.0,0.75555557,1.6666666,0.94444454,0.33333334,0.125,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,1.0999999,0.50000006,0.0,0.022222223,0.0,0.49166667,2.0222223,3.1833336,4.0444446,18.633335,25.844444,37.011112,42.11667,29.311111,10.341666,3.6888888,2.966667,0.7555556,0.3,0.09166667,0.10000001,0.0,0.0,0.0,0.0,0.074999996,1.8555555,7.6444445,25.858334,34.27778,6.9833336,6.755556,3.7416663,3.6999998,2.8111112,1.1083333,0.6555556,0.091666676,0.055555556,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.32222223,0.69166666,2.0,2.141667,1.888889,3.5333333,5.9888887,4.7,2.6833332,2.188889,4.5333333,7.744445,9.191668,11.966667,7.044445,1.3083334,0.18888889,0.09166667,0.022222223,0.13333334,0.0,0.0,0.0,0.0,0.0,0.12222223,0.6,1.9833333,2.688889,3.5777779,3.7416666,2.4666665,1.5833333,1.3111112,1.7666667,1.3000001,0.5888889,0.59999996,0.68888885,0.6916666,0.7444445,0.9583333,0.12222222,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.11666667,0.22222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,0.24444446,0.81666666,0.62222224,0.625,0.8999999,0.6,0.40833336,0.10000001,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.5833334,2.4,2.8,0.8666667,0.07777778,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,1.5888889,2.5583334,1.2,0.125,0.06666667,0.26666668,1.9222221,1.9555556,1.0916666,0.3,0.8666667,1.3333334,0.625,0.14444445,0.06666667,0.05,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.15833333,0.08888889,0.09166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,0.0,1.2111111,1.1583333,1.7444445,4.791667,6.8222218,12.750001,16.5,14.077777,9.891666,8.233333,12.408334,14.555555,8.183333,0.8000001,0.022222223,0.13333334,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11111111,0.5666667,2.4333334,6.9,6.425,4.8222227,4.5249996,6.2777777,4.055556,2.05,2.0666666,0.7916666,0.70000005,0.79999995,2.9222224,4.477778,3.2666664,1.4444444,0.51666665,0.1,0.40833336,1.1444445,0.96666664,4.288889,3.0444446,1.1,0.25555554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.79166675,0.0,0.0,0.0,0.16666669,0.3666667,1.8555557,1.7166667,7.922222,16.975002,14.455555,22.244444,31.583334,23.01111,3.45,4.3888893,1.4333334,0.099999994,0.6888889,0.48333335,0.31111112,0.0,0.0,0.0,0.0,0.0,0.78888893,4.7555556,17.358334,14.222221,18.091667,30.122223,19.208334,3.0555553,2.6333332,1.5666668,0.1,0.058333337,0.033333335,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333332,1.125,7.155556,8.158334,1.5666666,2.4416668,5.644445,8.911112,7.983333,3.6111114,5.4083333,9.644444,8.475,8.677778,10.177778,8.833334,3.6777778,0.96666664,0.9,0.78333336,0.6888889,0.4333333,0.31666663,0.033333335,0.0,0.0,0.0,4.175,2.4666667,1.2916667,0.62500006,0.4,0.28750002,1.0916667,1.44375,1.3,0.9,0.73125005,0.7583333,0.60625005,0.7916667,0.8875,1.2166667,1.1750001,1.1833334,1.0083333,1.2250001,0.5583334,0.33125,0.15,0.10000001,0.008333334,0.008333334,0.03125,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.13125001,0.19166666,0.087500006,0.29999995,0.70624995,0.6916667,0.66666675,0.33125,0.23333335,0.050000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45833334,3.625,3.875,1.85,0.18125,0.0,0.0,0.0,0.05,0.06666667,0.175,0.0,0.0,0.04375,0.0,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14375,0.24166667,0.05,0.075,0.083333336,0.075,0.16666667,0.4375,3.5333335,2.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17500001,0.5416666,1.10625,3.3666668,0.9499999,0.2,0.008333334,0.35000002,0.8000001,0.98125,10.616667,14.225,12.533334,15.299999,12.487499,7.5249996,3.99375,1.6333334,0.41250002,0.50000006,0.54999995,0.35000002,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.075,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,1.175,2.7083335,5.9312506,8.45,5.29375,2.7416666,3.8500001,2.7333336,4.05,3.6625004,1.575,0.68125,0.28333333,1.14375,2.641667,1.7,0.7500001,0.30833334,0.58750004,0.3083333,0.84375,0.575,4.68125,8.483333,8.683333,2.525,1.0583333,0.21875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.016666668,0.74375004,4.1083336,3.1375,13.775,20.562498,13.241666,7.5749993,7.7250004,8.599999,6.1,5.2666674,0.5625,0.56666666,1.1583334,2.08125,1.5500002,0.8937501,0.3416667,0.80625004,2.9583335,0.98749995,0.80833334,2.0416667,9.131251,8.716667,15.400001,13.416666,6.05625,1.0416667,1.3583333,0.44375,0.0,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333333,0.3125,3.266667,18.6875,25.366669,8.63125,2.6416667,5.4083333,9.65,10.666667,13.5625,27.2,24.143751,13.675001,12.725001,10.056251,6.3916674,5.33125,4.9750004,2.6999998,0.85833335,0.75,1.6062499,0.34166667,0.0,0.0,0.0,5.9666667,5.888889,4.722222,1.8083334,0.4333333,0.15000002,0.47777778,0.45833334,0.53333336,0.87777776,1.1916666,1.4777777,1.5250001,1.5444446,1.7750001,1.611111,1.1083333,0.7111111,0.43333334,0.52500004,0.5888889,0.5166667,0.4222222,0.36666667,0.49999997,0.15555556,0.083333336,0.122222215,0.25,0.18888889,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11111111,0.0,0.08888889,0.48333335,0.8333334,0.20833333,0.29999998,0.54444444,0.66666675,0.2,0.025,0.0,0.008333334,0.1,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,0.4111111,0.06666667,0.75555557,0.28333333,0.0,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2666667,0.48333335,0.33333337,0.6666667,2.2555556,12.2,26.177776,11.0,0.9777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8,0.64444447,3.2749999,3.6222222,3.2,4.6000004,4.155556,2.891667,1.1777776,0.3416667,0.033333335,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.033333335,0.08888889,0.24166667,0.3888889,0.26666665,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,0.88888896,2.9666665,5.4,4.6222224,3.7833333,1.5777777,2.1166666,4.2,4.8111115,3.2250004,1.4888889,0.1,0.18888888,0.5416666,0.23333335,0.14444444,0.041666668,0.0,0.26666665,0.6777778,0.2,2.9111114,5.3916664,7.6888885,10.944445,2.475,0.6333333,0.09166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46666664,0.099999994,1.1666667,3.1555557,3.4416664,8.98889,18.508333,19.322222,11.244444,5.1416674,4.6,2.2916667,0.2777778,0.1,0.28888887,0.35555556,0.57500005,1.1333334,1.0000001,0.42222226,1.35,5.4444447,8.125,4.622222,3.4333336,5.2333336,0.79999995,5.833333,3.7666664,6.6000004,0.13333334,0.0,0.0,0.2888889,1.8416667,0.40000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.44444445,0.0,0.9333333,0.0,0.75,1.288889,9.841667,19.555555,15.266668,6.7222223,5.4777775,3.1750002,2.7222223,2.4250002,5.0222225,9.666667,12.944444,12.322224,6.0666666,4.6333337,8.816667,10.244446,9.425001,5.4,2.7333333,2.6833336,1.3444445,0.025,0.0,0.0,6.5562496,4.208333,3.6583333,4.1187496,1.9500002,1.0812501,1.1916667,1.3874999,1.8666667,1.7333333,2.3375,2.3749998,3.6062498,3.7916667,4.76875,3.1833334,2.5187502,3.4916668,3.275,2.225,2.4416668,1.83125,1.675,1.1437501,0.5666667,0.8500001,1.0375001,0.71666664,0.36875,0.15833333,0.34375,0.325,0.19999999,0.375,0.033333335,0.025,0.0,0.0,0.0,0.0,0.0,0.10833333,0.09375,0.008333334,0.09375,0.041666668,0.575,0.45000002,0.49166667,0.1875,0.25833336,0.29375,0.21666667,0.1875,0.09166667,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.074999996,0.30624998,0.1,0.0,0.13333334,0.025,0.1,0.09375,0.09166666,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7437501,4.3333335,0.43125,0.0,0.0,0.0,0.0,0.0,0.0,0.16250001,2.5666666,6.2625003,2.8750002,1.0687501,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21666667,0.5375,0.05,0.083333336,0.13750002,3.1833334,11.743751,7.241667,7.937501,5.933333,4.4333334,1.93125,1.1166667,0.28125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.225,0.09166667,0.53125006,0.75000006,0.74375,0.35000002,0.03125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,1.3333334,3.9416664,2.59375,1.8,2.075,3.2416666,6.4125,3.9416664,2.7833333,2.6187499,0.6916667,0.27500004,0.21666667,0.28750002,0.05,0.09166666,0.025,0.11666667,0.41250005,0.108333334,1.34375,3.5583334,3.7437499,2.3833332,1.0333333,0.06875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08125,0.28333333,0.0,0.20625001,0.43333334,3.01875,20.583332,20.03125,18.408333,13.783333,5.6625,1.9583334,0.49374995,0.06666667,0.0,0.0,0.05,0.19375002,0.083333336,0.0,0.15,4.275,9.724999,11.91875,3.2833335,1.6916666,1.7125001,0.0,0.0,0.116666675,0.0125,0.0,0.0,0.26250002,3.6333337,2.5625002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.0,0.0,0.05,0.34375,1.1416667,1.6937501,5.116667,5.6062503,2.6666667,2.3000002,2.6875002,2.4666667,0.7625,0.54999995,1.6437498,3.875,3.7250004,1.86875,4.425,6.6687503,7.875,8.293751,5.6000004,5.316667,4.1687503,0.68333334,0.10625,0.0,0.0,4.8416667,6.5555553,8.233334,6.1083336,3.7111113,1.1750001,1.7111111,1.4416666,1.4777777,1.5888889,2.0166667,1.9777778,2.3666666,1.5888889,1.7166667,2.3444443,2.4500003,2.9222226,4.7555556,7.3999996,6.4666667,4.158333,2.4111114,2.1416667,2.0333333,0.9444444,1.4999999,1.5777779,0.7333334,0.34444442,0.12500001,0.31111112,0.31666666,0.5555556,0.6777778,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.074999996,0.23333335,0.05,0.0,0.033333335,0.375,0.31111112,0.11666667,0.10000001,0.20000002,0.11111112,0.050000004,0.0,0.0,0.0,0.0,0.041666668,0.07777778,0.125,0.05555556,0.18888888,0.06666667,0.0,0.0,0.06666667,0.17500001,0.3,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14166667,3.0777779,1.3000001,0.53333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9777778,2.175,2.277778,2.488889,2.0833335,5.2111115,17.55,15.17778,11.474999,4.8555555,1.7888889,0.39166668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.044444446,0.21666667,0.33333334,0.7111111,1.1666666,0.5888889,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.016666668,0.0,0.05,0.6666667,1.2333333,3.477778,2.9,0.6666667,0.96666676,3.8083334,8.733334,6.8,5.0666666,3.4111109,2.483333,0.9444445,0.39999998,0.36666664,0.19166666,0.44444442,0.5222223,0.041666668,0.044444446,0.058333337,0.8,2.2416668,2.3222225,1.0083333,0.14444445,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777777,0.6666667,1.2777778,9.258333,22.977777,23.849998,14.566667,8.944445,2.6166666,0.24444444,0.2666667,0.17777778,0.325,0.044444446,0.07777778,0.6166667,0.0,0.0,0.8888889,5.05,8.933333,3.9250002,0.0,0.044444446,0.9666667,0.37777779,0.0,0.0,0.0,0.0,0.0,0.05,2.1555555,1.425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.088889,0.9,0.22222222,0.30833334,0.9888889,1.3444444,0.68333334,0.81111115,0.79166675,0.055555556,0.033333335,0.13333334,0.48888886,0.95833325,3.7333336,6.1916666,6.4777775,7.4750004,8.111112,11.233335,9.75,5.4444447,1.7583334,0.1777778,0.0,1.9437499,4.1083336,3.8333333,3.6312501,2.1083333,1.73125,2.0583334,1.6812501,1.2166667,0.47500002,0.33749998,0.40000004,0.30625004,0.65000004,0.8812499,1.7,1.9312501,2.791667,4.8,7.98125,10.166667,8.8125,6.1583333,2.99375,1.1666666,0.9583334,0.9875001,0.9749999,0.9250001,0.59999996,0.30625,0.008333334,0.0,0.0,0.0,0.1,0.0,0.0,0.0,0.0,0.0,0.025,0.0625,0.0,0.0,0.0,0.00625,0.0,0.0,0.0,0.041666668,0.16250001,0.18333335,1.2375001,1.2416667,0.30624998,0.14999999,0.0,0.0,0.0,0.0,0.0,0.3375,0.5333333,1.075,0.64719653,1.0555556,0.6252778,0.35227272,0.15625,0.058333334,0.04375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6,0.38333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.716667,5.075,4.483333,3.8083332,3.79375,8.75,9.75625,7.4083343,1.35,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.2875,0.34166667,0.44374996,0.925,0.5916667,0.2375,0.15833333,0.050000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16874999,0.6416666,0.61249995,0.8,2.5125,5.625,4.76875,1.6750001,0.6,0.95624995,1.7083334,7.8187504,9.341667,8.01875,7.5166674,3.291667,1.81875,1.1333334,1.00625,1.2583334,0.52500004,1.1416668,0.25833336,0.0,0.05,0.875,2.0583332,1.7125,1.0500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5333333,1.85625,6.333334,11.36875,18.316668,16.81875,10.0,4.241667,0.63125,0.3416667,2.4625,11.366667,5.63125,2.3249998,1.3166666,0.70625,0.033333335,0.0125,2.9,13.1875,13.85,4.20625,0.25,0.058333337,0.47500002,1.9916667,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8000001,2.15,2.4666667,1.7187501,0.9583334,1.075,0.175,0.13333334,0.18125,0.0,0.0,0.008333334,0.21666668,1.3625001,2.125,5.74375,7.7833333,7.0624995,5.6833334,6.8333335,6.6687503,4.3583336,1.8000001,0.075,0.0,0.016666668,0.2777778,0.06666667,0.79166675,1.4000001,1.9833333,1.8666668,1.1750002,1.4222223,1.5444444,0.625,0.6222222,1.2333333,2.1222224,2.9833333,4.2222223,4.833334,4.9111114,3.577778,3.425,5.0,5.3,4.5222216,4.016667,3.3555555,3.4666665,3.3083336,2.222222,0.4,0.7666667,1.6416668,0.6888889,0.16666667,0.0,0.0,0.0,0.022222223,0.0,0.0,0.0,0.0,0.022222223,0.23333336,0.5333333,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8777778,4.841666,4.6333337,1.5,0.122222215,0.044444446,0.058333334,0.0,0.0,0.0,0.025,0.111111104,0.36666667,1.6999999,1.977778,3.325,3.2333333,1.5166667,0.37777779,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.51111114,2.8333333,2.8333333,0.5083334,0.0,0.0,0.0,1.888889,11.016666,5.8000007,1.2166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.9111111,0.45,1.0666667,0.3333333,2.4777777,4.6916666,5.9,4.833333,3.9,8.444445,13.224999,4.933334,0.375,0.022222223,0.0,0.0,0.0,0.058333334,0.022222223,0.0,0.0,0.0,0.0,0.0,0.05,0.45555556,0.65000004,0.2888889,0.6666666,0.36666667,0.044444446,0.65,0.34444442,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40000004,0.85555553,2.8416665,4.833334,6.500001,5.8,3.7916665,1.1444445,1.0333333,1.2750001,4.2222223,7.6500006,4.9111114,5.666667,5.5111113,0.9555556,0.6666667,0.67777777,0.89166665,0.32222223,0.80833334,0.44444448,0.0,0.0,0.8666667,1.5166667,1.3444444,0.84166664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.17777778,3.0166667,7.1,7.6250005,9.288889,12.058333,8.133334,4.366667,3.8833332,7.7333336,13.616667,23.122223,14.841666,7.5666666,4.233333,1.425,0.07777778,2.5416667,8.622222,14.416666,10.388888,5.1416664,5.333333,1.9333334,0.98333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22222222,0.8000001,1.0111111,3.4916666,2.9555557,6.9333334,14.444444,11.677777,5.258333,1.5111111,1.95,0.24444446,0.0,0.17777778,0.8777778,1.4250001,1.5888889,2.1583335,4.611111,7.308334,10.922222,10.0,4.858333,1.6333332,0.35833335,0.011111111,0.0,0.0,0.0,0.022222223,0.6416667,0.76666665,0.6750001,0.78888893,0.48333338,1.9333335,2.2,1.6333333,1.5444444,1.075,1.8,1.9749999,2.9333336,3.0583336,4.077778,3.1777778,2.8166666,2.1999998,1.5583334,1.4000001,0.45833334,0.95555544,2.4,3.766667,3.2000003,2.2250001,3.5777779,0.76666677,3.5444443,3.725,1.3222222,0.11111111,0.09166667,0.3888889,0.23333335,0.08888889,0.0,0.0,0.033333335,0.56666666,0.8222223,0.40833333,0.0,0.14166667,0.099999994,0.0,0.0,0.0,0.116666675,2.0111113,5.625001,6.577778,1.3916668,0.24444444,0.033333335,0.0,0.0,0.0,0.0,0.0,0.011111111,0.08888889,0.06666667,0.42222226,1.3666666,2.6555555,2.5833337,1.5777777,0.44166663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.025,0.14444445,0.24166667,0.044444446,0.0,0.0,4.2666664,13.683333,13.322223,2.3500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,1.5333334,2.0,5.044444,10.225,10.344444,4.4083333,5.2666664,4.5583334,4.088889,2.766667,2.6666663,3.1222222,3.6666667,0.31111112,0.025000002,0.0,0.0,0.1,1.0111111,1.2166667,0.0,0.0,0.0,0.0,0.0,0.0,0.275,0.44444445,0.3,0.2777778,0.65,0.055555556,0.46666664,1.175,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.025,0.0,0.0,0.14166668,1.4777778,3.2500002,5.822222,5.575,3.022222,2.3166666,1.1444445,1.0888889,3.1333332,7.9888887,6.316667,6.9444447,9.475,4.4444447,0.8888889,1.025,1.588889,0.5,0.32222223,0.26666668,0.044444446,0.0,0.075,0.90000004,0.85833335,1.2,0.21666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.125,0.0,0.0,0.0,0.0,0.022222223,0.0,0.44444445,0.36666667,3.1916666,4.0333333,3.0083332,4.7777777,7.691667,27.244446,18.944447,7.1500006,16.28889,23.341667,24.688889,24.200003,14.688889,11.322223,5.7666664,3.1333334,5.1833334,12.6888895,12.733334,7.4444447,5.1333337,7.6666665,1.8999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.0666668,6.0,3.1222222,4.1416664,7.0111113,8.911111,7.941666,1.3555557,1.4499999,1.4666667,1.0166667,0.62222224,0.4888889,0.09166667,0.23333332,1.9416668,5.8333335,7.791667,7.566667,6.277777,3.858333,1.6999999,0.7416667,0.17777778,0.0,0.0,0.016666668,0.083333336,0.5,0.30833334,0.25625002,0.16666667,1.1750001,1.6166668,0.7250001,0.40624994,0.5833333,0.53125,0.4833333,0.25000003,0.5083334,1.3687501,2.0083332,1.6833334,2.59375,3.175,2.65625,4.0833335,4.706249,2.825,3.0000002,4.025,1.9166669,0.95000005,0.76666665,0.59375,0.73333335,2.075,1.9583333,0.70000005,0.0625,0.15833333,1.14375,1.2,0.0125,0.0,0.0,0.125,0.8083333,2.2624998,0.9750001,0.90000004,0.32500002,0.23333335,0.0375,0.0,0.3,2.341667,3.875,3.7000003,1.5875001,0.8333334,0.49166664,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.28333336,1.3937501,1.6083333,0.54375005,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26875,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.16666667,0.78749996,1.1833334,1.23125,2.3833334,2.7833335,4.51875,6.133333,10.80625,13.516666,5.4875,1.7166667,2.8937502,2.0,1.0416667,0.49375,0.13333334,0.075,0.0,0.0,0.0,0.0,3.725,12.308333,3.7625,0.8833333,0.0125,0.0,0.0,0.0,0.0,0.087500006,0.175,0.0375,0.8166667,0.30624998,0.125,1.125,0.93125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19375,0.41666666,0.0375,0.0,0.0,0.0,0.46666667,4.4812503,7.3250003,3.64375,1.9000001,0.9499999,1.1666666,2.3,3.7125,3.1583333,4.7875,6.950001,4.6749997,3.0916667,2.3333335,1.2375001,0.55833334,0.2875,0.625,0.225,0.0,0.0,0.0,0.30000004,0.75624996,0.30833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0375,0.0,0.25,0.58124995,0.0,0.0,0.033333335,0.175,0.8666667,0.23750001,0.041666668,2.2666667,3.39375,3.6500006,3.6250002,3.2250004,5.86875,16.325,12.916666,24.181252,29.516668,30.13125,21.008333,26.406252,21.650002,12.083333,6.43125,4.875,6.60625,7.016667,14.18125,14.016666,6.48125,4.0166664,1.675,0.2875,0.0,0.043750003,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.5666666,1.5500001,1.5416667,4.525,3.225,1.7375,0.89166665,0.5,0.2,0.0,0.01875,0.22500001,0.25,1.425,0.30833334,0.13125,0.0,0.16874999,0.7083334,1.28125,2.5833335,3.7083335,3.76875,2.3083332,0.5375,0.05,0.175,0.0,1.6222222,1.7222223,0.5583334,0.42222226,0.79166675,1.4555556,0.9583333,0.6111111,0.3222222,0.55833334,0.5777778,0.275,0.34444442,0.3166667,0.2777778,1.2750001,1.2222222,0.6666667,1.5250001,2.1555555,2.1833334,2.5,3.8333333,6.3555555,7.611111,4.2083335,1.1111112,1.0,0.42222223,0.8916666,1.2111111,0.35000002,0.43333337,1.4111112,1.2166667,0.6111111,0.36666667,1.4555557,0.7666667,0.022222223,0.0,0.025000002,1.2555556,2.025,2.3777778,2.3916667,2.8222222,1.0444444,0.18333334,0.033333335,0.041666668,1.4,2.6,1.8555555,0.53333336,1.488889,1.7444444,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22500001,0.25555557,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,1.7500001,1.7000002,0.39166668,1.5666666,1.9333333,2.3333333,2.0333335,2.7083333,1.1111112,5.1583333,14.811111,25.95,13.544444,5.5499997,4.6888885,3.5000002,1.6166669,0.9111111,0.15,0.26666668,0.06666667,0.0,0.23333333,4.45,10.233334,8.808333,2.3888888,0.025,0.0,0.0,0.075,0.011111111,0.0,0.0,0.06666667,0.35555556,0.050000004,0.33333334,1.2222223,0.09166667,0.0,0.05,0.26666668,0.20833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,0.97499996,0.17777778,0.0,0.0,0.0,0.5083333,2.788889,5.358333,4.266667,1.825,0.32222223,1.0083333,2.5222223,1.4555556,0.9250001,1.0666667,4.4083333,4.466667,4.8166666,3.3555555,2.5333333,0.95,0.2777778,0.46666667,0.11111111,0.0,0.0,0.0,0.0,0.0,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31111112,0.1,0.0,0.15555555,0.23333333,0.07777778,0.0,0.22222224,0.76666665,1.9333334,1.0833334,0.5,3.7888887,4.491667,4.2777777,1.6916667,1.6555556,4.0083337,22.222223,25.122225,27.5,27.277779,19.075,9.711111,15.891666,27.311111,23.599998,13.333333,10.711111,15.933332,16.877777,12.375001,4.911111,3.65,1.3222222,1.2777777,0.275,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40000004,5.083334,3.3111112,0.39166668,0.61111116,0.033333335,0.93333334,0.8222222,0.05,0.0,0.26666668,0.7777778,0.0,0.0,0.0,0.033333335,0.044444446,0.24166667,0.5888889,0.36666667,0.21666667,0.6999999,0.06666667,0.0,0.38333333,1.26875,2.4416666,1.5916667,0.075,0.47500002,1.5625,2.7083333,2.4375,2.3750002,1.6083335,2.1,2.2166667,2.65,2.7583332,1.6,0.92499995,1.1187501,1.2416668,1.7166668,1.6750001,0.95,1.3499999,0.8416667,1.2624999,1.7250001,0.8166667,1.4875,3.6,8.075,3.9166667,0.78749996,1.2916666,1.475,1.275,0.87500006,1.3375,2.6666667,1.3249999,0.675,1.7875001,3.7083335,2.5666668,0.2875,0.22500001,1.2625,3.1416664,4.475,4.4999995,3.2833335,1.5999999,0.11666667,0.125,1.4583334,2.1437502,1.5500002,2.9375,3.0083332,1.175,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.48749998,0.35833332,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09375,0.5500001,0.525,0.081250004,0.6083334,1.5937501,2.1000001,2.20625,2.0916667,5.6666665,8.443749,6.375,8.225,15.050002,31.031248,22.791668,9.25,4.4249997,1.5333333,1.0125,1.0416667,0.4,0.125,0.05,0.0,0.0,1.21875,14.058332,15.19375,4.2333336,0.1375,0.041666668,0.525,0.39374998,0.008333334,0.0,0.0,0.00625,0.008333334,0.0125,0.23333335,0.2916667,0.70625,0.5833334,1.46875,1.4416666,0.95000005,1.7416667,0.69166666,0.0,0.0,2.63125,0.82500005,0.0,0.0,0.0,0.0,0.0,0.01875,0.21666667,0.55,0.033333335,0.0,0.3333333,0.42499998,1.0,2.0333333,1.7499998,1.1083333,0.43125004,0.60833335,2.7312503,1.3333331,0.34166667,0.19375001,2.4333336,4.0062504,4.6249995,3.5562499,1.9416665,1.8083334,0.59999996,0.05,0.056250002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.38333333,0.0,0.28333336,1.0333333,0.33124998,0.49166667,0.1875,0.40000004,1.30625,1.4666666,1.5749999,2.7,3.5666664,4.5875006,3.9499998,1.10625,1.6666667,5.2875,15.000001,24.633335,22.525002,14.941667,13.3375,15.141666,20.6375,28.425,31.933334,27.28125,19.883335,24.231249,21.841667,13.9375,7.591667,2.1999998,1.7333332,4.025,1.7437501,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.6166667,0.55,0.0,0.0,0.0,0.0,0.0,0.0,0.1,1.05,1.5,2.5874999,0.6416667,0.0,0.0,0.1,0.24166667,1.4124999,1.4166666,0.22500001,0.8375001,2.1083336,1.0187501,0.18333334,0.0,0.008333334,0.041666668,0.29999998,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.0125,0.0,0.0,0.38333333,0.7888889,0.23333332,0.083333336,0.3888889,0.87499994,1.3111112,2.4750001,1.8,2.6333334,2.7666667,2.2222223,2.575,2.6777778,1.2333333,0.81111115,2.1166668,1.7333335,1.2555556,1.1666666,1.0444444,1.1083333,1.1333334,2.5083332,1.9222223,1.4222221,1.5333333,2.5777779,0.9583334,0.4666667,1.2,2.788889,4.008333,4.522222,3.877778,2.1333332,1.1333333,3.0333333,3.2444444,1.2666667,1.7,5.133333,5.641667,0.6333333,0.041666668,0.4,1.6250001,3.1444442,4.733333,4.608333,5.1555552,2.1916666,1.4999999,1.0416666,1.9777777,5.2750006,3.3111112,0.46666667,0.11666667,0.08888889,0.1,0.9888889,0.23333335,0.0,0.0,0.083333336,0.5111111,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.0,0.0,0.0,0.0,0.016666668,0.06666667,0.3111111,1.4916668,4.2777777,2.3166666,0.111111104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9666667,0.73333335,2.266667,2.1000001,1.4444445,0.25,0.0,1.2750001,4.322222,7.422222,21.291668,18.311111,10.466667,6.477778,4.1333337,2.8333333,3.1333337,1.2555556,0.06666667,0.016666668,0.11111112,0.041666668,0.0,0.0,0.0,0.055555556,0.9916668,6.9333334,16.45,2.0333335,0.33333334,0.33333334,0.49999997,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.8111111,1.4666667,3.7444444,3.5416667,2.8777776,3.575,4.8444443,0.82222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.16666666,0.44166666,0.0,0.1,0.46666664,0.29999998,0.4666667,0.08888889,0.23333335,0.25555557,2.0333333,2.3333335,1.7,0.7777778,0.15555556,1.6,2.7444441,3.25,1.7888888,0.6,0.8333334,1.2666668,0.45833337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,0.32500002,0.32222223,0.05,0.24444447,0.43333334,0.5666667,0.64444447,0.6916667,0.44444445,2.125,0.8666668,1.2166667,1.4333334,2.7555554,4.616667,1.8333334,1.3916667,3.8,4.9333334,13.566667,20.9,22.55,12.233333,15.658333,15.811111,13.616667,16.366669,18.722221,22.275002,26.800001,27.883333,29.52222,16.2,5.1666665,1.9083335,9.433333,14.155556,3.7166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24444446,1.5416666,0.73333335,0.0,0.0,0.0,0.0,0.0,0.6,0.8,0.4,3.8333335,1.4777778,0.0,0.022222223,0.033333335,0.0,0.13333334,0.4888889,0.6666666,2.45,3.9444447,1.9416666,0.24444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.4562497,1.175,0.4333333,0.25625002,0.275,0.68125004,0.6,1.09375,1.75,3.0166667,1.6062499,1.5583334,2.75625,2.416667,2.3562498,3.1416664,4.7000003,3.891667,3.8583333,3.225,2.1666665,2.15625,1.9916666,2.575,2.5083337,2.8833332,4.35,4.875,3.6250002,3.5416667,3.7125,3.375,2.675,2.6000001,3.0166667,2.5125,1.9750001,1.5875001,3.1833334,3.675,1.8166667,1.2,3.40625,4.7416673,1.2249999,0.09166667,0.6625,2.7916665,6.9416676,7.10625,6.0249996,4.075,1.2916666,1.5062499,1.4666668,3.5437498,1.7083334,0.48333335,0.081250004,0.13333334,0.36875,2.175,3.1375,1.0666667,0.26666668,0.0,0.40833333,1.59375,0.35000002,0.0,0.275,0.6875,0.17500001,0.39999998,0.41875005,0.05,0.38125,0.1,0.00625,0.26666668,0.8666667,2.125,2.6166666,2.26875,0.41666666,0.95625,0.18333334,0.0,0.0,0.0,1.9000001,4.666667,0.0625,0.0,0.5125,2.025,6.541667,9.525,5.3083334,3.3937502,0.1,0.425,0.49166667,3.8666668,19.0,26.45,34.11875,19.858334,16.731249,10.483334,4.9812503,1.5583335,1.2583333,1.6000001,0.24999999,0.01875,0.0,0.44375,0.69166666,1.0583334,1.3999999,3.7,4.14375,3.0749998,2.3812501,0.425,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7,3.7833335,4.21875,15.791668,27.631248,29.858332,24.287502,7.5666666,1.7833333,0.3875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.34166667,0.5375,0.35000002,0.10625,0.0,0.10625,0.116666675,0.016666668,0.0375,0.17500001,0.6,2.916667,3.0000002,1.2333335,0.65,0.175,1.325,3.5249999,2.5583334,0.99375004,0.81666666,0.8250001,0.8666667,0.2916667,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.80833334,0.86249995,0.28333336,0.41250002,0.0,0.35,1.4875001,1.2666667,0.79999995,0.86666673,1.1937499,0.22500004,0.675,1.4000001,2.1,2.7875001,2.1583333,1.2375001,3.1916666,8.531251,20.850002,24.808332,20.2875,29.266668,17.7375,15.533333,13.931251,16.075,17.633333,20.95625,26.225,30.3875,26.166666,15.806252,5.9583335,2.8125,4.3083334,6.1083336,1.35625,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.112500004,0.0,0.0,0.0,0.0,0.95,1.8333334,0.0,0.0,0.0,0.0,0.0,1.7250001,3.8416667,3.4125004,0.375,0.025,0.058333337,0.0625,0.0,0.0,0.0,0.2916667,0.39374998,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.75,0.8333334,0.27777776,0.6333333,0.22222224,0.033333335,0.0,0.125,2.288889,6.755556,3.2500002,1.1555556,1.4749999,3.0555558,7.583334,9.966666,7.633333,7.077778,3.622222,2.3666668,1.8555557,1.5666666,2.0333333,2.3083334,1.6000001,4.211111,5.341667,4.9444447,4.366667,3.2222223,2.7250004,2.6,1.8583332,1.1777778,1.2111111,1.4833333,1.4555557,1.6416668,2.1555557,5.233333,7.077778,3.2,0.95000005,2.288889,4.408333,1.1666666,1.4666666,3.8333333,5.6888885,3.7999997,3.0000002,2.3,1.2333335,1.0333334,3.0888891,6.108333,6.633333,2.4666665,1.0666667,0.07777778,0.16666667,0.8,2.3000002,1.6777778,0.24444446,0.0,0.055555556,0.8833333,6.677778,12.150001,5.7444444,1.175,0.57777774,0.07777777,0.06666667,0.34444445,0.76666677,0.8333333,0.9833333,0.46666667,0.25555557,0.78333336,0.6333333,2.1583333,1.8444446,0.68333334,0.0,0.17777778,0.06666667,4.1555557,18.916668,22.400002,9.383333,0.0,1.6499999,7.2000003,8.044445,16.208332,33.11111,22.5,13.033333,6.15,6.033334,8.755556,26.133333,29.011112,31.791666,22.088888,24.25,29.122221,14.225,6.9666667,0.85,0.20000002,0.42222226,0.44166666,0.7444445,0.80833334,0.7888889,2.1333332,3.7499998,8.255556,9.141667,11.0222225,4.016667,0.25555557,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.8666667,0.8444445,2.3333333,2.022222,2.8083334,6.3111115,10.041668,16.244444,0.5777778,1.9333334,1.0666667,0.0,0.0,0.0,0.0,0.0,0.3333333,1.7222223,1.2916667,0.08888889,0.0,0.0,0.0,0.0,0.0,0.083333336,0.3666667,2.8833337,4.0111113,1.0999999,0.84444445,0.325,1.0333333,2.7111113,2.1916666,0.53333336,1.0083333,0.9777778,0.67499995,0.32222223,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,0.35555556,0.56666666,0.24444444,0.3333333,0.022222223,0.73333335,1.1583333,1.4444444,1.1916667,0.9999999,1.4000001,1.2222223,3.1083333,3.5222223,2.9555557,2.3666666,1.5888889,1.975,8.322223,15.433334,35.91111,34.31111,37.758327,47.433334,43.158337,24.777777,15.691668,20.099998,10.91111,11.591667,13.555555,20.875002,24.933334,15.425001,4.044445,2.2416668,3.1555557,2.0666666,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40000004,1.6916666,0.35555556,0.0,0.0,0.73333335,1.7111111,0.48888892,0.26666665,0.0,1.0666667,0.28888887,0.47499996,0.5666667,0.86666673,3.175,1.5666666,1.2166668,0.15555556,0.025,1.0111111,0.36666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26875,0.3,0.27500004,0.0375,0.0,0.0,0.0,0.46874997,3.191667,7.0166674,7.225,5.5916667,3.6937501,1.4416667,1.425,3.2,1.9749999,1.4083333,1.2333333,0.95625,0.35833332,0.38125,0.55,0.9375,2.1166668,2.9250002,4.56875,3.9083338,3.5187502,3.2416668,1.675,0.9333334,1.9125001,1.6583333,0.35000002,0.35624996,0.29999995,0.29999998,0.49999997,1.4437499,4.583334,6.5333333,4.2,1.1333333,1.86875,5.791667,6.7124996,5.6083336,3.7916672,2.0500002,0.9,0.75,1.0083332,1.6125001,2.5333335,3.8249998,6.5000005,9.5,8.88125,6.5000005,2.34375,1.4916667,1.06875,0.48333332,0.20833331,0.2875,0.116666675,0.58750004,7.491667,16.4625,9.925,4.58125,2.6999998,1.8833332,0.3,0.0,0.0,0.23333333,1.1625001,0.24166667,0.15,1.5749999,1.7,2.2875,0.82500005,0.26875,0.9000001,1.0083333,2.5062501,9.858335,22.48125,17.766666,10.3125,2.2166667,5.7437506,14.15,15.758334,30.43125,43.241665,42.893753,42.941666,26.70625,31.475,29.975004,31.062502,29.308334,21.006252,13.433333,12.043751,8.158335,8.412499,1.9333334,0.70075756,0.6329167,0.72121215,3.4401786,5.516667,8.21875,9.858334,9.008334,13.531251,9.658334,8.84375,4.8083334,1.1125001,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.16666667,0.2916667,0.675,0.35833335,1.10625,2.45,2.6625001,0.26666668,2.8,1.6437501,5.8500004,0.3875,0.075,0.0,0.0,0.03125,0.9166666,1.9166667,0.51875,0.05,0.0,0.0,0.0,0.0,0.016666668,0.13125,2.3000002,3.3625002,0.9333334,0.71875,0.30833334,0.74375,1.8333335,1.8833334,0.39999998,0.38333336,0.575,1.2833334,0.36875004,0.23333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37500003,0.4,0.10000001,0.041666668,0.11875,0.5833333,1.1583334,1.39375,2.4833333,1.48125,1.1250001,1.5,4.7083335,7.425,7.0666666,5.3416667,2.6062503,1.35,5.40625,21.525002,28.725002,34.225002,30.591667,22.112501,25.808336,24.75,19.25,11.650001,9.966667,7.366667,4.3875003,8.65,12.68125,15.133333,7.11875,0.125,1.0749999,1.0999999,0.6,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.075,0.0,0.0,0.0,0.0,0.18333334,0.0,0.275,0.8666667,0.1625,0.8416667,0.8062501,0.2,0.525,3.025,1.2916667,0.0,0.0,0.01875,0.35833335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4333333,0.1,0.18125,0.26666665,0.01875,0.0,0.0,0.18333332,0.2888889,0.17777778,0.05,0.0,1.0416666,1.4666667,1.2083334,3.5777779,7.488889,8.75,3.4666667,1.5333333,0.2777778,0.23333335,0.5666666,0.89166665,1.188889,1.2666665,2.7333336,1.8555557,1.2916667,1.3333334,2.125,2.411111,1.5444446,0.9833334,0.76666665,0.8416667,1.0111111,2.4916668,1.1,0.2166667,0.57777774,0.59999996,0.325,0.13333334,0.0,0.0,0.041666668,0.54444444,2.5444446,4.858333,3.755556,2.3750002,4.7555556,4.35,4.177778,2.0666666,1.8583333,1.2777779,0.9083334,1.6333333,1.5666668,1.0333334,0.8833334,1.0222224,4.277777,13.549999,27.155558,24.783335,15.500001,7.2,5.388889,1.3555557,0.5083334,0.6444445,0.36666667,0.4666667,2.15,3.5222228,3.033333,1.911111,1.5555556,0.60833335,0.044444446,0.0,0.0,0.46666664,0.0,0.3888889,2.375,2.3555555,1.25,1.0888889,0.97499996,1.9,3.333333,3.0249999,2.4222224,8.758333,11.055554,15.424999,12.6,23.725,34.055557,35.455555,54.758335,43.93333,31.100002,19.955557,20.025,29.922222,42.77778,37.075,26.233332,15.341667,22.122223,27.308336,15.377779,8.375,4.1333337,1.6111112,3.565,8.836112,14.128788,15.788889,22.308334,26.988888,28.21111,18.433334,5.244445,1.7416667,0.22222224,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.0,0.0,0.0,1.4416667,7.0111117,4.2833333,2.7666667,0.083333336,0.0,0.30833334,1.3555555,0.73333335,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.90833336,2.3,0.49166667,0.22222224,0.26666668,0.07777778,1.075,0.9111112,0.24444444,0.008333334,0.055555556,0.8000001,0.41111112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8333334,0.8666667,0.33333334,0.72222227,0.7166667,1.2777779,0.7555555,1.725,2.8333333,1.1,1.6444445,4.8916664,8.0222225,10.1,10.622223,6.977779,3.5750003,3.9333334,11.158334,23.41111,21.716665,14.088888,11.677778,8.333333,7.3444443,14.675,15.877779,14.366667,10.377778,6.455556,10.258333,13.155556,13.541668,11.611111,6.275,3.6333334,0.8416667,1.1000001,1.6,2.9,1.7333335,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.3333333,0.0,0.0,0.0,0.0,0.1,0.53333336,0.7,0.51111114,1.625,1.3444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333335,0.98888886,2.3,2.2666667,1.3222221,0.46666667,0.0,0.0,1.1500001,0.24444446,0.68888885,0.65000004,0.6888889,3.0,0.6666667,0.49999997,0.9555556,2.6222224,0.65,0.2888889,0.4,0.0,0.4,0.6888889,5.041667,2.9444444,4.7333336,6.633333,6.8222227,3.5416665,3.088889,3.1916666,2.6111112,1.2444445,0.2,0.2,0.041666668,0.033333335,0.29166666,0.4111111,0.025,0.0,0.7333334,1.175,0.11111111,0.033333335,0.23333332,0.52500004,0.28888887,0.5,1.9583334,4.7111115,4.1416664,2.0,0.9,0.6333333,0.73333335,2.8000002,1.9444445,0.59166664,1.6555556,1.275,0.79999995,0.09166667,2.888889,3.9999998,4.95,26.433334,35.583336,27.055557,10.791666,15.6,12.3,2.2833333,0.8555556,2.6333334,1.211111,0.29999998,0.9444444,2.6666667,3.588889,4.477778,3.2000003,1.1444446,0.38333338,0.4,0.1,0.0,0.43333334,1.8416666,2.8999999,3.2333333,1.4444444,0.29166666,0.9666667,3.1333332,3.2,2.1444445,4.608333,5.4,13.35,17.211113,23.4,32.633335,22.57778,38.541664,23.044445,20.508335,13.077779,18.7,18.822222,24.633335,36.51667,34.988888,23.750002,16.8,14.016666,10.1,8.6,7.322222,8.955555,15.341667,14.755557,13.112627,16.543056,12.408334,11.122222,11.48889,6.5583334,1.6555555,0.34999996,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,3.725,6.888889,0.21666668,0.0,0.43333337,0.8444444,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,1.1000001,0.34444445,0.108333334,0.25555557,0.0,0.011111111,0.53333336,0.8333334,0.0,0.0,0.033333335,0.4583333,0.07777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.1777778,0.06666667,0.45000002,0.62222224,0.3166667,0.35555556,1.225,0.41111112,0.4777778,0.6166667,0.8888889,1.0583334,2.811111,5.5583334,10.277779,11.266665,9.155556,6.2999997,2.575,4.6111107,10.133333,9.933333,10.966668,5.2444444,5.4,6.2000003,3.3777776,5.575,10.288889,12.900001,11.200001,11.566667,13.033333,18.633333,19.2,13.311112,14.750001,9.922222,4.125,1.5222223,0.54444444,1.5249999,0.64444447,0.13333334,0.07777778,0.016666668,0.0,0.099999994,0.6833334,0.11111112,0.0,0.0,0.13333333,0.0,0.0,0.0,0.0,0.0,0.0,0.4666667,1.3888888,3.2583332,3.1,1.5,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.1000001,3.4583335,0.2888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.25555557,0.6,1.3,2.7666671,2.3833332,3.2555556,4.625,0.15625,0.43333337,1.8166666,3.2375,7.5333333,9.325,4.2166667,0.8750001,0.13333334,5.191667,4.7687507,0.7833334,0.52500004,0.45000005,1.2750001,4.3083334,4.2000003,3.5083332,5.3166666,7.1937504,13.958334,9.85,7.7416663,4.425,1.4416667,0.008333334,0.0,0.0,0.0,0.0,0.0,0.116666675,0.043750003,0.0,0.9416666,2.2250001,1.9666666,1.16875,2.6750002,1.7062502,0.075,0.025,0.29999998,2.3916667,2.5625,0.5083333,0.05,0.23333333,0.55833334,2.5875,3.575,1.4875001,1.4583333,0.43125004,0.23333333,2.18125,4.683333,3.6749997,2.3374999,11.0,21.39375,19.933334,16.5625,15.341667,18.625,7.5125,1.3916668,3.94375,9.733334,6.7875004,4.7833333,0.85625005,2.35,5.0666666,8.181251,6.35,1.66875,0.70000005,0.1375,0.0,0.46666667,2.1999998,4.6583333,3.7437499,1.05,0.91249996,2.6166668,3.3916664,1.9375,0.45,2.2250001,1.4166667,1.625,3.791667,8.362499,5.541667,6.458333,6.6312504,5.2166667,4.4062505,10.916667,22.112501,28.916666,25.816666,30.50625,34.958332,36.39375,38.916668,25.325003,16.708334,11.3625,9.833334,8.883333,7.5875,6.5424247,6.1608334,7.3833327,5.19375,4.716666,3.5416667,1.44375,0.3,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22500002,1.4833333,2.5375,2.6166668,0.0,0.17500001,0.1,0.14166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.16875002,0.008333334,0.09375,0.075,0.0,0.0,0.43125004,0.0,0.0,0.0,0.20833336,0.18750001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.24375,0.5916667,0.25,0.15,0.4416667,0.08125,0.0,0.63124996,2.7583334,3.0999997,1.6874999,0.825,1.4937499,5.133333,6.24375,12.849999,16.756248,16.775002,7.566667,3.2187502,2.341667,4.0375004,3.1,9.1875,11.766666,7.1500006,9.18125,7.5333333,3.31875,5.133333,7.2562494,6.708333,8.875,11.818748,11.616667,12.118752,13.416667,19.525002,17.075,2.99375,2.05,1.8000001,1.1499999,1.2666667,0.64375,0.21666665,0.36874998,0.9833334,0.29166666,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.5625,1.7249998,1.925,1.2,1.8000001,0.9250001,0.0,1.5,3.3333335,3.0625002,3.25,0.01875,0.65000004,0.6,1.1625,0.9666667,1.925,2.4499998,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14375001,0.6666667,1.20625,3.1749997,3.8062496,0.19166668,0.15555556,0.7555555,2.5083332,5.1000004,9.974999,9.533334,1.7583332,0.36666667,3.6,2.8416667,1.1555556,2.141667,0.88888896,2.3750002,2.9999998,5.8833337,6.3666663,8.511111,8.591666,3.088889,5.933333,3.8222225,1.7083334,0.044444446,0.011111111,0.0,0.0,0.0,0.0,0.28333336,0.4888889,0.5083333,0.055555556,0.26666668,1.9583334,1.3333334,0.425,1.1444445,0.0,0.0,0.0,0.016666668,0.45555556,0.71666664,0.8222222,0.14166667,0.67777777,2.9333336,5.5249996,6.033334,3.5416665,1.2,0.3666667,0.6,1.8583336,1.6666667,3.3111112,6.375,9.388888,14.416667,14.000001,13.875,12.288889,8.388889,5.5750003,4.788889,7.6666665,11.733334,12.141668,10.633333,3.9,0.5777778,2.5222223,7.2500005,7.5222225,4.725,5.022222,2.3,0.41111112,0.044444446,5.141667,8.055555,5.1083326,2.611111,2.1666667,2.8222225,2.9666667,1.4916667,0.8777778,0.0,0.2,0.35833332,0.6888889,1.15,1.2888889,0.2,0.14166667,2.5444446,13.666667,26.822222,36.508335,47.511112,49.377777,62.733334,60.18889,47.408337,35.111115,18.008331,13.277777,9.450001,8.555555,7.377778,5.65,4.0111113,1.0916667,0.62222224,0.6416667,0.56666666,0.33333337,0.21666668,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,1.375,5.511111,2.4083333,0.22222222,0.0,0.4888889,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.325,0.0,0.0,0.041666668,0.12222224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17777778,0.05,0.11111111,0.06666667,0.06666667,0.12222223,0.058333337,0.0,0.50833327,1.3555555,2.466667,0.89166677,0.93333334,3.0916667,6.2111115,5.7,10.344445,15.5,20.300001,9.655556,8.166667,3.9555554,2.1416667,1.6111112,3.5083334,6.2222223,10.733335,11.183332,7.455555,5.0750003,5.1555557,4.925,3.1111112,2.3666666,8.475,11.500001,27.191666,18.377779,11.508333,7.622222,5.9333334,3.211111,1.0222223,1.625,1.8111111,1.4333334,0.8111111,0.108333334,0.53333336,0.22222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32222223,0.9666667,0.6666666,1.6083332,2.588889,1.2666667,1.1555556,0.0,0.0,0.0,0.0,0.0,1.5333333,0.22222224,0.0,0.0,0.11111111,0.3166667,0.08888889,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.25833333,1.2444444,4.2750006,1.3375,0.20833334,0.73333335,1.5062501,2.7416668,3.1375003,2.0416667,0.48125005,0.5,1.4583336,0.85625005,1.6,2.3375,2.9000003,3.7562501,3.6833334,5.81875,2.525,3.5,2.725,1.4583334,0.425,0.32500002,0.68125004,0.13333334,0.033333335,0.0,0.0,0.0,0.175,1.0062499,1.15,0.30624998,0.0,0.13333334,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.118750006,0.30833334,1.3125001,2.8500001,5.016667,4.49375,2.5333335,4.1875,4.8583336,2.0625,2.0833333,3.425,3.6583333,5.8333335,23.1875,19.04167,14.637501,5.966666,4.96875,6.5250006,6.6083336,7.3625,7.5833325,4.6562495,2.0916667,7.1125,9.7,9.84375,4.375,1.2166667,2.56875,4.1833334,4.28125,5.666666,5.7250004,2.725,2.591667,4.00625,6.808334,7.1687503,2.975,1.25,1.4166667,1.7666667,0.92499995,0.0,0.0,0.0,0.0,0.275,0.65625,0.9,0.05,1.65625,8.933333,14.293751,19.633333,24.7125,35.325005,61.216663,83.174995,63.45,42.822975,23.075003,12.73125,5.166667,2.5749998,1.3416667,0.81666666,0.60625,0.84166664,0.70000005,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.20000002,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.48333335,5.25,6.225001,1.6937499,0.0,0.0,0.0,0.5875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30625,0.0,0.0,0.10625,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.15,1.0416666,1.075,0.56875,0.23333335,0.36249998,0.041666668,0.47500002,0.7916667,1.5583335,0.70624995,1.0916667,3.4562497,5.033334,3.7000003,5.791667,10.1625,15.016667,11.366667,13.299999,7.55,4.10625,16.291668,10.2,6.0999994,13.816667,17.99375,17.558334,14.987499,11.191667,6.2625003,6.383333,6.2583337,7.90625,11.100001,22.7125,26.025,19.362501,7.175,2.3125,3.2583332,2.3083334,0.8999999,0.9,0.60625,0.35833332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333334,0.25625002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.71666664,0.8833334,1.75625,1.2583334,0.3625,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.63125,1.4749999,1.3555555,2.2444446,1.8666666,4.977778,8.633333,1.8111112,0.25000003,0.3,1.8555555,2.9,3.7000003,1.4749998,0.5111111,0.3,1.8555555,5.8583336,0.5111111,0.22222224,0.0,0.0,0.0,0.044444446,1.8,2.5555558,1.5111111,0.0,0.23333332,0.15833333,0.95555556,1.6916667,0.5555556,1.075,1.4444444,0.0,0.3166667,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19166668,0.24444446,0.65000004,1.7222223,1.9,3.075,1.8777778,5.5666656,12.044445,7.825,5.633333,7.4916663,6.3,18.688889,36.158337,23.344444,11.183333,1.8,1.025,3.1111114,4.277778,4.1499996,2.5555558,0.8083334,0.044444446,5.216667,7.0777774,6.916666,8.366668,6.588889,3.191667,4.0666666,3.4333334,2.1222222,3.716667,3.7888887,2.5555553,3.4833336,5.5444446,3.358333,2.6444447,1.3333335,0.3888889,0.15555556,0.22500001,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0666666,3.8333335,2.8416667,5.1444445,5.741667,10.48889,20.433334,20.475,13.622222,18.156818,22.2625,14.141666,2.9,0.7250001,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,1.825,0.17777778,0.0,0.0,0.0,0.09166667,0.011111111,0.0,0.18888889,0.9111112,4.566667,2.311111,0.35833332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.11666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22222222,0.5416667,0.7111112,0.82222223,1.0500002,0.33333337,0.40000004,0.14444445,0.15,0.7,0.9555555,0.46666667,0.18888889,1.7000002,2.1555557,1.9666667,2.6111112,3.0833333,4.9,13.422223,11.941667,8.155556,7.4833336,10.666667,8.633333,2.1999998,7.377778,9.616667,13.088888,16.125,19.333334,21.383335,12.777779,12.766666,12.35,14.377778,13.683333,20.911112,14.033333,6.8222227,2.7666671,3.6333334,3.088889,2.8333337,2.977778,0.61666673,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.0,0.33333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777778,0.6333333,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.35,4.0583334,6.3916664,2.18125,1.6916666,2.10625,0.975,0.7250001,0.6166667,0.7916667,6.8124995,7.9,4.2062507,0.38333336,0.0375,0.25,3.0374997,0.7750001,0.08333334,0.0,0.34166667,1.275,2.9083333,1.55,3.608333,3.9916668,0.6937501,0.48333335,1.2,3.6,0.79375005,0.18333334,1.29375,3.6000001,0.55,0.51875,1.6083333,0.9125,0.0,0.0,0.0,0.0,0.0,0.16666667,2.0125,0.083333336,0.14375,1.0916666,2.641667,3.5625,3.8500004,6.61875,12.45,12.549999,6.316667,6.5687504,7.7250004,39.216667,32.28125,14.283333,3.3125002,0.675,0.1,0.71666676,2.983333,4.8250003,2.4499998,1.2624998,0.9499999,3.0875,4.4,4.9125,5.0250006,7.008333,6.3625,4.7083335,4.46875,3.3083336,2.3999996,1.6583335,1.1833334,0.61875,0.041666668,1.33125,2.3333333,1.1687499,2.3500001,4.125,2.76875,0.5666666,0.0375,0.0,0.0,0.2,0.50000006,0.53333336,0.0,0.10625,0.48333335,1.8625,4.6,17.725002,27.10682,27.60394,23.543749,30.94167,34.968746,39.61333,24.899998,3.1083336,1.85,1.4166666,0.98333335,0.5875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2083334,0.54375,0.0,0.0,0.0,0.041666668,0.25625002,0.13333334,0.5125,1.0250001,1.5666666,2.45,0.7750001,0.075,0.16666667,0.55625004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14166668,0.2,0.33750004,0.725,0.50625,0.5,1.0625,1.2500002,0.41666666,0.38124996,0.49166667,0.86875,0.71666664,1.0750002,1.1916667,0.43125,2.5583334,7.2166667,5.7687497,7.2333336,10.5,7.9749994,3.18125,0.95,2.8916667,3.7062502,5.516667,12.437499,16.675,17.075,16.533333,19.575,15.793751,11.658334,5.14375,4.8083334,5.5,3.8083332,5.69375,2.6833334,3.1916668,1.5999999,0.6583334,0.04375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.49999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.55625,2.9,1.75,0.5625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.0833333,6.022222,10.077778,6.3999996,3.9777777,1.3000001,1.9111112,5.158334,2.6666665,1.1444443,4.6916666,9.622222,2.6999998,0.72222227,0.0,0.0,0.5,1.3111112,0.7777778,0.0,0.6111111,10.200001,10.788889,2.9333334,5.4222226,4.6666665,2.6583333,0.86666656,2.0083334,0.78888893,0.0,0.0,7.7,4.4222217,2.211111,1.0916667,2.0777779,0.7666667,0.0,0.0,0.0,0.0,0.050000004,0.43333334,1.3833333,0.05555556,0.20000002,1.3666668,3.066667,3.8416665,6.166667,6.6999993,6.7000003,10.058334,8.033334,13.625,27.144444,28.51111,20.508331,16.422222,17.775,7.0666666,5.6916666,8.177778,2.388889,7.158333,5.211111,3.6666667,1.9444444,1.5500001,2.1111112,4.3250003,4.566667,4.7000003,6.158334,5.8999996,4.3250003,3.9555557,2.9833333,1.5444446,0.43333334,0.0,0.0,0.65,1.5999999,3.2833335,10.800001,10.677778,4.4916663,1.4,0.05,0.0,0.525,1.5777779,0.06666667,0.0,0.0,0.6916667,3.2222223,2.0416667,6.866666,25.758333,35.09722,27.353016,48.825005,47.117065,60.433327,52.755558,21.816668,4.4888887,3.5083332,2.988889,3.2444444,3.25,1.0111111,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35833335,0.0,0.0,0.0,0.0,0.0,0.23333333,0.15833333,0.43333334,0.85833335,1.1222222,0.7111111,0.5166666,0.15555556,0.0,1.0444444,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12222222,0.31111112,0.0,0.0,0.1,0.17777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.3111111,0.18888889,0.56666666,0.9444444,0.60833335,1.1777778,1.7333333,1.4777777,0.23333333,0.19166669,0.87777776,1.225,0.7111111,0.375,0.36666667,0.06666667,1.0777777,1.0,1.3833334,3.711111,6.4000006,10.455556,13.641668,4.5222225,0.3555556,1.9416668,1.2555557,4.575,7.4111114,9.324999,16.4,16.88889,15.55,14.48889,11.483334,11.477777,10.941666,9.488889,8.716667,1.7222223,3.6333332,1.425,0.044444446,0.0,0.0,0.05,0.0,0.11111111,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,3.4,3.4777777,1.2166667,0.0,2.8249998,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31666666,4.0555553,6.711111,9.908333,8.5222225,3.3333333,0.53333336,4.825,6.577778,4.544444,4.258333,4.066667,0.26666668,0.0,0.19999999,0.24444444,5.0250006,6.5444446,4.1444445,4.225,4.4666667,7.325001,5.6555557,2.15,3.2000003,4.0,3.1833334,1.7777779,1.2666667,0.13333334,0.3,1.0444446,8.908334,4.8111115,2.0222223,0.34166667,0.41111112,0.0,0.0,0.0,0.0,0.0,0.15,1.2666668,1.2916666,1.1666667,1.2416667,2.511111,4.2333336,3.8333335,3.988889,7.2333336,5.7,5.0416665,7.6222215,18.325,23.444445,12.355556,17.983334,21.900002,41.48333,35.833336,24.458334,31.288889,12.1444435,6.4833336,8.344444,11.816668,13.4,7.3333335,3.1555557,3.7250004,5.266667,5.366667,4.508333,5.0111113,3.9166667,2.5222225,2.2916667,1.5222223,0.37777779,0.033333335,0.7111111,1.0833334,1.2333335,2.2583334,6.8111115,6.022222,1.8833332,0.7555556,0.0,0.93333334,1.4,0.51111114,0.1,0.14444445,2.6555557,15.641667,32.844444,27.699997,23.825,27.516668,40.03472,44.743053,49.4,49.444447,27.591667,18.055557,4.7166667,0.7777778,0.84166676,0.5222223,0.23333333,0.40833333,0.58888894,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333332,0.06666667,0.33333334,0.0,0.0,0.0,0.0,0.33333334,0.050000004,0.32222223,0.43333334,0.5333333,0.22222222,0.0,0.0,0.15833333,0.8444444,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1777778,0.51111114,0.0,0.0,0.4416666,0.36666667,0.0,0.08888889,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.05,0.022222223,0.57500005,1.4111112,0.5555556,0.425,1.1666669,0.9083333,0.43333334,0.9916667,1.3666667,0.23333333,0.033333335,0.17777778,0.36666667,0.4,0.3,0.3111111,0.041666668,0.3222222,0.3,0.25000003,0.95555556,2.8249998,6.3777776,19.191668,12.466665,3.4777777,0.16666667,0.32222223,2.0333333,3.5777776,3.8250003,7.433334,5.8999996,6.108333,9.422222,11.333334,15.055555,14.450001,7.577778,6.1166663,2.3777778,0.7,0.23333335,0.022222223,0.0,0.0,0.0,0.0,0.11111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,1.2,0.9083333,1.1777778,0.275,0.18888889,0.25833333,0.0,0.0,0.025,0.0,0.0,0.0,0.0,1.1562501,1.0,1.0,8.0375,14.991666,15.074999,1.8833333,0.5,4.016667,7.225,8.325001,6.8583336,3.7875001,0.008333334,0.3,1.7416668,11.687498,8.224999,6.091666,6.2999997,4.8250003,0.8812501,1.0916666,0.25,1.4083333,1.7083334,0.3125,0.0,0.10000001,0.25,0.6875,1.7833335,4.5,3.2916667,1.3083334,0.325,0.15833335,0.0,0.0,0.01875,0.18333334,0.44166666,1.85625,2.875,5.025,6.3083334,3.04375,2.4750001,2.991667,2.84375,3.5916665,4.09375,3.3333335,2.3812501,5.766667,16.15,19.85,28.008335,26.2,42.800003,40.356247,32.625,19.143751,9.641666,5.9666667,8.231251,10.891665,15.31875,20.45,19.48125,8.633333,5.3999996,4.458334,4.225,3.71875,2.8916667,2.75625,2.3999999,1.275,0.6750001,0.19166666,0.0,0.35000002,0.72499996,1.05,0.8375001,2.95,5.3666663,3.7937498,1.1916667,0.0625,0.0,0.31875,0.9916667,1.3874999,14.666668,32.475,45.225006,48.983334,45.4,42.71667,27.575003,25.258333,22.683334,17.956251,11.441667,4.05,2.8583333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.15625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43333334,0.0125,0.06666667,0.118750006,0.125,0.033333335,0.0,0.0,0.23124999,0.35833332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.081250004,0.10833334,0.43124998,0.35,0.20833334,0.22500001,0.033333335,0.05,0.083333336,0.0125,0.20833336,0.26250002,0.28333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.025,0.016666668,0.00625,0.0,0.0,0.0,0.0,0.15625,0.9916667,0.25,0.53333336,0.93750006,2.016667,0.8499999,1.325,1.0833334,1.13125,0.9916667,0.45000002,0.8833334,0.025,0.0,0.0,0.0125,0.058333337,0.14375,0.09166667,0.0625,0.40833333,0.125,0.0125,0.06666667,1.0374999,2.733333,7.2124996,6.3583336,2.0333333,2.25625,1.4166667,4.36875,5.7166667,2.6125,4.225,6.0333333,4.83125,3.4583335,7.668751,11.808334,8.606251,0.7916666,0.24375,0.15,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6583334,0.825,1.9124999,1.1750001,0.79375005,0.53333336,0.28750002,0.5833334,0.45833334,0.3,0.13333334,0.06875001,0.0,0.0,3.7166665,2.2444446,0.3888889,3.275,5.122222,5.766667,1.8222224,1.6416667,5.211111,17.544445,28.158335,29.944445,19.400002,9.133333,2.2,6.077778,9.625,9.255555,7.9666667,8.666666,5.5111113,1.5749999,0.055555556,5.7749996,7.933334,3.7555556,0.9583334,0.9333334,0.51666665,0.0,0.79166675,1.0333333,3.1333332,3.1222224,1.7666668,0.2916667,0.0,0.0,0.0,1.0916667,0.9666667,2.1777778,3.025,4.3111115,7.008333,6.122222,2.4333332,1.888889,3.1000001,1.875,0.9666666,2.125,1.5777777,6.941667,11.755555,42.15,67.53333,63.800003,52.233334,48.54445,24.366669,10.533334,6.0916667,1.5666666,1.1333334,3.1083336,9.733334,15.55,20.244446,18.633335,18.366667,10.25,5.5444446,3.9666667,2.4833333,1.7111112,0.8416666,1.1111112,0.7916667,0.9555556,1.0,0.6916667,0.4,0.17500001,1.2444446,2.0083334,4.4666667,7.455556,3.8333335,1.388889,1.05,0.56666666,1.3833333,1.588889,5.4999995,30.77778,44.45556,35.241665,21.977777,16.55,12.4777775,5.016667,4.511111,3.1444445,0.7416667,0.2888889,0.008333334,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.08888889,0.0,0.033333335,0.05,0.0,0.0,0.0,0.0,0.0,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,2.7583334,2.6222222,5.3444443,1.325,0.0,0.0,0.2888889,0.67499995,0.3111111,0.125,0.22222224,0.022222223,0.008333334,0.0,0.025,0.033333335,0.15833333,0.08888889,0.022222223,0.083333336,0.044444446,0.275,0.23333333,0.16666667,0.08888889,0.13333334,0.09166667,0.07777778,0.75,0.6111112,0.033333335,0.17777778,0.9416666,2.0666668,0.7,0.875,0.6888889,1.1583333,1.5666667,0.48333335,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.325,0.54444444,0.47777775,0.041666668,0.0,0.36666667,1.4666667,3.6166663,7.5000005,4.033334,1.4083334,1.9222223,1.1166667,3.488889,2.1583333,0.0,0.90000004,1.2916667,0.53333336,3.5416665,12.166666,13.000001,7.5222225,3.9416668,3.711111,2.6777778,1.3,1.2444445,0.9583333,0.70000005,0.35000002,0.07777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.77500004,0.36666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,1.0333333,2.0222223,1.6916667,0.08888889,0.0,0.0,0.125,0.5222223,0.22222224,0.016666668,0.022222223,0.050000004,0.0,0.2,5.8125,4.2250004,3.0333333,3.01875,3.4916668,3.6812503,3.291667,2.5125003,2.1583333,2.3416667,2.85,3.675,4.9437504,7.033334,16.675001,26.333334,24.525,17.949999,15.483333,13.368751,12.291667,8.79375,6.208334,7.3187494,7.408334,5.6166673,2.35,0.96666664,0.4125,0.16666667,0.46249998,1.3000001,2.16875,0.95000005,0.6,0.17500001,0.05,0.48749998,0.1,0.10000001,0.14166667,0.5833334,4.25,5.6833334,4.5624995,2.8749998,1.8937501,2.075,1.75,1.7062498,1.0333334,2.4125,5.191667,8.006249,24.333332,50.381252,54.333336,50.43334,42.41875,36.600002,29.8875,18.575003,11.95625,7.6833334,2.4583335,2.03125,3.8833334,9.200001,11.5,12.268749,12.741667,9.63125,3.491667,2.8833332,2.90625,0.56666666,0.40625,0.058333337,0.125,0.38333333,1.2750001,1.11875,0.26666668,0.05625,0.725,1.8500003,4.65,5.891667,3.3749998,1.525,0.36874998,0.95833325,1.2625003,1.6833335,8.65,20.299997,27.275,15.55,4.7833333,3.1750002,2.2333333,1.1687499,1.0833333,0.35833335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.075,0.025,0.0,0.18124999,0.125,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.4,3.6583338,7.716667,1.475,0.05,0.6374999,2.0083332,1.20625,0.6750001,0.54375,0.20833334,0.15833335,0.1125,0.083333336,0.29375,1.3666667,1.3375,0.25,0.40833333,0.51875,0.39166668,0.7624999,0.61666673,0.3875,0.34166667,0.47500002,0.35,0.27499998,0.30625,0.16666669,0.125,0.7,1.15,0.6333333,0.26666668,0.65000004,0.075,0.6625,0.62499994,0.26875,0.09166667,0.16666667,0.0,0.30833334,0.33125,0.0,0.0,0.0,0.2,0.041666668,0.0,0.0,0.0,0.0375,0.625,3.1000001,8.225,10.099999,1.2,0.94166666,3.0625002,7.0416665,5.83125,1.3333331,0.13333334,0.9812499,2.0,3.7125,7.2000003,11.300001,12.5,14.174999,17.166668,13.483333,5.84375,3.3999996,1.9562498,1.2416667,0.66875005,0.14166668,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.11666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.41666666,0.4625,0.0,0.82500005,2.0666666,2.4583335,4.3250003,1.0500001,0.05,0.0,0.22500001,0.45833334,0.2916667,0.21875001,0.0,0.0,0.0,0.0375,4.5333333,3.5111113,2.6888888,2.4583335,1.388889,1.775,2.211111,2.075,2.3666668,3.6777778,2.4416666,4.1666665,6.208334,10.4,19.741667,34.82222,39.050003,30.98889,27.300001,24.21667,19.066668,14.433334,6.8222227,3.2416668,2.577778,0.9666667,0.60833335,0.84444445,0.9083334,0.5888889,0.15833333,0.31111112,0.9499999,0.4888889,0.51111114,0.625,1.1,0.7583334,0.36666667,0.06666667,0.0,4.6555557,8.091665,8.700001,6.458334,2.8444445,2.5333333,1.7222223,0.5222223,0.14166667,0.6666667,3.2916665,5.2555556,11.675001,19.622223,21.791668,21.200003,20.944447,17.025002,24.755554,27.44167,13.077778,10.125001,8.5222225,3.611111,2.3583333,4.2444444,4.4666667,4.7000003,5.116667,4.922222,2.9666667,1.0555556,0.42222223,0.22500001,0.65555555,0.15833333,0.07777778,0.025,0.0,0.022222223,0.33333334,1.9444444,1.2333333,0.2111111,0.5083333,3.777778,4.0666666,1.8833333,0.07777778,0.0,0.0,0.49166664,1.8666668,4.3166666,9.0,6.2888894,3.2166667,0.32222223,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.0,0.53333336,0.23333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.2166667,15.777777,10.122223,0.058333334,0.35555556,0.8083333,0.7111112,0.46666667,0.47777778,0.6166667,0.2777778,0.2888889,0.15833335,0.6444445,0.89166665,1.7888889,0.68333334,0.45555556,1.5777779,1.4083333,1.2111112,0.9250001,0.8333334,0.6666667,0.8555556,0.62222224,0.4416667,0.3888889,0.40833336,0.6111111,1.6666666,1.0888889,0.5083333,0.13333334,0.0,0.0,0.17777778,0.13333334,0.2,0.17500001,0.044444446,0.011111111,0.0,0.6111111,0.3,0.0,0.0,0.0,0.18333335,0.055555556,0.0,0.0,0.0,0.25,0.13333334,0.39166665,4.011111,7.8555555,4.55,4.1000004,3.1916666,7.2111115,6.808333,2.6666667,1.7333332,0.31666666,0.0,0.06666667,0.15555556,1.0416667,4.4555554,11.091667,22.166668,21.97778,14.258333,7.666667,2.875,0.47777778,0.083333336,0.06666667,0.022222223,0.0,0.0,0.0,0.0,0.0,0.011111111,0.36666667,0.7,0.5222222,0.40000004,0.4888889,0.47500002,0.36666667,0.2916667,0.16666667,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.325,0.10000001,0.45833334,1.8111113,2.5000002,1.6777779,1.4888889,1.2,0.5555555,0.0,0.0,0.0,11.8625,6.5166664,4.166667,4.54375,5.8333335,6.3875,6.083333,7.3812504,7.183334,8.808334,10.362501,10.083334,10.087501,11.425,14.25625,12.35,13.11875,12.475,15.199999,19.21875,16.8,9.15625,4.641667,1.9187502,1.4000001,0.6333333,0.53125,0.29166666,0.24375,0.79166675,0.75000006,0.41666666,0.38750002,0.625,1.125,1.9875,2.1333334,1.53125,0.25,0.10625001,1.0666667,1.9583334,4.01875,5.266667,3.8375,3.6416667,2.6062498,0.26666665,0.15833333,1.15625,4.708334,3.7937503,4.05,6.35625,9.033334,9.062501,8.483334,5.925,5.4812503,11.900001,14.3,21.775,19.125,13.175001,5.5416665,2.5125,0.9666667,0.99375,0.97499996,1.09375,1.0416666,0.41875,0.13333333,0.44166666,1.7687502,1.9833332,1.1125,0.45,0.01875,0.0,0.033333335,0.087500006,0.43333337,0.59375,0.36666667,0.087500006,0.20833334,0.85,0.58750004,0.78333336,0.23125,0.0,0.05,1.2333333,4.2562494,5.4500003,0.3166667,0.38125002,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,1.0187501,1.1833334,0.6125,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.325,4.5666666,3.516667,0.23125,0.116666675,0.54375,0.425,0.53125006,0.70000005,0.56250006,0.425,0.30833337,0.6375,1.2166667,0.8375,0.8666666,0.375,0.8000001,1.5750002,1.89375,1.1666667,0.80625,0.725,0.99375004,0.8416667,0.69166666,0.80625004,1.9166667,2.3249998,3.266667,3.03125,0.875,0.5500001,0.3416667,0.0,0.0,0.0,0.0125,0.008333334,0.0125,0.008333334,0.0,0.0,0.21666667,0.26250002,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.17500001,0.9,0.9166666,1.8083334,3.00625,2.8666666,3.90625,6.266667,3.25625,2.1,2.1999998,1.3125,0.60833335,0.17500001,0.15000002,0.8812499,1.3583332,3.2749999,7.3916664,9.525001,9.3125,7.1083336,5.05625,3.9250002,2.15625,0.8666667,0.6666667,0.9625001,1.1333333,1.4250001,1.15,0.5625,0.73333335,0.58124995,0.18333334,0.025,0.28125,1.0749999,0.3625,0.041666668,0.21875,0.175,0.09166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.31875,0.9583334,1.03125,2.4250002,2.9812503,3.1000004,3.4916668,2.5562503,0.90000004,0.32500002,0.041666668,0.0,20.133333,20.666668,17.322224,9.933333,7.644444,7.4666677,8.822223,10.416667,8.088889,7.888889,8.550001,8.8,7.45,6.3777785,5.8583336,4.455556,3.5166671,3.666667,6.1444445,9.558333,8.044444,2.8166666,2.0888891,3.9333334,3.4333334,4.4666667,6.3,7.2111115,5.558333,4.766667,2.7833333,1.4888889,1.475,1.188889,0.11111111,0.2,0.0,0.0,0.0,0.016666668,0.044444446,0.76666665,2.65,4.3555555,3.6916666,1.4111111,0.39166665,0.6555556,3.3111112,6.2833333,9.622221,12.141666,4.666667,1.0333334,2.0333333,5.383333,8.255556,7.722222,11.266666,17.422222,15.883333,31.011112,29.458332,17.233335,10.211112,7.133334,1.2555556,0.7916667,0.0,0.008333334,0.0,0.7083334,1.2888889,1.5444444,1.8916667,1.3444445,1.65,1.0,0.0,0.22222222,0.22222222,0.25,1.1888889,0.8666667,0.41111112,0.33333334,0.31111112,0.8333334,1.125,1.7111113,1.225,0.0,0.48333335,2.4444444,1.6250001,1.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.3333333,0.07777777,1.5333334,0.34444445,0.0,0.0,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.20833334,0.12222222,0.16666667,0.0,0.11111111,1.1833334,1.0666667,0.7916666,1.5111111,0.5833333,0.6,0.8333334,1.5833334,1.0111111,0.87500006,0.5777778,1.95,2.1333334,1.9111112,1.5083333,0.88888884,0.975,1.2333333,1.4416666,1.3666667,0.94444454,2.175,5.666667,5.825001,6.2777777,4.8416667,2.3666666,0.825,0.41111115,0.6,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.28333336,0.7111112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3333333,0.0,0.0,0.0,0.033333335,1.2,1.225,0.5555556,0.24166667,0.3,0.65555555,0.525,0.5555556,0.39166665,0.033333335,0.13333334,0.32222223,0.8833333,3.7999997,4.5222216,4.8916664,4.066667,2.8500001,3.0666666,3.3416667,2.2666667,1.1333334,0.35833335,0.35555556,0.53333336,1.2444445,2.275,2.7222223,1.6916668,0.36666667,0.3888889,0.675,1.5111113,2.025,0.4888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.20000002,1.5749999,4.3333335,4.7666664,4.3888893,3.8555558,2.9333334,0.77777785,0.575,0.32222223,0.14999999,9.1,15.811111,9.033334,9.425,7.7333336,5.408334,5.466667,5.55,3.7444446,4.0333333,4.275,4.711111,3.6750002,3.3333335,3.816667,3.8333333,4.6000004,9.111113,15.911112,22.35,15.477777,8.875001,9.944444,11.174999,11.222222,11.933334,9.375,6.133333,3.7666671,2.1222222,0.70000005,0.20000002,0.26666665,0.21111111,0.0,0.0,0.0,0.0,0.044444446,0.09166667,0.62222224,1.0555556,1.1416667,2.1999998,2.2083333,2.6222222,3.2333333,5.7000003,8.677778,9.516666,8.711111,7.625,5.6555557,6.1916666,12.900001,21.45,23.122223,18.533333,16.533333,14.933334,13.958334,26.388887,34.358334,24.177776,16.699999,10.658334,3.477778,4.791667,0.13333334,0.0,0.0,0.16666667,1.1777779,1.2444445,2.0916667,1.4555556,0.625,0.15555556,0.0,0.44444445,0.6666667,0.5833334,0.5555556,0.69166666,0.12222223,0.98333335,3.0444443,3.1222224,4.0583334,3.1333334,0.425,0.0,0.65000004,0.9333334,1.1416667,0.70000005,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17777778,1.125,0.73333335,0.0,0.75555557,0.6666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.025,0.0,0.2,0.0,0.22222222,1.5916666,1.0666667,1.475,0.8555556,0.61666673,0.5555555,1.7777779,1.6166667,1.2222222,0.925,2.1111112,2.6166666,2.966667,1.8555558,1.5333334,1.3444445,1.2500001,1.5222223,1.8083334,1.4888889,2.2333336,5.2,7.622222,8.091667,7.811111,3.7000003,1.2888889,0.40833336,0.022222223,0.78888893,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43333337,3.2888892,3.8222225,4.6,5.8555555,5.891667,6.0111117,6.766667,5.911112,4.6444445,3.1416667,2.8777778,3.241667,3.888889,4.4833336,4.6222224,3.5833335,1.8333334,1.7444447,1.2500001,1.0333333,2.1583333,1.3111112,0.14166668,0.08888889,0.0,0.0,0.0,0.35,0.5888889,0.14166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15555555,0.7083334,3.1111112,4.1833334,3.4222221,2.6444447,0.68333334,0.16666667,0.5083333,0.4111111,0.29999998,5.6249995,5.633333,3.55,4.2375,2.7416666,1.2312502,1.3250002,1.125,1.0166667,1.1,0.38750002,0.29166663,0.38125002,0.5666667,0.97499996,1.6999999,2.6875,3.641667,5.591667,6.8687506,6.566667,6.00625,6.991667,8.23125,7.975,6.5916667,3.58125,1.4916667,0.4,0.55833334,1.26875,0.9166667,0.106249996,0.0,0.0,0.0,0.058333334,0.56875,0.76666665,0.50624996,0.21666667,0.06666667,0.8125,3.891667,4.5437503,3.008333,2.3750005,3.8999999,4.4333334,4.88125,10.783332,15.950002,18.425001,22.33125,25.525002,19.900002,17.541668,13.433334,10.5625,8.95,10.349999,14.45,25.725,25.716667,17.883335,9.95625,6.5583344,1.4625,0.05,0.0,0.0,0.0,0.18333334,0.275,0.375,0.083333336,0.20625,0.0,0.0,0.0,0.0,0.0,0.06666667,0.33749998,0.34166667,0.21875,0.6916667,0.6916667,1.2,0.875,1.3562498,0.77500004,0.66875,0.5833334,0.775,1.2666668,0.65,0.275,0.0,0.24375,0.9166667,0.25,0.33333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.21666667,0.31666666,0.0,0.0,0.0,0.0,0.15625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20625,0.85530305,0.17500001,0.0,0.0,0.0375,0.9416667,1.4562501,1.2916666,1.4625,1.125,0.8000001,1.0083333,2.6083333,1.59375,1.4,2.9875002,3.8583338,3.5625,1.5416667,1.5916667,1.63125,1.4916666,1.475,1.7583334,2.275,3.6499996,4.3166666,4.71875,5.5249996,5.6937494,4.766667,2.60625,0.55833334,0.118750006,0.05,0.11666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.1,0.52500004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40000004,0.0,0.0,0.0,0.0,0.5625,0.5333333,0.0,0.0,0.112500004,1.5166667,1.6166668,2.25,3.2000005,3.9000003,5.2000003,6.1000004,5.0750003,3.9750001,3.2375002,2.516667,0.89375,0.925,4.1000004,7.491667,8.40625,7.1083336,5.633333,6.7875004,6.9166665,6.6937504,3.7250001,3.8312502,2.7666664,1.2583333,0.87500006,0.875,0.25625,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.725,1.7062502,1.6166668,1.0999999,0.3,0.0,0.29999998,0.35000002,0.41875002,9.258333,8.4,5.811111,6.208333,7.911112,3.2749999,2.3111112,1.1166667,1.0555556,1.0222222,0.26666668,0.23333335,0.3166667,0.3888889,1.0,1.3555554,1.8833334,2.2555559,3.3222222,4.833333,5.1222224,3.1000001,2.5888886,1.0749999,0.6888889,0.29999998,0.20833334,0.22222224,0.28333333,0.8333334,1.4999999,0.75555557,0.0,0.011111111,0.35555556,1.7583334,1.4444443,0.35,0.15555555,0.0,0.0,0.011111111,0.7833334,1.5999999,1.6166667,0.29999998,0.17500001,7.3333335,10.788889,8.333334,8.322222,9.266667,8.066667,8.241667,6.7555556,5.8916664,5.433334,5.2111115,5.8,7.255555,9.2,12.833333,18.408333,18.722221,13.5222225,7.566667,5.8333335,0.92499995,0.0,0.0,0.0,0.0,0.0,0.16666667,0.0,0.0,0.0,0.11111112,0.05,0.13333334,0.11111111,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.9666667,0.9416666,0.8777778,0.48333332,0.19999999,0.76666665,0.0,0.0,0.0,0.5888889,0.675,1.3,1.9416666,3.8444448,3.4222224,1.5250001,0.7111111,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14444445,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.75,0.7222222,0.0,0.0,0.0,0.40833333,1.6888888,1.3500001,2.5555558,1.875,1.4444445,1.4916667,2.0,2.611111,1.7583332,3.0777779,4.6833334,4.4666667,2.525,2.2555556,2.0222223,0.9833334,2.3888888,2.3999999,3.2555556,4.558333,4.9777775,4.3333335,4.4750004,4.611111,3.0083332,2.688889,0.92,0.35555556,0.1507576,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,0.44444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.075,1.2777779,0.0,0.0,0.0,0.0,0.0,0.050000004,0.23333332,0.15833333,1.3222222,2.4666662,2.6555552,2.6333332,3.1416664,3.2444448,2.2166667,1.8555555,2.8333335,5.7555556,7.15,6.711112,6.900001,11.3,13.322223,12.158334,8.800001,8.225,5.8444448,3.7777777,3.0333333,3.1666665,2.05,0.25555557,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22222222,1.8416667,2.2444444,0.85555553,0.6166666,0.25555554,0.7333334,0.8000001,1.6666667,13.025001,14.658333,16.866667,15.643751,14.200001,10.85625,10.008334,8.30625,10.258334,10.641667,11.606251,8.133333,8.93125,4.2,2.5874999,0.5,0.3,0.26666668,1.0583334,2.4,5.083334,7.10625,7.2750006,6.7249994,5.683334,4.7500005,2.8687503,1.9,1.21875,0.8333334,2.0875,3.0666666,1.7874999,0.825,0.82500005,1.18125,0.24166667,0.0,0.0,0.0,0.0,0.016666668,0.087500006,0.14166668,0.08125001,0.0,0.89375,3.3416667,3.1749997,2.08125,1.0583333,0.43125004,0.69166666,0.9,1.2,1.96875,2.7833333,3.6166668,4.86875,5.8583336,8.9375,12.9,13.656252,9.625,6.333333,3.0125,1.9583333,0.55625004,0.15,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.35,0.0375,0.0,0.0,0.375,6.666667,4.8750005,0.0,0.0,0.0,0.16666667,0.48125,0.70000005,1.1937499,0.975,1.2562499,1.3916667,0.60625,0.6916667,0.7333334,1.475,4.6083336,3.8187504,3.241667,2.5937498,1.3416667,1.0583333,0.8312501,1.0250001,1.06875,0.8000001,0.88124996,0.7,0.45,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06875,0.083333336,0.075,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.025,0.0,0.0,0.15,0.775,0.13333334,0.0,0.0,0.14166667,0.7875,1.1166668,1.4625001,2.9166665,2.6625001,2.7583332,2.875,3.0749998,2.0916667,2.4624999,3.575,4.2437496,5.166667,4.8312507,3.883333,3.6033332,2.0125,2.937879,4.65625,6.166667,5.83125,5.0833335,5.658333,5.625,3.525,2.8125,2.709091,1.9875,0.33000004,0.04375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06875,0.12500001,0.0,0.00625,0.1,0.00625,0.0,0.0,0.0,0.0,0.15,0.5833333,0.0,0.13333334,0.55,0.0,0.0,0.0,0.0,0.675,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.65833324,1.3875,1.3750001,1.7500001,2.5437503,1.7666667,1.63125,3.1916666,4.425,4.516667,5.08125,8.933333,11.974999,9.962501,8.691667,8.56875,5.683333,4.8375,4.366667,3.3333333,4.0249996,3.1499999,0.6062499,0.075,0.06875,0.2,0.15,0.0,0.083333336,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28750002,0.925,0.7916666,0.78125,0.26666668,0.75625,0.5916667,1.4000001,22.016665,21.977777,25.222221,26.216667,21.233334,20.241667,19.866667,15.491668,15.2,17.677776,17.05,10.5222225,11.791666,3.9333332,4.191666,1.6333334,0.0,0.011111111,0.011111111,0.6916667,2.711111,4.5250006,4.277777,3.1666665,3.711111,3.7444444,2.9916666,2.2666667,1.9083332,1.6777779,1.1416667,0.66666675,0.06666667,0.1777778,0.033333335,0.0,0.25555557,0.25,0.11111112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10833334,0.13333334,0.15555556,0.075,0.0,0.0,0.033333335,0.06666667,0.12222223,0.44166666,0.8000001,1.2888889,2.0833335,2.6,3.7000003,4.166667,2.4833336,1.0,1.0666666,0.35833335,0.3,0.05,0.0,0.39999998,0.4888889,0.0,0.0,0.0,0.0,0.0,0.008333334,0.21111111,0.15,0.17777778,0.0,2.733333,19.811111,16.441666,2.3000002,0.89166665,0.5333333,0.54444444,0.65,0.5,0.525,0.36666667,0.15833333,0.0,0.7166667,2.4444444,3.677778,6.7,14.51111,9.391666,5.8444443,5.8666663,5.722222,5.1,3.8333335,2.2222223,1.3583333,1.1555556,0.28333333,0.0,0.26666668,0.70000005,0.21111113,0.0,0.0,0.0,0.0,0.0,0.35555556,0.6,0.25,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.2888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.0,0.0,0.016666668,0.54444444,0.5,0.23333332,0.15833333,0.11111111,0.41111112,0.625,1.7444444,2.75,3.2333333,2.2666664,3.0333333,2.9166665,0.75555557,1.6999999,5.8250003,3.9444444,4.9500003,5.666667,8.400001,6.0222216,3.577778,3.5083334,5.6777773,7.233333,7.377778,6.708334,7.066667,5.722223,4.7083335,3.766667,4.9666667,5.7,3.4416666,0.43333334,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.05,0.022222223,0.0,0.0,0.033333335,0.022222223,0.0,0.016666668,0.13333334,0.016666668,0.0,0.016666668,0.044444446,0.0,0.0,0.044444446,0.016666668,0.06666667,2.2166667,1.111111,0.11111111,0.13333334,0.3777778,1.0666666,0.6666667,0.09166667,0.0,0.0,0.0,0.0,0.0,0.06666667,0.1,0.7444444,1.8166667,2.1444445,2.488889,2.8666668,2.2666667,1.5083334,1.6111112,3.1166668,5.111111,5.5,5.3666673,4.888889,5.5249996,6.4000006,8.233334,8.611111,5.6250005,7.233334,8.655556,7.0166664,3.6444445,1.3499999,0.25555554,0.30833334,0.37777779,0.083333336,0.16666667,0.19999999,0.39166665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.5888889,2.1166668,2.0666666,0.9333333,0.6,0.89166665,18.3375,20.158333,25.883333,25.28125,24.008333,19.24375,16.766668,12.19375,9.616666,8.358334,6.6062503,6.683334,3.60625,0.60833335,0.0375,0.008333334,0.0125,0.0,0.0,0.03125,0.20833333,0.66875005,0.7833333,0.39999998,0.91666657,1.125,2.975,4.833333,3.7,2.65,2.2375002,1.6083333,0.50625,0.725,1.1416667,0.94375,0.4416667,0.0625,0.10833334,0.21875,0.025000002,0.06666667,0.06875,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.225,0.59999996,0.95625013,1.4499999,3.341667,2.7437499,0.7750001,1.23125,2.1000001,2.0625,1.6,0.8833334,0.5125,0.5083334,0.7625,0.4416667,0.3375,0.24166667,0.081250004,0.0,0.0,0.0,0.0,0.09375001,0.3083333,0.33124998,0.44166672,2.975,6.05625,5.633333,4.1250005,2.2416666,1.8125,4.35,3.8083332,2.75,2.9333334,1.48125,0.51666665,0.25625002,0.45833337,2.9250002,9.025,7.2833333,8.71875,15.908333,13.950001,9.933334,9.018749,9.516666,9.949999,11.937499,11.533334,7.0875006,3.225,2.2125,1.2166667,1.44375,0.24166667,0.06666667,0.0,0.0,0.075,0.52500004,1.6250002,1.175,0.23333335,0.0125,0.016666668,0.0,0.0,0.0,0.0,0.0,0.025,0.24166667,1.0562501,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18333334,0.05,0.0,0.0,0.23125002,0.89166677,0.57500005,0.9250001,1.3624998,2.9166667,2.5333335,3.85625,4.1583333,4.78125,4.8333335,3.8500004,3.1666667,3.21875,2.7083333,4.883333,8.243751,12.691666,12.900001,10.791667,10.15625,7.875,4.116667,4.9625006,6.3833337,7.75,9.008333,8.3125,6.0,5.125,4.4625,4.625,4.0062504,3.75,3.3125,1.5916667,0.60625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41250002,0.38333333,0.3375,0.083333336,0.0,0.0,0.14374998,0.033333335,0.0,0.20625001,0.083333336,0.0,0.0,0.4375,0.5500001,0.325,0.075,0.24166667,0.03125,0.0,0.0,0.0,0.025000002,0.23124999,0.10000001,0.0375,0.0,0.0,0.0,0.0,0.016666668,0.375,0.58125,1.4499999,2.2624998,3.25,4.66875,5.2916665,5.908334,7.018749,4.625,2.4562502,1.6500001,2.2625003,3.15,3.0312502,3.7416668,4.133333,3.4999998,2.9916668,3.9125,3.0416665,4.05,6.7083335,6.558333,6.1125,4.0416665,1.5312501,0.30833334,0.35625002,0.40833336,0.17500001,0.0,0.125,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.1,0.68125004,2.0,1.5222223,3.411111,4.7749996,5.788889,6.55,8.166666,8.225,6.8444448,5.5,6.0000005,3.488889,2.5749998,2.8333333,2.45,2.1222224,2.3416667,2.0777776,1.4555557,1.3916668,1.3888888,1.1333333,2.0222223,1.9250001,3.9666667,5.6888885,6.7833333,8.055555,10.608334,8.844444,5.850001,4.6777782,2.0833333,2.1555557,2.1666665,1.6666666,2.6777775,3.2333336,1.6666667,1.625,0.73333335,0.8888889,0.30833334,0.10000001,0.0,0.0,0.0,0.044444446,0.23333332,1.4333334,3.4777777,5.1,2.4444447,2.3,4.4888887,10.366667,17.533335,21.088888,16.350002,7.0,6.8250003,6.8444443,7.625,6.622223,5.1000004,4.05,4.844445,4.0250006,2.4666667,2.5166667,1.6111112,0.37500003,0.011111111,0.0,0.0,0.0,0.0,0.0,0.47500002,4.0444446,7.2222223,15.858334,26.244446,16.716667,6.211111,7.3083334,11.922222,9.788889,6.7083325,2.5222223,0.80833334,0.32222223,0.14166668,0.4,1.7916666,5.2222223,5.4666667,6.0583334,10.044444,12.758333,14.41111,15.250001,8.966667,9.422222,15.333334,19.011112,15.266666,7.922222,3.825,1.8444445,0.425,0.17777778,0.12222222,0.0,0.2888889,1.8083335,2.9222226,2.25,1.1222222,0.9666667,0.85833335,0.9666667,0.8999999,0.0,0.0,0.0,0.0,0.0,0.06666667,0.3416667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15833333,0.07777777,0.0,0.011111111,0.18888889,0.35000002,0.36666667,0.45000005,1.188889,2.875,3.9444447,4.7555556,5.441666,3.8111115,3.8333337,3.5666668,3.1,2.9555554,3.975,6.4888887,8.788889,15.374999,16.488888,17.108334,15.133334,11.566666,6.7555556,4.6777782,6.1749997,8.288888,8.433333,7.4333334,5.3166676,4.311111,3.6222224,4.008333,5.633333,6.541667,6.588889,5.466667,1.6333334,0.0,0.0,0.0,0.0,0.7888889,0.19166666,0.0,0.0,0.0,0.0,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17777778,0.20833334,0.07777778,0.23333332,0.0,0.30833334,0.4222222,0.6888889,0.5666666,0.33333334,0.0,0.0,0.0,0.0,0.0,0.12500001,0.35555553,0.25,0.24444446,0.075,0.11111111,0.5083334,0.6111111,1.2222222,1.05,1.9,3.1499999,4.5444446,6.525,7.8444443,7.5111113,8.349999,8.133333,5.933333,4.3,3.3333333,3.4222224,5.408333,5.366667,5.6888895,6.1833334,4.922222,3.1,2.1444445,2.4666667,2.388889,1.7444446,1.2916667,0.6,0.61666673,2.8555555,3.3083334,1.488889,0.1,0.0,0.8111111,0.9083333,0.88888896,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29166666,5.1749997,6.441667,8.133333,12.0375,16.383333,14.943749,15.066667,16.26875,15.650001,13.308333,9.168751,5.3583336,7.4937506,9.016668,12.25625,12.883334,10.806251,8.066667,7.516668,6.549999,5.866667,5.3875,4.983333,5.6625,5.2333336,5.116667,4.10625,3.5583334,2.6062503,2.1666665,1.625,1.4666667,0.9,1.6333334,3.1750002,2.8125,3.5666668,2.375,1.9666666,2.6875,4.0916667,2.4416668,0.5625,0.13333334,0.025,0.09166667,0.6875,2.2416668,4.491667,7.2499995,10.450001,12.887499,14.866667,19.26875,27.591667,32.831253,33.858334,33.95,27.043753,19.833334,16.63125,18.733334,24.16875,22.233332,17.575,15.48125,12.458334,6.387501,3.9250002,2.8812504,1.1916666,0.5500001,0.26666665,0.25,0.04375,0.0,0.0,0.15,1.4125,3.5666673,6.6166673,9.687499,18.616667,14.181252,7.2666674,1.64375,3.7416668,4.583333,2.5875,0.35,0.13750002,0.06666667,0.10625001,0.38333336,0.61875004,1.3083334,2.625,5.2437506,6.983333,10.525,13.408333,12.53125,11.45,13.983333,15.875,15.691667,11.275001,4.3916664,1.0250001,0.65833336,0.28125,0.0,0.0,0.50624996,1.3416668,1.75,2.2416668,2.3500004,2.6916668,2.3250003,1.6937501,1.0,0.36875,0.0,0.0,0.0,0.0,0.0,0.16666667,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21666668,0.0,0.13333334,0.0375,0.0,0.26250002,0.19166666,0.20833334,1.0749999,1.0583333,1.4,2.666667,2.6375,3.283333,3.741667,2.30625,1.7166668,1.6249999,1.7499998,1.5125,1.5500001,4.6312504,8.908334,14.199999,16.3625,17.208332,15.606251,11.866667,9.15625,5.25,3.3083334,4.5687504,6.083333,5.5937505,4.3250003,2.9687502,1.8833334,1.525,1.3687501,3.7250001,4.9500003,5.666667,5.5249996,2.125,0.01875,0.0,0.0,0.0,0.033333335,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.13125,0.0,0.0,0.0,0.0,0.0,0.0,0.69375,1.95,1.0375,0.075,0.025,0.70000005,0.6833334,1.5062501,0.6333333,0.15,0.1,0.1,0.3,0.65,1.66875,1.8083333,1.05625,0.5,0.3125,1.25,1.9499999,2.4916668,2.1166668,1.7125,2.025,1.9875,1.9833333,3.1562498,4.6499996,6.3,9.11875,11.650001,12.3125,10.966666,9.400001,9.783334,10.450001,9.625001,10.15,11.06875,10.308333,8.28125,6.7333336,4.2125,2.0,1.9166667,1.8437499,1.4166665,0.9,1.0916667,1.2375002,0.5916667,0.34375,0.3,1.1916666,1.8249999,0.425,0.04375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,11.1,13.211112,12.355555,12.716667,12.922223,12.083332,11.322222,14.475002,13.166666,13.055556,13.833335,13.666667,10.775001,10.544445,8.116667,5.8333335,4.6833334,1.4777777,2.1666667,2.4250002,1.7777779,1.5416667,0.85555553,1.9833336,3.3999999,4.2,3.8166673,2.511111,1.3999999,0.7444445,0.44166672,0.16666669,0.06666667,0.32222223,0.32222223,0.71666664,1.3666668,2.2833335,3.6111112,3.2166667,1.3666668,1.0555556,2.9416666,4.4,3.125,2.5555556,3.1666665,5.377778,8.444445,13.416666,20.033333,26.341667,30.922222,37.666668,37.81111,44.408333,46.17778,52.08889,40.983334,31.855556,34.200005,37.4,35.425003,30.355555,19.222221,8.566667,2.477778,3.2500005,4.433334,2.2500002,2.1000001,1.5083333,0.7444445,0.2777778,0.025000002,0.0,0.0,0.055555556,0.72499996,2.0111113,2.7444444,4.691666,10.677778,13.225,8.5,0.2,0.022222223,0.033333335,0.9083334,0.9666667,1.5250001,2.4777777,3.5416667,3.7444446,5.375,6.355556,6.1888895,5.258333,4.1,4.9083333,4.611111,6.7250004,8.233335,8.51111,8.191667,8.566667,2.816667,0.71111107,0.2,0.8666667,0.25,0.0,0.23333335,0.52500004,0.72222227,0.2916667,0.5444445,2.3333333,1.0888889,0.5888889,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15833335,0.7888889,0.19166668,0.0,0.0,1.1888889,1.4833333,0.7777778,1.1666666,1.3083334,1.6555556,1.8749999,2.188889,2.3500001,2.5888886,1.7222221,1.9833333,1.7222222,1.3499999,1.9555557,2.2083333,6.1222224,13.150001,16.899998,17.400002,15.558334,14.222223,11.483333,9.8,6.6833334,2.9444444,1.977778,2.6416664,2.3111112,2.408333,1.6888889,0.94166666,0.35555556,0.57777774,1.2666667,1.3111111,1.3166666,2.2555554,2.2666667,0.7,0.6500001,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333334,0.5333333,0.9666666,2.875,3.1,1.0500001,0.45555553,0.116666675,0.26666668,1.6000001,2.55,2.0444446,0.6916667,0.6333333,0.61666673,0.62222224,0.75555557,0.64166677,1.1111112,0.6166667,0.42222226,1.4916667,3.5111113,2.625,1.1444445,0.17777778,0.29166666,0.8555556,1.0083333,0.7888889,1.7583334,3.911111,3.8777776,4.2,6.2999997,8.208333,9.833333,11.025,12.511111,13.658333,12.533334,12.2,12.208334,11.644444,10.858333,8.977778,7.925,8.0,8.988889,8.491667,6.4111114,4.891667,4.2333336,2.2000003,0.5777778,0.5833333,1.4,2.0,3.0500002,2.1222222,0.575,0.0,0.041666668,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,11.858334,17.31111,19.155558,18.150002,14.177778,10.908334,8.644444,9.041667,7.3,7.811112,7.341666,10.066667,9.600001,11.355557,14.466667,17.433334,21.408333,20.511112,16.11111,11.908333,8.711112,5.45,5.544444,4.316667,3.8666668,3.1333334,1.9833333,1.2444445,0.5416667,0.23333332,0.34166667,0.7777778,1.1083333,2.1444445,2.5,3.6916666,4.0555553,3.475,3.9333334,7.0583334,13.666667,17.011112,18.175,13.499999,4.983333,5.0444455,8.216666,11.177777,14.644445,19.883333,25.811111,30.249998,33.044445,43.058334,43.355556,43.525,43.166668,35.41111,32.074997,27.17778,19.650002,21.233332,23.158333,19.58889,13.011112,4.125,2.6222222,1.925,0.9888889,0.5833333,0.7222222,0.75,1.7444445,0.16666667,0.016666668,0.0,0.016666668,0.48888892,2.025,3.9777777,1.8222222,1.2166667,1.7555556,2.15,3.788889,0.7833333,0.0,0.0,4.2166667,13.677776,20.116669,24.244444,20.808332,20.511112,14.15,10.255556,5.5888886,3.9083333,2.0777779,2.0750003,2.7222223,2.3333335,0.95555556,1.4777777,0.5916667,1.1,0.4166667,0.12222223,1.0,0.41111112,0.0,0.022222223,0.06666667,0.13333334,0.8777778,1.65,3.7111113,0.70000005,0.22222222,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.20000002,0.083333336,0.0,0.8333333,2.4111114,1.9250001,1.3555555,1.8444445,2.1666665,2.6555555,3.4250002,2.688889,2.075,1.2777777,1.0666666,1.4583333,1.1777778,2.6249998,4.744445,10.941668,13.977778,17.025002,18.255556,18.0,16.191666,10.933334,8.883334,8.622223,5.291667,1.6444445,1.0666666,0.45000002,0.26666668,0.30833334,0.055555556,0.0,0.13333334,0.2666667,0.4166667,0.46666667,0.65,0.6666667,0.5833334,0.77777785,0.6166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24166667,2.3000002,3.811111,3.2916667,1.3888888,0.9250001,1.7333333,1.075,0.0,1.3222222,1.5666668,1.2444445,0.6750001,1.3444445,2.2083333,1.7777779,1.1777778,0.4166667,2.222222,1.9416668,2.6000001,2.1916666,1.5777779,1.1916667,0.0,0.0,0.0,0.0,0.0,0.0,0.23333335,0.8777778,1.4222223,3.5833333,5.711111,6.7,5.8999996,5.9083333,7.3888893,8.5,8.588889,7.544444,4.991667,3.8888888,4.083333,4.5111113,6.3166666,7.1000004,7.344445,8.616668,10.688889,11.983334,10.166667,5.916667,2.488889,2.0500002,2.4222224,2.988889,3.7833335,2.711111,0.7166667,0.8,0.47500002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,9.443749,13.341666,18.633333,22.650002,26.191664,29.2875,32.283333,32.84375,35.633335,22.541668,22.375,21.741667,21.13125,19.641666,22.449999,23.466665,31.325,34.4,30.233335,17.96875,14.5,8.68125,4.791667,4.0,5.033334,6.924999,6.95,6.5166664,3.45,1.9750001,2.9562502,2.9916668,2.6312501,3.2583334,4.3250003,5.1875,6.2583337,8.43125,12.983334,16.5,21.775002,22.216667,18.018753,11.1,12.600001,10.525001,10.51875,12.708332,15.066666,20.362501,29.958332,33.90625,39.791664,41.674995,36.76667,30.675,23.150002,26.766666,21.2125,16.958334,10.793749,14.975,10.975,9.716667,7.408333,4.26875,1.4666666,0.425,1.3333334,2.2312498,1.3,1.3125,1.1916666,0.425,0.29375,0.48333335,1.3687501,2.7833333,10.21875,12.55,9.85,9.74375,4.675,2.7187502,4.0333333,4.1874995,3.3333335,3.466667,7.4187503,21.458336,31.256247,41.175003,41.3125,28.933332,13.787499,6.008333,1.9666667,0.6812501,1.1833333,1.9437501,3.258333,2.0187502,4.825,3.3333335,1.9437501,1.075,0.4,0.8916667,0.5125,0.0,0.0,0.0,0.06666667,0.43125004,0.83333325,1.8,3.2583337,1.05,0.28333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11666667,0.14375001,0.025,0.1875,0.6166667,1.9125,1.325,1.4875002,2.0916667,2.1916666,2.7812505,3.1666663,2.7312498,2.4833333,1.79375,1.1166666,1.0916667,1.525,3.8750002,6.1437497,11.783333,13.706249,14.133335,16.8125,19.666666,18.19167,14.4937525,11.775,9.58125,6.0750003,3.0437503,1.1166668,0.25,0.36875004,0.40833336,0.4,0.25,0.050000004,0.0,0.0,0.043750003,0.3166667,0.8437501,0.92500013,0.675,0.3,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.1,1.7416667,2.0666666,1.6812501,1.0083333,2.6437502,5.1000004,3.6375003,0.108333334,0.40000004,0.55,1.2166667,1.3812501,1.5916668,2.8875003,2.1666665,0.7083334,0.8624999,1.1666666,0.725,0.058333337,0.17500001,0.075,0.0,0.0,0.0,0.056250002,0.6666667,0.34374997,0.15,0.25625,0.225,0.5833333,1.325,2.266667,2.96875,2.891667,2.275,1.8750001,2.5375,4.075,5.2833333,5.1125,3.5,4.25,3.525,3.3500001,3.7750003,4.2,5.887501,9.258334,14.424998,16.408333,11.95,7.0666666,5.8125,3.975,2.7583332,3.2625,3.6583333,1.7937499,0.55833334,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.658333,4.1555557,5.0666666,7.183334,13.7,23.941668,30.911112,33.100002,31.744446,29.888891,28.825,28.222223,27.758335,30.111113,32.975002,34.944447,40.63333,32.72222,24.444445,19.099998,12.777778,10.974999,8.28889,11.691667,21.122221,26.077776,40.274998,44.7,33.066666,25.122223,12.583334,8.4777775,5.3499994,2.3666666,1.8,2.3249998,1.3444445,3.3249998,4.9222217,8.566668,12.322223,14.900001,14.983335,14.077778,13.524999,7.8555555,9.458335,16.733334,26.455555,32.658333,39.977776,38.35,35.9,30.150002,26.61111,23.216667,17.988888,13.044445,8.891666,8.166666,10.333333,9.400002,9.175001,9.644444,8.444445,3.6749997,1.0777777,0.28333336,0.70000005,0.8416667,0.7,1.0000001,2.277778,1.888889,3.35,3.4222226,3.8833334,6.0,21.766666,28.266668,29.08889,23.599998,19.633335,9.341667,8.644444,3.4916666,4.1111107,6.5000005,6.091667,10.533334,11.541668,13.18889,9.6,5.8555555,3.1749997,1.6222223,0.9555556,0.6000001,0.08888889,0.8583334,1.6000001,3.1666667,4.688889,1.9666667,1.1166667,0.39999998,0.09166667,0.12222223,0.075,0.0,0.0,0.0,0.7,2.85,5.1888895,5.316667,1.7,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.23333333,0.28333333,0.0,0.31111112,0.11666667,0.12222222,0.35,1.7,3.9333336,2.6444445,2.108333,1.6555555,1.6555557,1.1583333,0.7888889,0.85833335,1.4444444,2.2833333,2.788889,2.377778,4.608333,8.077778,10.025,11.544445,11.283334,16.755554,19.383335,22.222223,19.433334,16.058334,12.566668,10.091667,5.322222,2.1999998,1.0333334,1.011111,1.1166666,1.3555555,1.4416667,1.2666667,0.25,0.36666664,0.32222223,0.57500005,1.0111111,0.6166666,0.24444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,0.2777778,0.0,0.022222223,0.11111111,0.16666667,0.6888889,1.35,4.2666664,2.8250003,0.5222222,0.8333333,1.7166666,4.366667,3.0666668,1.588889,1.5500002,1.0888889,0.45555556,3.7166667,9.5,6.8250003,1.4222221,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.22222224,0.59166664,1.1777779,1.4777778,1.3416666,1.1999999,1.4916667,2.588889,3.8083334,4.5222225,2.725,1.277778,0.98888886,1.1583333,2.1444447,4.9750013,5.6,6.566666,7.8333335,7.2777777,8.183333,12.533334,16.925,18.655558,17.308334,18.544443,18.691668,14.355556,9.355556,5.325,4.055556,3.0416667,1.6666666,0.37500003,0.0,0.0,0.008333334,0.07777778,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.7500005,5.7916665,5.5416665,3.1750002,3.666667,6.74375,11.700002,18.64375,30.275003,30.208334,33.74375,34.600002,34.29375,35.65,37.287502,39.533333,44.156254,40.766666,33.916668,23.406252,20.258335,12.831251,8.241667,11.225,17.791666,22.383331,22.493752,18.133335,11.762499,9.683334,4.7375007,2.1583333,0.66249996,0.22500001,0.0,0.7062501,1.6166667,3.4687502,7.233333,13.787499,17.333334,20.658335,24.256248,19.958332,17.33125,13.866667,21.637503,30.474998,39.491665,45.468754,45.366665,35.8375,26.55,20.875,17.491667,14.900001,11.925,5.7250004,7.33125,8.791667,7.387501,7.758334,6.0687504,4.741667,4.408334,4.5249996,2.1083336,0.55,0.45,0.53125,0.9166666,0.66249996,0.875,1.4416667,1.0312499,1.7833333,8.5375,10.508333,20.768751,28.691666,29.391668,20.362501,15.533333,8.550001,5.3000007,1.93125,1.6416667,2.1083336,6.3875003,13.141667,12.299999,5.525,3.3062499,2.7583332,1.6687499,0.625,0.9,0.25,0.0,0.04375,0.3666667,0.14375,0.0,0.05,0.01875,0.0,0.0,0.0,0.0,0.0,0.2,1.1083333,3.0750003,4.6124997,3.591667,1.09375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.058333334,0.24375,0.19166668,0.10000001,0.13333334,0.26666668,0.075,0.09166667,0.3125,1.2583333,2.0499997,1.8416665,1.55,1.325,1.5666667,0.65,0.65,1.7750001,3.2416663,3.2,2.2,2.5083334,4.8812494,7.575,9.243749,7.5416665,6.381251,6.075,10.76875,14.558333,15.875001,14.431251,13.3583355,10.593751,7.175,4.1812506,2.416667,2.266667,2.8499997,3.5083337,3.2062502,2.1583335,1.98125,1.1750001,0.98333335,0.83125,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.10833334,0.081250004,2.2833333,1.7625,1.7333333,2.0500002,3.0625,3.9250002,2.075,0.575,0.05625,0.06666667,0.0,0.425,2.1,2.4,0.8833334,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.056250006,0.3,0.70625,1.3666666,1.4333332,1.1937499,0.7583333,0.46875003,0.67499995,1.15625,1.8416668,2.15,1.35,1.0749999,1.3125002,1.1250001,0.95625,0.8833334,1.875,4.4416666,5.4916663,6.9249997,9.833333,13.84375,19.358334,21.275,22.833334,24.931252,22.125,17.933334,11.125001,5.416667,3.3125,2.8583338,1.43125,0.16666667,0.033333335,0.3625,1.5333334,1.825,0.38333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0;
 } 
