netcdf ecmwf_r24_2018072300_f096 {
dimensions: 
 lat = 601; 
 lon = 701; 
variables:  
float lat(lat) ; 
   lat:long_name = "latitude" ;
   lat:units = "degrees_north" ;
   lat:standard_name = "latitude" ;
float lon(lon) ;
   lon:long_name = "longitude" ;
   lon:units = "degrees_east" ;
   lon:standard_name = "longitude" ;
float APCP_24(lat, lon) ;
   APCP_24:name = "APCP_24" ;
   APCP_24:long_name = "Total Precipitation" ;
   APCP_24:level = "A24" ;
   APCP_24:units = "kg/m^2" ;
   APCP_24:_FillValue = -9999.f ;
   APCP_24:init_time = "20180723_000000" ;
   APCP_24:init_time_ut = "1532304000.0" ;
   APCP_24:valid_time = "20180727_000000" ;
   APCP_24:valid_time_ut = "1532649600.0" ;
   APCP_24:accum_time = "240000" ;
   APCP_24:_FillValue = 65535 ;
   APCP_24:accum_time_sec = 86400 ;
 // global attributes: 
 :_NCProperties = "version=1|netcdflibversion=4.4.1.1" ;
	:FileOrigins = "ECMWF_HR_APCP24" ; 
	:MET_version = "V7.0" ;
	:Projection = "LatLon" ;
	:lat_ll = "0.0 degrees_north" ; 
	:lon_ll = "70.0 degrees_east" ; 
	:delta_lat = "0.10 degrees" ;
	:delta_lon = "0.10 degrees" ;
	:Nlat = "601 grid_points" ; 
	:Nlon = "701 grid_points" ; 
data:
lat = 0.0,0.1,0.2,0.3,0.4,0.5,0.6,0.7,0.8,0.90000004,1.0,1.1,1.2,1.3000001,1.4,1.5,1.6,1.7,1.8000001,1.9,2.0,2.1000001,2.2,2.3,2.4,2.5,2.6000001,2.7,2.8,2.9,3.0,3.1000001,3.2,3.3,3.4,3.5,3.6000001,3.7,3.8,3.9,4.0,4.1,4.2000003,4.3,4.4,4.5,4.6,4.7000003,4.8,4.9,5.0,5.1,5.2000003,5.3,5.4,5.5,5.6,5.7000003,5.8,5.9,6.0,6.1,6.2000003,6.3,6.4,6.5,6.6,6.7000003,6.8,6.9,7.0,7.1,7.2000003,7.3,7.4,7.5,7.6,7.7000003,7.8,7.9,8.0,8.1,8.2,8.3,8.400001,8.5,8.6,8.7,8.8,8.900001,9.0,9.1,9.2,9.3,9.400001,9.5,9.6,9.7,9.8,9.900001,10.0,10.1,10.2,10.3,10.400001,10.5,10.6,10.7,10.8,10.900001,11.0,11.1,11.2,11.3,11.400001,11.5,11.6,11.7,11.8,11.900001,12.0,12.1,12.2,12.3,12.400001,12.5,12.6,12.7,12.8,12.900001,13.0,13.1,13.2,13.3,13.400001,13.5,13.6,13.7,13.8,13.900001,14.0,14.1,14.2,14.3,14.400001,14.5,14.6,14.7,14.8,14.900001,15.0,15.1,15.2,15.3,15.400001,15.5,15.6,15.7,15.8,15.900001,16.0,16.1,16.2,16.300001,16.4,16.5,16.6,16.7,16.800001,16.9,17.0,17.1,17.2,17.300001,17.4,17.5,17.6,17.7,17.800001,17.9,18.0,18.1,18.2,18.300001,18.4,18.5,18.6,18.7,18.800001,18.9,19.0,19.1,19.2,19.300001,19.4,19.5,19.6,19.7,19.800001,19.9,20.0,20.1,20.2,20.300001,20.4,20.5,20.6,20.7,20.800001,20.9,21.0,21.1,21.2,21.300001,21.4,21.5,21.6,21.7,21.800001,21.9,22.0,22.1,22.2,22.300001,22.4,22.5,22.6,22.7,22.800001,22.9,23.0,23.1,23.2,23.300001,23.4,23.5,23.6,23.7,23.800001,23.9,24.0,24.1,24.2,24.300001,24.4,24.5,24.6,24.7,24.800001,24.9,25.0,25.1,25.2,25.300001,25.4,25.5,25.6,25.7,25.800001,25.9,26.0,26.1,26.2,26.300001,26.4,26.5,26.6,26.7,26.800001,26.9,27.0,27.1,27.2,27.300001,27.4,27.5,27.6,27.7,27.800001,27.9,28.0,28.1,28.2,28.300001,28.4,28.5,28.6,28.7,28.800001,28.9,29.0,29.1,29.2,29.300001,29.4,29.5,29.6,29.7,29.800001,29.9,30.0,30.1,30.2,30.300001,30.4,30.5,30.6,30.7,30.800001,30.9,31.0,31.1,31.2,31.300001,31.4,31.5,31.6,31.7,31.800001,31.9,32.0,32.100002,32.2,32.3,32.4,32.5,32.600002,32.7,32.8,32.9,33.0,33.100002,33.2,33.3,33.4,33.5,33.600002,33.7,33.8,33.9,34.0,34.100002,34.2,34.3,34.4,34.5,34.600002,34.7,34.8,34.9,35.0,35.100002,35.2,35.3,35.4,35.5,35.600002,35.7,35.8,35.9,36.0,36.100002,36.2,36.3,36.4,36.5,36.600002,36.7,36.8,36.9,37.0,37.100002,37.2,37.3,37.4,37.5,37.600002,37.7,37.8,37.9,38.0,38.100002,38.2,38.3,38.4,38.5,38.600002,38.7,38.8,38.9,39.0,39.100002,39.2,39.3,39.4,39.5,39.600002,39.7,39.8,39.9,40.0,40.100002,40.2,40.3,40.4,40.5,40.600002,40.7,40.8,40.9,41.0,41.100002,41.2,41.3,41.4,41.5,41.600002,41.7,41.8,41.9,42.0,42.100002,42.2,42.3,42.4,42.5,42.600002,42.7,42.8,42.9,43.0,43.100002,43.2,43.3,43.4,43.5,43.600002,43.7,43.8,43.9,44.0,44.100002,44.2,44.3,44.4,44.5,44.600002,44.7,44.8,44.9,45.0,45.100002,45.2,45.3,45.4,45.5,45.600002,45.7,45.8,45.9,46.0,46.100002,46.2,46.3,46.4,46.5,46.600002,46.7,46.8,46.9,47.0,47.100002,47.2,47.3,47.4,47.5,47.600002,47.7,47.8,47.9,48.0,48.100002,48.2,48.3,48.4,48.5,48.600002,48.7,48.8,48.9,49.0,49.100002,49.2,49.3,49.4,49.5,49.600002,49.7,49.8,49.9,50.0,50.100002,50.2,50.3,50.4,50.5,50.600002,50.7,50.8,50.9,51.0,51.100002,51.2,51.3,51.4,51.5,51.600002,51.7,51.8,51.9,52.0,52.100002,52.2,52.3,52.4,52.5,52.600002,52.7,52.8,52.9,53.0,53.100002,53.2,53.3,53.4,53.5,53.600002,53.7,53.8,53.9,54.0,54.100002,54.2,54.3,54.4,54.5,54.600002,54.7,54.8,54.9,55.0,55.100002,55.2,55.3,55.4,55.5,55.600002,55.7,55.8,55.9,56.0,56.100002,56.2,56.3,56.4,56.5,56.600002,56.7,56.8,56.9,57.0,57.100002,57.2,57.3,57.4,57.5,57.600002,57.7,57.8,57.9,58.0,58.100002,58.2,58.3,58.4,58.5,58.600002,58.7,58.8,58.9,59.0,59.100002,59.2,59.3,59.4,59.5,59.600002,59.7,59.8,59.9,60.0;
lon = 70.0,70.1,70.2,70.3,70.4,70.5,70.6,70.7,70.8,70.9,71.0,71.1,71.2,71.3,71.4,71.5,71.6,71.7,71.8,71.9,72.0,72.1,72.2,72.3,72.4,72.5,72.6,72.7,72.8,72.9,73.0,73.1,73.2,73.3,73.4,73.5,73.6,73.7,73.8,73.9,74.0,74.1,74.2,74.3,74.4,74.5,74.6,74.7,74.8,74.9,75.0,75.1,75.2,75.3,75.4,75.5,75.6,75.7,75.8,75.9,76.0,76.1,76.2,76.3,76.4,76.5,76.6,76.7,76.8,76.9,77.0,77.1,77.2,77.3,77.4,77.5,77.6,77.7,77.8,77.9,78.0,78.1,78.2,78.3,78.4,78.5,78.6,78.7,78.8,78.9,79.0,79.1,79.2,79.3,79.4,79.5,79.6,79.7,79.8,79.9,80.0,80.1,80.2,80.3,80.4,80.5,80.6,80.7,80.8,80.9,81.0,81.1,81.2,81.3,81.4,81.5,81.6,81.7,81.8,81.9,82.0,82.1,82.2,82.3,82.4,82.5,82.6,82.7,82.8,82.9,83.0,83.1,83.2,83.3,83.4,83.5,83.6,83.7,83.8,83.9,84.0,84.1,84.2,84.3,84.4,84.5,84.6,84.7,84.8,84.9,85.0,85.1,85.2,85.3,85.4,85.5,85.6,85.7,85.8,85.9,86.0,86.1,86.2,86.3,86.4,86.5,86.6,86.7,86.8,86.9,87.0,87.1,87.2,87.3,87.4,87.5,87.6,87.7,87.8,87.9,88.0,88.1,88.2,88.3,88.4,88.5,88.6,88.7,88.8,88.9,89.0,89.1,89.2,89.3,89.4,89.5,89.6,89.7,89.8,89.9,90.0,90.1,90.2,90.3,90.4,90.5,90.6,90.7,90.8,90.9,91.0,91.1,91.2,91.3,91.4,91.5,91.6,91.7,91.8,91.9,92.0,92.1,92.2,92.3,92.4,92.5,92.6,92.7,92.8,92.9,93.0,93.1,93.2,93.3,93.4,93.5,93.6,93.7,93.8,93.9,94.0,94.1,94.2,94.3,94.4,94.5,94.6,94.7,94.8,94.9,95.0,95.1,95.2,95.3,95.4,95.5,95.6,95.7,95.8,95.9,96.0,96.1,96.2,96.3,96.4,96.5,96.6,96.7,96.8,96.9,97.0,97.1,97.2,97.3,97.4,97.5,97.6,97.7,97.8,97.9,98.0,98.1,98.2,98.3,98.4,98.5,98.6,98.7,98.8,98.9,99.0,99.1,99.2,99.3,99.4,99.5,99.6,99.7,99.8,99.9,100.0,100.1,100.2,100.3,100.4,100.5,100.6,100.7,100.8,100.9,101.0,101.1,101.2,101.3,101.4,101.5,101.6,101.7,101.8,101.9,102.0,102.100006,102.2,102.3,102.4,102.5,102.600006,102.7,102.8,102.9,103.0,103.100006,103.2,103.3,103.4,103.5,103.600006,103.7,103.8,103.9,104.0,104.100006,104.2,104.3,104.4,104.5,104.600006,104.7,104.8,104.9,105.0,105.100006,105.2,105.3,105.4,105.5,105.600006,105.7,105.8,105.9,106.0,106.100006,106.2,106.3,106.4,106.5,106.600006,106.7,106.8,106.9,107.0,107.100006,107.2,107.3,107.4,107.5,107.600006,107.7,107.8,107.9,108.0,108.100006,108.2,108.3,108.4,108.5,108.600006,108.7,108.8,108.9,109.0,109.100006,109.2,109.3,109.4,109.5,109.600006,109.7,109.8,109.9,110.0,110.100006,110.2,110.3,110.4,110.5,110.600006,110.7,110.8,110.9,111.0,111.100006,111.2,111.3,111.4,111.5,111.600006,111.7,111.8,111.9,112.0,112.100006,112.2,112.3,112.4,112.5,112.600006,112.7,112.8,112.9,113.0,113.100006,113.2,113.3,113.4,113.5,113.600006,113.7,113.8,113.9,114.0,114.100006,114.2,114.3,114.4,114.5,114.600006,114.7,114.8,114.9,115.0,115.100006,115.2,115.3,115.4,115.5,115.600006,115.7,115.8,115.9,116.0,116.100006,116.2,116.3,116.4,116.5,116.600006,116.7,116.8,116.9,117.0,117.100006,117.2,117.3,117.4,117.5,117.600006,117.7,117.8,117.9,118.0,118.100006,118.2,118.3,118.4,118.5,118.600006,118.7,118.8,118.9,119.0,119.100006,119.2,119.3,119.4,119.5,119.600006,119.7,119.8,119.9,120.0,120.100006,120.2,120.3,120.4,120.5,120.600006,120.7,120.8,120.9,121.0,121.100006,121.2,121.3,121.4,121.5,121.600006,121.7,121.8,121.9,122.0,122.100006,122.2,122.3,122.4,122.5,122.600006,122.7,122.8,122.9,123.0,123.100006,123.2,123.3,123.4,123.5,123.600006,123.7,123.8,123.9,124.0,124.100006,124.2,124.3,124.4,124.5,124.600006,124.7,124.8,124.9,125.0,125.100006,125.2,125.3,125.4,125.5,125.600006,125.7,125.8,125.9,126.0,126.100006,126.2,126.3,126.4,126.5,126.600006,126.7,126.8,126.9,127.0,127.100006,127.2,127.3,127.4,127.5,127.600006,127.7,127.8,127.9,128.0,128.1,128.2,128.3,128.4,128.5,128.6,128.7,128.8,128.9,129.0,129.1,129.2,129.3,129.4,129.5,129.6,129.7,129.8,129.9,130.0,130.1,130.2,130.3,130.4,130.5,130.6,130.7,130.8,130.9,131.0,131.1,131.2,131.3,131.4,131.5,131.6,131.7,131.8,131.9,132.0,132.1,132.2,132.3,132.4,132.5,132.6,132.7,132.8,132.9,133.0,133.1,133.2,133.3,133.4,133.5,133.6,133.7,133.8,133.9,134.0,134.1,134.20001,134.3,134.4,134.5,134.6,134.70001,134.8,134.9,135.0,135.1,135.20001,135.3,135.4,135.5,135.6,135.70001,135.8,135.9,136.0,136.1,136.20001,136.3,136.4,136.5,136.6,136.70001,136.8,136.9,137.0,137.1,137.20001,137.3,137.4,137.5,137.6,137.70001,137.8,137.9,138.0,138.1,138.20001,138.3,138.4,138.5,138.6,138.70001,138.8,138.9,139.0,139.1,139.20001,139.3,139.4,139.5,139.6,139.70001,139.8,139.9,140.0;
APCP_24 = 7.4627824,6.5950966,6.4064693,6.094377,5.2987127,4.0880685,3.6868064,3.4021509,2.9322972,2.369845,2.2120838,1.8108221,1.7833855,1.8142518,1.8382589,2.0440342,1.8965619,1.9239986,1.9514352,1.9720128,2.1674993,2.1057668,1.8965619,1.6496316,1.5090185,1.6770682,1.4335675,1.5090185,1.6496316,1.6770682,1.4953002,1.6667795,2.0646117,1.9239986,1.2620882,0.8848336,0.6036074,0.45956472,0.37039545,0.28122616,0.18176813,0.25721905,0.45613512,0.6276145,0.8745448,1.5707511,1.8519772,2.8945718,3.998899,4.9214582,5.874883,4.8494368,5.381023,6.948344,8.594546,8.9100685,9.472521,10.6488695,11.7086115,12.840376,15.138199,15.858413,14.555169,14.126471,15.254805,16.403717,16.513464,15.954441,15.71094,15.988737,16.21852,14.54831,13.807519,13.4474125,13.680624,15.488017,15.097044,14.586036,14.225929,14.476289,15.9921665,17.075916,17.487467,17.021042,15.704081,13.762935,12.908967,13.063298,13.9481325,14.918706,14.953001,14.856973,15.014734,15.282242,15.868701,17.333136,19.483486,20.128248,19.94648,19.819586,20.858751,19.95677,17.772121,17.171944,18.632948,20.217419,21.37662,21.93221,22.261452,22.223726,21.150267,19.257133,18.28999,18.1288,18.44432,18.677534,18.44432,18.28656,18.608942,19.54179,20.920483,21.20171,21.150267,21.12283,21.4555,22.491234,22.223726,21.266872,20.303158,19.675543,19.394318,20.224277,21.28402,22.069395,22.096832,20.889618,20.53637,19.843594,19.390888,19.847023,21.956219,23.568125,22.011093,19.589804,18.169954,19.1954,17.988186,17.71382,17.254255,16.112202,14.404267,13.903547,13.999576,15.79325,18.482046,19.346302,18.70154,17.412016,17.134218,17.669235,16.997036,15.107333,15.172495,16.064188,16.45516,14.832966,13.4645605,12.425395,11.670886,11.201033,11.077567,10.48082,11.317638,13.125031,14.3974085,12.603734,10.81006,11.595435,13.049581,14.016724,14.112752,14.164196,13.279363,12.30193,12.048141,13.306799,13.169616,13.200482,14.037301,15.357693,15.88242,13.749216,12.747777,12.71691,13.275933,13.824667,15.885849,16.101913,16.252815,17.007324,17.899017,18.386019,18.132229,18.327715,19.716698,22.597551,22.43979,22.638706,22.70044,22.316326,21.37662,22.53582,23.173723,23.235455,22.741594,21.78817,21.067955,21.723007,22.20315,22.19286,22.583834,21.78817,20.821026,20.96164,21.815605,21.314886,21.28059,22.52553,23.146286,22.77932,22.583834,23.69502,23.496103,23.35549,23.828773,24.658733,22.412354,21.476076,21.328604,20.817596,18.142517,18.680964,18.320856,17.885298,17.995045,19.058218,18.557497,18.478617,18.838724,19.421753,19.775002,18.87302,18.351723,17.741257,17.168514,17.364002,18.231688,19.11652,20.073376,20.402617,18.646667,20.649546,21.815605,21.901346,21.1194,20.141968,20.179693,20.443771,20.913624,22.041958,24.76505,24.751333,24.291767,23.554407,22.587263,21.314886,21.013083,18.656956,16.715809,16.108772,16.21852,14.778092,14.208781,13.481709,12.185325,10.515115,9.23245,10.593996,12.079007,12.607163,12.55915,15.035312,16.588915,16.009314,13.684054,11.595435,8.189855,6.2864337,5.9160385,8.872343,18.722118,17.21996,11.5645685,8.498518,9.403929,10.268185,8.875772,8.868914,6.2555676,2.393852,3.9680326,6.1286726,5.552502,5.195825,6.358455,8.666568,11.365653,13.63261,14.750656,13.978998,10.573419,7.2775846,6.4098988,7.0786686,8.934075,12.144169,9.716022,7.891481,5.2747054,2.5481834,2.486451,3.4776018,2.3972816,1.704505,2.2155135,3.083199,4.1326528,5.192395,5.147811,4.1463714,3.5873485,2.5241764,1.8176813,1.4164196,1.1420527,0.70306545,0.21263443,0.06516216,0.041155048,0.048014224,0.12346515,0.17147937,0.26407823,0.33952916,0.39440256,0.5041494,0.6379033,0.9911508,1.5536032,2.2909644,3.1586502,3.0866287,3.4055803,3.8342788,4.0229063,3.5702004,3.2409601,2.819121,2.4590142,2.16064,1.7696671,2.2223728,2.3801336,2.0646117,1.4267083,0.9602845,1.155771,1.3169615,1.4815818,1.5090185,1.0837497,1.155771,1.430138,1.5398848,1.5364552,1.8931323,2.5138876,3.1277838,3.8925817,4.8117113,5.751418,3.82399,3.865145,3.99204,3.6319332,3.508468,3.5839188,3.5290456,3.5770597,3.7005248,3.6147852,3.8720043,3.433017,2.5619018,2.1332035,3.6456516,2.5619018,2.2600982,2.719663,3.4535947,3.5393343,4.3349986,4.15666,3.5530527,2.8156912,1.9994495,1.4507155,1.2312219,1.4369972,1.8965619,2.1503513,2.311542,2.2841053,2.9254382,4.280125,5.6005163,5.562791,3.2649672,1.9239986,2.2052248,2.2429502,2.8911421,2.4212887,2.5550427,3.40901,3.4947495,2.884283,3.8308492,6.142391,10.052121,16.204802,14.3974085,10.823778,10.079557,11.47197,9.016385,9.445084,9.259886,7.764586,6.135532,7.431916,6.125243,8.131552,10.31277,11.478829,12.421966,5.778855,5.8508763,6.667118,5.9983487,5.3398676,5.377593,4.746549,4.9351764,5.9571934,6.3481665,2.9185789,4.1463714,5.15467,4.705394,5.219832,4.4859004,6.526505,7.1884155,5.3398676,2.8980014,2.7882545,3.275256,3.566771,3.525616,3.6456516,3.292404,3.4707425,3.340418,2.867135,2.7916842,3.782835,3.2135234,2.6167753,2.3904223,1.8142518,2.0474637,2.095478,1.7250825,1.1934965,1.2655178,1.2792361,0.88826317,1.1934965,2.2498093,3.0660512,2.2258022,2.1332035,1.8691251,1.2586586,0.85396725,0.939707,1.1523414,1.3306799,1.3032433,0.90198153,2.452155,2.1160555,1.9137098,2.3046827,2.1812177,2.4761622,2.4487255,2.301253,2.1640697,2.0920484,3.690236,5.206114,5.3090014,4.280125,4.012617,2.095478,2.1743584,3.0866287,3.2889743,0.8848336,0.32238123,0.12003556,0.082310095,0.12346515,0.24350071,0.7442205,1.1454822,1.0597426,0.6001778,0.3806842,0.37039545,0.65848076,0.85396725,0.7613684,0.39783216,0.89855194,0.8196714,0.85739684,1.2243627,1.6633499,2.627064,2.1640697,1.6084765,1.786815,3.0214665,3.532475,2.8122618,2.3767042,2.6133456,2.7470996,2.8328393,3.292404,3.7313912,3.998899,4.180667,5.0346346,4.8734436,5.147811,5.768566,5.096367,5.7925735,5.5079174,4.787704,4.1429415,4.057202,3.192946,5.4736214,7.301592,6.90033,4.3487167,3.8960114,3.4535947,3.7039545,3.940596,2.061182,1.7319417,1.9411465,1.8382589,1.5158776,2.0303159,2.8945718,2.5173173,2.1503513,2.0920484,1.6770682,1.2517995,1.3272504,1.2723769,0.84367853,0.18176813,0.12346515,0.061732575,0.030866288,0.08573969,0.30523327,0.32924038,0.6207553,3.5016088,7.3530354,6.6225333,1.6290541,1.1694894,2.836269,5.305572,8.347616,7.9086285,7.164408,6.1149545,5.3227196,5.919468,4.540774,3.3987212,3.1723683,3.5153272,3.0523329,2.7470996,2.4590142,2.4658735,2.884283,3.6765177,5.6073756,6.958633,5.5902276,2.767677,3.1586502,5.8200097,8.224151,9.139851,8.827758,9.047252,8.913498,7.689135,6.0737996,4.7499785,4.3933015,4.9694724,6.5950966,8.669997,9.716022,7.3839016,7.8503256,8.405919,7.953213,6.5642304,5.4770513,5.137522,5.288424,4.8734436,3.7553983,2.7162333,2.7539587,1.8999915,1.7971039,3.0043187,5.020916,4.616225,5.3330083,5.977771,5.9983487,5.446185,5.130663,5.2335505,4.911169,4.2766957,4.4104495,4.6779575,4.5819287,4.5270553,4.6093655,4.6093655,4.15666,3.642222,3.2272418,3.2855449,4.4104495,4.7499785,4.2698364,4.122364,4.4927597,4.5784993,5.2747054,6.0154963,6.5230756,6.591667,6.1046658,6.9346256,8.515666,8.783174,7.349606,5.4941993,7.1061053,6.125243,5.377593,4.588788,3.7759757,3.2581081,2.5138876,2.2635276,2.1640697,2.07833,2.0646117,2.0234566,1.8382589,1.6873571,1.6256244,1.5810398,1.670209,1.6667795,1.611906,1.5844694,1.704505,1.5536032,1.4781522,1.6530612,1.8588364,1.4815818,1.4335675,1.471293,1.5193073,1.4541451,1.1043272,1.0014396,0.99801,0.83681935,0.53501564,0.37382504,0.23664154,0.18176813,0.14404267,0.1097468,0.1097468,0.23321195,0.45270553,0.77508676,1.1900668,1.6804979,2.2635276,3.3952916,4.4275975,4.9214582,4.65395,4.8117113,5.6005163,6.869464,8.06639,8.22758,8.985519,10.624862,11.921246,13.248496,16.588915,17.28169,16.173935,15.673215,16.311117,16.746675,16.317978,15.858413,15.570327,15.446862,15.268523,15.265094,14.987297,14.634049,14.754086,16.269962,15.234227,14.908417,15.769243,17.508043,19.041069,18.907316,18.235117,17.19938,15.947581,14.592895,13.495427,13.4474125,13.872682,14.369971,14.7095,14.699212,15.62863,16.856422,18.12194,19.517782,21.637268,21.795029,20.86561,19.847023,19.871029,18.235117,16.568336,16.269962,17.415445,18.77699,19.750994,20.340883,20.913624,21.297739,20.76958,19.023922,18.650097,19.058218,19.843594,20.78673,20.604961,19.668684,18.687822,18.217968,18.650097,19.740705,20.231136,20.361462,20.382038,20.550089,20.94449,20.61182,20.131678,19.78529,19.565796,19.03764,19.360022,20.323736,21.393766,21.719578,20.995934,20.560377,20.183123,20.03908,20.724997,22.412354,22.847912,21.78474,20.172834,20.135109,19.171394,17.837284,17.055338,17.000465,17.075916,15.748666,15.275383,15.560039,16.774113,19.349733,18.917604,17.353712,16.431154,16.47231,16.338554,14.788382,14.712931,15.357693,15.947581,15.71094,13.708061,12.205902,11.540562,11.482259,11.211322,11.38623,10.916377,11.835506,13.88983,14.555169,13.337666,12.950122,13.070158,13.54687,14.393978,15.1862135,15.642348,15.721229,15.584045,15.601193,13.982429,12.30193,13.536582,16.877,17.703531,16.20137,15.518884,15.450292,15.820687,16.496315,17.302269,17.748116,18.145947,18.571217,18.886738,19.003344,18.811287,18.852442,19.716698,22.048819,22.60441,23.098272,22.889067,21.94936,20.851892,20.03908,20.402617,20.567236,20.176264,19.898466,20.03565,20.135109,20.237995,20.388897,20.642687,19.771572,19.603521,20.131678,20.841602,20.742146,20.999365,21.400625,21.671564,21.928782,22.679861,23.811626,23.60242,23.324625,23.681301,24.806206,23.70188,22.69701,21.716148,20.553518,18.87645,18.934752,18.094503,17.676094,17.95389,18.166525,17.442883,17.28512,17.384579,17.799559,18.945042,18.451181,18.396307,18.296848,17.95389,17.425734,18.320856,19.102802,19.901896,20.265432,19.171394,19.726988,20.234566,20.954779,21.44521,20.556948,20.896477,21.836184,21.839613,21.157125,21.846472,21.20171,20.433481,19.8676,19.613811,19.596663,18.547209,17.003895,16.249386,16.269962,15.755525,15.018164,13.855534,12.6586075,11.736049,11.293632,12.240198,16.194511,17.504614,15.752095,15.7795315,16.684942,15.364552,12.507706,10.2921915,12.367092,9.438225,8.944365,8.179566,7.840037,11.996697,15.896138,16.986746,13.193623,7.699424,8.927217,4.1772375,5.874883,5.5593615,3.316411,7.798882,6.6705475,7.5416627,8.48137,9.22216,11.156448,11.657167,12.072148,11.866373,10.4533825,7.191845,6.4544835,7.14726,8.7317295,10.960961,13.87954,10.72775,7.56567,4.5990767,2.7402403,3.5873485,4.9248877,2.7916842,2.16064,3.6044965,3.2889743,4.6127954,4.496189,3.9851806,3.5221863,2.9494452,2.270387,1.6530612,1.3272504,1.3478279,1.5913286,0.42183927,0.116605975,0.09602845,0.08573969,0.1097468,0.216064,0.28122616,0.32581082,0.37039545,0.42869842,0.72021335,1.4129901,2.07833,2.5070283,2.719663,2.7059445,2.843128,3.093488,3.2889743,3.117495,3.1620796,3.000889,2.942586,2.8396983,2.0886188,1.9925903,2.3149714,2.0165975,1.1900668,1.0460242,1.2826657,1.4781522,1.6599203,1.6393428,1.0460242,1.3341095,1.6839274,1.9171394,1.9445761,1.7833855,2.1229146,2.760818,3.6147852,4.623084,5.7274113,5.1066556,4.4996185,3.6216443,2.585909,1.8862731,1.7456601,2.5310357,3.2272418,3.9474552,5.9126086,4.4584637,4.0229063,3.6285036,3.2375305,3.7553983,3.3061223,3.9028704,4.383013,4.413879,4.5270553,4.180667,3.5633414,3.2615378,3.1895163,2.5961976,2.1263442,1.8142518,1.6873571,1.8073926,2.2978237,4.125794,3.0626216,2.4727325,3.4673128,4.90431,2.417859,4.2869844,6.0566516,6.2144127,6.2212715,6.420188,7.9600725,9.908078,9.72288,3.2855449,3.74168,6.893471,8.968371,8.947794,8.577398,11.866373,9.414218,8.64942,11.317638,13.474849,7.3187394,8.100685,8.368194,6.3001523,5.7102633,4.033195,7.589677,9.73317,9.191295,10.052121,7.4353456,5.778855,5.4804807,6.012067,5.9400454,5.9469047,4.664239,4.314421,4.945465,4.420738,3.6559403,3.9611735,4.012617,3.6010668,3.6559403,4.2698364,3.450165,3.806842,5.0003386,3.74168,2.585909,2.5550427,2.8122618,3.0900583,3.6696587,3.4844608,3.7759757,3.7313912,3.3987212,3.6970954,3.7176728,3.083199,2.4212887,2.136633,2.4144297,2.2463799,2.3492675,2.1915064,1.7388009,1.4610043,0.91569984,0.85739684,2.8054025,5.411889,4.420738,1.8313997,1.5810398,1.9342873,1.9342873,1.4164196,1.6873571,2.07833,2.8911421,3.426158,1.9857311,2.9700227,2.3835633,2.170929,2.6853669,2.6716487,2.0063086,2.5756202,3.0729103,3.4192986,4.763697,5.0929375,5.1512403,4.9077396,4.6436615,4.9420357,2.2429502,1.5193073,1.6564908,1.8005334,1.3478279,1.0494537,0.58988905,0.65505123,1.1283343,1.0734608,1.2723769,1.1934965,0.9911508,0.78194594,0.65162164,0.6276145,0.9945804,1.1866373,1.0151579,0.6790583,0.8471081,0.6344737,0.6962063,1.1489118,1.5913286,2.3286898,2.5070283,2.4487255,2.551613,3.2649672,4.108646,3.57363,2.8705647,2.7916842,3.6970954,4.2835546,4.866585,5.305572,5.528495,5.535354,6.0875177,6.0052075,5.960623,5.9126086,5.096367,5.576509,5.0483527,4.4721823,4.1943855,3.974892,2.7642474,6.1492505,8.934075,8.39563,4.262977,4.0949273,3.350707,3.532475,4.1943855,2.9391565,1.9548649,1.978872,2.3629858,2.6887965,2.760818,3.1106358,3.1072063,2.8945718,2.5207467,1.9582944,1.3066728,1.4815818,1.3443983,0.66876954,0.14747226,0.09602845,0.06516216,0.041155048,0.18862732,0.8676856,1.2998136,1.3478279,1.7490896,2.4075704,2.3972816,2.218943,3.059192,4.705394,6.7528577,8.591117,7.613684,6.9792104,6.169828,5.188966,4.5647807,4.6127954,4.4550343,4.2355404,3.758828,2.503599,2.2669573,2.253239,2.4007113,2.702515,3.2135234,3.0900583,2.7813954,3.415869,4.8494368,5.662249,6.125243,7.5862474,8.508806,8.855195,10.062409,8.988949,7.6205435,6.715132,6.2247014,5.284994,5.693115,7.4456344,8.4093485,7.9017696,6.715132,7.459353,7.7885933,6.931196,5.4599032,5.271276,5.144381,4.7431192,4.331569,3.6765177,2.0337453,2.020027,2.8054025,4.2046742,5.641671,6.142391,5.377593,5.336438,5.720552,6.0223556,5.5319247,5.2644167,5.394741,5.4770513,5.381023,5.302142,5.442755,4.996909,4.705394,4.5784993,3.923448,3.940596,3.8205605,3.542764,3.391862,3.957744,4.046913,3.9337368,3.7862647,3.683377,3.6147852,4.7774153,5.562791,5.693115,5.470192,5.7754254,6.8763227,8.39563,8.995808,8.169277,6.2247014,5.3707337,4.437886,3.8857226,3.3850029,2.8637056,2.5207467,2.1023371,2.0646117,1.9891608,1.8073926,1.8176813,1.8828435,1.7765263,1.6942163,1.6770682,1.6016173,1.6839274,1.7559488,1.6530612,1.471293,1.5673214,1.3478279,1.2792361,1.4198492,1.5227368,1.0323058,1.0014396,0.9568549,0.881404,0.7579388,0.548734,0.5624523,0.4938606,0.37039545,0.23664154,0.16119061,0.09945804,0.082310095,0.072021335,0.072021335,0.1097468,0.22978236,0.41840968,0.7442205,1.2860953,2.1194851,2.8328393,3.4227283,3.9371665,4.273266,4.184097,4.6436615,5.56965,6.90033,8.107545,8.2310095,8.903209,10.299051,11.334786,12.229909,14.500296,15.848124,16.21166,16.283682,16.352274,16.300829,15.875561,15.614912,15.597764,15.549749,14.829536,14.956431,14.846684,15.055889,15.728088,16.582056,15.13134,15.385129,16.475739,17.857862,19.301718,19.418324,18.406595,17.000465,15.7795315,15.158776,15.405707,15.525743,15.724659,16.05733,16.45173,16.033321,16.578627,18.025911,20.03908,22.007662,22.998814,22.77932,22.083115,21.28059,20.37175,18.197392,16.846134,16.475739,16.925014,17.71382,20.296299,21.939072,22.806757,22.844482,21.764162,19.644676,18.938183,18.9519,19.411465,20.4472,21.37319,21.664703,20.697561,19.106232,18.759844,19.641247,19.819586,19.963629,20.361462,20.899906,20.814167,20.19341,19.500635,19.05136,19.013634,18.674105,18.176813,18.344864,19.288,20.406046,20.937632,20.7833,20.666695,20.762722,20.728426,21.592682,22.127699,21.956219,21.270302,20.810738,19.915615,18.756414,17.820137,17.62122,18.725548,18.20425,18.269413,17.569777,16.702091,18.20425,17.562918,16.86671,16.386568,16.177364,16.108772,15.429714,14.942713,14.904987,15.103903,14.867262,14.054449,12.452832,11.818358,12.257345,12.205902,12.836946,11.808069,11.729189,13.190193,14.778092,14.027013,13.934414,13.834956,13.96185,15.409137,15.995596,17.446312,18.269413,17.761833,15.981877,14.520873,13.601744,14.191633,15.803539,16.499744,16.482597,17.103354,17.333136,17.099922,17.29541,17.110212,17.463459,18.053349,18.656956,19.143957,19.123379,19.871029,20.382038,20.526081,21.033659,21.860191,22.336903,22.052248,20.94449,19.312008,18.248835,18.506054,18.62609,18.310568,18.427174,18.327715,18.430603,18.800999,19.263992,19.432043,18.855871,18.814716,19.085653,19.713268,21.002794,21.170843,21.03709,21.03023,21.410915,22.28546,23.911083,24.295198,24.140865,24.041409,24.473536,24.329493,23.256033,21.633839,19.987637,18.986197,18.478617,17.974468,17.96761,18.060207,16.945591,17.28512,17.315987,16.973028,16.79126,17.912735,18.12537,17.826996,17.398296,17.096493,17.04848,18.344864,19.010202,19.46291,19.829874,19.932762,18.773561,18.331144,19.027351,20.179693,20.001354,20.189981,20.673553,20.711279,20.128248,19.322296,19.03078,18.804428,18.180243,17.302269,16.921585,16.575195,16.266533,16.575195,16.911295,15.522313,14.606613,13.588025,13.173045,13.406258,13.660047,14.033872,16.901007,17.350283,15.223939,15.110763,15.611482,13.817808,14.116182,16.979887,18.95533,13.042721,11.718901,10.360784,8.31332,8.89635,9.774324,10.244178,10.089847,9.057541,6.869464,3.5873485,6.6293926,7.222711,5.178677,8.906639,5.288424,6.094377,8.724871,11.067279,11.506266,12.253916,10.940384,9.482809,8.539673,7.4936485,8.457363,9.321619,10.405369,11.523414,11.986408,10.484249,7.1232533,4.417309,3.4604537,3.9063,3.6799474,2.0714707,1.9445761,3.4535947,4.0366244,4.214963,4.0846386,3.707384,3.1380725,2.417859,1.9480057,1.4095604,1.2209331,1.4987297,2.054323,0.548734,0.13032432,0.11317638,0.12346515,0.09602845,0.23321195,0.34638834,0.4355576,0.4972902,0.5041494,0.7442205,1.3684053,2.0749004,2.6064866,2.7745364,2.6922262,2.527606,2.7059445,3.1586502,3.316411,3.2889743,3.1826572,3.0111778,2.7402403,2.2841053,1.978872,2.095478,1.7765263,1.1111864,1.1317638,1.2826657,1.5433143,1.7902447,1.7662375,1.0734608,1.3855534,1.8656956,2.2566686,2.3904223,2.1469216,2.3664153,3.1655092,3.9097297,4.48933,5.329579,5.7102633,5.06893,3.9680326,2.7128036,1.3786942,2.0474637,3.1106358,4.232111,5.6245236,8.05953,5.3878818,4.1600895,3.875434,4.187526,4.8734436,4.513337,4.482471,4.3452873,4.3178506,5.2609873,5.4599032,4.482471,3.6593697,3.433017,3.340418,3.2135234,2.6750782,2.8259802,3.3712845,2.6167753,3.083199,3.0660512,2.7059445,2.6990852,4.3178506,2.5070283,7.133542,9.911508,8.995808,8.97523,7.9257765,10.398509,12.47341,10.981539,3.5359046,4.6882463,9.352485,10.415657,6.711703,3.0351849,6.807731,6.4098988,5.8337283,7.4936485,12.205902,4.846007,7.160979,8.378482,6.046363,6.0395036,6.101236,7.390761,8.182996,7.7611566,6.4133286,7.0478024,6.989499,6.8145905,6.7219915,6.5470824,6.2967224,5.288424,4.2355404,3.7005248,4.091498,3.2615378,3.3266997,3.4467354,3.5118976,4.1155047,4.57164,2.8877127,2.5893385,3.666229,2.568761,1.4164196,1.4575747,2.0028791,2.6647894,3.3747141,3.8720043,3.7176728,3.3026927,3.059192,3.4638834,3.083199,3.1552205,2.74367,2.0989075,2.6819375,2.3904223,2.585909,2.5996273,2.2120838,1.6564908,0.89169276,0.7305021,2.4075704,4.73969,4.1120753,1.8519772,1.1454822,1.2003556,1.371835,1.1523414,1.1180456,1.2312219,1.7662375,2.3218307,1.8176813,1.9720128,1.5364552,1.4232788,1.7422304,1.7765263,1.5021594,1.646202,2.1674993,3.2443898,5.284994,6.001778,5.2815647,4.787704,5.0586414,5.5113473,1.9514352,1.0357354,1.7799559,2.702515,1.8313997,1.1900668,1.2209331,3.2203827,5.977771,5.7754254,6.944915,7.1952744,7.233,6.625963,3.8308492,1.9685832,1.4507155,1.2929544,1.0048691,0.61046654,0.75450927,0.64133286,0.6344737,0.89169276,1.3512574,1.8245405,2.1674993,2.7951138,3.415869,3.0420442,3.940596,4.1189346,3.8925817,3.7931237,4.5682106,5.518206,5.381023,5.7068334,6.5779486,6.615674,6.6225333,6.6293926,6.4579134,6.0497923,5.442755,5.7308407,5.0757895,4.32471,3.765687,3.1380725,2.9288676,5.0655007,7.7268605,8.4093485,3.9303071,4.2286816,3.5221863,3.2443898,3.782835,4.4756117,4.588788,3.5599117,3.1963756,3.7725463,4.0057583,3.9268777,3.7553983,3.1586502,2.2600982,1.6633499,1.2277923,1.1900668,0.9842916,0.51100856,0.14747226,0.08916927,0.06859175,0.06516216,0.3018037,1.2346514,3.3609958,3.5702004,3.0283258,2.6304936,2.9906003,3.1586502,3.625074,5.2506986,7.4799304,8.323608,7.116394,6.468202,6.0875177,5.7068334,5.079219,4.7191124,4.0777793,3.8617156,3.8857226,3.0797696,2.6990852,2.020027,1.8382589,2.3424082,3.1346428,3.5530527,4.3590055,5.0757895,5.6176643,6.3035817,7.0478024,8.992378,10.6317215,11.561139,12.504276,10.508256,9.191295,8.22758,7.239859,5.802862,5.809721,6.7700057,7.3564653,6.8626046,5.192395,6.252138,6.5299344,5.844017,4.804852,4.835718,4.496189,4.400161,4.2595477,3.6765177,2.153781,2.020027,3.0969174,4.98662,6.7940125,7.130112,6.8454566,6.4098988,6.118384,5.909179,5.3432975,5.593657,6.0154963,6.3721733,6.3035817,5.3398676,5.7136927,5.2335505,4.647091,4.2595477,3.9097297,4.15323,3.9131594,3.5942078,3.5016088,3.8171308,3.4398763,3.450165,3.3747141,3.2066643,3.3815732,4.064061,4.770556,5.535354,6.39961,7.4113383,7.970361,8.683716,8.803751,8.323608,7.9909387,3.7176728,3.000889,2.7951138,2.644212,2.3629858,2.0337453,1.8999915,1.8965619,1.8073926,1.5981878,1.3924125,1.471293,1.5364552,1.5158776,1.430138,1.371835,1.4644338,1.611906,1.5193073,1.2346514,1.1489118,0.94999576,0.91569984,0.9328478,0.864256,0.548734,0.52815646,0.47671264,0.38754338,0.29837412,0.25721905,0.32238123,0.274367,0.18862732,0.12346515,0.08916927,0.061732575,0.0548734,0.061732575,0.09602845,0.18862732,0.36353627,0.52815646,0.91227025,1.5570327,2.3218307,3.0557625,3.4878905,3.8377085,4.2183924,4.636802,5.127233,6.183546,7.346176,8.176137,8.217292,8.64942,9.678296,10.467101,10.971251,11.955542,13.742357,14.990726,15.553179,15.642348,15.817257,15.059319,14.843254,15.21365,15.642348,15.055889,14.994157,14.38369,14.517444,15.570327,16.602633,15.896138,16.45859,17.031332,17.412016,18.423744,19.301718,19.020493,17.744686,16.13278,15.354263,16.05733,16.232237,16.331696,16.636929,17.257685,17.082775,17.230247,18.197392,20.045938,22.426073,22.823904,22.885637,22.834194,22.43979,21.04395,18.71526,17.566347,17.288551,17.525192,17.87158,20.467777,22.710728,23.972816,23.983105,22.789608,21.45893,19.881319,18.917604,18.897026,19.603521,20.834743,22.158566,21.908205,20.334024,19.596663,20.107672,19.888178,19.936192,20.60839,21.62012,21.335464,20.52951,19.641247,18.927893,18.46147,18.313997,17.569777,17.192522,17.597214,18.643238,19.823015,20.20027,20.711279,21.325174,21.074816,21.150267,21.211998,21.43835,21.654415,21.328604,20.749004,20.183123,19.188541,18.348293,19.274282,20.21056,21.074816,20.351171,18.434032,17.61779,16.45859,16.564907,16.70895,16.383139,15.810398,15.683503,15.254805,14.832966,14.483148,14.044161,14.339106,13.46799,12.864383,12.905538,12.922686,13.526293,12.655178,12.30193,13.066729,14.171056,14.568888,14.496866,14.315098,14.778092,17.000465,17.278261,18.499195,19.312008,18.735836,16.160215,15.608052,16.0539,15.892709,15.097044,15.189643,15.830976,16.743246,17.171944,17.144508,17.466888,16.770683,16.743246,17.086205,17.549198,17.916164,18.95533,19.94305,20.344313,20.159115,19.905325,20.53637,20.742146,20.594673,19.963629,18.530062,17.031332,17.055338,17.271402,17.233677,17.364002,17.267973,17.54234,18.025911,18.485476,18.602083,18.807858,18.883308,18.855871,19.353163,21.575535,21.685282,21.393766,21.486366,22.065966,22.546108,23.890507,24.339783,24.394655,24.27119,23.893936,23.94195,22.841053,21.215427,19.665255,18.752985,18.001905,17.751545,17.854433,17.682953,16.108772,17.562918,17.645227,16.931873,16.276823,16.80155,17.350283,17.137648,16.640358,16.359133,16.828985,18.166525,18.663815,18.787281,18.979338,19.658396,17.87158,17.271402,17.655516,18.550638,19.20912,19.648108,19.44576,19.486916,19.565796,18.37916,18.36887,18.595222,17.744686,16.0539,15.29253,15.6526375,15.834405,16.352274,16.660936,15.12448,14.064738,13.63261,14.284232,15.337115,14.96672,14.627191,15.745236,15.827546,14.616901,14.081886,13.471419,12.648318,14.699212,18.073925,16.616352,12.614022,14.061309,15.302819,13.831526,10.281903,5.2026844,4.180667,6.2487082,8.220721,4.7019644,6.1321025,8.282454,8.1212635,6.540223,8.3922,4.856296,6.509357,10.686595,14.081886,12.737488,12.22648,10.542552,9.081548,8.419638,8.303031,10.131001,10.679735,11.2593355,11.526843,9.496528,9.211872,6.56766,5.178677,5.2472687,3.5873485,2.253239,1.6016173,1.7010754,2.6304936,4.465323,4.1326528,3.8274195,3.4707425,2.959734,2.1434922,1.7525192,1.2826657,1.1660597,1.5501735,2.3286898,0.6824879,0.17490897,0.13032432,0.15090185,0.116605975,0.2469303,0.40126175,0.53158605,0.59331864,0.53501564,0.8676856,1.2929544,1.845118,2.411,2.719663,2.7368107,2.4144297,2.5584722,3.1895163,3.5187566,3.3747141,3.350707,3.1243541,2.7093742,2.452155,2.085189,1.9754424,1.6667795,1.214074,1.1454822,1.2380811,1.5330256,1.8382589,1.8656956,1.2277923,1.471293,2.0131679,2.452155,2.6167753,2.551613,2.8225505,3.6319332,4.245829,4.465323,4.650521,5.2335505,5.0895076,4.3178506,3.1723683,2.0749004,3.199805,3.9954693,5.206114,6.742569,7.706283,6.0566516,4.8597255,4.8288593,5.5833683,5.6793966,5.5559316,5.003768,4.482471,4.496189,5.6039457,5.7411294,4.8837323,4.0263357,3.7348208,4.170378,4.6608095,3.899441,3.957744,4.523626,2.8980014,3.0489032,3.841138,3.340418,2.452155,4.9420357,3.6559403,6.4990683,7.805741,6.6739774,6.9723516,6.108095,7.5588107,8.707723,7.5416627,2.6407824,6.029215,10.545981,9.873782,4.314421,0.78194594,5.8165803,5.9571934,4.633373,5.1238036,10.590566,4.2355404,6.8797526,7.7371492,5.271276,7.1884155,9.112414,7.7748747,7.486789,8.196714,5.501058,6.025785,7.486789,8.889491,9.462232,8.656279,6.3961806,7.1712675,6.258997,3.6387923,3.9646032,3.0797696,3.4981792,3.9714622,4.245829,5.051782,4.8322887,3.4707425,3.059192,3.7176728,3.6113555,1.5124481,1.2003556,2.1400626,3.350707,3.4124396,4.0846386,3.9680326,3.4055803,2.959734,3.3850029,2.5996273,3.0248961,2.9974594,2.4041407,2.6887965,2.4315774,2.551613,2.5584722,2.2292318,1.6153357,0.9431366,0.59674823,1.7079345,3.532475,3.457024,2.0234566,0.9294182,0.5041494,0.64476246,0.83681935,0.7373613,0.607037,0.7990939,1.2998136,1.7147937,1.8313997,1.6290541,1.5981878,1.6633499,1.1660597,1.4815818,2.0406046,2.7779658,3.8034124,5.4187484,6.941485,6.7528577,6.094377,5.7377,5.9640527,3.1689389,2.3218307,2.603057,2.8637056,1.605047,0.97400284,2.9871707,5.411889,6.8866115,6.931196,9.002667,10.576848,11.609154,10.916377,6.1801167,5.809721,5.7068334,4.4516044,2.2635276,0.9945804,0.7613684,0.64476246,0.5761707,0.6310441,1.0288762,1.430138,1.8519772,2.719663,3.4947495,2.6750782,3.8137012,4.3658648,4.5647807,4.619654,4.722542,5.2644167,5.336438,5.8508763,6.6739774,6.6053853,6.7322803,6.8626046,6.667118,6.2041235,5.895461,5.857735,5.164959,4.3590055,3.6765177,3.0454736,2.976882,5.0243454,6.9037595,6.9792104,4.249259,4.7362604,4.057202,3.7039545,4.15666,4.887162,6.0806584,4.852866,3.9714622,4.307562,4.8322887,4.602506,4.057202,3.2306714,2.2978237,1.546744,1.1454822,0.922559,0.72364295,0.47328308,0.18176813,0.09259886,0.072021335,0.08573969,0.34981793,1.3512574,3.9783216,4.8494368,4.602506,4.0434837,4.15666,4.0023284,3.8720043,5.0483527,7.058091,7.658269,6.625963,6.3001523,6.2247014,5.9880595,5.2438393,5.1100855,4.2698364,3.782835,3.8479972,3.8171308,2.9734523,1.99602,1.5947582,1.99602,2.9391565,4.1943855,5.06893,5.2781353,5.312431,6.4407654,8.158989,10.203023,11.540562,11.856084,11.55771,11.135871,10.593996,9.582268,8.347616,7.723431,7.1026754,6.9723516,6.944915,6.509357,5.0620713,5.429037,5.3158607,4.8940215,4.4550343,4.40702,4.273266,3.782835,3.5221863,3.3884325,2.6167753,2.0165975,2.9322972,5.1066556,7.455923,8.073249,7.8126,7.3839016,6.90033,6.3618846,5.693115,6.341307,6.4304767,6.5710897,6.6465406,5.8337283,5.6142344,5.003768,4.4584637,4.1600895,4.0263357,4.249259,3.7108135,3.2203827,3.1209247,3.2855449,2.9871707,3.1037767,3.1586502,3.1312134,3.450165,3.7931237,4.5682106,5.857735,7.39762,8.573969,8.597976,8.7317295,8.553391,8.31332,8.968371,2.750529,2.2738166,2.2635276,2.2258022,1.9925903,1.7079345,1.605047,1.4472859,1.3958421,1.3546871,0.9534253,1.0288762,1.1934965,1.1351935,0.89512235,0.84024894,0.9774324,1.1351935,1.0734608,0.78194594,0.4698535,0.3806842,0.4115505,0.3806842,0.2709374,0.21263443,0.24007112,0.24007112,0.22978236,0.22292319,0.24350071,0.20920484,0.15433143,0.10288762,0.06859175,0.061732575,0.0548734,0.061732575,0.10288762,0.1920569,0.35324752,0.6001778,0.82996017,1.3889829,2.1126258,2.335549,3.0214665,3.8342788,4.513337,5.0449233,5.662249,6.108095,7.2878733,8.035523,8.097256,8.14527,8.423067,9.098696,9.72631,10.196163,10.714031,12.360233,13.37882,14.027013,14.555169,15.223939,13.828096,13.663476,14.376831,15.251375,15.223939,15.402277,14.157337,13.498857,14.239647,15.978448,16.616352,17.21653,17.45317,17.511473,18.073925,19.233126,19.908754,19.164536,17.185663,15.254805,15.145059,15.179354,15.155347,15.313108,16.328266,17.412016,17.885298,18.163095,18.835295,20.680412,20.94449,21.37662,21.77102,21.767591,20.851892,18.910746,17.988186,18.019053,18.54035,18.684393,19.435472,21.085104,22.44322,22.87192,22.264881,22.738165,20.78673,19.058218,18.62609,19.013634,19.648108,20.968498,21.476076,20.882757,20.104242,20.436913,20.220848,20.162544,20.604961,21.53781,21.654415,21.067955,20.388897,19.70641,18.574646,17.947031,17.250826,16.79126,16.763824,17.243965,17.916164,18.773561,19.94648,21.019941,21.04395,21.04395,20.913624,21.067955,21.421204,21.37319,21.28059,21.239435,20.574095,19.521212,19.236557,21.013083,22.501524,22.686722,21.19485,18.28656,16.571766,16.763824,17.264544,17.058767,15.707511,15.37827,15.289101,14.977009,14.476289,14.30481,14.977009,15.1862135,14.517444,13.450842,13.365103,13.718349,13.502286,13.666906,14.147048,13.872682,15.584045,15.055889,14.634049,15.6697855,18.499195,19.102802,19.380598,19.637817,19.346302,17.134218,17.158226,18.495766,18.005335,15.782962,15.155347,15.927004,16.04018,16.04018,16.287111,16.96274,16.365992,15.9750185,15.817257,15.851553,15.954441,18.406595,18.883308,18.694681,18.636377,18.989626,19.11652,18.807858,18.893597,19.243416,18.77699,16.71238,16.37971,16.6335,16.846134,16.88043,17.141079,17.4566,17.778982,18.04649,18.197392,19.167965,19.582945,19.596663,19.87446,21.592682,21.69214,21.939072,22.642136,23.492674,23.557837,23.756752,23.537258,23.715597,24.003683,22.995384,22.669573,21.650986,20.526081,19.504065,18.392878,17.689812,17.247395,17.027903,16.753534,15.927004,17.593784,17.545769,16.79126,16.03675,15.704081,16.071047,16.486027,16.496315,16.317978,16.846134,17.652086,17.988186,18.053349,18.12194,18.533491,17.425734,17.398296,17.463459,17.562918,18.581505,19.305147,18.825006,18.773561,19.202261,18.584934,18.45804,18.547209,17.586924,15.9613,15.690363,16.108772,15.944152,15.738377,15.440002,14.387119,13.701202,14.085316,15.429714,16.503176,14.918706,14.870691,15.0078745,15.237658,15.155347,14.05102,11.952112,12.4802685,13.015285,11.835506,8.1487,10.6145735,15.87899,19.408035,18.746124,13.516005,3.9474552,2.8911421,4.540774,5.2301207,3.433017,9.050681,8.81747,8.14527,8.580828,7.795452,5.8474464,9.084977,14.040731,17.28169,15.419425,11.712041,10.494537,9.9869585,9.301042,8.450503,10.264755,10.264755,10.662587,10.943813,7.8777623,7.394191,5.9434752,6.2830043,7.1129646,3.0797696,1.8108221,1.9925903,1.920569,1.8554068,4.0366244,4.3590055,3.6525106,3.1072063,2.867135,2.0131679,1.6496316,1.2655178,1.138623,1.4815818,2.469303,0.8025235,0.23664154,0.15433143,0.16804978,0.14747226,0.28122616,0.44927597,0.607037,0.6790583,0.5555932,1.0254467,1.255229,1.5433143,1.9582944,2.3458378,2.6579304,2.3972816,2.5378947,3.1792276,3.5564823,3.3644254,3.415869,3.3061223,2.976882,2.702515,2.2600982,2.0097382,1.786815,1.4987297,1.1283343,1.255229,1.5330256,1.8382589,1.9411465,1.4987297,1.5638919,2.085189,2.4830213,2.6304936,2.8396983,3.2066643,3.9097297,4.4550343,4.513337,3.9165888,4.1326528,4.6402316,4.3933015,3.4878905,3.1620796,4.1463714,4.616225,5.669108,6.715132,5.4496145,6.447624,6.334448,6.444195,6.7322803,5.7651367,5.744559,5.4633327,5.2609873,5.336438,5.761707,4.99005,4.479041,4.149801,4.122364,4.7499785,5.9880595,5.0449233,4.496189,4.5990767,3.2649672,4.273266,4.629943,3.4535947,2.417859,5.7479887,4.5613513,3.07634,1.937717,1.5536032,2.0989075,4.0880685,3.059192,2.435007,2.7093742,1.4575747,7.599966,10.377932,7.98408,2.7333813,1.0425946,8.076678,7.781734,5.960623,6.217842,9.97324,5.346727,7.425057,7.332458,4.7088237,7.682276,10.487679,8.412778,7.6033955,8.690575,6.773435,5.096367,6.924337,10.412228,12.88496,10.816919,5.857735,8.357904,8.471081,4.770556,4.2218223,3.532475,4.3178506,4.955754,5.079219,5.576509,4.9934793,4.108646,3.9954693,5.007198,6.756287,2.7333813,1.6359133,2.8019729,4.4550343,3.7005248,4.3452873,4.5167665,3.899441,3.117495,3.7382503,2.6545007,2.7162333,2.8465576,2.6750782,2.5207467,2.3629858,2.3046827,2.1983654,1.9068506,1.3409687,0.88826317,0.48357183,1.2963841,2.8259802,2.901431,2.7059445,1.3752645,0.4389872,0.3806842,0.64133286,0.83338976,0.77508676,1.0425946,1.6599203,2.0680413,2.4487255,2.417859,2.49331,2.4898806,1.5398848,1.6736387,2.983741,4.105216,4.822,6.0635104,7.8126,8.237869,7.3358874,6.001778,6.0086374,5.3913116,4.712253,3.4535947,1.920569,1.2483698,1.0048691,4.386442,5.394741,3.5290456,3.782835,6.0978065,8.580828,10.7757635,11.118723,6.927767,9.448513,10.6145735,8.453933,4.166949,2.1297739,1.0117283,0.64133286,0.5418748,0.53501564,0.7305021,1.2037852,1.8485477,2.5653315,2.9803114,2.452155,3.9268777,4.3761535,4.650521,4.8425775,4.307562,4.0023284,5.0312047,5.9400454,6.1046658,5.7239814,6.691125,6.914048,6.684266,6.307011,6.101236,5.7136927,5.223262,4.5819287,3.9131594,3.5221863,3.0797696,6.5710897,7.514226,5.288424,5.130663,5.56965,4.5853586,4.506478,5.267846,4.417309,5.099797,4.8837323,4.5682106,4.6402316,5.2747054,5.0449233,4.1772375,3.3884325,2.784825,1.8416885,1.1729189,0.89512235,0.7613684,0.58302987,0.24350071,0.1097468,0.08573969,0.09602845,0.34638834,1.3581166,3.2272418,4.7191124,5.209543,4.7774153,4.2252517,4.448175,4.3624353,4.8768735,6.0052075,6.869464,6.433906,6.591667,6.5470824,5.926327,4.7945633,5.40503,5.0620713,4.2355404,3.5873485,3.9646032,2.9185789,2.2635276,1.8965619,1.937717,2.7128036,3.782835,3.6696587,3.923448,5.1512403,7.0203657,8.820899,9.9801,10.220171,9.4862385,7.949784,10.199594,10.628291,10.028113,9.421077,10.041832,8.766026,7.874333,7.0615206,6.3378778,6.0532217,5.164959,4.482471,4.2183924,4.214963,3.9680326,4.2423997,3.0386145,2.5721905,3.1689389,3.2855449,1.937717,2.609916,4.962613,7.682276,8.512236,7.9737906,7.7783046,7.658269,7.3530354,6.6053853,7.023795,6.3961806,6.0978065,6.3790326,6.3721733,5.3432975,4.4996185,4.1429415,4.1635194,4.0537724,4.064061,3.3815732,2.760818,2.5070283,2.4761622,2.7402403,2.935727,3.0866287,3.3061223,3.7794054,4.3041325,5.195825,6.2864337,7.3290286,7.9737906,7.9943686,8.2653055,8.2481575,8.1384115,8.851766,2.2120838,1.7353712,1.7559488,1.670209,1.3684053,1.2209331,1.1489118,1.0117283,0.90541106,0.8779744,0.91569984,0.96371406,0.9568549,0.823101,0.64476246,0.65505123,0.6207553,0.7099246,0.6001778,0.31209245,0.21263443,0.20234565,0.20920484,0.18862732,0.15090185,0.15090185,0.18862732,0.17147937,0.13375391,0.1097468,0.12346515,0.09602845,0.072021335,0.0548734,0.048014224,0.061732575,0.072021335,0.13032432,0.25378948,0.42869842,0.61046654,0.7682276,1.2483698,2.037175,2.784825,2.8225505,3.3850029,4.413879,5.4084597,6.0875177,6.392751,6.478491,7.7097125,8.296172,8.097256,8.621983,9.23245,9.22902,9.441654,10.179015,11.214751,12.312219,12.809509,13.179905,13.540011,13.625751,12.247057,12.689473,13.591455,14.078457,13.749216,14.870691,14.273943,13.169616,12.682614,13.855534,14.356253,15.405707,17.106783,18.975908,19.929333,19.87789,19.692692,19.418324,18.36887,15.121051,14.620332,14.651197,14.284232,13.862392,14.983868,17.912735,19.78186,20.111101,19.363451,18.934752,17.765263,16.95931,16.969599,17.813278,19.058218,18.142517,17.658945,17.816708,18.279701,18.159666,18.060207,17.943602,18.248835,18.71526,18.3723,19.70298,19.548649,18.468328,17.511473,18.217968,19.047928,19.86074,20.478067,20.604961,19.836735,20.03222,20.419764,20.412905,20.097382,20.217419,20.570665,20.2037,20.2037,20.515793,19.94305,18.36887,16.811838,15.933864,15.854982,16.160215,16.280252,16.732958,17.765263,19.13024,20.080235,21.153696,21.496655,21.174273,20.52951,20.186552,20.176264,20.4472,21.143406,21.472647,19.713268,20.189981,22.093403,23.60928,23.252604,19.898466,18.019053,17.501184,18.04992,18.502625,16.828985,15.525743,14.942713,14.904987,15.29596,16.050468,16.96617,17.178804,16.098484,14.538021,14.7095,15.247946,15.810398,16.578627,16.901007,15.289101,16.619781,16.486027,16.071047,16.47231,18.708399,20.941061,21.434921,21.479506,21.126259,19.20912,18.149376,19.678972,19.377169,16.96274,16.266533,18.903887,18.948471,17.264544,15.165636,14.435134,14.582606,14.424845,14.280802,14.503725,15.501736,17.079346,17.765263,17.916164,17.998474,18.584934,18.255693,17.130789,17.28169,18.605513,18.814716,18.056778,17.53891,17.086205,16.856422,17.319416,17.161655,17.20281,17.63494,18.296848,18.660385,19.270851,20.056227,20.587814,20.567236,19.823015,19.589804,21.626978,23.410364,24.058556,24.3535,23.633287,22.721018,22.762173,23.129137,21.407484,21.150267,20.382038,19.552078,18.821575,18.04992,17.21996,16.307688,15.758954,15.755525,16.21852,16.55119,16.503176,16.259674,15.752095,14.678635,14.7026415,15.707511,16.341984,16.369421,16.660936,16.688372,17.003895,17.604073,18.190533,18.20425,18.190533,18.262554,18.163095,17.995045,18.20425,17.61779,17.655516,17.837284,17.926455,17.912735,17.669235,16.969599,16.516893,16.80155,18.080786,18.03277,17.689812,16.37285,14.445422,13.337666,13.629181,14.891269,16.204802,16.702091,15.580616,16.45859,16.21166,15.96816,15.697222,14.222499,12.754636,13.855534,12.737488,10.467101,13.944703,18.36544,17.511473,12.596875,8.244728,12.466551,3.199805,1.7010754,3.6216443,5.446185,4.4721823,7.8023114,7.034084,10.220171,15.097044,9.078118,6.368744,9.14328,13.361672,16.520323,17.655516,11.9040985,9.716022,9.3764925,9.438225,8.742019,9.561689,8.419638,8.207003,8.793462,7.034084,5.7891436,5.3227196,6.090947,6.5470824,3.1277838,2.1503513,3.0969174,2.9254382,1.6942163,2.5481834,3.6593697,3.5599117,3.1415021,2.6373527,1.6496316,1.3786942,1.1489118,1.0425946,1.3101025,2.335549,0.78537554,0.2503599,0.17147937,0.18176813,0.12346515,0.35324752,0.53844523,0.7888051,0.9945804,0.823101,0.9328478,0.97057325,1.1592005,1.5158776,1.845118,2.4212887,2.3424082,2.534465,3.175798,3.7382503,3.4192986,3.2135234,3.1346428,3.1552205,3.2032347,2.4967396,2.0646117,1.99602,1.9720128,1.2517995,1.4335675,1.6530612,1.8965619,2.037175,1.8142518,1.4610043,1.9582944,2.435007,2.6819375,3.1586502,3.3781435,4.2218223,4.7499785,4.4996185,3.4638834,3.7211025,4.3692946,4.3281393,3.5290456,2.9288676,4.0880685,5.0929375,6.0532217,6.3893213,4.852866,7.160979,7.9737906,7.133542,5.6313825,5.6313825,4.3487167,4.8254294,5.7411294,6.310441,6.2864337,5.6039457,4.7259717,4.3349986,4.4550343,4.4550343,6.2487082,5.1238036,4.201245,4.3521466,4.180667,3.4124396,2.386993,1.4815818,1.4850113,3.5873485,4.7808447,3.542764,2.4144297,2.136633,1.6496316,9.386781,6.341307,2.8499873,2.7402403,3.3266997,8.796892,9.338767,6.6533995,2.9734523,1.0666018,5.363875,7.1712675,8.659708,9.668007,7.689135,5.6999745,8.700864,9.006097,5.936616,5.813151,8.279024,8.4093485,6.632822,4.588788,5.127233,4.307562,6.6122446,10.587136,12.950122,8.604835,3.9303071,4.3933015,5.4599032,5.672538,6.636252,4.122364,4.2183924,4.650521,4.756838,5.4770513,5.501058,3.9611735,3.4227283,4.839148,7.5382333,2.5584722,1.2655178,2.1400626,3.4810312,3.433017,5.4839106,4.695105,3.1449318,2.4555845,3.799983,3.309552,2.6853669,2.1983654,2.0337453,2.287535,2.2292318,2.201795,2.1469216,1.8759843,1.0837497,0.6310441,0.33609957,0.6173257,1.3752645,1.9994495,4.880303,3.2546785,1.3752645,0.7510797,0.15433143,0.48357183,0.8676856,1.7525192,2.6922262,2.3492675,1.2758065,1.3649758,1.7559488,2.1160555,2.6407824,1.0048691,0.53158605,1.3546871,3.57363,7.2467184,7.881192,5.926327,4.3590055,4.262977,4.835718,5.65539,5.2918534,3.8274195,2.2841053,2.6407824,2.2600982,1.4164196,1.845118,3.0386145,2.2600982,4.297273,4.266407,6.2144127,9.3936405,8.268735,6.036074,6.1732574,5.56965,3.9371665,3.8137012,1.6427724,0.7888051,0.66533995,0.75450927,0.59674823,0.91227025,2.0165975,2.9391565,3.1586502,2.609916,3.8925817,4.3590055,4.547633,4.5990767,4.256118,3.9646032,4.5682106,5.453044,5.9331865,5.2506986,6.958633,7.1026754,6.6876955,6.1972647,5.6005163,5.223262,5.4667625,4.972902,3.6559403,2.7162333,4.266407,8.014946,8.433355,5.6656785,5.5079174,6.1904054,4.3041325,3.998899,5.552502,5.3707337,2.527606,3.5016088,5.099797,5.919468,6.3481665,5.7994323,4.856296,3.8925817,3.0523329,2.2566686,1.4027013,1.0700313,0.9568549,0.78194594,0.30523327,0.17147937,0.12003556,0.106317215,0.4046913,1.6016173,3.8102717,4.7019644,5.0757895,5.055212,4.105216,4.3349986,5.2266912,5.720552,5.7822843,6.392751,6.9071894,6.8969,6.6396813,6.1972647,5.4153185,4.6127954,4.5030484,3.957744,3.0351849,2.976882,3.2683969,2.7573884,2.369845,2.5310357,3.1277838,2.6647894,4.307562,6.0875177,7.3255987,8.604835,8.189855,8.114404,8.601405,9.0369625,7.949784,8.707723,8.7317295,9.102125,9.650859,8.940934,7.4044795,6.691125,6.0532217,5.4187484,5.3707337,4.5784993,4.029765,3.8788633,3.8445675,3.234101,2.8568463,2.952875,3.4673128,4.105216,4.3487167,2.393852,2.5927682,4.383013,6.5813785,7.4010496,7.936065,7.798882,7.881192,8.097256,7.3393173,6.447624,6.0806584,6.025785,5.8337283,4.822,5.1992545,4.3795834,3.6147852,3.5290456,4.0880685,3.7965534,3.4467354,3.059192,2.6579304,2.3046827,2.7573884,2.7402403,2.7882545,3.340418,4.746549,5.6005163,6.169828,6.245279,5.8988905,5.5079174,6.2418494,7.3839016,7.579388,7.298162,8.851766,1.5055889,1.430138,1.5913286,1.646202,1.488441,1.2312219,0.90541106,0.66876954,0.5590228,0.5555932,0.5624523,0.7373613,0.6756287,0.5555932,0.48357183,0.48357183,0.44927597,0.41498008,0.31895164,0.20234565,0.21263443,0.1920569,0.16462019,0.1371835,0.11317638,0.10288762,0.09259886,0.08916927,0.08916927,0.07545093,0.048014224,0.072021335,0.06859175,0.08573969,0.13375391,0.19548649,0.16804978,0.31209245,0.45270553,0.6207553,1.039165,1.2826657,1.8142518,2.417859,2.9391565,3.2855449,4.0229063,4.7808447,5.960623,7.1884155,7.298162,7.0889573,7.579388,7.915488,7.9189177,8.083538,8.471081,8.98209,9.465661,9.746887,9.654288,10.779194,11.729189,12.21962,12.147599,11.588576,12.103014,12.668896,13.087306,13.21763,12.953552,13.433694,13.025573,12.521424,12.408247,12.867812,12.898679,13.831526,15.083325,16.482597,18.241976,18.320856,18.694681,18.8593,18.091074,15.440002,15.251375,15.12448,14.808959,14.363112,14.167625,15.357693,16.37285,16.78783,16.760393,17.055338,16.95931,16.969599,17.065628,17.20624,17.350283,16.317978,15.656067,15.697222,16.736387,19.03764,19.994495,19.884748,19.408035,18.506054,16.359133,16.986746,17.226818,17.20281,17.072487,17.04848,17.905876,18.907316,19.750994,20.111101,19.654966,19.44919,19.692692,19.857311,19.833303,19.925903,19.94648,19.421753,18.972477,18.828436,18.831865,18.53692,17.394867,16.21852,15.477728,15.306249,15.251375,15.71094,16.427725,17.350283,18.602083,20.262003,21.390337,21.589252,20.920483,19.905325,20.138538,20.61182,21.465788,22.017952,20.738716,20.28944,21.256582,22.450079,22.841053,21.582394,20.12139,19.86417,19.871029,19.62753,19.041069,18.005335,16.050468,15.282242,15.896138,16.173935,17.000465,17.315987,16.616352,15.525743,15.782962,15.608052,16.029892,17.027903,18.02934,17.902447,18.265984,18.344864,17.995045,17.741257,18.742695,20.498644,21.585823,22.076254,21.805317,20.35803,18.828436,19.668684,20.237995,19.246845,16.753534,19.078794,20.992504,20.910194,18.831865,16.352274,15.422854,15.752095,16.321407,16.722668,17.175373,17.391438,18.406595,18.886738,18.722118,19.023922,19.339443,17.899017,17.405157,18.430603,19.401176,18.495766,17.96418,17.802988,17.95046,18.259123,16.94902,16.732958,17.243965,18.012194,18.4649,18.71526,19.13024,20.100813,20.810738,19.246845,19.250275,20.899906,22.371199,23.070835,23.657295,23.35549,22.316326,21.70929,21.503513,20.457489,20.141968,19.723558,18.989626,18.084215,17.501184,17.072487,16.317978,15.772673,15.635489,15.769243,15.05246,15.193072,15.367981,14.953001,13.505715,14.088745,14.822677,15.71094,16.671225,17.54234,17.487467,17.04505,17.178804,17.919594,18.351723,18.28999,17.799559,17.607502,17.744686,17.532051,16.359133,17.086205,17.70696,17.748116,18.241976,18.938183,18.389448,18.118511,18.602083,19.277712,17.62808,16.650646,14.030442,10.899229,11.859513,13.869251,15.066177,15.556609,15.498305,15.079896,15.196502,15.271953,15.618341,15.542891,13.341095,11.46854,11.238758,13.337666,16.674654,18.427174,14.2533655,11.050131,8.995808,8.327039,9.366203,3.1072063,1.8828435,4.108646,6.3618846,3.3712845,7.641121,7.6274023,11.180455,15.964729,9.469091,8.272165,8.7145815,10.593996,13.591455,17.264544,12.960411,12.751206,12.840376,11.293632,8.049242,8.378482,7.881192,8.124693,8.268735,5.0929375,5.9297566,5.8062916,5.809721,5.3878818,2.3595562,3.0523329,4.8185706,4.338428,2.1915064,2.8396983,3.6113555,3.2718265,2.6373527,2.054323,1.4164196,1.2072148,1.039165,0.91227025,1.0631721,1.9823016,0.72364295,0.22635277,0.14061308,0.1920569,0.17147937,0.32581082,0.5418748,0.8848336,1.1934965,1.0940384,1.3786942,1.2895249,1.3375391,1.6153357,1.7971039,1.9411465,2.2052248,2.510458,2.942586,3.7382503,3.3815732,3.1209247,2.9734523,2.8637056,2.6304936,2.5961976,2.2566686,2.2498093,2.3664153,1.5673214,1.6256244,1.7765263,2.0406046,2.2498093,2.061182,1.6290541,1.8999915,2.2463799,2.5001693,2.9871707,3.5016088,3.9337368,4.2766957,4.2389703,3.2203827,3.8171308,3.9440255,3.6765177,3.1106358,2.3561265,3.0454736,3.532475,5.0620713,6.6431108,5.0346346,6.8626046,7.9463544,7.281014,6.0497923,7.630832,6.869464,5.31929,4.870014,5.6176643,5.895461,5.857735,4.8494368,4.7431192,5.6245236,5.809721,5.377593,5.137522,5.038064,4.695105,3.3987212,2.5241764,1.8588364,1.7456601,2.1297739,2.5481834,2.3389788,3.8377085,3.5633414,1.5707511,1.4541451,4.681387,5.003768,3.3438478,1.6667795,2.983741,4.166949,5.754848,7.208993,6.8728933,1.9720128,2.1469216,5.6348124,7.8503256,7.6925645,7.531374,7.699424,8.56025,8.220721,6.186976,3.3609958,8.64942,7.1198235,4.513337,3.9851806,6.1149545,5.0929375,6.2384195,6.9552035,6.550512,6.2384195,4.3349986,3.981751,3.882293,3.9200184,5.147811,4.705394,5.038064,5.6793966,5.8645945,4.5270553,5.2438393,4.3658648,4.396731,6.025785,8.134981,6.759717,3.4604537,2.2841053,3.7279615,4.763697,4.7362604,3.7485392,3.069481,3.0043187,2.9322972,2.7470996,2.3732746,1.961724,1.7113642,1.862266,2.0337453,1.9068506,1.8862731,1.7765263,0.77851635,0.5796003,0.4355576,0.50757897,1.6221949,5.2815647,10.000677,6.725421,4.420738,4.6265135,1.4575747,1.6427724,2.4795918,3.3747141,3.5873485,2.2395205,3.5599117,6.667118,6.7974424,3.649081,1.430138,1.6804979,2.5927682,3.2135234,3.6559403,5.1238036,7.8091707,9.280463,7.6033955,5.627953,10.978109,4.48933,8.855195,10.590566,6.1561093,1.9685832,2.6236343,2.7711067,3.07634,3.2718265,2.1469216,2.253239,4.996909,6.252138,5.302142,4.852866,5.2266912,3.707384,4.9591837,7.040943,1.4095604,1.3375391,0.94999576,0.66533995,0.6001778,0.5590228,0.7476501,1.704505,2.527606,2.7951138,2.5481834,3.525616,4.2046742,4.5339146,4.389872,3.5599117,3.5221863,4.029765,4.880303,5.579939,5.3330083,5.813151,6.3310184,6.3138704,5.7651367,5.2335505,4.846007,5.1100855,5.0655007,4.046913,1.6907866,4.1017866,6.824879,6.23156,3.865145,6.461343,4.389872,4.245829,3.8617156,2.8156912,2.417859,2.335549,3.2375305,4.866585,6.324159,6.0806584,5.802862,5.675967,4.9831905,3.799983,2.9665933,1.9651536,1.3238207,1.0288762,0.88826317,0.548734,0.2503599,0.17147937,0.18176813,0.5727411,2.054323,3.590778,4.3692946,4.557922,4.5167665,4.8254294,5.4084597,5.874883,5.871454,5.610805,5.8817425,6.276145,6.025785,5.562791,5.3090014,5.662249,5.3913116,4.712253,3.940596,3.4433057,3.6353626,3.5359046,3.1620796,2.7711067,2.726522,3.4810312,4.2081037,4.619654,4.9214582,5.3878818,6.3481665,7.486789,8.008087,8.1212635,7.6376915,5.98463,5.638242,6.3378778,7.332458,7.7371492,6.550512,5.693115,5.3707337,5.336438,5.2438393,4.6402316,4.6745276,4.3349986,3.6765177,3.0626216,3.1723683,2.3252604,2.2326615,2.9906003,4.040054,4.1772375,2.2360911,2.2738166,3.6525106,5.658819,7.5210853,7.7851634,7.1369715,7.016936,7.675417,8.158989,6.944915,6.691125,6.7357097,6.478491,5.394741,4.73969,4.1360826,3.5050385,3.1620796,3.8205605,3.4981792,3.192946,2.9494452,2.8568463,3.0489032,3.3232703,3.1552205,3.2889743,3.99204,5.0620713,5.586798,6.0154963,6.2041235,6.310441,6.776865,6.8557453,7.5210853,7.7851634,7.8777623,9.253027,1.0700313,1.196926,1.2998136,1.1934965,0.91569984,0.7133542,0.50757897,0.42183927,0.4046913,0.4081209,0.40126175,0.5041494,0.4629943,0.42869842,0.44584638,0.45956472,0.33609957,0.25721905,0.20920484,0.18862732,0.19548649,0.14747226,0.1097468,0.082310095,0.06859175,0.06516216,0.048014224,0.048014224,0.044584636,0.041155048,0.048014224,0.08573969,0.14061308,0.22978236,0.33952916,0.42183927,0.42183927,0.6344737,0.881404,1.1729189,1.6942163,2.07833,2.6613598,3.100347,3.426158,4.0537724,4.4104495,5.3432975,6.619104,7.6651278,7.5862474,7.7885933,8.604835,8.820899,8.289313,7.922347,8.7145815,9.630281,9.97324,9.647429,9.14328,9.962952,10.600855,11.30049,11.770344,11.197603,11.849225,12.418536,12.792361,12.950122,12.984418,12.644889,12.517994,12.79922,13.183334,12.895248,12.6757555,13.581166,14.747226,16.067617,18.180243,18.999914,19.6241,19.6241,18.890167,17.63151,17.1205,15.6526375,14.788382,14.925565,15.278812,15.7795315,16.05733,15.971589,15.6526375,15.515453,15.621771,15.951012,16.688372,17.669235,18.406595,17.350283,16.37285,15.580616,15.662926,17.902447,19.497204,19.322296,18.663815,17.820137,16.12935,15.395418,15.704081,16.444872,17.051908,16.993607,17.154797,17.61779,18.410025,19.003344,18.317427,18.471758,19.229696,19.654966,19.596663,19.70641,19.263992,18.684393,18.317427,18.12537,17.686382,17.813278,17.497755,16.96617,16.335125,15.604623,14.781522,15.13134,15.854982,16.588915,17.439453,19.353163,20.577524,21.009653,20.752434,20.100813,20.803877,21.304598,21.736725,21.939072,21.4555,21.524092,21.585823,21.969936,22.467228,22.350622,21.85333,21.664703,20.95135,19.871029,19.582945,19.342873,17.69667,16.894148,17.12393,16.506605,16.088194,16.606062,16.901007,16.6335,16.263103,15.367981,15.536031,16.208231,17.086205,18.142517,18.945042,18.962189,18.44432,18.0362,18.752985,20.001354,21.527521,22.5221,22.210009,19.840164,18.653526,18.95876,20.148827,20.656404,17.95732,18.307138,19.967058,21.19485,21.047379,19.411465,18.420315,18.324286,18.680964,19.243416,19.963629,19.740705,19.79901,19.709839,19.54179,19.87446,20.104242,19.065077,18.639809,19.308577,20.159115,19.243416,18.687822,18.471758,18.37573,18.008764,16.842705,16.7844,17.388008,18.193962,18.728977,18.351723,18.61923,19.634388,20.649546,20.073376,20.107672,20.591244,21.297739,21.86362,21.798458,22.415783,22.062536,21.328604,20.560377,19.843594,19.490345,19.161106,18.804428,18.307138,17.484037,17.04505,16.993607,16.671225,15.88242,14.904987,14.586036,14.829536,14.915276,14.555169,13.872682,14.404267,14.459141,14.822677,15.71437,16.80155,17.655516,17.346853,16.986746,17.343424,18.825006,18.862732,18.180243,17.864721,18.101362,18.187103,17.154797,17.322845,17.700102,17.857862,17.923023,17.78927,17.425734,17.346853,17.679523,18.166525,16.599203,14.1299,10.912948,8.694004,10.786053,11.907528,13.145609,14.30138,15.21365,15.769243,14.568888,15.522313,16.345413,15.385129,11.622872,11.63659,10.357354,12.545431,16.352274,13.320518,9.6645775,8.56368,9.4862385,11.074138,11.163307,6.3618846,5.1066556,5.5490727,6.042933,5.130663,8.361334,9.071259,11.173596,13.6086035,10.353925,9.836057,9.321619,9.47595,11.06042,14.915276,12.120162,12.80608,12.857523,10.854645,8.056101,7.8606143,7.3118806,8.114404,9.019815,5.8337283,4.8082814,4.9523244,5.144381,4.7191124,3.457024,4.122364,3.9886103,3.117495,2.2223728,2.668219,3.1449318,2.9117198,2.3664153,1.7662375,1.2312219,1.2758065,1.4061309,1.2998136,1.196926,1.920569,0.9911508,0.4081209,0.18519773,0.21263443,0.274367,0.3806842,0.5144381,0.7956643,1.097468,1.0871792,1.4815818,1.4404267,1.3821237,1.5021594,1.7593783,1.7936742,2.170929,2.3595562,2.4418662,3.0969174,3.4433057,3.3712845,3.0420442,2.6819375,2.5961976,2.5550427,2.3561265,2.4590142,2.6373527,1.99602,1.8656956,1.8965619,2.1434922,2.3458378,1.920569,1.6290541,1.8245405,2.136633,2.4144297,2.726522,3.5461934,3.998899,4.1326528,3.8034124,2.6647894,3.8960114,3.6799474,3.275256,2.9494452,1.9651536,2.860276,3.525616,4.2835546,4.6608095,3.3952916,4.887162,5.926327,6.121814,6.142391,7.740579,8.203573,6.444195,5.3844523,5.861165,6.632822,6.7322803,5.5079174,4.972902,5.3090014,4.8940215,4.629943,4.996909,5.7754254,5.892031,3.4227283,2.702515,3.0214665,3.3129816,3.1277838,2.644212,2.085189,3.292404,3.1277838,1.4369972,1.039165,1.8416885,2.3252604,1.8656956,1.214074,2.4967396,2.7539587,3.6456516,5.4941993,6.667118,3.5804894,4.7774153,7.486789,7.3255987,4.7671266,5.1409516,5.312431,5.754848,7.15069,8.186425,5.5387836,7.8777623,6.355026,5.3158607,5.9571934,6.307011,8.498518,7.9120584,5.6965446,3.6456516,4.180667,3.7279615,3.532475,3.8102717,4.6916757,6.2418494,4.249259,4.7088237,5.9126086,6.5539417,5.7239814,4.99005,3.9611735,4.2046742,5.826869,7.4696417,7.881192,4.506478,2.5378947,3.1586502,3.549623,4.187526,4.139512,4.2218223,4.2595477,3.0900583,3.3198407,3.4638834,3.0351849,2.2395205,2.0097382,2.170929,1.7456601,1.6084765,1.6427724,0.7373613,0.59674823,0.432128,0.5418748,1.2758065,3.0283258,6.385892,9.349055,10.257896,8.968371,6.8385973,3.5804894,3.083199,5.6039457,8.3922,5.662249,4.650521,5.4667625,6.8797526,6.7185616,1.879414,3.0454736,3.2203827,2.8877127,3.1689389,5.830299,9.194724,9.918367,7.0718093,4.5956473,11.276484,5.90575,5.7925735,5.5902276,3.566771,1.5913286,6.5196457,4.822,2.5721905,1.9651536,1.3341095,12.240198,10.175586,6.118384,4.5682106,3.549623,3.3952916,2.1126258,3.5359046,5.7411294,1.0563129,0.77508676,0.9911508,1.0666018,0.864256,0.7510797,0.75450927,1.5158776,2.411,3.083199,3.4467354,3.450165,4.07435,4.341858,4.0229063,3.6353626,3.8274195,4.0263357,4.4516044,5.0483527,5.4941993,5.8680243,6.0635104,5.7068334,5.038064,4.9214582,4.523626,4.681387,4.180667,2.702515,0.8128122,2.5070283,5.0346346,5.6245236,5.130663,8.035523,9.112414,5.7891436,3.1895163,2.8739944,2.8396983,3.7725463,3.9474552,4.6402316,5.73427,5.7377,5.456474,5.6073756,5.2815647,4.40359,3.7279615,2.867135,1.8485477,1.097468,0.7373613,0.6001778,0.31895164,0.1920569,0.26407823,0.823101,2.386993,3.3129816,4.616225,5.15467,4.928317,5.1066556,6.3035817,6.3173003,5.8543057,5.4496145,5.4770513,5.7136927,5.675967,5.6073756,5.5833683,5.528495,4.6848164,4.0366244,3.5702004,3.3301294,3.433017,3.4295874,3.2889743,2.877424,2.633923,3.5530527,3.7211025,4.2115335,4.8768735,5.5559316,6.077229,7.390761,7.4010496,6.9792104,6.619104,6.427047,5.658819,5.689686,6.1458206,6.4716315,5.9434752,4.914599,5.0140567,5.6793966,6.125243,5.3432975,5.120374,4.7362604,4.232111,3.6147852,2.884283,2.527606,2.6613598,2.935727,3.450165,4.729401,2.9734523,2.7333813,3.5016088,4.887162,6.608815,6.7631464,7.31531,7.5690994,7.64798,8.498518,7.7611566,6.931196,6.6396813,6.7665763,6.444195,5.8062916,4.914599,4.1635194,3.758828,3.7176728,3.4021509,3.3781435,3.2855449,3.093488,3.069481,3.199805,3.1586502,3.450165,4.1943855,5.1238036,5.5250654,5.768566,5.7308407,5.7822843,6.7665763,6.9792104,7.349606,7.6514096,7.9292064,8.47451,0.83338976,0.9294182,0.8848336,0.6790583,0.42183927,0.32924038,0.31895164,0.34981793,0.39097297,0.42526886,0.47328308,0.47671264,0.4629943,0.4698535,0.47671264,0.41840968,0.26750782,0.18862732,0.16804978,0.17490897,0.14747226,0.09945804,0.06859175,0.048014224,0.034295876,0.041155048,0.024007112,0.020577524,0.0274367,0.05144381,0.12689474,0.18862732,0.35324752,0.5041494,0.58988905,0.6241849,0.7990939,1.0254467,1.3375391,1.8279701,2.644212,2.9391565,3.40901,3.8617156,4.3109913,4.972902,5.1066556,6.1046658,7.1541195,7.723431,7.5931067,7.98065,9.081548,9.657719,9.205012,7.939495,8.800322,9.897789,10.185875,9.571979,8.9100685,9.417647,9.650859,10.405369,11.574858,12.175035,12.336226,12.339656,12.377381,12.562579,12.922686,11.561139,11.64345,12.511135,13.327377,13.070158,13.018714,13.516005,14.068168,14.750656,16.21509,17.45317,18.358582,18.416885,17.778982,17.243965,17.37429,16.12935,15.145059,15.031882,15.371411,16.105343,16.324837,16.45173,16.37285,15.443433,15.0250225,15.402277,16.489456,17.960749,19.239986,17.919594,16.585485,15.5085945,15.169065,16.266533,17.302269,16.928444,16.341984,15.995596,15.597764,14.438563,14.637479,15.601193,16.698662,17.267973,17.53891,17.384579,17.446312,17.573206,16.839275,16.527182,17.53891,18.492336,18.886738,19.099373,18.44775,18.12194,18.166525,18.272842,17.79613,17.741257,17.78927,17.724108,17.343424,16.441442,15.6252,15.752095,16.12249,16.46888,16.955881,18.434032,19.37031,19.967058,20.327166,20.443771,21.191422,21.849901,22.134558,22.052248,21.911634,22.312897,22.186,22.330044,22.85477,23.170294,23.125708,22.624989,21.517231,20.28258,19.997925,20.018501,18.996485,18.187103,17.754974,16.750105,15.978448,16.112202,16.777542,17.439453,17.384579,15.985307,15.29253,15.350834,16.091625,17.326277,18.293419,18.37573,17.95046,17.576635,18.001905,19.099373,21.35947,23.304047,23.382927,19.967058,18.45804,18.03277,19.140528,20.60839,19.634388,18.406595,18.533491,19.432043,20.303158,20.107672,20.889618,20.845032,20.79016,21.019941,21.301168,21.554956,21.393766,20.872469,20.430052,20.872469,20.827885,20.440342,20.141968,20.138538,20.430052,19.387459,19.11309,19.03078,18.62266,17.405157,17.405157,17.401728,17.995045,19.006773,19.473198,19.164536,19.157675,19.740705,20.670124,21.150267,21.356041,20.94449,20.965069,21.19828,20.152256,20.954779,21.260014,20.824455,19.932762,19.414894,19.102802,18.866161,18.759844,18.54378,17.689812,17.401728,17.7927,17.593784,16.496315,15.141628,15.011304,14.928994,14.671775,14.315098,14.208781,14.349394,14.459141,14.764374,15.237658,15.597764,17.312557,17.929884,17.480608,16.938732,18.214539,17.802988,17.79613,18.070496,18.37916,18.348293,17.665806,17.518333,18.070496,18.79757,18.471758,17.401728,17.233677,16.993607,16.568336,16.719238,15.275383,12.079007,10.103564,9.856634,9.379922,11.2421875,13.083877,14.390549,15.230798,16.263103,14.774663,16.047039,16.523752,14.915276,12.199042,13.1593275,10.48082,10.031544,11.135871,6.5642304,5.5387836,7.3393173,10.275044,12.130451,10.175586,5.754848,5.1409516,5.31929,5.267846,5.98463,8.114404,10.64201,12.792361,13.354814,10.679735,9.585697,8.06639,8.069819,9.753747,11.485688,11.537132,11.849225,11.201033,9.537683,7.9600725,7.8331776,6.989499,7.548522,8.803751,7.2192817,5.0757895,4.8322887,4.3178506,3.5599117,4.804852,4.2286816,2.9803114,2.153781,2.2326615,3.0866287,2.750529,2.3904223,2.0131679,1.6564908,1.3958421,1.7833855,2.0234566,1.7388009,1.3272504,1.9548649,1.2277923,0.6344737,0.28808534,0.216064,0.32924038,0.48357183,0.5796003,0.69963586,0.823101,0.82996017,1.1832076,1.3409687,1.3581166,1.4061309,1.762808,1.8039631,2.1503513,2.3561265,2.435007,2.8225505,3.4364467,3.357566,2.9494452,2.585909,2.633923,2.4761622,2.301253,2.4555845,2.6853669,2.16064,2.0508933,2.0440342,2.1674993,2.201795,1.6942163,1.5021594,1.7010754,2.0337453,2.3629858,2.6647894,3.690236,4.2218223,3.899441,3.018037,2.5241764,3.6936657,3.3198407,2.884283,2.6819375,1.8245405,3.059192,3.450165,3.3232703,3.0900583,3.2512488,5.627953,6.711703,6.866034,6.8111606,7.610255,8.320179,6.7940125,5.5113473,5.4016004,5.8817425,5.7411294,5.171818,4.8768735,4.787704,4.046913,4.256118,4.856296,5.761707,6.029215,3.8445675,4.057202,4.770556,4.4756117,3.275256,2.884283,3.5393343,3.7211025,2.9082901,1.4644338,0.6276145,0.5624523,0.9945804,1.0151579,0.8676856,1.9548649,2.2909644,2.2086544,4.033195,6.866034,6.574519,6.6122446,6.9552035,5.8200097,4.046913,5.103226,4.201245,3.625074,5.0929375,7.0958166,4.90431,4.870014,5.0140567,6.9209075,9.270175,7.8331776,9.537683,8.189855,6.3893213,5.535354,5.8165803,6.217842,4.695105,4.187526,5.6039457,7.8331776,5.5147767,5.0826488,5.813151,6.5367937,5.638242,5.086078,4.6402316,4.5647807,4.712253,4.5099077,6.001778,5.6005163,3.8274195,1.9445761,1.9754424,4.2046742,4.7774153,5.2644167,5.5319247,3.7451096,4.3521466,4.3487167,3.7005248,2.6545007,1.7422304,2.1297739,1.5227368,1.1351935,1.1729189,0.83681935,0.52472687,0.3566771,0.5727411,1.0940384,1.5330256,2.1332035,6.433906,8.337327,6.8900414,6.279575,3.8274195,4.822,8.186425,11.067279,8.838047,7.936065,7.4696417,7.291303,6.245279,2.177788,3.7759757,4.7602673,4.057202,3.3472774,7.085528,7.3084507,7.1266828,5.2815647,3.7759757,7.8777623,6.81802,3.1312134,0.88826317,1.0048691,1.2243627,6.2692857,8.40249,9.469091,8.848335,3.433017,14.894698,9.654288,5.096367,5.5319247,2.2052248,2.726522,3.1415021,5.31929,7.208993,2.8259802,1.1729189,0.89169276,1.2072148,1.546744,1.5433143,1.1489118,1.5981878,2.170929,2.6990852,3.5770597,3.8617156,4.15323,4.170378,3.9508848,3.841138,3.957744,4.016047,4.3281393,4.8837323,5.353586,6.036074,6.0875177,5.3878818,4.5099077,4.722542,4.4859004,4.2869844,3.4295874,1.9411465,0.5693115,1.255229,3.093488,4.4859004,5.312431,6.924337,9.033533,5.178677,2.7745364,3.6696587,4.1360826,4.6573796,4.4584637,4.557922,5.130663,5.528495,4.8322887,4.98662,4.98662,4.513337,3.9371665,3.4364467,2.3835633,1.3581166,0.7133542,0.5453044,0.32581082,0.25721905,0.45956472,1.2312219,3.0454736,2.8122618,4.4241676,5.5113473,5.3741636,5.0140567,6.492209,6.341307,5.610805,5.1855364,5.7754254,5.528495,5.007198,5.188966,5.7582774,5.1100855,4.2252517,3.690236,3.5804894,3.666229,3.3952916,3.8171308,3.782835,3.2546785,2.750529,3.3198407,3.292404,4.0606318,5.1752477,5.977771,5.593657,6.2864337,6.447624,6.252138,6.094377,6.56766,5.7136927,5.2506986,5.195825,5.4941993,6.0154963,4.914599,5.254128,6.252138,6.831738,5.6485305,5.07236,4.7191124,4.413879,3.8925817,2.8225505,2.6476414,2.767677,2.8156912,3.1140654,4.6676683,3.981751,3.642222,3.865145,4.5647807,5.360445,6.619104,7.9086285,8.416207,8.320179,8.762596,8.591117,7.6376915,6.944915,6.8866115,7.164408,6.591667,5.4804807,4.6127954,4.180667,3.8102717,3.3781435,3.3266997,3.3781435,3.3609958,3.223812,3.1380725,3.292404,3.782835,4.496189,5.0929375,4.8768735,5.07236,5.127233,5.188966,6.118384,6.773435,7.1061053,7.281014,7.3393173,7.1987042,0.65162164,0.58988905,0.45270553,0.33609957,0.28465575,0.28465575,0.38754338,0.44927597,0.4972902,0.5555932,0.64133286,0.6001778,0.6001778,0.5693115,0.4698535,0.30866286,0.2194936,0.16119061,0.1371835,0.12346515,0.07545093,0.058302987,0.044584636,0.030866288,0.017147938,0.024007112,0.006859175,0.024007112,0.06859175,0.15090185,0.29837412,0.4046913,0.65848076,0.8265306,0.85396725,0.89169276,1.2758065,1.4472859,1.7730967,2.5070283,3.8171308,3.9714622,4.190956,4.6779575,5.346727,5.802862,6.0086374,6.756287,7.3839016,7.6445503,7.7440085,7.8777623,8.851766,10.076128,10.494537,8.573969,8.652849,9.3936405,9.716022,9.314759,8.656279,8.882631,8.889491,9.417647,10.755186,12.751206,12.71691,12.048141,11.5645685,11.660598,12.298501,10.9541025,11.022695,11.7086115,12.428825,12.812939,13.077017,12.943263,12.566009,12.22648,12.319078,13.296511,14.507155,15.004445,14.575747,13.756075,15.151917,15.782962,15.505165,14.658057,14.030442,15.076467,15.549749,16.29397,16.95931,15.988737,15.29596,15.745236,16.777542,17.936743,18.87302,17.466888,16.108772,15.433144,15.412566,15.3302555,14.973578,14.29452,13.776653,13.776653,14.531162,14.095605,14.325387,15.247946,16.63007,17.971039,19.013634,18.595222,17.576635,16.62321,16.191082,15.038741,15.649208,16.983316,18.190533,18.605513,18.118511,18.145947,18.512913,18.897026,18.849012,18.28313,18.145947,18.145947,17.984756,17.333136,17.168514,17.04162,16.842705,16.70552,17.021042,17.689812,18.214539,18.900457,19.744135,20.443771,20.94792,21.935642,22.583834,22.62156,22.309467,22.354052,22.631847,23.118849,23.671013,24.007113,23.907654,23.132568,22.141417,21.301168,20.903336,20.584383,19.833303,18.948471,18.077356,17.21996,17.075916,16.496315,16.664366,17.720678,18.77699,17.418875,15.539461,14.791811,15.395418,16.12935,16.657507,16.969599,16.96617,16.825556,17.014183,18.176813,20.94449,23.753323,24.648445,21.287449,18.838724,17.549198,17.778982,19.092514,20.265432,19.161106,17.878439,17.261114,17.53891,18.317427,21.479506,22.326614,22.216867,21.825895,21.133118,21.849901,22.371199,22.038528,21.222288,21.332033,21.469217,21.60983,21.184563,20.37175,20.104242,18.849012,18.989626,19.267422,18.814716,17.151367,18.691252,18.677534,19.109661,20.217419,20.45406,20.766151,20.594673,20.567236,20.982216,21.825895,22.213438,21.668133,21.404055,21.242865,19.62067,19.884748,20.179693,20.063087,19.603521,19.387459,19.061647,18.866161,18.667244,18.389448,18.02934,18.060207,18.231688,17.96761,17.20624,16.410576,15.724659,15.076467,14.658057,14.445422,14.188204,13.893259,14.71636,15.621771,15.892709,15.127911,16.969599,18.324286,18.087645,16.808409,16.698662,15.920145,17.04505,18.21111,18.509483,17.991615,17.29198,17.185663,18.228258,19.634388,19.277712,18.012194,18.022482,17.61779,16.47231,15.621771,14.040731,10.940384,11.029553,12.734058,8.220721,12.88839,15.114192,15.484588,15.244516,16.300829,15.662926,16.393429,15.981877,14.359683,13.893259,14.723219,10.707172,7.0135064,5.055212,2.5310357,2.9117198,5.8508763,8.98209,9.668007,4.979761,1.4472859,1.8897027,3.4844608,4.8185706,5.885172,7.689135,12.583157,16.311117,16.276823,11.543991,8.718011,6.252138,6.8043017,9.277034,8.793462,11.413667,10.748327,9.304471,8.303031,7.6925645,8.06296,7.0032177,6.8145905,7.8537555,8.512236,6.9860697,5.3432975,3.275256,2.1503513,5.0243454,3.4227283,2.7059445,2.301253,2.3664153,3.782835,2.4967396,1.7902447,1.5193073,1.5364552,1.6804979,2.2600982,2.3732746,1.8965619,1.4164196,2.2223728,1.5810398,0.90198153,0.4046913,0.216064,0.3566771,0.5727411,0.67219913,0.6379033,0.53844523,0.48700142,0.66533995,1.0494537,1.2792361,1.3889829,1.7902447,1.786815,2.0680413,2.49331,2.8705647,2.9563043,3.1860867,2.8739944,2.568761,2.469303,2.4075704,2.3801336,2.1983654,2.3321195,2.5824795,2.0714707,2.1023371,2.1400626,2.085189,1.8862731,1.5776103,1.3512574,1.5330256,1.8828435,2.2909644,2.784825,3.8308492,4.262977,3.4604537,2.2223728,2.767677,3.2478194,2.9460156,2.6716487,2.6064866,2.3149714,3.4913201,2.9803114,2.620205,3.350707,5.2164025,8.388771,9.578837,9.280463,8.423067,8.354475,7.963502,6.307011,4.8905916,4.297273,4.1943855,3.7759757,4.2081037,4.623084,4.6402316,4.3590055,4.629943,5.0243454,5.2918534,5.113515,4.0880685,5.470192,5.8165803,4.722542,3.0454736,2.9117198,4.9248877,4.482471,2.9734523,1.4129901,0.42526886,0.36696586,1.2895249,1.3752645,0.7613684,1.5604624,1.670209,1.2758065,3.8617156,8.834618,11.526843,6.6431108,4.341858,4.6093655,6.619104,8.735159,5.288424,3.069481,2.884283,3.415869,1.2072148,1.7388009,3.6799474,7.514226,11.201033,10.172156,7.3598948,6.7459984,7.3701835,8.224151,8.2653055,10.30591,7.366754,5.422178,6.358455,7.966932,7.4524937,6.8214493,6.420188,5.844017,3.9337368,6.5367937,7.239859,6.2144127,3.9268777,1.1626302,2.7642474,6.1046658,5.7068334,1.9582944,1.1249046,3.9646032,5.5319247,6.3001523,6.125243,4.232111,5.8988905,5.4770513,4.064061,2.4418662,1.0734608,1.7147937,1.1763484,0.64476246,0.6207553,0.9259886,0.3806842,0.28465575,0.53501564,1.1454822,2.253239,0.91569984,0.47671264,0.53501564,0.6790583,0.45956472,2.4041407,6.447624,8.748878,8.711152,8.964942,10.957532,11.451392,8.368194,3.4433057,2.2326615,3.5153272,6.4236174,6.012067,3.6525106,7.0203657,3.7485392,3.2375305,3.4947495,3.5942078,3.7005248,5.3227196,2.5001693,0.42869842,0.58988905,0.7442205,2.6133456,10.189304,16.599203,16.46545,5.9126086,6.831738,3.192946,2.9906003,5.353586,0.5144381,2.6887965,4.557922,8.038953,10.748327,6.0052075,5.0929375,2.1674993,1.1626302,2.469303,2.9151495,1.8897027,1.7696671,1.7388009,1.7971039,2.7573884,4.2526884,4.2046742,3.9886103,4.07435,4.0057583,3.724532,3.8925817,4.4721823,5.086078,5.0312047,5.73427,5.9880595,5.3673043,4.4104495,4.6127954,4.698535,4.046913,3.2443898,2.3972816,1.1146159,0.9774324,1.4747226,2.3904223,3.457024,4.3624353,3.841138,3.6147852,3.8548563,4.4584637,5.0449233,4.5682106,4.372724,4.4413157,4.73969,5.2335505,4.1017866,4.108646,4.307562,4.180667,3.6353626,3.542764,2.8499873,1.8931323,0.9945804,0.4629943,0.3018037,0.36010668,0.78537554,1.821111,3.8205605,2.7059445,3.940596,5.1580997,5.3673043,4.955754,5.888602,5.802862,5.195825,4.9420357,6.2692857,5.48734,4.280125,4.40359,5.411889,4.6402316,4.341858,3.9097297,3.9611735,4.232111,3.566771,4.280125,4.2355404,3.6627994,3.0420442,3.1072063,3.542764,4.1943855,5.171818,5.778855,4.523626,4.756838,5.586798,6.0497923,5.90232,5.6142344,4.9660425,4.7431192,4.7979927,5.171818,6.090947,5.267846,5.5902276,6.392751,6.715132,5.2987127,4.7979927,4.557922,4.139512,3.4913201,2.959734,2.5756202,2.3904223,2.702515,3.415869,4.033195,5.1100855,4.7774153,4.557922,4.787704,4.633373,7.7131424,8.381912,8.594546,9.023245,9.050681,9.074688,8.604835,7.720001,6.992929,7.466212,6.7048435,5.5319247,4.5784993,4.0880685,3.9063,3.4021509,3.1655092,3.3369887,3.683377,3.6044965,3.3884325,3.707384,4.262977,4.7328305,4.7774153,3.8445675,4.187526,4.65395,4.9077396,5.456474,6.276145,6.783724,6.869464,6.574519,6.0840883,0.31895164,0.22292319,0.24350071,0.26750782,0.2709374,0.31895164,0.45613512,0.6173257,0.70649505,0.6893471,0.5796003,0.5693115,0.58302987,0.47328308,0.2709374,0.19891608,0.1371835,0.10288762,0.07888051,0.05144381,0.01371835,0.0274367,0.020577524,0.01371835,0.01371835,0.0,0.01371835,0.07888051,0.20920484,0.3841138,0.5796003,0.7133542,0.90198153,1.0254467,1.1489118,1.5261664,1.8313997,1.8965619,2.294394,3.316411,4.99005,5.610805,5.686256,5.7582774,5.9983487,6.193835,6.3310184,6.6739774,7.160979,7.781734,8.573969,8.501947,9.3079,10.72432,11.797781,10.8958,9.283894,8.597976,8.573969,8.766026,8.546532,8.275595,8.100685,8.117833,8.539673,9.674867,10.429376,10.39165,10.127572,10.185875,11.077567,13.2862215,13.015285,11.979549,11.362224,11.825217,11.825217,11.588576,11.293632,10.868362,9.962952,10.209882,11.4033785,12.199042,11.924676,10.604284,11.595435,13.1593275,14.225929,14.284232,13.38225,13.248496,12.984418,12.850664,13.169616,14.328816,15.402277,16.338554,17.497755,18.516342,18.310568,18.214539,17.802988,17.223389,16.585485,15.9750185,14.87755,13.924125,13.289652,13.323947,14.555169,14.812388,15.700651,17.165085,18.849012,20.093952,20.766151,20.61525,19.236557,17.446312,17.288551,17.436022,17.096493,17.638369,18.996485,19.668684,19.569225,19.456049,19.425184,19.360022,18.921034,17.809847,17.658945,18.008764,18.310568,17.943602,17.408587,17.171944,17.130789,17.130789,16.983316,17.494326,17.69667,18.142517,18.879879,19.456049,20.35803,21.599543,22.755312,23.36921,22.978235,22.624989,22.985096,23.35206,23.533829,23.849352,24.226606,24.27805,23.725885,22.758743,22.004232,21.674994,20.875898,20.310017,19.905325,18.845583,18.45461,18.025911,17.569777,17.46003,18.44775,18.104792,15.803539,13.96871,13.663476,14.603184,15.103903,15.46744,15.858413,16.475739,17.562918,18.344864,19.901896,22.035099,23.60928,22.583834,20.141968,18.351723,17.178804,16.691803,17.04505,18.30028,17.717249,16.61292,16.143068,17.302269,20.183123,22.093403,22.669573,22.258022,21.925352,21.20514,21.647556,22.035099,21.623549,20.172834,21.637268,21.921923,21.157125,20.008213,19.654966,18.358582,18.437462,18.804428,18.725548,17.823566,20.251715,20.766151,20.906765,21.19828,21.150267,21.404055,22.007662,21.839613,21.229147,21.973368,21.897917,21.94593,21.921923,21.585823,20.646116,20.889618,20.052797,19.589804,19.901896,20.340883,19.630959,19.044498,18.38259,17.96761,18.6158,18.578075,17.881868,17.480608,17.46003,17.04505,15.666355,14.918706,15.13134,15.62863,14.723219,14.284232,15.199932,16.482597,17.226818,16.616352,17.521763,17.545769,17.189093,16.698662,16.0539,16.942162,18.338005,19.11309,19.068506,18.921034,17.175373,16.19794,16.722668,17.960749,17.593784,16.921585,17.03819,17.532051,17.243965,14.267084,13.337666,9.6645775,9.489669,11.96926,9.184435,15.374841,15.741806,14.935853,15.275383,16.739817,16.739817,16.602633,16.026463,14.479718,11.183885,13.810948,9.952662,6.2418494,4.557922,2.0303159,2.9082901,3.758828,4.6573796,4.383013,0.42869842,0.9774324,1.371835,2.8225505,5.4976287,8.498518,10.477389,16.13278,19.709839,19.174824,16.21852,11.118723,9.355915,8.464222,8.011517,9.599416,10.014396,9.266746,8.258447,7.6685576,7.949784,8.292743,7.250148,7.3118806,8.879202,10.268185,8.40249,4.197815,1.6907866,1.9239986,2.959734,2.9220085,2.6133456,2.369845,2.452155,3.0351849,2.037175,1.3649758,1.0837497,1.1317638,1.3272504,1.5844694,1.6393428,1.5536032,1.7833855,3.1723683,2.7093742,1.3855534,0.4389872,0.28465575,0.5041494,0.5658819,0.53501564,0.4972902,0.4629943,0.36696586,0.37725464,0.7579388,1.1043272,1.3512574,1.7559488,1.5364552,1.8656956,2.452155,2.8705647,2.5790498,2.5070283,2.1400626,2.037175,2.1263442,1.7250825,2.2120838,2.3081124,2.4487255,2.5721905,2.1194851,1.9754424,1.9925903,1.8759843,1.6496316,1.6633499,1.3581166,1.3821237,1.6633499,2.136633,2.7470996,3.5873485,3.6696587,3.0248961,2.2669573,2.609916,2.9151495,2.9631636,3.1963756,3.683377,4.1360826,4.341858,3.1209247,3.4707425,5.65539,7.2158523,7.3530354,8.282454,9.6817255,10.81006,10.528833,8.673427,6.2692857,4.5956473,4.280125,5.295283,5.099797,4.914599,4.695105,4.7362604,5.675967,6.262427,5.9880595,5.6142344,5.0655007,3.4192986,4.602506,4.695105,4.746549,4.619654,3.0214665,3.1792276,2.469303,1.646202,1.0460242,0.59674823,0.59674823,1.08032,1.5261664,1.6942163,1.6324836,0.9259886,1.3066728,4.5099077,10.782623,18.87302,9.499957,6.0395036,7.517656,11.495977,14.081886,4.756838,2.5550427,2.9254382,2.9665933,1.4027013,3.8102717,4.629943,5.610805,7.5245147,10.1481495,5.2644167,6.368744,5.7274113,2.428148,2.3801336,8.875772,9.692014,9.373062,8.721441,4.791134,5.206114,9.3936405,9.345626,4.8254294,3.3712845,11.012405,11.550851,8.903209,5.4976287,2.2738166,1.3958421,3.5359046,6.351596,6.7665763,0.9911508,1.4678634,7.2158523,8.865483,5.31929,3.7691166,8.738589,9.366203,6.0326443,1.5261664,1.039165,1.0254467,0.78537554,0.6859175,0.7888051,0.84024894,0.36353627,0.34638834,0.4664239,0.7990939,1.8005334,1.99602,1.155771,1.1694894,1.8142518,0.77851635,1.8039631,3.2855449,2.8156912,1.5570327,4.2423997,5.4016004,5.2335505,5.4976287,5.809721,3.6627994,2.8945718,4.2835546,3.673088,1.7696671,4.149801,6.444195,3.6216443,1.7010754,2.2600982,2.4418662,0.6962063,0.12346515,0.017147938,0.037725464,0.18176813,4.6882463,2.719663,0.4664239,0.16462019,0.07545093,0.6756287,0.4389872,0.12346515,0.024007112,0.0,0.037725464,0.15433143,3.1346428,7.8126,9.095266,16.45516,7.8674736,1.7525192,3.292404,4.4413157,2.6956558,1.4987297,1.3649758,2.0097382,2.3664153,3.4021509,3.5976372,3.549623,3.7142432,4.4104495,3.690236,4.0023284,4.6436615,5.1169443,5.1409516,4.887162,5.1409516,5.1238036,4.722542,4.5167665,4.8940215,4.1017866,3.391862,3.0317552,2.2738166,1.1489118,0.66876954,0.6310441,1.8485477,6.135532,4.2526884,7.2535777,8.090397,5.813151,5.56965,4.8494368,4.064061,3.789694,4.0263357,4.197815,3.525616,3.2272418,3.4673128,3.865145,3.525616,3.6113555,3.3472774,2.6407824,1.5741806,0.42869842,0.35324752,0.42869842,1.1763484,2.5378947,3.8445675,4.417309,4.479041,4.5099077,4.846007,5.675967,4.870014,4.6402316,4.770556,5.0586414,5.3398676,4.804852,4.8425775,5.007198,4.9694724,4.5167665,3.9543142,3.9714622,3.9646032,3.642222,3.0043187,3.1037767,3.1826572,3.0489032,2.9494452,3.5702004,3.5942078,3.6936657,4.3590055,5.07236,4.3041325,5.5730796,5.5319247,5.5079174,5.6039457,4.698535,4.773986,5.147811,5.9400454,6.6053853,5.919468,5.2747054,5.3673043,5.6245236,5.7239814,5.6142344,5.6519604,5.312431,4.386442,3.2272418,2.7779658,2.9117198,2.6785078,3.2409601,4.3281393,4.2423997,6.684266,6.012067,5.2781353,5.4633327,5.4633327,9.002667,8.093826,7.281014,8.124693,9.184435,8.820899,8.573969,7.8949103,7.222711,7.98065,7.1987042,5.703404,4.4996185,3.9200184,3.6010668,3.5633414,3.8205605,4.0949273,4.105216,3.5564823,3.690236,4.1635194,4.3281393,4.029765,3.6147852,3.3952916,4.0023284,4.537344,4.822,5.3707337,5.4084597,6.1321025,6.7185616,6.660259,5.768566,0.2709374,0.33952916,0.4389872,0.45956472,0.42183927,0.48014224,0.41840968,0.47328308,0.548734,0.5761707,0.4938606,0.42526886,0.3806842,0.29837412,0.1920569,0.1371835,0.07545093,0.05144381,0.030866288,0.01371835,0.01371835,0.017147938,0.017147938,0.01371835,0.017147938,0.024007112,0.106317215,0.26407823,0.45956472,0.65505123,0.8128122,0.9568549,1.1249046,1.3341095,1.5810398,1.8416885,2.7230926,3.2718265,3.6113555,4.0777793,5.2335505,5.9743414,5.9743414,5.754848,5.675967,5.9400454,6.200694,6.509357,7.0443726,7.8194594,8.711152,9.253027,9.414218,9.877212,10.542552,10.528833,9.873782,9.259886,8.89635,8.700864,8.275595,8.299602,8.299602,7.8674736,7.2364297,7.257007,8.30646,8.707723,8.889491,9.342196,10.6145735,12.325937,12.867812,12.511135,11.794352,11.495977,12.140739,12.13731,11.893809,11.369082,10.086417,9.949233,10.5597,11.327928,11.760056,11.447963,11.430815,12.3911,13.430264,14.05102,14.164196,14.243076,13.762935,13.63604,14.092175,14.706071,14.150477,14.291091,15.278812,16.400288,16.064188,15.440002,15.638919,15.697222,15.440002,15.46401,15.145059,14.760944,14.490007,14.71636,16.047039,16.62321,16.955881,17.672665,18.718689,19.339443,20.049368,20.851892,20.755863,19.435472,17.226818,16.45516,16.362562,17.178804,18.739265,20.474638,21.294308,21.057667,20.406046,19.840164,19.70298,18.423744,17.641798,17.37429,17.367432,17.089634,16.767254,16.160215,15.892709,16.156786,16.715809,17.089634,17.29541,17.418875,17.583494,17.95389,18.584934,20.234566,21.832754,22.868488,23.406935,23.022821,23.046827,22.967947,22.86163,23.372639,23.304047,23.554407,23.677872,23.403505,22.638706,21.517231,20.773012,20.62897,20.683842,19.905325,18.948471,18.879879,18.8593,18.482046,17.751545,17.926455,16.540901,14.819247,13.598314,13.310229,13.526293,14.102464,14.856973,15.899568,17.658945,18.567787,19.630959,20.502073,20.899906,20.61868,19.53493,18.434032,17.521763,16.750105,15.824117,17.353712,16.986746,15.71094,14.805529,15.837835,18.845583,22.223726,24.27119,24.662163,24.442669,22.480946,20.416334,19.579515,19.895037,19.8676,20.845032,20.917053,20.323736,19.61724,19.654966,19.219408,19.03078,18.547209,17.63494,16.564907,20.2037,21.77788,22.196291,22.168854,22.19972,22.02481,22.391777,22.10712,21.27716,21.287449,22.017952,21.939072,21.294308,20.502073,20.155685,20.478067,19.260563,18.341434,18.427174,19.082224,19.010202,18.79757,18.71526,19.065077,20.189981,18.639809,17.257685,16.671225,16.571766,15.724659,14.970149,14.942713,15.241087,15.391989,14.870691,14.832966,15.254805,16.098484,17.257685,18.581505,17.590355,18.056778,18.739265,18.718689,17.408587,17.010754,17.436022,17.724108,17.494326,16.955881,16.21509,16.077906,16.53747,17.106783,16.78783,16.146498,15.916716,15.21022,14.29452,14.596324,9.928656,7.0478024,6.831738,8.721441,10.710602,13.2690735,14.044161,15.090185,16.527182,16.554619,16.527182,16.732958,15.885849,13.443983,9.623423,10.518545,10.755186,8.875772,5.8200097,4.9351764,5.178677,3.1552205,1.7525192,1.8005334,2.0749004,5.425607,4.040054,4.880303,8.628842,9.657719,14.30138,17.508043,20.131678,21.434921,19.075365,14.754086,9.513676,6.914048,7.4627824,8.608265,8.447074,8.663138,8.416207,7.870903,8.169277,6.5985265,7.157549,8.035523,8.001227,6.4236174,4.3109913,4.2595477,3.450165,2.4658735,5.2781353,3.9337368,2.9151495,2.784825,2.9734523,1.7902447,1.786815,1.3203912,0.9945804,1.1351935,1.7799559,1.3512574,1.2860953,1.7490896,2.760818,4.2115335,2.3904223,1.1660597,0.5212973,0.35324752,0.45613512,0.42869842,0.34638834,0.32924038,0.36696586,0.32924038,0.37039545,0.5007198,0.72021335,1.0357354,1.4369972,1.4438564,1.7696671,2.153781,2.3767042,2.2498093,2.527606,2.153781,1.8656956,1.8108221,1.5638919,2.0337453,2.2566686,2.270387,2.194936,2.2292318,1.8588364,1.8588364,1.7422304,1.5055889,1.6153357,1.4541451,1.4369972,1.4781522,1.7422304,2.6373527,2.9906003,2.7093742,2.287535,2.1469216,2.633923,2.6750782,2.9803114,3.3232703,3.7382503,4.4996185,3.4192986,2.8808534,4.7671266,8.056101,8.827758,8.083538,8.083538,8.961512,10.024684,9.784613,8.008087,5.885172,4.4859004,4.098357,4.232111,4.1943855,3.7759757,3.2032347,3.292404,5.4324665,4.698535,4.314421,4.1155047,3.8308492,3.100347,3.1895163,2.9185789,3.2786856,3.6593697,1.8245405,2.4144297,2.2360911,1.6873571,1.7216529,3.8171308,1.9994495,1.7971039,2.1915064,2.4830213,2.3046827,6.7048435,4.3487167,2.8808534,5.3330083,10.134431,11.698323,10.405369,8.711152,8.371623,10.4705305,4.249259,2.750529,4.064061,5.4599032,3.3815732,3.724532,2.7642474,3.0043187,5.7891436,11.293632,15.405707,12.0138445,7.284444,4.1292233,2.1983654,7.764586,12.771784,13.197053,10.319629,10.72432,7.7680154,8.7283,8.467651,5.895461,3.9337368,8.724871,7.720001,5.8474464,5.2506986,5.288424,5.579939,5.871454,5.844017,4.852866,1.920569,3.2855449,3.6525106,5.346727,6.975781,3.450165,6.866034,4.7499785,2.8088322,2.527606,1.1729189,1.3066728,1.0563129,0.939707,1.039165,1.0117283,0.5727411,0.66876954,0.75450927,0.805953,1.2895249,1.5021594,1.1077567,1.0425946,1.1797781,0.33952916,1.0014396,1.2106444,3.923448,7.099246,3.6936657,7.9772205,6.7528577,5.5319247,5.0174866,1.1111864,0.8093826,5.195825,8.268735,7.2775846,2.7333813,2.4795918,1.3786942,0.7888051,1.0117283,1.2929544,0.45613512,0.116605975,0.23664154,0.58988905,0.7579388,1.4335675,1.4747226,1.0528834,0.44584638,0.041155048,0.94999576,1.0494537,0.64476246,0.22292319,0.45270553,0.09602845,0.030866288,2.335549,8.100685,17.418875,8.069819,2.952875,1.255229,1.6221949,2.1332035,1.5193073,1.1489118,1.1763484,1.5536032,2.0234566,3.275256,3.4295874,3.2718265,3.3712845,4.057202,3.7759757,4.2423997,4.6402316,4.8322887,5.3741636,5.0895076,5.336438,5.377593,4.9523244,4.2835546,4.9077396,4.4104495,3.5599117,2.6545007,1.5158776,2.8156912,1.6564908,0.53501564,1.0082988,3.6936657,3.542764,3.6353626,5.4084597,7.3358874,4.9351764,5.844017,4.180667,3.1243541,3.357566,3.0626216,3.3369887,2.867135,2.6647894,2.959734,3.1826572,3.199805,3.1037767,2.760818,2.037175,0.78194594,0.34638834,0.53501564,1.7010754,3.1483612,3.1380725,4.482471,4.866585,4.746549,4.513337,4.5030484,4.2252517,4.245829,4.383013,4.5682106,4.839148,4.537344,4.636802,4.6916757,4.5201964,4.187526,3.8685746,4.1155047,4.331569,4.1155047,3.2375305,3.5804894,3.7931237,3.7622573,3.782835,4.57164,4.2526884,4.1635194,4.3933015,4.756838,4.7774153,5.0140567,4.6848164,4.636802,5.195825,6.1766872,5.977771,5.206114,4.9694724,5.212973,4.722542,5.0243454,4.822,4.633373,4.8254294,5.6039457,4.9077396,4.8254294,4.3624353,3.4810312,3.117495,2.7951138,2.6373527,3.3301294,4.623084,5.329579,6.0497923,5.6828265,5.4804807,5.8371577,6.2555676,8.604835,9.352485,9.102125,8.916927,10.319629,8.05953,7.0546613,6.550512,6.186976,5.967482,5.302142,4.122364,3.2546785,2.884283,2.527606,2.9185789,3.0797696,3.3129816,3.6147852,3.6525106,3.2992632,3.3266997,3.210094,2.7779658,2.2360911,2.5927682,3.2683969,4.029765,4.5201964,4.2595477,4.297273,4.8151407,5.2301207,5.2815647,5.0346346,0.24007112,0.3566771,0.4629943,0.4629943,0.39783216,0.4355576,0.40126175,0.39097297,0.3806842,0.35324752,0.30866286,0.3018037,0.30523327,0.23321195,0.116605975,0.07545093,0.037725464,0.024007112,0.017147938,0.006859175,0.006859175,0.006859175,0.010288762,0.030866288,0.06859175,0.14061308,0.36353627,0.61046654,0.77165717,0.8711152,1.097468,1.2895249,1.5810398,1.9480057,2.3389788,2.6819375,3.940596,4.7945633,4.9934793,4.8734436,5.3398676,6.0223556,6.7871537,7.133542,6.9209075,6.385892,6.358455,6.3447366,6.5779486,7.2021337,8.2481575,8.958082,8.748878,8.800322,9.445084,10.179015,10.477389,10.13786,9.650859,9.119273,8.255017,8.344186,8.299602,7.7097125,6.9723516,7.257007,7.750868,8.05953,8.464222,9.06097,9.746887,10.528833,11.358793,11.979549,12.421966,12.9981365,13.526293,13.203912,12.490558,11.540562,10.199594,10.405369,10.820349,11.595435,12.408247,12.47341,12.006986,12.240198,13.087306,14.256795,15.275383,15.752095,14.781522,13.944703,13.834956,14.078457,13.817808,13.732068,14.30481,15.182784,15.182784,14.527733,14.29452,14.071597,14.009865,14.822677,15.9613,16.462019,16.2974,15.930434,16.328266,16.993607,18.115082,19.006773,19.243416,18.674105,19.29143,20.015072,20.512363,20.310017,18.79414,17.4566,16.63007,16.859852,18.070496,19.558937,21.019941,21.177702,20.337454,19.281141,19.257133,18.554068,17.669235,16.743246,15.9578705,15.549749,15.755525,15.858413,16.050468,16.348843,16.582056,16.667795,16.732958,16.767254,16.839275,17.082775,17.309128,18.591793,19.980776,21.139977,22.333473,22.36091,22.237446,22.144846,22.179142,22.374628,22.470657,22.566685,22.803328,22.94051,22.384918,21.236006,20.515793,20.124819,19.843594,19.339443,19.054789,19.510923,19.823015,19.480057,18.355152,17.641798,17.03819,15.951012,14.668345,14.339106,13.46799,13.440554,14.352823,15.820687,16.979887,18.053349,19.003344,19.469769,19.346302,18.770132,18.386019,17.854433,17.583494,17.161655,15.3817,16.832415,16.729528,15.9750185,15.453721,16.023033,16.928444,19.648108,22.18943,23.547548,23.69845,22.53925,20.478067,19.480057,19.836735,20.165974,20.652975,20.659836,20.220848,19.53836,18.975908,19.569225,19.476627,18.910746,17.998474,16.80155,19.380598,20.773012,21.218857,21.222288,21.565247,21.53095,21.157125,20.697561,20.3546,20.28601,21.980227,21.901346,20.574095,19.095943,19.12681,18.965618,18.358582,17.79613,17.62808,18.073925,18.742695,18.752985,18.993055,19.750994,20.70442,18.643238,17.521763,16.63007,15.697222,14.928994,14.867262,15.169065,15.563468,15.6869335,15.090185,14.750656,14.760944,15.501736,16.979887,18.845583,17.840714,17.813278,18.20425,18.276272,17.106783,16.70552,16.79126,16.780972,16.585485,16.609491,16.21852,15.769243,15.608052,15.707511,15.642348,15.536031,15.738377,15.673215,15.227368,14.760944,9.105555,8.158989,8.690575,9.719451,12.504276,13.666906,14.613472,15.758954,16.582056,15.621771,16.427725,16.722668,15.549749,13.224489,11.327928,10.693454,9.338767,6.824879,4.1600895,3.8034124,3.5153272,2.3252604,1.4267083,1.5364552,2.8808534,5.07236,4.5647807,5.9743414,9.856634,12.686044,19.143957,18.115082,18.3723,21.4555,21.647556,16.578627,10.203023,6.5127864,6.773435,9.534253,8.628842,8.700864,8.594546,8.131552,8.1041155,6.0326443,6.433906,7.8194594,8.375052,5.9743414,4.979761,4.5853586,4.0434837,3.6319332,4.650521,4.098357,2.901431,2.435007,2.5824795,1.7353712,1.5501735,1.2243627,1.0494537,1.1351935,1.4164196,1.3169615,1.1249046,1.4027013,2.4144297,4.149801,2.1434922,1.08032,0.5727411,0.35324752,0.29494452,0.30523327,0.23664154,0.23664154,0.30866286,0.31895164,0.42183927,0.45613512,0.5178677,0.72021335,1.2037852,1.4678634,1.9548649,2.2223728,2.1297739,1.845118,2.2052248,2.0131679,1.821111,1.7353712,1.4267083,1.728512,2.1503513,2.2223728,2.0097382,2.0920484,1.762808,1.646202,1.4850113,1.3272504,1.5570327,1.529596,1.5776103,1.5364552,1.6016173,2.3149714,2.644212,2.3321195,2.020027,1.99602,2.2360911,2.335549,2.8637056,3.4364467,3.9200184,4.4104495,3.841138,3.7691166,5.9914894,9.561689,10.789482,9.626852,9.0644,8.865483,8.536243,7.346176,6.2830043,4.6265135,3.9268777,4.029765,3.0900583,2.7951138,2.8945718,3.0626216,3.4398763,4.629943,2.9906003,2.49331,2.4624438,2.5378947,2.6750782,3.2066643,2.3664153,2.6785078,3.765687,2.3492675,3.1620796,2.4007113,1.5604624,1.7353712,3.5976372,3.3061223,2.5996273,2.0303159,1.8656956,2.095478,5.2815647,4.681387,3.2512488,3.1140654,5.5319247,7.596536,6.8557453,5.5902276,5.0586414,5.5113473,5.178677,5.137522,7.966932,10.960961,6.135532,4.57507,4.5647807,4.057202,3.5118976,5.90575,13.138749,13.265644,9.349055,4.482471,1.7765263,5.120374,11.574858,13.642899,11.489118,12.956982,8.803751,8.580828,8.656279,7.4936485,5.675967,6.4133286,6.601956,5.3261495,3.940596,6.060081,6.2212715,6.2830043,5.3432975,3.666229,2.6716487,3.4192986,4.0057583,4.887162,6.307011,8.289313,4.540774,2.784825,2.1091962,1.6907866,0.77508676,1.5261664,1.5124481,1.4061309,1.3546871,0.99801,0.8505377,0.7613684,0.8093826,0.9774324,1.1317638,1.7388009,1.471293,1.214074,1.1420527,0.72364295,0.7339317,0.4698535,3.2443898,8.052671,9.541112,10.302481,6.56766,3.9165888,3.2272418,0.6824879,0.5212973,2.4555845,4.040054,3.9028704,1.7662375,1.3752645,0.84367853,0.72021335,0.9294182,0.7888051,0.5796003,0.23664154,0.1371835,0.29837412,0.36010668,0.32924038,0.72364295,0.7373613,0.34638834,0.34295875,0.9431366,0.9568549,0.9294182,0.89169276,0.37382504,0.12689474,0.106317215,0.9602845,3.549623,8.971801,5.56965,2.633923,1.1454822,0.96714365,0.86082643,0.6859175,0.7339317,0.9328478,1.1832076,1.3615463,2.6236343,2.7779658,2.843128,3.1689389,3.4364467,3.426158,4.0846386,4.7671266,5.212973,5.5319247,6.1321025,6.3173003,6.0497923,5.2918534,4.0057583,4.506478,3.9063,3.4055803,3.3232703,3.093488,4.2286816,3.216953,1.8279701,1.196926,1.8108221,2.201795,4.619654,6.39961,6.8454566,7.2295704,4.6676683,2.5996273,1.961724,2.3972816,2.2738166,2.5138876,2.3801336,2.2395205,2.2738166,2.4658735,2.5310357,2.6750782,2.609916,2.0920484,0.90541106,0.36010668,0.7579388,2.1091962,3.5050385,3.1243541,4.1943855,4.5167665,4.523626,4.417309,4.184097,4.081209,4.3178506,4.396731,4.3007026,4.496189,4.32471,4.170378,4.0434837,4.012617,4.214963,4.139512,4.496189,4.5030484,3.99204,3.3952916,4.012617,3.8548563,3.6627994,3.8137012,4.3349986,4.928317,4.729401,4.4584637,4.3109913,3.9371665,3.9063,4.4927597,5.192395,5.6656785,5.7479887,5.751418,5.0483527,4.8117113,5.1855364,5.295283,5.144381,4.8254294,4.846007,5.329579,6.029215,5.3501563,4.962613,4.420738,3.6456516,2.9391565,2.8054025,3.000889,3.690236,4.756838,5.7925735,5.6245236,5.5079174,5.874883,6.6293926,7.140401,7.589677,7.8777623,7.7851634,7.7542973,8.8929205,8.495089,7.1952744,6.15268,5.5593615,4.6573796,4.125794,3.5221863,2.942586,2.49331,2.294394,2.5378947,2.7093742,3.0797696,3.549623,3.6216443,3.000889,2.7985435,2.4761622,1.9754424,1.7079345,2.0406046,2.4007113,2.8088322,3.1620796,3.2409601,3.1895163,3.4981792,3.9543142,4.338428,4.413879,0.28465575,0.3806842,0.42526886,0.42183927,0.37725464,0.31552204,0.33609957,0.34981793,0.31895164,0.25721905,0.22978236,0.23321195,0.2194936,0.15433143,0.06516216,0.034295876,0.01371835,0.010288762,0.010288762,0.006859175,0.0,0.0,0.05144381,0.14061308,0.2469303,0.34638834,0.72707254,0.9602845,1.0597426,1.1249046,1.3375391,1.6290541,2.1640697,2.819121,3.4433057,3.8479972,5.0483527,6.108095,6.478491,6.15268,5.669108,6.420188,7.881192,8.868914,8.755736,7.4936485,7.0923867,6.6225333,6.4373355,6.8111606,7.9257765,8.577398,8.498518,8.498518,8.824328,9.156999,9.832627,10.017825,9.774324,9.201583,8.450503,8.48137,8.594546,8.189855,7.490219,7.56224,7.747438,8.1041155,8.628842,9.283894,9.983529,9.935514,10.268185,11.156448,12.590015,14.390549,15.031882,14.191633,12.850664,11.55771,10.429376,10.624862,11.015835,11.893809,12.926115,13.179905,12.644889,12.284782,12.740917,13.903547,14.932424,15.494876,14.507155,13.564018,13.347955,13.639469,14.754086,14.812388,14.723219,14.805529,14.778092,14.970149,14.270514,13.615462,13.653188,14.750656,16.321407,16.976458,17.075916,16.945591,16.88386,16.86671,18.20425,19.353163,19.52807,18.70497,19.078794,19.425184,19.87446,20.217419,19.901896,18.818146,17.826996,17.487467,17.895588,18.71183,20.076805,20.419764,19.661825,18.495766,18.413456,17.971039,17.353712,16.348843,15.127911,14.249936,14.534592,15.179354,15.999025,16.616352,16.462019,16.564907,16.842705,16.815268,16.578627,16.798119,16.925014,17.665806,18.684393,19.819586,21.112541,21.061096,20.776442,20.587814,20.659836,20.995934,21.671564,22.065966,22.295748,22.316326,21.897917,21.143406,20.19684,19.342873,18.636377,17.892159,17.96761,19.178253,20.066517,19.936192,18.862732,17.778982,17.641798,17.014183,15.906426,15.7795315,14.356253,13.516005,14.13676,15.717799,16.362562,17.412016,18.30028,18.53692,18.097933,17.436022,17.147938,17.12393,17.442883,17.412016,15.594335,16.184223,16.417435,16.403717,16.444872,17.027903,16.647217,17.974468,19.222837,19.816156,20.364891,20.858751,20.340883,20.100813,20.347742,20.2037,20.79016,20.992504,20.766151,20.066517,18.866161,20.056227,19.884748,19.476627,19.12681,18.307138,18.564358,18.982767,19.181683,19.288,19.95334,20.320305,19.490345,19.05136,19.349733,19.497204,21.160555,20.930773,19.428614,17.929884,18.348293,18.399736,18.303709,17.981327,17.71382,18.163095,19.253704,19.456049,19.713268,20.183123,20.220848,18.142517,17.312557,16.338554,15.206791,15.29596,15.309678,15.46744,15.964729,16.307688,15.316538,14.778092,14.661487,15.073037,16.095055,17.78927,18.03963,17.679523,17.4566,17.559488,17.610931,17.093063,16.660936,16.146498,15.673215,15.659496,15.241087,14.435134,13.927555,13.934414,14.198492,14.452282,15.258235,15.676644,15.498305,15.268523,9.774324,9.729739,10.916377,11.838936,13.7526455,14.874121,16.115631,16.80498,16.678083,15.87899,17.312557,16.94902,15.12448,12.9638405,12.370522,9.729739,6.5059276,3.6868064,1.9582944,1.6976458,1.4198492,1.4027013,1.2998136,1.3615463,2.452155,4.108646,6.6225333,8.735159,10.635151,13.975569,19.281141,16.671225,15.12448,17.412016,20.100813,15.717799,11.036412,7.3358874,6.1629686,9.325048,8.083538,8.381912,8.961512,9.088407,8.532814,6.526505,6.725421,8.591117,9.925226,6.8591747,6.8591747,5.5422134,4.7774153,4.7774153,4.125794,3.8925817,2.9288676,2.3595562,2.277246,1.7353712,1.4815818,1.2689474,1.2380811,1.3409687,1.3443983,1.3615463,1.2175035,1.2209331,1.728512,3.1380725,1.6976458,0.9568549,0.5658819,0.32238123,0.15433143,0.21263443,0.17147937,0.18519773,0.26407823,0.2777966,0.41840968,0.4046913,0.3806842,0.52815646,1.08032,1.3615463,1.8382589,2.061182,1.9171394,1.6324836,1.8108221,1.8279701,1.8348293,1.7696671,1.3512574,1.4987297,1.8931323,2.0406046,1.9102802,1.9274281,1.7319417,1.5055889,1.2517995,1.1214751,1.4404267,1.5364552,1.6084765,1.5261664,1.4438564,1.8039631,2.2292318,2.0406046,1.8416885,1.8382589,1.8588364,2.1640697,2.5756202,3.0043187,3.426158,3.9028704,4.057202,4.184097,6.0223556,9.541112,12.922686,10.432805,8.81404,7.798882,6.7357097,4.5853586,5.086078,3.998899,3.82399,4.2938433,2.3732746,2.0920484,2.6716487,3.3678548,3.7142432,3.532475,1.8656956,1.5261664,1.6496316,1.845118,2.1983654,3.1826572,2.6990852,3.2546785,4.3624353,2.534465,3.0866287,2.4898806,2.620205,3.5804894,3.6970954,4.180667,3.642222,2.510458,1.6839274,2.534465,4.8151407,4.8322887,3.5221863,2.4967396,4.0846386,4.629943,5.4941993,5.439326,4.4996185,3.99204,4.90431,7.082098,11.533703,14.726648,8.584257,4.5819287,5.5559316,5.744559,3.8274195,2.9220085,7.0272245,10.755186,10.683165,6.6705475,1.8554068,2.5173173,7.699424,11.177026,11.345076,11.201033,8.971801,7.963502,7.7097125,7.284444,5.3158607,5.295283,5.353586,4.386442,3.2546785,4.791134,5.8474464,5.689686,5.2987127,4.7362604,3.1552205,2.983741,5.9434752,6.9689217,6.036074,8.162418,3.3472774,2.3081124,1.7902447,0.86082643,0.89169276,1.8348293,1.8656956,1.8519772,1.8691251,1.1797781,1.0563129,0.84024894,0.922559,1.2209331,1.1694894,1.7525192,1.8039631,1.605047,1.2895249,0.84024894,0.82996017,0.48014224,1.6873571,4.7328305,8.279024,6.9654922,3.899441,1.9994495,1.6530612,0.72021335,0.99801,1.605047,1.961724,1.9720128,2.0406046,1.7525192,1.1283343,1.1180456,1.5741806,1.2860953,1.3306799,0.5693115,0.041155048,0.07888051,0.34295875,0.26064864,0.37039545,0.38754338,0.3806842,0.7888051,1.3341095,0.99801,0.9911508,1.214074,0.24350071,0.12003556,0.17490897,0.16804978,0.32581082,1.3546871,3.8891523,2.6476414,1.1797781,0.7510797,0.34295875,0.26750782,0.4664239,0.7305021,0.91569984,0.9534253,1.8691251,2.0817597,2.301253,2.6853669,2.843128,3.059192,3.8720043,4.972902,5.8508763,5.7891436,6.7459984,6.931196,6.420188,5.3090014,3.7211025,3.9440255,3.292404,3.0420442,3.3369887,3.216953,4.7945633,5.394741,4.214963,2.0577524,1.3341095,1.371835,5.1409516,6.2864337,4.7259717,6.636252,4.664239,3.57363,2.4658735,1.4610043,1.7010754,1.6427724,1.821111,1.8691251,1.7525192,1.7525192,1.8554068,2.1126258,2.2120838,1.8862731,0.90198153,0.45270553,0.922559,2.1674993,3.5221863,3.7725463,4.338428,4.461893,4.417309,4.297273,3.9954693,4.1017866,4.341858,4.386442,4.2218223,4.15323,4.4413157,4.029765,3.8137012,4.0091877,4.1360826,4.184097,4.245829,3.9440255,3.5118976,3.7794054,4.434457,3.99204,3.7142432,4.0057583,4.4104495,5.2609873,4.9420357,4.40702,4.0846386,3.882293,3.6044965,4.386442,5.4599032,6.1046658,5.6210938,5.7068334,5.3913116,5.4153185,5.885172,6.2898636,5.6348124,5.4496145,5.6142344,5.9469047,6.193835,5.4016004,4.9488945,4.341858,3.5153272,2.8465576,2.8808534,3.3438478,3.923448,4.5956473,5.627953,5.130663,5.147811,5.813151,6.869464,7.671987,7.3221693,7.174697,7.099246,7.099246,7.3255987,8.385342,7.0718093,5.7274113,5.0174866,3.9200184,3.4604537,3.1586502,2.8225505,2.5207467,2.5756202,2.4727325,2.534465,2.8294096,3.192946,3.2272418,2.668219,2.3972816,2.054323,1.7250825,1.9411465,2.095478,1.9720128,1.8485477,1.9068506,2.2326615,2.1297739,2.3492675,3.083199,3.998899,4.2286816,0.36353627,0.39097297,0.3841138,0.40126175,0.4046913,0.2503599,0.29494452,0.33609957,0.32924038,0.274367,0.23664154,0.17833854,0.09602845,0.044584636,0.034295876,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.0034295875,0.0274367,0.15776102,0.32924038,0.5041494,0.65162164,1.0666018,1.2380811,1.3409687,1.4575747,1.5638919,2.037175,2.784825,3.7382503,4.616225,4.931747,5.796003,6.941485,7.6925645,7.582818,6.3653145,6.9963584,8.532814,9.757176,9.942374,8.862054,8.399059,7.613684,7.0718093,7.1678376,8.100685,8.450503,8.803751,8.838047,8.4264965,7.654839,7.9292064,8.56025,8.827758,8.680285,8.738589,8.748878,8.995808,8.831187,8.162418,7.438775,7.699424,8.3922,9.019815,9.6817255,11.063849,10.504827,10.134431,10.64201,12.151029,14.222499,15.079896,14.171056,12.7272,11.444533,10.491108,10.261326,10.597425,11.526843,12.668896,13.21763,13.049581,12.442543,12.500846,13.176475,13.272504,13.282792,12.795791,12.569438,12.864383,13.433694,15.693792,16.21166,15.752095,14.959861,14.321958,15.402277,14.750656,14.064738,14.085316,14.599753,15.515453,15.827546,16.37285,17.20624,17.586924,16.925014,17.566347,18.674105,19.459478,19.188541,19.263992,19.384027,19.408035,19.387459,19.565796,19.068506,18.581505,18.193962,18.073925,18.478617,19.013634,19.140528,18.602083,17.761833,17.61779,16.993607,16.54433,15.810398,14.706071,13.478279,13.392539,13.975569,15.189643,16.417435,16.462019,16.811838,17.45317,17.370861,16.722668,16.839275,17.04848,17.484037,18.317427,19.356592,20.076805,19.69955,19.325726,18.907316,18.746124,19.46634,20.649546,21.678423,22.137987,22.004232,21.647556,21.308027,20.02193,18.79757,17.826996,16.46888,16.317978,18.03963,19.469769,19.675543,18.965618,18.344864,18.279701,17.689812,16.702091,16.640358,15.659496,14.435134,14.46943,15.659496,16.2974,17.031332,17.63494,17.610931,16.94902,16.13278,15.947581,16.479168,17.161655,17.336565,16.232237,15.618341,16.11906,16.63007,17.014183,18.104792,18.46147,18.732407,17.78927,16.335125,16.897577,18.344864,19.473198,20.334024,20.749004,20.327166,21.397196,21.843042,21.839613,21.297739,19.843594,20.773012,20.296299,20.052797,20.382038,20.313446,18.320856,17.487467,17.195951,17.29198,18.104792,18.739265,18.11165,17.95732,18.62266,19.061647,19.77843,19.281141,18.193962,17.384579,17.96418,18.756414,18.948471,18.831865,18.831865,19.476627,20.361462,20.831314,20.95135,20.62211,19.565796,17.864721,16.87357,16.002455,15.518884,16.55119,15.999025,15.6869335,16.05733,16.499744,15.37827,15.227368,15.340545,15.278812,15.268523,16.194511,17.78927,17.737827,17.38115,17.586924,18.722118,17.144508,16.208231,15.433144,14.664916,14.044161,13.570878,12.79922,12.439114,12.672326,13.145609,13.317088,14.267084,14.308239,13.72178,14.740367,10.7586155,10.854645,12.38424,13.80409,14.699212,16.026463,17.446312,17.737827,17.110212,17.20967,18.37573,17.065628,14.678635,12.308789,10.755186,6.615674,3.8960114,2.1091962,1.0014396,0.53501564,0.5212973,0.69963586,0.67219913,0.6344737,1.3478279,3.6868064,8.567109,10.7586155,10.367643,12.867812,14.637479,13.169616,11.273054,11.108434,14.201921,12.38767,10.847785,8.237869,5.885172,7.7851634,6.9209075,7.870903,9.297611,9.97324,8.796892,7.2775846,8.014946,10.196163,11.451392,7.864044,8.224151,6.941485,5.8680243,5.425607,4.5956473,3.8617156,3.2032347,2.7470996,2.393852,1.821111,1.7319417,1.8073926,1.8176813,1.7422304,1.7593783,1.4781522,1.4987297,1.3752645,1.2380811,1.8005334,1.1249046,0.78194594,0.5418748,0.3018037,0.1097468,0.16462019,0.14061308,0.16462019,0.23664154,0.22978236,0.34981793,0.31209245,0.28808534,0.432128,0.90198153,1.0014396,1.2826657,1.5398848,1.6530612,1.605047,1.5776103,1.7525192,1.9068506,1.8519772,1.4404267,1.4575747,1.6221949,1.7319417,1.7490896,1.7833855,1.728512,1.4232788,1.0666018,0.91569984,1.3032433,1.4335675,1.5021594,1.4027013,1.2312219,1.2826657,1.6804979,1.6770682,1.670209,1.7765263,1.8416885,2.2223728,2.2429502,2.201795,2.3595562,2.952875,3.549623,3.649081,4.8014226,7.689135,12.133881,8.937505,6.8145905,5.8645945,5.1580997,2.702515,4.5922174,4.15666,4.2286816,4.6882463,2.4452958,2.2360911,2.8945718,3.5804894,3.6696587,2.7470996,1.646202,1.4953002,1.762808,2.2052248,2.860276,3.666229,3.99204,4.6848164,5.007198,2.6476414,2.5619018,2.719663,4.0229063,5.6005163,4.7945633,4.1943855,4.1429415,3.433017,2.5413244,3.6182148,6.217842,4.8082814,2.9254382,2.510458,3.8925817,4.698535,7.6274023,8.165848,5.977771,4.90431,3.083199,7.191845,12.103014,13.917266,9.983529,4.372724,5.4839106,6.8145905,5.7925735,3.7622573,2.9906003,6.550512,9.47938,8.851766,3.789694,2.9563043,5.7136927,8.3922,9.115844,7.8126,8.282454,6.6431108,5.662249,5.456474,3.4981792,4.8734436,3.3815732,3.0248961,4.2835546,4.105216,5.586798,4.8940215,5.271276,6.200694,3.4295874,3.2992632,7.589677,9.2153015,6.5024977,3.1723683,2.9185789,1.961724,1.0048691,0.66876954,1.5021594,2.1846473,2.16064,2.3492675,2.609916,1.7147937,1.371835,1.1420527,1.2998136,1.6359133,1.4472859,1.5021594,1.821111,1.8348293,1.3409687,0.52472687,0.9294182,0.6379033,0.2777966,0.17490897,0.35324752,0.29494452,0.44584638,0.67219913,0.805953,0.6207553,1.2929544,2.819121,3.6010668,3.2958336,2.7882545,2.2120838,1.4164196,1.4369972,2.1572106,2.311542,2.0817597,0.97400284,0.22292319,0.2777966,0.7888051,0.52472687,0.37039545,0.490431,0.8162418,1.0597426,1.7559488,1.2209331,0.91227025,1.0254467,0.5212973,0.274367,0.24007112,0.19891608,0.18176813,0.48357183,1.6907866,2.0714707,1.9720128,1.704505,1.529596,0.4629943,0.34981793,0.5212973,0.6756287,0.8505377,1.2758065,1.5638919,1.8416885,2.1572106,2.486451,2.9254382,3.7759757,5.0346346,6.135532,5.960623,6.6636887,6.708273,6.060081,4.8734436,3.4878905,3.4021509,2.942586,2.702515,2.6613598,2.177788,4.602506,7.517656,6.7665763,3.0351849,1.8554068,1.1900668,3.3644254,4.2423997,3.433017,4.290414,6.029215,5.8988905,3.724532,1.1146159,1.4644338,1.2072148,1.3581166,1.4164196,1.2689474,1.1797781,1.2998136,1.5055889,1.646202,1.5193073,0.88826317,0.58302987,0.96714365,1.961724,3.2889743,4.4859004,4.8425775,4.852866,4.557922,4.108646,3.7794054,4.0777793,4.105216,4.1429415,4.187526,3.9371665,4.7808447,4.389872,4.262977,4.5647807,4.1120753,4.0194764,3.5804894,3.1106358,3.1106358,4.256118,4.7088237,4.331569,4.187526,4.5853586,5.07236,5.305572,5.0346346,4.530485,4.1943855,4.57164,4.149801,4.307562,5.147811,6.1321025,6.0875177,6.1046658,5.9812007,6.2144127,6.8111606,7.267296,6.5882373,6.591667,6.526505,6.210983,6.012067,5.1169443,4.7808447,4.1360826,3.223812,3.0043187,2.884283,3.3266997,3.7348208,4.1155047,5.0929375,4.8082814,4.804852,5.377593,6.4098988,7.4113383,7.4284863,7.6376915,7.8331776,7.7611566,7.1198235,7.610255,6.3173003,5.1580997,4.5956473,3.6216443,3.2272418,2.8225505,2.585909,2.5961976,2.8465576,2.4761622,2.2978237,2.301253,2.4212887,2.5653315,2.3286898,2.0817597,1.8554068,1.8416885,2.3904223,2.4315774,2.1229146,1.8485477,1.7490896,1.7182233,1.6187652,1.8965619,2.836269,4.057202,4.513337,0.34981793,0.25378948,0.32924038,0.39097297,0.3841138,0.39783216,0.48357183,0.3566771,0.20920484,0.12689474,0.09259886,0.041155048,0.01371835,0.006859175,0.01371835,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.1371835,0.30523327,0.4629943,0.66533995,1.0666018,1.1900668,1.4781522,1.728512,1.8691251,1.9685832,2.7128036,3.3850029,4.341858,5.2987127,5.3090014,6.1149545,7.1232533,7.874333,8.025234,7.3530354,6.7459984,7.56224,8.429926,8.961512,9.764035,9.997248,9.403929,8.7283,8.443645,8.772884,8.323608,8.766026,8.519095,7.421627,6.773435,6.0052075,6.3173003,7.0135064,7.822889,8.89635,9.153569,8.601405,8.152129,7.9737906,7.5210853,7.425057,8.371623,9.139851,9.647429,10.940384,10.096705,10.233889,10.871792,11.485688,11.537132,11.427385,11.873232,11.880091,11.067279,9.674867,9.599416,9.637141,10.216741,11.30049,12.373952,13.3033695,12.96727,13.032433,13.430264,12.343085,11.039842,10.8958,11.327928,11.907528,12.360233,13.7526455,15.134769,15.683503,15.103903,13.625751,13.615462,13.612033,13.622321,13.392539,12.3911,13.111313,14.105893,14.935853,15.635489,16.70895,17.600643,17.86815,18.684393,19.70298,19.044498,18.969048,19.171394,18.852442,18.11165,17.929884,16.914726,16.204802,16.438013,17.429163,18.173384,17.576635,17.436022,17.178804,16.811838,16.921585,16.496315,15.343974,14.153908,13.306799,12.878101,12.744347,13.032433,14.123041,15.741806,16.938732,17.1205,17.384579,17.439453,17.192522,16.753534,16.523752,17.113642,18.169954,18.989626,18.54035,18.989626,18.986197,18.612371,18.159666,18.11165,18.941612,19.919044,21.071384,22.011093,21.925352,21.561817,20.323736,18.969048,17.689812,16.12935,16.153357,17.147938,18.166525,18.855871,19.456049,18.831865,18.430603,17.658945,16.774113,16.859852,16.88386,16.352274,16.05733,16.307688,16.907866,17.065628,16.931873,16.907866,16.338554,13.519434,14.606613,15.885849,16.78783,17.099922,16.952452,16.12249,16.520323,16.928444,17.264544,18.571217,21.085104,21.37319,19.901896,17.936743,17.532051,17.350283,18.320856,19.582945,20.79016,22.11055,23.060547,23.235455,23.304047,23.11542,21.699,21.270302,20.687271,20.676983,21.20514,21.482935,18.993055,17.20967,16.256245,16.153357,16.80155,17.079346,17.288551,17.549198,17.988186,18.708399,18.927893,18.37916,17.87158,17.672665,17.501184,17.940172,19.041069,20.207129,21.050808,21.393766,21.270302,22.155134,22.350622,21.44521,20.310017,19.723558,18.056778,17.04505,17.134218,17.501184,16.355703,15.645778,15.193072,14.949572,15.001016,15.951012,16.619781,16.681513,16.12249,15.244516,16.523752,17.29541,17.892159,18.183672,17.562918,13.780083,13.519434,14.027013,14.057879,13.886399,13.71492,13.1593275,13.066729,13.526293,13.855534,13.622321,13.564018,12.977559,11.664027,9.918367,10.81006,12.9809885,15.001016,16.191082,16.616352,17.093063,17.71382,17.703531,17.233677,17.439453,17.12393,15.9921665,14.232788,11.399949,6.4098988,3.9303071,3.998899,3.8137012,2.5001693,1.0837497,0.58302987,0.6962063,0.548734,0.28808534,1.0666018,1.9239986,3.4364467,4.616225,6.3961806,11.657167,10.803201,8.868914,7.8983397,7.997798,7.3393173,7.888051,7.689135,6.852316,6.258997,7.5519514,7.822889,8.519095,8.985519,8.601405,6.8043017,6.7322803,8.608265,10.377932,10.635151,8.621983,9.208443,8.052671,6.4716315,5.2781353,4.791134,4.6436615,3.8034124,2.952875,2.627064,3.1895163,2.4452958,3.3369887,3.2958336,2.1160555,1.9685832,1.7730967,1.786815,1.4815818,1.0185875,1.2517995,0.8471081,0.7305021,0.59674823,0.36696586,0.18176813,0.17147937,0.15090185,0.16804978,0.22978236,0.29151493,0.3018037,0.34295875,0.31209245,0.24350071,0.30523327,0.40126175,0.6207553,0.99801,1.3992717,1.4953002,1.704505,2.0028791,2.1126258,1.9891608,1.8313997,1.6221949,1.7079345,1.587899,1.3169615,1.5261664,1.5981878,1.2243627,0.8265306,0.75450927,1.2655178,1.1934965,1.4129901,1.4061309,1.1489118,1.097468,1.1832076,1.4267083,1.704505,2.0097382,2.4247184,2.3767042,2.1469216,1.9068506,1.7079345,1.4644338,2.8328393,2.8088322,3.3198407,4.040054,2.3801336,3.5393343,4.417309,4.856296,4.482471,2.702515,3.566771,3.8857226,4.32471,4.605936,3.4947495,2.3458378,2.7299516,3.5290456,3.8925817,3.234101,2.2326615,1.5707511,2.0063086,3.8479972,6.9723516,7.239859,6.759717,5.994919,5.3844523,5.3090014,4.6882463,3.99204,2.7230926,1.9857311,4.5030484,2.8156912,2.3767042,2.9322972,3.789694,3.8137012,3.1792276,2.061182,2.054323,2.8328393,2.136633,4.1635194,5.7308407,6.276145,5.1100855,1.4507155,1.670209,5.3227196,7.4284863,7.579388,9.932085,6.989499,8.333898,7.7851634,4.372724,2.335549,4.2869844,4.170378,3.3781435,4.1463714,9.551401,10.844356,13.155897,9.9869585,4.1635194,7.8126,6.0532217,5.147811,4.787704,4.729401,4.791134,2.935727,2.3252604,4.180667,7.4970784,9.047252,5.178677,4.5784993,3.9131594,2.784825,3.724532,5.895461,7.5107965,7.394191,5.6485305,3.6456516,0.9259886,0.20920484,0.22635277,0.53844523,1.5261664,2.3081124,2.767677,3.2546785,3.4844608,2.534465,2.277246,1.937717,2.0714707,2.4830213,2.2292318,1.8725548,1.4095604,1.2209331,1.1592005,0.548734,0.4629943,0.31552204,0.17490897,0.1097468,0.18176813,0.37725464,0.37382504,0.36696586,0.4972902,0.84024894,0.5453044,0.8848336,1.1180456,1.1797781,1.6770682,1.3238207,0.9534253,0.96371406,1.5158776,2.5173173,1.3341095,1.0460242,0.90541106,0.65162164,0.5178677,0.8128122,0.7476501,1.1454822,1.646202,0.71678376,0.77851635,0.8848336,0.8162418,0.8265306,1.6324836,0.97400284,0.5144381,0.3566771,0.44584638,0.5796003,1.3478279,3.3266997,4.98662,5.874883,6.6053853,1.5776103,0.15433143,0.12003556,0.3018037,0.59674823,0.9602845,1.2346514,1.8142518,2.5001693,2.486451,3.1209247,3.7931237,4.5613513,5.2644167,5.5079174,6.632822,5.8508763,4.8322887,4.170378,3.4021509,3.0248961,2.8945718,2.7402403,2.9117198,4.3624353,4.4241676,8.182996,7.915488,3.357566,1.7079345,0.7682276,0.70649505,3.4192986,7.500508,8.268735,5.778855,2.9254382,1.7388009,2.1469216,1.9514352,1.587899,1.2586586,0.922559,0.65505123,0.65505123,0.8505377,0.9911508,1.0597426,1.0597426,1.0220171,0.6207553,0.9568549,1.8725548,3.069481,4.1189346,4.7774153,4.9523244,4.5990767,4.033195,3.9371665,3.923448,3.673088,3.649081,3.9371665,4.2423997,4.852866,5.0312047,5.161529,5.2506986,4.945465,4.273266,3.7931237,3.426158,3.4021509,4.256118,4.513337,4.513337,4.671098,5.0483527,5.3398676,5.535354,5.9126086,5.5593615,4.523626,3.8137012,4.2423997,4.715683,5.3741636,5.90575,5.5387836,5.8680243,5.593657,6.1321025,7.5725293,8.683716,8.182996,7.9909387,7.4010496,6.464772,6.012067,6.169828,5.212973,4.040054,3.2478194,3.1140654,2.6133456,2.6887965,2.9220085,3.3952916,4.715683,5.3878818,5.206114,5.3707337,5.9571934,5.919468,5.7754254,6.543653,7.8126,8.903209,8.865483,7.658269,6.1286726,5.1752477,4.7088237,3.6456516,3.4776018,2.819121,2.311542,2.2120838,2.3972816,2.0063086,1.670209,1.5536032,1.7113642,2.0920484,2.1743584,1.9411465,1.786815,1.8656956,2.061182,2.0234566,2.5447538,3.2272418,3.525616,2.7299516,2.620205,3.0146074,3.4433057,3.9268777,4.99005,0.37382504,0.36696586,0.35324752,0.28808534,0.22292319,0.32238123,0.34981793,0.20920484,0.09945804,0.06516216,0.017147938,0.017147938,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.006859175,0.017147938,0.06516216,0.22292319,0.39440256,0.61046654,0.8162418,1.039165,1.371835,1.7799559,2.07833,2.2120838,2.2258022,2.2841053,3.2272418,4.098357,4.839148,5.4016004,5.785714,6.2418494,6.948344,7.610255,7.922347,7.56224,7.1678376,7.582818,8.172707,8.796892,9.825768,9.530824,9.115844,8.951223,8.889491,8.261876,8.289313,8.683716,8.615124,7.915488,7.0923867,5.579939,5.48734,6.0326443,6.711703,7.298162,7.699424,7.390761,7.0958166,7.0546613,7.034084,7.1129646,7.449064,7.9463544,8.525954,9.146709,9.417647,10.110424,10.796341,11.207891,11.266195,12.456262,12.349944,11.585147,10.772334,10.504827,10.508256,10.329918,10.549411,11.2421875,11.982979,12.325937,12.020704,11.914387,11.941824,11.0981455,10.456812,10.319629,10.449953,10.700313,11.005547,11.537132,12.668896,13.687484,13.96871,12.977559,11.873232,11.612583,11.862943,11.986408,11.022695,11.410237,11.986408,12.826657,13.708061,14.109323,14.911846,15.525743,16.650646,17.909306,17.833855,18.221397,19.065077,19.582945,19.510923,19.11309,18.187103,17.484037,17.511473,18.087645,18.344864,17.638369,17.412016,17.243965,17.089634,17.274832,17.326277,16.54433,15.666355,14.898128,13.903547,13.330807,13.083877,13.485138,14.579176,16.108772,17.29541,17.580065,17.36057,16.96274,16.619781,16.575195,16.808409,17.63151,18.571217,18.392878,18.36544,18.71526,18.728977,18.303709,17.940172,18.12537,18.746124,19.62067,20.388897,20.498644,20.749004,20.025362,18.986197,17.977898,17.021042,15.9613,16.208231,16.914726,17.669235,18.492336,17.63494,17.099922,16.979887,17.010754,16.568336,16.877,16.96274,17.21996,17.55263,17.357141,17.466888,17.189093,17.03819,16.602633,14.544881,14.438563,15.265094,16.252815,17.069057,17.830425,16.835844,17.343424,17.785841,17.947031,18.962189,21.815605,22.748453,22.371199,21.270302,19.997925,19.668684,20.36832,20.917053,21.229147,22.292318,23.139427,23.35206,23.647005,23.818485,22.734735,21.342323,20.159115,19.658396,19.853882,20.299728,18.44432,16.986746,16.160215,16.060759,16.63007,16.753534,17.243965,17.717249,18.067066,18.475187,18.224829,17.844143,18.025911,18.660385,18.831865,18.550638,18.550638,19.401176,20.941061,22.309467,22.69358,22.306036,20.958208,19.514353,19.881319,19.37374,18.46147,17.768692,17.405157,16.938732,15.71437,15.361122,15.011304,14.654627,15.134769,15.549749,15.71094,15.9750185,15.954441,14.500296,14.246507,15.028452,15.402277,14.812388,13.584596,13.011855,13.416546,13.248496,12.583157,13.104454,13.101024,12.343085,11.856084,11.914387,12.048141,13.320518,13.433694,13.207341,13.032433,12.847235,13.035862,14.46257,15.340545,15.350834,15.6526375,16.568336,16.698662,16.355703,15.96816,16.098484,15.889278,15.237658,12.281353,7.48336,3.6147852,7.0443726,6.0669403,4.787704,5.3878818,8.152129,4.2423997,2.2566686,1.99602,2.6990852,3.069481,1.2895249,1.0871792,1.4164196,2.7711067,7.2021337,6.036074,6.5127864,7.466212,7.421627,4.5922174,6.667118,8.069819,7.73372,6.375603,6.468202,7.222711,10.278474,9.80862,6.492209,7.490219,7.3290286,7.599966,8.4093485,9.342196,9.47595,8.615124,8.399059,8.412778,7.905199,5.754848,5.9126086,4.448175,3.0351849,2.7059445,3.8720043,3.1586502,3.8034124,3.9611735,3.1380725,2.201795,2.9803114,2.6785078,1.6873571,0.8196714,1.2758065,0.72707254,0.51100856,0.42183927,0.34295875,0.26750782,0.17833854,0.18862732,0.19548649,0.18862732,0.22978236,0.38754338,0.45613512,0.42526886,0.33609957,0.28122616,0.36010668,0.44584638,0.6962063,1.0254467,1.0940384,1.3478279,1.8348293,2.054323,1.9480057,1.9171394,1.6393428,1.605047,1.471293,1.2620882,1.3924125,1.6324836,1.2758065,0.89855194,0.7682276,0.8505377,1.1797781,1.2346514,1.1592005,1.0837497,1.1214751,1.0631721,1.4918705,1.8176813,1.8828435,1.9754424,1.5055889,1.3512574,1.430138,1.488441,1.0871792,2.726522,2.2223728,2.037175,2.6133456,2.369845,4.7191124,4.8014226,3.923448,3.0489032,2.7985435,2.8637056,3.2821152,3.6182148,3.7176728,3.7005248,2.8088322,2.702515,2.609916,2.3629858,2.417859,2.1194851,2.0268862,2.6236343,4.2183924,6.9723516,6.4407654,5.4496145,4.3281393,3.6147852,4.0880685,5.147811,3.192946,2.0063086,2.5207467,2.8294096,2.0131679,1.8999915,1.978872,1.9480057,1.7388009,1.8279701,2.1332035,2.194936,1.9445761,1.6976458,1.3512574,1.646202,2.1674993,2.3972816,1.6942163,6.601956,8.97866,9.537683,9.078118,8.491658,7.7680154,7.438775,5.7822843,3.309552,2.7745364,6.574519,5.761707,3.415869,2.0920484,3.841138,11.7257595,11.458252,7.531374,4.9934793,9.434795,6.2727156,7.0923867,5.9434752,3.223812,5.7068334,5.3158607,3.3301294,4.197815,7.208993,6.4716315,5.9126086,4.537344,4.012617,4.091498,2.5996273,2.6236343,2.836269,3.0043187,2.7539587,1.5707511,0.5178677,0.4389872,0.5590228,0.83338976,1.9411465,2.8396983,3.3952916,3.7211025,3.7313912,3.1312134,3.2855449,2.867135,2.3664153,2.054323,1.9823016,2.4212887,2.1469216,1.6736387,1.3375391,1.2929544,0.7407909,0.61046654,0.42869842,0.13032432,0.08573969,0.1920569,0.28122616,0.52815646,1.155771,2.4247184,2.4555845,2.3321195,2.760818,3.4810312,3.2786856,2.5927682,2.369845,2.061182,2.428148,5.56965,3.0077481,1.9445761,1.5844694,1.4164196,1.2037852,0.66533995,0.5555932,0.8848336,1.4507155,1.8519772,1.670209,1.3546871,1.097468,1.0666018,1.4129901,0.65505123,0.40126175,0.37382504,0.5007198,0.89855194,2.3595562,2.153781,2.952875,4.698535,4.5819287,2.7059445,0.922559,0.06516216,0.14747226,0.34981793,0.6001778,0.881404,1.5193073,2.393852,2.9391565,3.2889743,3.8308492,4.383013,4.7774153,4.887162,5.4736214,5.470192,5.360445,5.0895076,4.0846386,3.0248961,2.74367,2.8980014,2.901431,1.9239986,2.6373527,3.865145,4.5510626,3.9371665,1.587899,0.75450927,1.0631721,1.7593783,2.49331,3.350707,4.355576,3.2889743,2.6819375,3.0146074,2.7230926,2.4452958,1.6599203,1.0082988,0.7305021,0.6927767,0.8505377,0.9362774,1.0185875,1.0837497,1.0460242,0.5658819,0.7099246,1.5261664,2.877424,4.4241676,4.6848164,4.4927597,4.314421,4.2766957,4.170378,3.82399,3.6387923,3.666229,3.9543142,4.523626,4.98662,5.4016004,5.377593,4.9180284,4.417309,3.532475,3.0729103,2.8499873,2.884283,3.426158,4.249259,4.57507,4.8905916,5.40503,6.060081,6.667118,5.9400454,5.1512403,4.5784993,3.508468,3.974892,4.605936,5.336438,5.857735,5.6005163,5.0312047,5.90232,6.7494283,7.438775,9.146709,7.394191,6.8283086,6.3618846,5.7479887,5.5593615,6.5882373,6.169828,5.099797,3.8925817,2.7711067,2.7573884,2.9117198,2.9117198,3.100347,4.506478,4.5922174,4.098357,4.173808,5.0826488,6.1904054,5.3501563,5.2266912,5.717122,6.7219915,8.169277,6.9209075,5.353586,4.273266,3.8308492,3.5016088,3.0660512,2.4830213,2.2463799,2.2635276,1.8691251,1.5673214,1.4815818,1.5364552,1.6084765,1.529596,1.7113642,1.605047,1.9925903,2.7951138,3.0489032,3.1483612,3.2718265,3.3198407,3.2203827,2.9254382,3.391862,3.4398763,3.6387923,4.3349986,5.662249,0.2709374,0.30523327,0.24350071,0.16119061,0.12003556,0.17833854,0.16119061,0.08573969,0.034295876,0.020577524,0.0,0.0034295875,0.006859175,0.0034295875,0.0034295875,0.010288762,0.010288762,0.030866288,0.09259886,0.22635277,0.45613512,0.8093826,1.0425946,1.2037852,1.4369972,1.978872,2.352697,2.702515,2.8156912,2.760818,2.867135,3.6970954,4.6848164,5.446185,5.878313,6.1801167,6.2898636,6.7048435,7.160979,7.473071,7.514226,6.8728933,6.691125,7.1884155,8.069819,8.532814,8.323608,8.4093485,8.553391,8.340756,7.1884155,7.689135,8.330468,8.275595,7.5450926,7.006647,5.5730796,5.103226,5.3981705,6.012067,6.2555676,6.5710897,6.7391396,6.831738,6.869464,6.800872,7.459353,7.9772205,8.162418,8.083538,8.076678,9.071259,9.918367,10.323058,10.600855,11.667457,13.502286,13.780083,12.9638405,11.592006,10.264755,10.052121,10.041832,10.446524,10.995257,10.943813,11.842365,11.712041,11.485688,11.4376745,11.201033,10.717461,10.583707,10.662587,10.88551,11.231899,11.4205265,12.133881,12.854094,13.176475,12.843805,11.818358,11.05699,10.792912,10.984968,11.321068,11.032983,11.293632,12.277924,13.491997,13.797231,14.174485,14.445422,15.083325,15.937293,16.221949,16.29054,17.573206,19.243416,20.522652,20.663265,19.70298,18.77699,18.547209,18.79071,18.396307,17.254255,16.756964,16.777542,17.233677,18.077356,17.662374,17.288551,16.719238,15.858413,14.747226,13.906977,13.543441,13.677195,14.315098,15.450292,16.942162,17.412016,17.185663,16.592344,15.981877,16.026463,16.105343,16.846134,18.008764,18.492336,18.516342,19.11309,19.322296,18.77699,17.70696,17.37772,17.782412,18.413456,18.831865,18.629519,18.893597,18.989626,18.821575,18.320856,17.436022,16.242527,15.9921665,16.37971,17.106783,17.87501,16.695232,15.728088,15.604623,16.115631,16.20137,16.750105,16.904436,17.137648,17.346853,16.86671,16.856422,17.364002,17.586924,17.04505,15.580616,15.12448,14.990726,15.409137,16.45173,18.03277,17.288551,17.470318,17.943602,18.492336,19.315437,20.893047,22.244305,22.978235,22.868488,21.832754,21.568676,21.77102,21.839613,21.699,21.798458,21.94936,22.5221,23.18744,23.554407,23.170294,22.258022,20.841602,19.579515,18.917604,19.099373,17.768692,16.582056,16.002455,16.047039,16.273392,16.609491,17.144508,17.487467,17.63151,17.96761,17.662374,17.638369,18.139088,19.03078,19.805868,19.847023,19.020493,18.886738,20.186552,22.8582,23.427511,22.563255,20.738716,19.020493,19.071936,17.741257,16.973028,16.6335,16.341984,15.481158,15.049029,14.730078,14.555169,14.647768,15.21365,14.79867,14.730078,14.997586,15.062748,13.838386,13.320518,13.433694,13.245067,12.641459,12.360233,12.600305,12.517994,12.459691,12.710052,13.485138,13.193623,12.662037,12.397959,12.63803,13.354814,14.452282,13.972139,13.310229,13.05301,12.977559,13.070158,13.488567,13.87954,14.404267,15.748666,16.45173,15.728088,14.983868,14.613472,14.013294,13.677195,12.020704,8.440215,4.2389703,2.620205,4.5201964,5.223262,5.1992545,5.4599032,7.548522,8.879202,5.0655007,2.4761622,2.6750782,2.417859,2.1126258,1.9994495,2.1812177,3.6285036,8.165848,6.1286726,7.0718093,7.2432885,5.641671,4.016047,5.7822843,7.407909,7.8503256,7.0135064,5.7377,6.351596,7.997798,8.014946,6.8591747,8.080108,7.671987,7.5245147,7.641121,8.189855,9.496528,9.462232,9.784613,10.14472,9.554831,6.3618846,6.2144127,4.914599,3.9783216,3.9268777,4.273266,3.8720043,4.6093655,5.171818,4.7945633,3.2649672,3.6456516,3.6182148,2.386993,0.78537554,1.2449403,0.5796003,0.36353627,0.32238123,0.29494452,0.25378948,0.22292319,0.25721905,0.2709374,0.25378948,0.26750782,0.3841138,0.41840968,0.4424168,0.4355576,0.29151493,0.32924038,0.42526886,0.61046654,0.83681935,0.96371406,1.0288762,1.4610043,1.7765263,1.8176813,1.7833855,1.5261664,1.546744,1.5947582,1.5398848,1.3958421,1.5947582,1.2792361,1.0323058,0.97400284,0.764798,1.097468,1.1934965,1.1317638,1.0082988,0.94656616,0.980862,1.4644338,1.8691251,1.9857311,1.9171394,1.8759843,1.5433143,1.3341095,1.3272504,1.2380811,2.3389788,2.8088322,2.7333813,2.2909644,1.7422304,3.350707,3.474172,3.0146074,2.7745364,3.4638834,3.5187566,3.6970954,4.0709205,4.4996185,4.623084,3.7279615,3.2718265,2.8328393,2.3664153,2.201795,1.8897027,2.719663,3.6593697,3.9886103,3.3129816,3.1723683,2.5550427,1.9651536,1.8176813,2.4212887,2.5927682,1.7353712,2.1880767,3.8171308,4.012617,3.100347,3.0111778,2.9151495,2.5893385,2.4384367,2.2669573,2.5550427,2.8877127,2.6785078,1.1763484,2.0508933,2.4590142,4.0263357,5.9914894,5.223262,7.0032177,6.999788,7.407909,8.2653055,7.48336,7.208993,8.615124,9.225591,8.073249,5.703404,6.2212715,5.6793966,4.1463714,2.4075704,1.9720128,6.1732574,6.807731,5.130663,4.3349986,9.530824,8.594546,6.2830043,4.6127954,4.290414,4.7362604,5.8405876,3.415869,3.2718265,5.778855,5.892031,5.7891436,5.593657,4.3590055,2.4247184,1.4232788,1.0494537,0.82996017,0.8265306,0.85739684,0.5041494,0.23664154,0.548734,0.89512235,1.3546871,2.620205,3.3061223,4.249259,4.588788,4.0949273,3.1723683,3.2203827,3.2855449,3.0077481,2.5447538,2.5619018,2.6922262,2.4658735,2.1057668,1.821111,1.8005334,0.9534253,0.7339317,0.70649505,0.59674823,0.29151493,0.18519773,0.4046913,0.77851635,1.2620882,1.9342873,2.3389788,2.8225505,3.8171308,4.6882463,3.7313912,3.4021509,3.4433057,4.0194764,5.1752477,6.8283086,4.4927597,3.2615378,2.7128036,2.393852,1.8313997,1.3855534,1.1317638,1.2620882,1.9857311,3.508468,2.0577524,1.587899,1.4575747,1.371835,1.4129901,0.9534253,0.7133542,0.59674823,0.5761707,0.7099246,1.7182233,1.845118,2.5996273,4.431027,6.728851,2.6167753,0.6859175,0.061732575,0.07545093,0.23664154,0.4389872,0.6824879,1.3238207,2.3801336,3.5187566,3.7931237,4.262977,4.6573796,4.7808447,4.5030484,4.5339146,4.756838,4.928317,4.8425775,4.331569,3.3541365,2.7539587,2.6819375,2.6853669,1.7147937,2.3904223,2.7951138,4.166949,5.003768,1.0631721,0.5796003,1.1592005,2.0028791,2.4727325,2.1194851,2.5447538,2.0886188,2.095478,2.8122618,3.3712845,3.415869,2.3835633,1.4095604,0.97057325,0.8848336,0.91569984,0.94656616,0.9568549,0.9362774,0.91569984,0.5693115,0.6207553,1.255229,2.5207467,4.307562,4.928317,4.619654,4.125794,3.8479972,3.8788633,3.508468,3.4467354,3.5016088,3.7862647,4.722542,5.4187484,5.686256,5.535354,5.0929375,4.5819287,3.765687,3.3472774,3.1620796,3.2409601,3.8137012,4.99005,5.302142,5.545643,5.8337283,5.5902276,6.9209075,6.2144127,5.4496145,5.079219,4.029765,3.5873485,3.7313912,4.1017866,4.48933,4.8288593,3.9680326,4.7842746,5.778855,6.557371,7.8434668,6.9071894,6.029215,5.2026844,4.647091,4.7979927,5.7274113,5.693115,4.9934793,3.957744,2.9494452,2.6785078,2.8739944,2.9871707,3.1415021,4.108646,4.383013,3.82399,3.899441,5.0140567,6.48535,5.98463,5.7891436,5.8234396,6.2247014,7.363324,6.6053853,4.996909,3.5393343,2.8225505,3.0351849,2.2841053,1.937717,1.8965619,1.9445761,1.7216529,1.3306799,1.3443983,1.4164196,1.3581166,1.1420527,1.3066728,1.471293,2.0440342,2.8980014,3.3884325,3.923448,3.8205605,3.6627994,3.7553983,4.1120753,4.383013,4.0023284,3.8342788,4.15666,4.6402316,0.17490897,0.18519773,0.12003556,0.06516216,0.05144381,0.0548734,0.034295876,0.017147938,0.006859175,0.0,0.006859175,0.006859175,0.0274367,0.034295876,0.020577524,0.0274367,0.037725464,0.09602845,0.22978236,0.4355576,0.70306545,1.2826657,1.4129901,1.5673214,1.9857311,2.644212,2.8534167,3.1895163,3.3884325,3.426158,3.508468,4.166949,5.1169443,5.7891436,6.0635104,6.2658563,6.2418494,6.5470824,6.684266,6.5985265,6.6636887,5.8817425,5.689686,6.186976,6.9792104,7.2021337,7.517656,7.9292064,7.9120584,7.2638664,6.121814,6.433906,7.2775846,7.500508,6.9723516,6.560801,5.6313825,5.1100855,5.360445,6.060081,6.200694,6.416758,6.660259,6.697984,6.6225333,6.831738,7.747438,8.56368,8.453933,7.64798,7.459353,8.752307,9.482809,9.774324,10.199594,11.770344,13.38568,13.985858,13.54687,12.157887,10.017825,9.788043,9.945804,10.449953,10.878652,10.405369,11.540562,11.646879,11.489118,11.454823,11.571428,11.146159,11.039842,10.909517,10.844356,11.348505,10.813489,11.173596,11.921246,12.614022,12.88839,12.0309925,11.111863,10.700313,11.159878,12.651748,12.504276,12.493987,12.994707,13.762935,13.937843,14.452282,14.476289,14.760944,15.488017,16.276823,15.80011,16.516893,18.070496,19.771572,20.62554,20.53294,19.984205,19.62753,19.360022,18.317427,16.79469,15.724659,15.549749,16.269962,17.463459,17.487467,17.508043,17.278261,16.763824,16.13621,15.001016,14.387119,14.267084,14.538021,15.0250225,16.170506,16.828985,16.952452,16.61292,16.012743,15.933864,15.927004,16.407146,17.28512,17.96418,18.608942,19.579515,19.915615,19.318867,18.145947,17.470318,17.525192,17.775553,17.813278,17.38115,17.28169,17.477179,17.885298,18.197392,17.885298,16.811838,16.280252,16.331696,16.7844,17.21996,16.252815,15.079896,14.634049,15.028452,15.542891,16.180794,16.143068,15.999025,15.927004,15.700651,15.927004,17.195951,18.0362,17.864721,16.990177,16.012743,15.018164,14.706071,15.450292,17.305698,17.480608,17.655516,18.180243,18.979338,19.569225,19.733847,21.12283,22.648996,23.564695,23.468666,23.214878,23.019392,22.810186,22.309467,21.016512,21.225718,22.172283,22.988525,23.393215,23.681301,23.074265,21.843042,20.268862,18.924463,18.677534,17.305698,16.221949,15.810398,15.971589,16.108772,16.527182,16.993607,17.099922,16.96617,17.223389,17.247395,17.401728,17.885298,18.735836,19.823015,20.2037,19.318867,18.900457,19.843594,22.223726,22.799898,22.017952,20.69413,19.45262,18.739265,16.911295,15.933864,15.484588,15.13134,14.328816,14.315098,13.982429,14.184773,14.79524,14.706071,14.081886,13.824667,13.594885,13.371962,13.471419,12.922686,12.531713,12.164746,11.910957,12.061859,12.295071,12.089295,12.1921835,12.672326,12.912396,12.127021,12.185325,12.445972,12.823228,13.783512,14.05102,13.173045,12.614022,12.644889,12.377381,12.466551,12.4974165,13.210771,14.575747,15.830976,16.21852,15.062748,13.543441,12.103014,10.419086,10.179015,8.385342,5.703404,3.309552,2.9082901,3.1415021,4.5956473,5.768566,6.001778,5.4907694,10.007536,6.842027,3.9063,3.5530527,2.5756202,2.5756202,3.1243541,3.9131594,5.171818,7.6616983,6.210983,7.239859,6.341307,3.7039545,4.139512,5.8062916,7.48336,7.870903,7.1678376,7.0923867,8.330468,6.8385973,7.0306544,9.14328,9.208443,8.687145,8.4093485,8.134981,8.213862,9.599416,10.045261,10.360784,9.935514,8.471081,5.970912,5.5730796,4.7328305,4.417309,4.7088237,4.7774153,4.7945633,5.2987127,6.0737996,6.2075534,4.0880685,4.2835546,3.9646032,2.5927682,0.97400284,1.2449403,0.58988905,0.33609957,0.29494452,0.31552204,0.2777966,0.33609957,0.4081209,0.42183927,0.39097297,0.44584638,0.39783216,0.37039545,0.4081209,0.4389872,0.28122616,0.32581082,0.42183927,0.58988905,0.77165717,0.83681935,0.7888051,1.138623,1.4575747,1.5776103,1.5741806,1.4644338,1.5707511,1.7559488,1.8039631,1.4129901,1.5776103,1.3341095,1.1592005,1.1111864,0.8265306,1.0288762,1.1626302,1.1214751,0.94656616,0.82996017,0.9362774,1.3924125,1.7971039,1.9857311,2.0508933,2.201795,2.0268862,1.670209,1.3478279,1.3375391,2.085189,3.199805,3.5016088,2.8808534,2.2909644,2.7230926,2.843128,2.9322972,3.2203827,3.8925817,4.0777793,4.15666,4.557922,5.1238036,5.1169443,4.5990767,3.625074,2.877424,2.5173173,2.1743584,2.335549,3.1449318,3.9714622,3.8377085,1.4267083,2.277246,1.8519772,1.6804979,2.3458378,3.4947495,1.3478279,0.89512235,3.3712845,6.776865,5.861165,3.8514268,2.9803114,2.620205,2.935727,4.880303,2.7745364,2.2978237,2.5001693,2.3561265,0.7613684,2.4212887,3.216953,4.8734436,6.6636887,5.394741,4.2595477,3.4810312,3.9268777,5.06893,4.976331,4.955754,8.8929205,11.619442,11.177026,8.81747,6.200694,4.8151407,4.2698364,3.8479972,2.5070283,2.1023371,4.4927597,5.9880595,6.433906,9.239308,7.3530354,4.0537724,3.1826572,4.3521466,2.942586,5.802862,5.302142,4.3487167,4.4687524,5.7891436,6.0806584,5.7925735,3.9200184,1.3375391,0.77508676,0.39097297,0.1920569,0.10288762,0.082310095,0.1371835,0.13375391,0.5418748,1.0528834,1.845118,3.590778,4.0777793,4.9831905,5.2335505,4.5510626,3.457024,3.2992632,3.625074,3.5873485,3.1517909,3.117495,3.175798,2.8499873,2.4795918,2.1503513,1.7216529,1.214074,0.82996017,0.7476501,0.86082643,0.77851635,0.33609957,0.432128,0.7133542,0.9877212,1.2277923,1.6942163,2.8019729,4.046913,4.804852,4.307562,4.695105,4.822,5.5147767,6.694555,7.3564653,4.897451,4.057202,3.4021509,2.6545007,2.6716487,2.633923,2.3904223,2.452155,3.0351849,4.0880685,2.2223728,1.7696671,1.7971039,1.7353712,1.3958421,1.8931323,1.2517995,0.6824879,0.59674823,0.61389613,1.0185875,1.4575747,1.9857311,3.117495,5.8337283,1.8176813,0.3841138,0.061732575,0.05144381,0.19891608,0.66191036,0.881404,1.3169615,2.1983654,3.5050385,4.07435,4.6882463,5.103226,5.120374,4.5922174,4.016047,3.9851806,4.081209,4.0229063,3.6765177,3.433017,2.6785078,2.386993,2.5584722,2.2292318,2.177788,2.3218307,3.865145,4.931747,0.5693115,0.4115505,1.3032433,2.5584722,3.3369887,2.6407824,2.0577524,1.611906,1.8313997,2.7230926,3.7622573,4.1326528,3.1826572,2.095478,1.4232788,1.0734608,0.97057325,0.922559,0.8848336,0.864256,0.939707,0.607037,0.58302987,1.0357354,2.0749004,3.7553983,4.5682106,4.40702,3.8205605,3.309552,3.3301294,3.175798,3.2546785,3.5221863,4.1292233,5.442755,5.871454,6.0086374,5.950334,5.675967,5.0312047,4.4996185,4.07435,3.7794054,3.8137012,4.547633,5.5490727,5.717122,6.042933,6.4887795,5.9812007,7.0032177,6.948344,6.4064693,5.627953,4.4996185,3.2889743,3.0660512,3.3061223,3.806842,4.695105,3.457024,3.7519686,4.8082814,5.8645945,6.1766872,5.7308407,4.938606,4.122364,3.7211025,4.314421,4.465323,4.5922174,4.3487167,3.765687,3.2443898,2.6956558,2.6956558,2.8705647,3.100347,3.5221863,4.0434837,3.8857226,4.122364,5.0449233,6.1801167,5.7822843,5.6519604,5.6039457,5.6073756,5.813151,5.4941993,4.4275975,3.1037767,2.136633,2.2635276,1.5913286,1.4404267,1.5433143,1.6496316,1.5364552,1.2209331,1.3101025,1.3478279,1.1660597,0.89169276,1.2003556,1.5981878,2.0714707,2.6167753,3.223812,3.882293,3.865145,3.882293,4.2081037,4.6779575,4.9523244,4.431027,3.9028704,3.7348208,3.858286,0.1097468,0.072021335,0.037725464,0.020577524,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.017147938,0.017147938,0.017147938,0.061732575,0.07545093,0.0548734,0.06516216,0.09259886,0.22978236,0.4355576,0.6927767,1.0151579,1.6290541,1.646202,1.8519772,2.4418662,3.0489032,3.1620796,3.474172,3.8205605,4.07435,4.15323,4.6402316,5.288424,5.720552,5.888602,6.108095,6.090947,6.3893213,6.228131,5.645101,5.5079174,4.9214582,5.192395,5.545643,5.7582774,6.1458206,6.9826403,7.606825,7.431916,6.48535,5.4187484,5.06893,5.90575,6.4819202,6.293293,5.768566,5.40503,5.1855364,5.562791,6.3378778,6.6533995,6.927767,6.701414,6.2212715,5.98463,6.7391396,7.675417,8.608265,8.323608,7.181556,7.1061053,8.30646,8.920357,9.290752,9.80519,10.8958,11.753197,12.445972,12.600305,11.931535,10.261326,10.055551,10.268185,10.618003,10.813489,10.539123,11.283342,11.660598,11.852654,11.952112,11.986408,11.578287,11.321068,10.703742,10.103564,10.816919,9.6645775,9.746887,10.690024,11.88352,12.487128,11.760056,11.194174,11.4033785,12.504276,14.143619,14.637479,14.493437,14.246507,14.164196,14.2533655,15.148488,15.251375,15.481158,16.208231,17.240536,16.61292,16.568336,17.027903,17.926455,19.21255,20.53637,20.800447,20.467777,19.692692,18.348293,16.486027,14.79524,14.153908,14.63062,15.453721,16.743246,17.144508,17.254255,17.388008,17.573206,16.311117,15.422854,14.994157,14.898128,14.79524,15.090185,15.79325,16.46545,16.808409,16.674654,16.475739,16.341984,16.348843,16.585485,17.137648,18.358582,19.61724,20.02193,19.5315,18.95876,18.358582,18.0362,17.826996,17.556059,17.024471,16.492886,16.060759,16.403717,17.394867,18.108221,17.439453,16.87357,16.684942,16.808409,16.856422,16.39,15.316538,14.544881,14.4317045,14.791811,15.412566,15.21022,14.688923,14.29795,14.441993,15.29939,16.811838,18.04306,18.437462,17.820137,16.331696,15.066177,14.284232,14.393978,15.971589,17.20967,17.909306,18.560926,19.250275,19.651537,19.006773,20.052797,21.86705,23.68473,24.888515,24.658733,24.243753,23.917942,23.228596,20.975357,21.575535,22.679861,23.424082,23.719027,24.254042,23.310905,22.477516,21.098822,19.469769,18.818146,17.38115,16.506605,16.21166,16.311117,16.427725,16.417435,16.595774,16.61292,16.47231,16.554619,17.130789,17.315987,17.586924,18.173384,19.05136,19.377169,19.140528,19.360022,20.162544,20.762722,20.896477,20.495214,20.080235,19.62753,18.571217,17.106783,15.933864,15.035312,14.3974085,14.040731,13.807519,13.522863,14.030442,14.754086,13.71492,13.570878,13.097594,12.250486,11.80464,13.337666,12.627741,12.329367,12.349944,12.38424,11.914387,12.0138445,12.068718,11.910957,11.509696,10.984968,10.583707,11.47197,12.168177,12.38767,13.029003,11.962401,11.032983,11.30735,12.360233,12.291641,12.46998,12.80265,14.057879,15.62863,15.542891,15.505165,14.020154,11.458252,8.546532,6.385892,8.512236,8.128122,6.2247014,4.15323,3.6353626,4.3692946,4.770556,6.166398,7.8023114,6.848886,7.596536,6.632822,6.042933,5.90232,4.2698364,2.510458,3.2855449,4.513337,4.98662,4.372724,4.6676683,6.018926,5.0586414,2.7573884,4.420738,6.5196457,8.515666,8.193284,6.989499,10.014396,11.633161,7.997798,7.9463544,11.664027,10.659158,10.131001,9.836057,9.654288,9.671436,10.179015,9.493098,9.088407,7.6788464,5.65539,5.0757895,4.705394,4.547633,4.7808447,5.3330083,5.871454,5.8337283,5.3878818,6.0737996,6.989499,4.7945633,4.6608095,3.4913201,2.1263442,1.2312219,1.3169615,0.6962063,0.36696586,0.29837412,0.37382504,0.37725464,0.490431,0.6241849,0.6207553,0.548734,0.7099246,0.4972902,0.39440256,0.37039545,0.3566771,0.2503599,0.3566771,0.39783216,0.5418748,0.72364295,0.64476246,0.61389613,0.9259886,1.1626302,1.2346514,1.371835,1.4472859,1.5776103,1.7765263,1.8485477,1.3889829,1.587899,1.4575747,1.2929544,1.1592005,0.90884066,0.96714365,1.0700313,1.0185875,0.84367853,0.7990939,0.9362774,1.3272504,1.6221949,1.7971039,2.1674993,2.1332035,2.3458378,2.1229146,1.5021594,1.2312219,1.937717,2.877424,3.4878905,3.625074,3.5599117,3.2272418,3.1895163,3.4433057,3.789694,3.8514268,4.2183924,4.3178506,4.5339146,4.852866,4.863155,5.0620713,3.6627994,2.6853669,2.5927682,2.277246,3.0077481,2.9048605,3.275256,3.707384,2.0817597,3.7142432,3.5050385,3.350707,4.0606318,5.353586,1.8039631,0.8471081,4.0263357,8.23444,5.7239814,3.0454736,1.8142518,1.4815818,2.5824795,6.7391396,2.6167753,1.4027013,1.4472859,1.5398848,0.89855194,1.7971039,2.620205,3.1277838,3.0351849,2.0063086,1.3032433,1.4232788,1.546744,1.4987297,1.7353712,2.2120838,6.958633,9.767465,9.331907,9.22902,7.116394,5.857735,6.478491,7.641121,5.6313825,2.352697,4.8288593,7.822889,8.803751,7.9429245,3.069481,2.201795,2.9940298,3.3850029,1.6016173,5.2164025,7.222711,5.9812007,3.8479972,7.174697,7.6205435,5.4599032,3.3472774,2.0886188,0.6310441,0.17147937,0.09259886,0.14061308,0.18519773,0.22292319,0.24350071,0.5761707,1.1832076,2.2463799,4.15323,4.712253,5.2301207,5.3673043,4.98662,4.139512,3.8479972,4.081209,4.0366244,3.6044965,3.3541365,3.789694,3.3952916,2.8396983,2.270387,1.3203912,1.5776103,1.1317638,0.764798,0.7990939,1.1077567,0.5453044,0.45956472,0.50757897,0.61389613,0.9602845,1.2483698,2.4830213,3.5804894,4.273266,5.099797,5.967482,5.8165803,5.7102633,6.2487082,7.5690994,4.386442,4.012617,3.590778,2.8225505,3.9337368,4.1429415,4.0949273,4.3590055,4.8425775,4.763697,3.4124396,2.4658735,2.0337453,1.8725548,1.371835,2.6716487,1.704505,0.85396725,0.8745448,0.89855194,0.9602845,0.939707,1.0117283,1.3512574,2.1263442,1.3615463,0.64476246,0.1920569,0.11317638,0.40126175,1.1729189,1.3546871,1.4267083,1.7971039,2.8054025,3.8205605,4.729401,5.288424,5.3913116,5.038064,4.201245,3.7108135,3.4913201,3.2855449,2.6373527,3.1140654,2.503599,2.270387,2.6545007,2.6545007,1.6736387,1.4781522,2.5481834,3.350707,0.31552204,0.39097297,1.5776103,2.8225505,3.5873485,3.8445675,3.1860867,2.3664153,2.2909644,3.0454736,3.8685746,4.4687524,3.8308492,2.8705647,2.0406046,1.3169615,1.097468,0.91912943,0.84367853,0.90541106,1.1283343,0.66533995,0.5555932,0.85739684,1.6564908,3.0523329,3.5942078,3.7108135,3.40901,2.935727,2.7813954,2.8637056,3.0317552,3.6319332,4.8288593,6.5813785,6.351596,6.5470824,6.728851,6.5162163,5.593657,5.353586,4.8768735,4.389872,4.2835546,5.0895076,5.994919,5.994919,6.3790326,7.1884155,7.222711,7.0032177,7.5382333,7.2604365,5.9434752,4.705394,3.1346428,2.7230926,3.0420442,3.7931237,4.8151407,3.6147852,3.3644254,4.07435,5.099797,5.164959,4.396731,3.8720043,3.415869,3.2272418,3.875434,3.192946,3.3232703,3.4673128,3.3712845,3.3301294,2.8465576,2.5550427,2.6304936,2.935727,3.0386145,3.4604537,3.7691166,4.1600895,4.65395,5.099797,4.5167665,4.461893,4.5510626,4.48933,4.081209,3.8720043,3.6627994,2.959734,1.9582944,1.5227368,1.214074,1.1523414,1.3169615,1.4918705,1.2826657,1.155771,1.3649758,1.4335675,1.2106444,0.8471081,1.371835,1.7696671,1.9823016,2.16064,2.651071,3.1963756,3.4913201,3.8342788,4.2183924,4.3349986,4.791134,4.4721823,3.8171308,3.3850029,3.8308492,0.0,0.0,0.0,0.01371835,0.0274367,0.01371835,0.01371835,0.01371835,0.041155048,0.06859175,0.030866288,0.030866288,0.020577524,0.041155048,0.08916927,0.1371835,0.18519773,0.44584638,0.7373613,1.0528834,1.5398848,1.5776103,1.786815,1.978872,2.2052248,2.7916842,3.1209247,3.5873485,4.046913,4.4584637,4.897451,5.0826488,5.0277753,5.31929,5.90232,6.0737996,5.8405876,5.90232,5.720552,5.3741636,5.56965,5.422178,5.597087,5.3158607,4.681387,4.6676683,5.329579,6.6636887,7.548522,7.2158523,5.2506986,4.7602673,5.4153185,5.6176643,5.0346346,4.6093655,4.557922,4.73969,5.038064,5.4804807,6.2247014,6.824879,5.9400454,5.120374,5.0895076,5.7377,7.349606,8.272165,8.1212635,7.274155,6.8969,7.7268605,8.621983,8.841476,8.515666,8.635701,9.074688,10.2921915,11.129011,11.201033,10.8958,9.966381,10.285333,10.504827,10.333347,10.528833,11.115293,11.818358,12.672326,13.330807,13.059869,12.329367,11.348505,10.127572,9.325048,10.254466,10.449953,10.158438,10.041832,10.316199,10.741467,10.912948,10.984968,12.257345,14.2533655,14.695783,14.5243025,14.644339,14.846684,15.193072,16.03675,16.012743,16.170506,16.0539,15.676644,15.518884,15.848124,17.230247,17.816708,17.676094,18.79757,20.323736,20.714708,20.409475,19.750994,18.982767,16.407146,14.654627,14.027013,14.147048,13.975569,15.343974,16.163645,16.516893,16.719238,17.302269,16.70552,16.300829,15.769243,15.110763,14.647768,13.831526,14.284232,15.275383,16.221949,16.722668,16.955881,16.582056,16.187653,16.331696,17.576635,18.005335,18.825006,19.143957,18.883308,18.79757,19.164536,18.907316,18.506054,18.015623,17.075916,16.414005,15.62863,15.440002,16.033321,17.058767,17.864721,17.607502,17.487467,17.768692,17.806417,17.03819,15.985307,15.172495,14.767803,14.572317,15.230798,15.230798,14.791811,14.232788,13.975569,15.4914465,16.71238,17.442883,17.319416,15.79325,15.196502,14.606613,13.958421,13.725209,14.908417,16.081335,17.480608,18.44432,18.917604,19.456049,18.636377,19.109661,20.683842,23.019392,25.619019,25.85223,25.214327,24.86108,24.68617,23.331484,22.477516,23.36921,24.164873,24.226606,24.154585,22.971376,22.271742,20.971928,19.1954,18.279701,18.279701,18.406595,18.44432,18.183672,17.439453,16.21852,15.577187,15.892709,16.678083,16.554619,17.580065,18.101362,18.214539,18.173384,18.416885,18.526632,19.013634,19.87446,20.567236,20.018501,18.578075,18.54035,18.392878,17.689812,17.04505,16.654078,15.830976,14.867262,14.225929,14.5414505,14.150477,13.917266,13.982429,13.972139,12.9707,13.227919,12.603734,12.109874,12.264205,13.107883,12.373952,12.840376,13.416546,13.341095,12.205902,11.828648,11.084427,10.014396,9.054111,9.016385,11.80121,13.557159,14.143619,14.064738,14.479718,10.854645,9.537683,10.439664,12.3911,13.121602,14.013294,14.575747,15.275383,15.848124,15.275383,14.116182,10.984968,7.5931067,5.23698,4.822,15.22051,16.79469,11.327928,4.0503426,3.6456516,4.341858,3.765687,5.0312047,9.170717,15.151917,6.0840883,4.804852,6.4990683,7.5416627,5.4770513,3.415869,3.1655092,2.760818,2.0303159,2.5790498,3.1655092,4.722542,4.90431,4.0674906,5.2644167,6.910619,9.153569,8.954653,7.805741,11.749766,10.076128,8.707723,9.530824,11.646879,11.369082,10.573419,10.926665,11.681175,12.034423,11.108434,7.7748747,5.7719955,4.897451,4.866585,5.295283,5.0140567,6.108095,7.301592,7.970361,8.117833,6.6053853,4.386442,4.863155,7.2707253,6.697984,3.7794054,2.393852,1.6187652,1.1797781,1.4507155,0.607037,0.28808534,0.23664154,0.31895164,0.48700142,0.61046654,0.805953,0.78194594,0.65162164,0.9294182,0.6859175,0.4972902,0.3806842,0.32238123,0.274367,0.4081209,0.41498008,0.45270553,0.53501564,0.53501564,0.4355576,0.6859175,0.8196714,0.83681935,1.1900668,1.2758065,1.3238207,1.488441,1.6324836,1.3272504,1.5364552,1.5673214,1.5021594,1.3238207,0.94656616,0.8471081,0.88826317,0.77851635,0.5693115,0.64133286,0.9842916,1.3169615,1.4678634,1.5673214,2.0440342,2.2635276,2.2566686,1.9994495,1.587899,1.2209331,1.4267083,2.1846473,2.9185789,3.216953,2.8396983,2.3492675,2.6750782,3.2821152,3.7279615,3.6936657,4.7534084,4.4721823,4.029765,4.0091877,4.3624353,4.914599,3.9886103,3.457024,3.5461934,2.8396983,2.2395205,1.6976458,2.1297739,2.8122618,1.371835,2.5584722,4.0537724,3.99204,2.3389788,0.8848336,0.432128,0.65848076,0.97057325,0.9774324,0.48700142,0.47671264,2.277246,3.391862,3.4913201,4.3933015,2.0508933,0.980862,2.1880767,4.046913,2.287535,2.6922262,3.0317552,2.5893385,1.6153357,1.2963841,2.627064,2.7402403,2.2566686,1.6496316,1.2346514,1.7593783,3.1655092,3.7862647,3.4535947,3.4810312,7.226141,13.29994,17.46003,17.487467,13.152468,4.715683,3.1483612,2.8808534,2.2086544,3.2821152,2.4384367,2.9974594,4.3452873,4.9214582,2.2120838,2.7985435,2.9254382,2.2909644,3.806842,13.594885,10.799771,7.2364297,4.976331,3.6353626,0.34981793,0.20577525,0.15776102,0.32238123,0.5761707,0.5658819,0.5761707,0.96371406,1.7833855,2.6750782,2.884283,3.9714622,4.588788,5.0174866,5.188966,4.698535,4.32128,4.619654,4.650521,4.1463714,3.525616,3.9028704,3.8137012,3.3266997,2.5173173,1.4815818,2.0303159,1.9274281,1.4335675,0.8265306,0.4115505,0.6310441,0.9877212,0.91569984,0.5212973,0.59674823,0.9602845,1.8485477,2.9185789,3.9886103,5.051782,5.2815647,4.417309,4.256118,5.394741,7.2021337,4.187526,3.4433057,4.033195,5.0826488,5.751418,5.7274113,5.830299,6.64997,8.107545,9.47595,7.840037,4.6127954,2.0920484,1.2277923,1.6187652,1.6667795,1.6599203,1.8965619,2.1332035,1.5707511,1.3272504,1.1283343,1.4232788,2.2600982,3.309552,2.860276,1.8039631,0.7613684,0.35324752,1.2209331,1.611906,1.6187652,1.4095604,1.3409687,1.937717,2.9631636,3.998899,4.633373,4.9180284,5.3570156,5.4667625,4.7774153,3.9851806,3.3438478,2.6853669,2.6853669,2.428148,2.5378947,2.9494452,2.8980014,1.704505,0.9911508,0.9568549,1.1077567,0.29151493,0.6310441,1.862266,3.1792276,4.32128,5.552502,4.7979927,3.0523329,2.417859,3.1723683,3.782835,4.540774,4.1429415,3.3987212,2.6716487,1.8759843,1.5227368,1.1420527,0.90198153,0.90884066,1.1900668,0.72707254,0.5658819,0.7339317,1.3924125,2.8088322,2.9288676,3.1620796,3.093488,2.7299516,2.486451,2.4624438,2.5653315,3.2855449,4.8734436,7.3393173,7.1678376,7.5382333,7.7577267,7.4010496,6.3001523,6.0223556,5.521636,4.9523244,4.6745276,5.2506986,7.6651278,7.473071,7.143831,7.407909,7.2467184,6.392751,6.601956,6.550512,5.8645945,5.096367,3.059192,1.9720128,1.8485477,2.386993,2.959734,3.8891523,3.2409601,2.4590142,2.819121,5.4324665,4.9694724,4.1017866,3.4844608,3.1312134,2.411,1.8245405,2.0165975,2.3458378,2.5961976,2.976882,2.901431,2.6922262,2.6990852,2.9665933,3.234101,3.1483612,2.9254382,3.0729103,3.5016088,3.525616,3.6353626,4.091498,4.197815,3.9200184,3.9200184,3.5187566,3.3644254,2.952875,2.2052248,1.4507155,1.1317638,1.1249046,1.2312219,1.3066728,1.2826657,1.0494537,1.4129901,1.7113642,1.6290541,1.1900668,1.5193073,1.4918705,1.4369972,1.5158776,1.7250825,2.6887965,3.175798,3.57363,3.9543142,4.0880685,3.9440255,3.8891523,3.649081,3.3781435,3.6456516,0.0,0.030866288,0.020577524,0.01371835,0.017147938,0.01371835,0.01371835,0.024007112,0.030866288,0.037725464,0.030866288,0.030866288,0.09602845,0.16119061,0.22292319,0.31895164,0.6241849,1.0323058,1.2483698,1.2998136,1.5536032,1.6873571,1.8348293,1.9685832,2.153781,2.534465,3.0420442,3.7142432,4.2835546,4.6127954,4.6916757,4.8254294,4.846007,4.9660425,5.178677,5.2301207,5.1066556,4.8940215,4.866585,5.0243454,5.0929375,4.8185706,4.7431192,4.4756117,3.974892,3.532475,4.0949273,5.130663,5.796003,5.6965446,4.8837323,4.4241676,4.7431192,4.73969,4.32128,4.413879,4.1292233,4.3692946,4.722542,5.113515,5.809721,5.970912,6.2487082,6.186976,5.857735,5.857735,6.48535,7.425057,7.9772205,8.100685,8.433355,8.971801,9.740028,9.716022,8.97523,8.697433,9.31133,10.0041065,10.72775,11.283342,11.31078,11.074138,10.923236,10.5597,10.065839,9.870353,9.966381,10.607714,12.072148,13.725209,14.013294,13.670336,12.065289,10.329918,9.585697,10.912948,11.80121,11.794352,11.159878,10.532263,10.899229,11.571428,12.240198,13.745787,15.844694,17.21996,17.021042,16.016174,15.29253,15.542891,17.03819,16.29054,15.4914465,15.333686,15.6697855,15.529172,14.531162,14.997586,16.20137,17.665806,19.140528,20.217419,21.146837,21.589252,21.335464,20.313446,17.892159,15.896138,14.771234,14.586036,15.001016,15.316538,15.810398,16.204802,16.304258,16.023033,15.549749,15.446862,15.073037,14.352823,13.783512,13.190193,13.581166,14.205351,14.771234,15.46744,15.621771,15.580616,15.3302555,15.110763,15.415996,16.54776,17.141079,17.597214,17.943602,17.857862,18.410025,18.492336,18.54378,18.506054,17.820137,16.914726,16.486027,16.11906,15.930434,16.53404,17.144508,17.309128,17.549198,17.87501,17.79613,17.600643,17.38115,17.024471,16.568336,16.194511,16.269962,16.225378,15.923574,15.453721,15.148488,15.422854,15.433144,15.745236,16.317978,16.499744,15.844694,15.073037,14.387119,14.157337,14.918706,16.12249,16.636929,16.695232,16.914726,18.28313,19.085653,19.099373,19.54179,20.968498,23.27661,25.413242,25.52985,24.905664,24.315775,24.013971,23.2869,23.34863,23.623,23.69159,23.27661,21.966507,20.817596,19.634388,18.488907,17.730967,17.768692,18.595222,19.339443,19.239986,17.63494,16.153357,15.5085945,15.865272,16.715809,16.897577,17.532051,18.674105,19.288,19.288,19.54179,18.732407,19.11995,20.27915,21.1194,19.884748,18.327715,17.593784,17.171944,16.877,16.825556,16.47231,16.03675,15.289101,14.428274,14.040731,13.522863,14.054449,14.335675,14.150477,14.349394,14.068168,13.231348,13.035862,13.320518,12.583157,12.816368,14.037301,14.339106,13.272504,11.852654,11.698323,11.485688,11.38623,11.506266,11.897239,11.742908,11.506266,11.756626,12.360233,12.504276,11.30049,10.97468,10.593996,10.545981,12.535142,13.437123,14.712931,15.549749,15.251375,13.224489,11.30049,8.268735,7.2535777,8.371623,8.7283,8.405919,8.443645,11.314209,14.712931,11.55771,8.766026,7.1849856,8.155559,10.017825,8.107545,5.90232,4.863155,4.3178506,3.806842,3.0626216,2.1812177,3.0660512,3.0660512,2.201795,3.199805,3.3781435,3.1963756,3.4433057,4.5647807,6.680836,8.1041155,7.7577267,7.8091707,9.074688,11.015835,8.220721,8.759167,10.864933,12.699762,12.367092,12.960411,12.240198,11.72233,10.998687,7.7268605,6.1046658,6.121814,6.6568294,7.1952744,7.846896,8.375052,8.090397,7.267296,6.701414,7.6788464,7.5416627,5.0655007,4.166949,4.90431,3.5016088,1.862266,1.488441,1.4335675,1.3752645,1.6324836,0.6241849,0.2777966,0.2194936,0.26750782,0.42869842,0.45270553,0.6962063,0.83338976,0.8265306,0.9431366,0.77851635,0.5555932,0.42183927,0.4046913,0.432128,0.37382504,0.38754338,0.42869842,0.48700142,0.59674823,0.58645946,0.59331864,0.64476246,0.7373613,0.83681935,1.1077567,1.1866373,1.2792361,1.4232788,1.4987297,1.3924125,1.3546871,1.3924125,1.3821237,1.08032,0.97400284,0.96714365,0.84024894,0.66876954,0.7990939,0.85739684,1.1729189,1.371835,1.4335675,1.6530612,1.9514352,2.2463799,2.2738166,2.0303159,1.7833855,1.7456601,2.1400626,2.8534167,3.3438478,2.644212,2.867135,2.6990852,2.784825,3.3301294,4.0949273,4.5510626,4.372724,4.201245,4.3041325,4.557922,4.3761535,3.450165,3.7794054,4.633373,2.568761,2.3904223,3.1895163,3.4810312,2.7162333,1.2758065,2.07833,1.8382589,1.2895249,0.8779744,0.7613684,2.4590142,2.9871707,2.8980014,2.5481834,2.0989075,2.4967396,2.0131679,3.2581081,5.1100855,2.7230926,1.3341095,1.6324836,5.1992545,8.7283,4.0229063,3.8891523,2.4967396,1.5330256,1.762808,3.018037,2.8637056,2.644212,3.1209247,5.2575574,10.196163,6.5127864,8.042382,9.654288,9.263316,7.8126,9.674867,12.47341,13.749216,12.881531,11.077567,5.2609873,2.8739944,5.079219,9.31133,9.273604,7.06495,7.4113383,7.5519514,6.252138,3.82399,4.7499785,3.069481,2.1194851,3.350707,6.2967224,4.1635194,6.800872,7.7885933,5.103226,1.0940384,0.7442205,0.5521636,0.6036074,0.83681935,1.039165,0.9259886,1.4644338,2.5310357,3.4535947,3.018037,3.9303071,4.605936,4.9420357,5.209543,6.0806584,4.6265135,4.3281393,4.2938433,3.9200184,2.877424,3.000889,3.1655092,3.3198407,3.0557625,1.5913286,1.4644338,1.3203912,1.2655178,1.1866373,0.7407909,1.0014396,1.08032,0.96371406,0.7442205,0.6310441,0.8128122,1.1763484,1.9102802,2.760818,3.0626216,4.249259,4.273266,4.2766957,4.791134,5.7479887,4.540774,4.650521,5.144381,5.878313,7.486789,6.464772,6.2041235,7.4353456,8.769455,6.680836,5.4941993,3.8720043,2.2978237,1.4987297,2.435007,1.5947582,1.4198492,1.5981878,1.8588364,1.9514352,1.8142518,1.5981878,1.4850113,1.5810398,1.9068506,2.0817597,1.8691251,1.2792361,0.77508676,1.2826657,1.5844694,1.5981878,1.5227368,1.5261664,1.7559488,2.585909,3.5564823,4.262977,4.6779575,5.137522,5.871454,5.1512403,4.2526884,3.5804894,2.6476414,2.6476414,2.6579304,2.6716487,2.8259802,3.3644254,2.0989075,1.5330256,1.529596,1.937717,2.585909,1.3238207,3.5839188,5.120374,4.756838,4.3590055,4.256118,3.5016088,3.4776018,4.266407,4.650521,4.8322887,4.3933015,3.923448,3.5118976,2.767677,2.177788,1.6427724,1.2449403,1.0768905,1.2380811,0.7956643,0.5796003,0.70649505,1.2483698,2.2326615,2.767677,3.1140654,3.1517909,2.9494452,2.8054025,2.1743584,2.5721905,3.5050385,4.8117113,6.691125,6.893471,7.442205,7.6033955,7.267296,6.9620624,5.977771,5.645101,5.4084597,5.195825,5.4084597,6.632822,6.1801167,5.6828265,5.8405876,6.392751,7.1198235,7.298162,6.6636887,5.5387836,4.8288593,3.6079261,2.719663,2.5207467,2.6922262,2.2395205,2.5927682,3.1277838,3.4433057,3.707384,4.650521,3.5050385,2.860276,2.4247184,2.0646117,1.8142518,1.3924125,1.5158776,1.9480057,2.4247184,2.6579304,2.6236343,2.6133456,2.5413244,2.5207467,2.8568463,2.8019729,2.2978237,2.0646117,2.2360911,2.3767042,2.4007113,3.100347,3.450165,3.2375305,3.0420442,3.1586502,3.8479972,3.9371665,3.1449318,2.085189,1.4918705,1.3101025,1.196926,1.1214751,1.3443983,1.2003556,1.3786942,1.605047,1.6324836,1.2517995,1.3958421,1.6359133,1.8245405,2.0440342,2.603057,3.2066643,3.2615378,3.3061223,3.5461934,3.858286,3.6525106,3.8102717,3.6319332,3.1860867,3.316411,0.0,0.030866288,0.034295876,0.11317638,0.1920569,0.024007112,0.017147938,0.020577524,0.020577524,0.0274367,0.048014224,0.11317638,0.22978236,0.36696586,0.53844523,0.7956643,1.1180456,1.3958421,1.471293,1.4095604,1.5021594,1.6530612,1.7559488,1.9651536,2.2806756,2.534465,3.018037,3.4913201,4.0229063,4.420738,4.2183924,4.201245,4.413879,4.633373,4.7191124,4.616225,4.636802,4.633373,4.7945633,4.9831905,4.7259717,4.523626,4.431027,4.256118,3.957744,3.642222,3.9028704,4.7019644,5.099797,4.791134,4.105216,3.7485392,3.9680326,4.2081037,4.32471,4.6127954,4.0057583,4.1772375,4.695105,5.2438393,5.597087,5.830299,6.3138704,6.4133286,6.0223556,5.56965,5.7582774,6.5230756,7.2638664,7.922347,8.985519,9.499957,10.343636,10.628291,10.326488,10.268185,10.38479,10.683165,11.351934,11.986408,11.561139,11.345076,11.369082,11.080997,10.436234,9.914937,9.6988735,10.690024,12.157887,13.450842,13.996146,13.193623,11.417097,10.017825,9.89436,11.499407,11.96926,11.8115,11.276484,10.659158,10.30934,11.1393,11.941824,13.660047,15.577187,15.306249,15.385129,14.514014,13.989287,14.565458,16.482597,16.835844,16.739817,16.37971,15.885849,15.350834,14.613472,14.596324,15.350834,16.71238,18.28313,19.737276,21.232576,22.326614,22.676432,22.04539,19.336014,17.017612,15.385129,14.603184,14.7095,15.035312,15.29596,15.539461,15.638919,15.306249,14.911846,14.802099,14.606613,14.349394,14.452282,13.783512,13.975569,14.407697,14.791811,15.169065,14.901558,14.534592,14.2533655,14.191633,14.445422,15.854982,16.403717,16.434584,16.410576,16.88386,17.532051,17.700102,17.782412,17.895588,17.895588,17.288551,16.88386,16.345413,15.896138,16.29397,16.489456,16.698662,17.024471,17.357141,17.370861,17.761833,18.156237,18.20768,17.778982,16.938732,16.448301,16.355703,16.143068,15.752095,15.587475,15.265094,14.836395,14.894698,15.484588,16.101913,15.275383,14.928994,14.994157,15.2033615,15.12448,16.143068,16.410576,16.400288,16.438013,16.719238,18.101362,18.595222,18.629519,18.746124,19.603521,22.919933,24.308916,24.240324,23.52354,23.2869,22.12427,21.959648,22.511812,23.060547,22.453508,20.968498,19.637817,18.416885,17.525192,17.418875,16.94902,17.477179,18.231688,18.54378,17.86815,17.058767,16.47231,16.321407,16.616352,17.158226,17.278261,17.748116,18.156237,18.38259,18.629519,17.892159,18.149376,18.814716,19.250275,18.752985,17.466888,16.973028,16.684942,16.516893,16.87014,16.21509,15.494876,14.832966,14.225929,13.577737,13.21763,14.037301,14.30481,13.965281,14.658057,14.016724,13.227919,13.077017,13.21763,12.175035,12.987847,13.605173,13.773223,13.471419,12.891819,11.64345,11.447963,11.567999,11.495977,10.933525,11.749766,12.46312,13.207341,13.80409,13.776653,13.505715,13.176475,12.439114,11.97269,13.498857,13.917266,15.145059,14.493437,12.13731,11.0981455,12.6929035,10.930096,9.445084,9.115844,8.038953,5.6005163,4.8117113,8.635701,14.112752,12.363663,11.835506,10.096705,8.858624,8.165848,6.385892,5.9983487,4.5201964,3.2375305,2.6545007,2.4658735,1.4472859,2.3972816,2.767677,2.3321195,3.1655092,3.875434,3.690236,4.3281393,6.0395036,7.5931067,7.157549,7.949784,9.328478,10.556271,10.789482,9.373062,10.405369,12.140739,13.077017,11.952112,11.622872,10.319629,8.460793,6.8969,6.927767,7.431916,7.8846216,8.31332,8.536243,8.189855,9.129561,8.453933,6.948344,5.9126086,7.191845,6.615674,5.4153185,4.1463714,3.3781435,3.6696587,1.8999915,1.5398848,1.4164196,1.2277923,1.5398848,0.58645946,0.24007112,0.15433143,0.14747226,0.2194936,0.2777966,0.48357183,0.7613684,1.0151579,1.1008976,0.881404,0.6790583,0.5453044,0.48014224,0.42869842,0.36696586,0.38754338,0.38754338,0.42526886,0.72021335,0.6962063,0.6001778,0.61389613,0.6893471,0.5658819,0.89512235,1.1592005,1.1729189,1.0940384,1.4129901,1.3032433,1.1660597,1.1832076,1.313532,1.2895249,1.1111864,1.0940384,0.9328478,0.6962063,0.8128122,0.97400284,1.0528834,1.1523414,1.3306799,1.5844694,1.6290541,2.0817597,2.2635276,2.1126258,2.170929,1.9925903,2.2052248,2.8877127,3.4776018,2.767677,3.1346428,2.8637056,2.74367,3.100347,3.8034124,4.0194764,4.081209,4.2252517,4.4756117,4.6265135,4.588788,4.040054,3.8548563,3.8514268,2.784825,2.4727325,2.836269,2.9254382,2.4795918,1.9548649,3.2066643,2.5413244,2.5310357,3.6559403,4.2835546,5.7994323,6.0223556,5.4324665,4.695105,4.6436615,2.551613,1.6599203,3.5599117,5.785714,1.8382589,1.1592005,2.620205,7.997798,11.993267,2.2498093,3.4021509,2.860276,2.2360911,2.1915064,2.4418662,2.7299516,3.2649672,3.649081,4.547633,7.6925645,6.831738,8.80718,9.849775,9.112414,8.683716,11.094715,14.140189,13.845244,10.316199,7.740579,4.5030484,4.8151407,8.779744,13.015285,10.662587,5.1821065,6.0703697,6.725421,4.839148,2.3972816,3.0489032,2.2909644,2.2978237,3.957744,6.869464,4.8734436,6.992929,9.366203,8.958082,3.5599117,1.7525192,0.91912943,0.90541106,1.2963841,1.4061309,1.5981878,1.845118,2.651071,3.6456516,3.6113555,3.2683969,3.858286,4.48933,5.0346346,6.1046658,5.305572,4.773986,4.341858,3.7622573,2.726522,2.8808534,3.1037767,3.1723683,2.8637056,1.9480057,1.8656956,1.670209,1.5810398,1.5090185,1.0357354,0.9602845,0.823101,0.7407909,0.70306545,0.59674823,0.85396725,1.1214751,1.7113642,2.4212887,2.5173173,3.6593697,4.2595477,4.633373,5.003768,5.4770513,4.6848164,5.4667625,6.3001523,6.8763227,8.083538,7.233,6.324159,6.914048,8.008087,6.0737996,6.23499,5.171818,3.5564823,2.3629858,2.8499873,1.9582944,1.920569,2.0577524,2.1023371,2.218943,2.1812177,2.1194851,1.8073926,1.5364552,2.0886188,2.6236343,2.49331,2.136633,1.8279701,1.6633499,1.8039631,1.845118,1.8313997,1.7422304,1.4815818,2.3561265,3.0351849,3.5839188,4.1189346,4.7774153,5.305572,5.0757895,4.4584637,3.673088,2.7951138,2.5447538,2.6236343,2.6545007,2.726522,3.3952916,2.5550427,1.9685832,1.6427724,1.6873571,2.335549,1.4129901,2.2909644,3.9783216,4.8254294,2.503599,2.6819375,2.9494452,3.5942078,4.389872,4.602506,5.1580997,4.976331,4.413879,3.7451096,3.1723683,2.5996273,2.1160555,1.6427724,1.2620882,1.214074,0.9362774,0.6927767,0.6790583,1.0425946,1.862266,2.4898806,2.9631636,3.1449318,3.0420442,2.8019729,2.218943,2.750529,3.6044965,4.6676683,6.5127864,6.8557453,7.1129646,7.4181976,7.795452,8.169277,7.332458,6.3207297,5.796003,5.7994323,5.768566,6.636252,6.1801167,5.813151,6.0669403,6.608815,7.14726,7.4284863,6.7185616,5.2781353,4.386442,3.5633414,2.8328393,2.5001693,2.4830213,2.2806756,2.1126258,2.3904223,2.750529,2.9460156,2.836269,2.2120838,1.9480057,1.845118,1.7353712,1.5090185,1.0631721,1.097468,1.4232788,1.8142518,2.0097382,2.095478,2.2463799,2.1057668,1.7696671,1.762808,2.0234566,1.8039631,1.6153357,1.6770682,1.9068506,2.0817597,2.651071,2.9906003,2.9048605,2.6304936,2.8980014,3.5461934,3.8445675,3.4947495,2.6373527,1.920569,1.5536032,1.2620882,1.0323058,1.138623,1.2449403,1.2209331,1.2620882,1.3272504,1.1283343,1.3821237,1.7936742,2.0920484,2.3664153,3.0797696,3.525616,3.4227283,3.3850029,3.5976372,3.789694,3.3952916,3.532475,3.532475,3.2718265,3.1723683,0.09259886,0.061732575,0.044584636,0.12003556,0.19548649,0.017147938,0.017147938,0.020577524,0.0274367,0.061732575,0.14747226,0.31895164,0.4938606,0.6859175,0.97057325,1.4815818,1.3684053,1.5158776,1.5810398,1.5021594,1.4815818,1.6290541,1.7490896,2.0440342,2.469303,2.726522,3.0900583,3.234101,3.4947495,3.789694,3.5770597,3.6044965,3.9714622,4.2252517,4.2286816,4.170378,4.3041325,4.437886,4.7671266,5.099797,4.8494368,4.557922,4.4516044,4.355576,4.190956,3.9440255,3.8788633,4.3761535,4.5647807,4.149801,3.4227283,3.1346428,3.3266997,3.707384,4.0846386,4.3795834,3.8308492,4.0229063,4.616225,5.2026844,5.2747054,5.720552,6.3790326,6.691125,6.4716315,5.9228973,5.9297566,6.3173003,6.8557453,7.5245147,8.539673,9.499957,10.618003,11.293632,11.523414,11.910957,11.838936,11.941824,12.370522,12.696333,11.89038,11.513125,11.55428,11.31078,10.683165,10.179015,9.97324,10.690024,11.712041,12.679185,13.488567,12.346515,11.070708,10.240748,10.299051,11.537132,11.993267,12.113303,11.948683,11.595435,11.218181,11.982979,12.322508,13.437123,14.733508,13.824667,13.615462,13.430264,13.618892,14.335675,15.542891,16.39,16.62321,16.19794,15.446862,15.076467,15.155347,15.350834,15.6526375,16.04018,16.513464,18.080786,20.124819,21.815605,22.683292,22.60098,20.395756,18.02934,16.105343,14.863832,14.184773,14.448852,14.421415,14.5243025,14.79867,14.904987,14.908417,14.685493,14.565458,14.743796,15.251375,14.589465,14.726648,15.2033615,15.566897,15.37827,15.0456,14.459141,14.05102,14.05102,14.476289,15.700651,16.400288,16.139639,15.436573,15.789821,16.273392,16.54433,16.602633,16.616352,16.918156,16.859852,16.808409,16.63007,16.46545,16.726099,16.6335,16.678083,16.852993,17.093063,17.254255,17.394867,17.96418,18.269413,17.929884,16.859852,15.827546,15.635489,15.594335,15.46058,15.415996,14.815818,14.664916,14.654627,14.7197895,15.0456,14.356253,14.421415,15.21365,16.163645,16.173935,16.890718,17.04162,17.027903,16.897577,16.352274,17.062197,17.857862,17.86815,17.21653,17.024471,19.78186,21.908205,22.655855,22.213438,21.726437,20.406046,20.138538,20.749004,21.52066,21.218857,19.819586,18.739265,17.778982,17.110212,17.247395,16.846134,16.897577,17.333136,17.833855,17.854433,17.38115,17.099922,16.811838,16.63007,16.986746,16.997036,16.746675,16.70895,16.897577,16.856422,16.63007,17.017612,17.29541,17.288551,17.367432,16.753534,16.671225,16.602633,16.45173,16.523752,15.621771,14.79524,14.260224,13.992717,13.728639,13.594885,13.992717,13.951562,13.629181,14.308239,13.749216,13.419975,13.138749,12.699762,11.869802,12.507706,12.596875,12.950122,13.437123,12.9809885,11.530273,12.260776,13.574307,13.776653,11.091286,12.72034,13.186764,13.708061,14.38369,14.198492,13.865822,13.756075,13.540011,13.516005,14.589465,14.640909,14.160767,12.545431,11.351934,14.273943,15.367981,13.025573,10.659158,9.167287,6.927767,5.610805,3.957744,5.967482,9.760606,7.5725293,9.945804,9.729739,10.501397,11.756626,8.916927,5.113515,4.389872,4.4275975,4.187526,3.9131594,2.1126258,3.2683969,3.6799474,3.1586502,5.0312047,5.2164025,5.120374,5.4839106,6.3035817,6.8557453,6.5950966,8.573969,10.707172,11.619442,10.618003,10.88894,11.873232,12.991278,13.13189,10.669447,8.745448,7.8091707,6.186976,4.756838,6.9209075,9.465661,9.441654,8.940934,8.639131,7.8194594,7.716572,6.931196,5.7239814,4.866585,5.6485305,5.4324665,5.5422134,4.931747,3.9474552,4.2938433,2.5653315,1.903421,1.5261664,1.1866373,1.155771,0.4698535,0.19548649,0.10288762,0.072021335,0.08573969,0.16804978,0.30866286,0.6001778,0.980862,1.2483698,0.9842916,0.8505377,0.7305021,0.5761707,0.42183927,0.40126175,0.40126175,0.3566771,0.36353627,0.6893471,0.70306545,0.58302987,0.61389613,0.7407909,0.5521636,0.7373613,1.0666018,1.0768905,0.89169276,1.2003556,1.2175035,1.1180456,1.0837497,1.1729189,1.3306799,1.1832076,1.1832076,1.0425946,0.77851635,0.7133542,1.0425946,1.0048691,1.0425946,1.2860953,1.5638919,1.5913286,2.0097382,2.2326615,2.2120838,2.452155,2.16064,2.294394,2.836269,3.333559,2.9151495,3.3232703,3.1380725,3.1037767,3.4192986,3.7279615,3.8720043,4.0537724,4.273266,4.5099077,4.705394,4.928317,4.046913,3.6559403,3.8479972,3.2066643,2.9563043,2.4898806,2.1332035,2.1023371,2.510458,3.1860867,3.175798,3.74168,4.7979927,4.8940215,6.591667,7.3873315,6.776865,5.394741,4.979761,2.4967396,2.2292318,4.07435,5.5833683,1.9720128,2.3081124,4.256118,8.025234,9.729739,1.4129901,4.629943,5.65539,5.4804807,4.629943,3.1552205,4.033195,4.290414,3.8617156,3.3438478,3.981751,4.7362604,6.0875177,6.5642304,6.3824625,7.459353,9.73317,12.55915,11.773774,7.840037,5.8543057,5.3707337,6.5813785,10.069269,13.841815,13.317088,5.7994323,4.822,4.911169,3.508468,0.9431366,1.3581166,1.3101025,1.8039631,3.3850029,6.166398,4.396731,6.2898636,8.48137,8.460793,4.5922174,2.1846473,1.08032,1.0940384,1.6496316,1.7799559,2.3321195,2.469303,2.9254382,3.6970954,4.0366244,3.0214665,3.391862,4.0606318,4.6127954,5.284994,5.4976287,5.1683884,4.6265135,3.9783216,3.0900583,3.1415021,3.199805,3.1723683,3.0043187,2.6990852,2.469303,2.301253,2.1160555,1.8519772,1.4438564,1.039165,0.7373613,0.6173257,0.6276145,0.59674823,1.0254467,1.2860953,1.786815,2.4144297,2.5310357,3.0317552,3.8377085,4.705394,5.429037,5.826869,5.3261495,6.1149545,6.7048435,6.824879,7.407909,6.608815,5.7239814,5.953764,6.8797526,6.4887795,7.0375133,5.8200097,4.190956,3.0420442,2.7779658,2.311542,2.4761622,2.6407824,2.5721905,2.4212887,2.1846473,2.335549,2.3218307,2.1091962,2.2086544,2.6956558,2.5893385,2.6545007,2.8259802,2.2258022,1.9720128,1.9514352,2.0097382,1.8931323,1.2620882,2.170929,2.6407824,2.9700227,3.3850029,4.040054,4.173808,4.4721823,4.2766957,3.5393343,2.8122618,2.3218307,2.411,2.5447538,2.6613598,3.1723683,3.0866287,2.5447538,1.8725548,1.4438564,1.7010754,1.430138,1.1763484,2.8877127,4.791134,1.4164196,3.7279615,3.333559,3.1517909,3.9063,4.139512,5.1340923,5.3844523,4.8151407,3.806842,3.1860867,2.6853669,2.2806756,1.8382589,1.4095604,1.2380811,1.0151579,0.7990939,0.7579388,1.0323058,1.7456601,2.2909644,2.644212,2.8328393,2.843128,2.6476414,2.386993,2.9048605,3.4913201,4.2835546,6.262427,6.893471,7.2535777,7.689135,8.213862,8.48137,8.008087,6.835168,6.0154963,5.895461,6.0737996,6.468202,5.9297566,5.689686,6.0806584,6.5196457,6.8591747,7.0478024,6.4544835,5.2335505,4.307562,3.4776018,2.9185789,2.5001693,2.253239,2.352697,2.3149714,2.2566686,2.2978237,2.2841053,1.821111,1.5947582,1.587899,1.6804979,1.6907866,1.3684053,0.9534253,0.89169276,1.039165,1.2483698,1.3889829,1.4747226,1.6427724,1.5913286,1.3306799,1.1763484,1.4164196,1.5055889,1.5398848,1.6256244,1.8588364,2.1160555,2.469303,2.74367,2.7745364,2.3732746,2.74367,3.1586502,3.4844608,3.4878905,2.8499873,2.201795,1.7250825,1.3649758,1.0940384,0.90541106,1.0357354,0.980862,0.91569984,0.94999576,1.1420527,1.4232788,1.8725548,2.2463799,2.609916,3.3472774,3.3781435,3.4535947,3.6559403,3.8514268,3.6627994,3.3198407,3.4947495,3.57363,3.3644254,3.0969174,0.18176813,0.09602845,0.044584636,0.024007112,0.020577524,0.0034295875,0.017147938,0.041155048,0.09602845,0.19548649,0.34638834,0.6001778,0.83681935,1.0631721,1.3958421,2.0508933,1.4987297,1.6153357,1.7490896,1.6736387,1.587899,1.6942163,1.8828435,2.201795,2.603057,2.9322972,3.1243541,3.0660512,3.0111778,3.0283258,3.0043187,3.2409601,3.6182148,3.7931237,3.7862647,3.9646032,4.180667,4.2046742,4.557922,5.120374,5.144381,4.712253,4.5442033,4.4447455,4.2389703,3.758828,3.532475,3.758828,3.865145,3.590778,2.959734,2.7745364,2.8499873,3.0420442,3.2512488,3.433017,3.4055803,3.7725463,4.338428,4.8014226,4.773986,5.3158607,6.461343,7.3118806,7.4524937,6.9380555,6.9037595,6.989499,7.291303,7.6685576,7.7714453,9.177576,10.645439,11.574858,12.010415,12.655178,12.771784,12.80608,12.97413,13.056439,12.38424,11.667457,11.393089,11.173596,10.882081,10.676306,10.686595,10.549411,10.998687,12.085866,13.169616,12.020704,11.485688,11.026124,10.679735,11.046701,12.171606,13.169616,13.509145,13.38568,13.71492,14.21564,13.834956,13.684054,13.999576,14.140189,13.258785,13.653188,14.565458,15.271953,15.100473,15.309678,15.100473,14.7095,14.452282,14.7095,15.518884,16.441442,16.907866,16.660936,15.745236,16.523752,18.28656,20.018501,21.236006,21.980227,21.054237,19.095943,17.20281,15.734947,14.318527,14.102464,13.858963,13.941273,14.373401,14.832966,15.326826,15.100473,14.970149,15.21022,15.594335,15.114192,15.309678,15.841265,16.180794,15.6252,15.662926,15.343974,14.932424,14.7369375,15.12448,15.7966795,16.513464,16.335125,15.395418,14.928994,15.0456,15.556609,15.7966795,15.676644,15.707511,15.892709,16.37285,16.87014,17.230247,17.436022,17.388008,17.343424,17.29198,17.29198,17.46003,16.780972,17.03819,17.357141,17.19938,16.352274,15.0250225,14.647768,14.685493,14.822677,14.932424,14.342535,14.712931,14.757515,14.311668,14.308239,13.9138365,13.954991,14.922135,16.54433,17.772121,18.471758,18.440891,18.156237,17.833855,17.405157,16.859852,17.264544,17.322845,16.777542,16.441442,17.422304,19.219408,20.423193,20.508932,19.826445,18.938183,18.509483,18.62609,19.089085,19.411465,18.667244,18.104792,17.61779,17.271402,17.29884,17.549198,17.315987,17.243965,17.350283,17.027903,16.503176,16.750105,16.849564,16.561478,16.321407,16.499744,16.071047,15.758954,15.659496,15.247946,15.594335,16.249386,16.53747,16.434584,16.564907,16.516893,16.540901,16.479168,16.20137,15.608052,14.675205,14.123041,13.821238,13.749216,14.016724,14.095605,13.828096,13.529722,13.416546,13.612033,13.450842,13.697772,13.22106,12.113303,11.691463,11.732618,11.996697,12.655178,13.13189,12.089295,11.856084,13.900118,16.047039,16.424294,13.481709,13.708061,12.569438,12.610593,13.776653,13.395968,12.71691,13.395968,14.119612,14.579176,15.470869,15.529172,12.922686,12.089295,15.223939,22.275171,17.305698,12.80265,10.213311,9.0644,6.992929,6.3138704,4.5853586,6.193835,8.464222,1.670209,4.619654,7.6445503,13.584596,18.763273,13.008426,3.7176728,5.0312047,6.7974424,5.953764,6.5539417,4.1360826,5.2335505,5.2747054,4.5922174,8.4264965,7.5210853,7.1369715,6.4064693,5.4941993,5.593657,7.425057,9.194724,10.861504,11.732618,10.443094,11.732618,12.672326,12.9638405,12.0138445,8.958082,6.2212715,6.7974424,6.615674,5.5559316,7.473071,10.827208,10.501397,8.875772,7.5759587,7.4696417,5.7377,5.1169443,4.307562,3.2786856,3.2512488,4.4721823,5.086078,5.576509,5.638242,4.173808,3.1552205,2.287535,1.6942163,1.2860953,0.7476501,0.36696586,0.18176813,0.09602845,0.058302987,0.06859175,0.12003556,0.216064,0.4115505,0.7613684,1.3032433,1.0700313,0.99801,0.88826317,0.6927767,0.5178677,0.45270553,0.4081209,0.36010668,0.3566771,0.50757897,0.6173257,0.5453044,0.6344737,0.8505377,0.7682276,0.7579388,0.922559,0.96371406,0.8848336,0.9877212,1.0631721,1.0940384,1.0563129,1.0185875,1.1454822,1.1454822,1.1900668,1.138623,0.94656616,0.66191036,0.9911508,1.0700313,1.1283343,1.2723769,1.4987297,1.8039631,2.0680413,2.2292318,2.3218307,2.469303,2.194936,2.3218307,2.6236343,2.867135,2.8328393,3.275256,3.216953,3.40901,3.8720043,3.8788633,4.0674906,4.2423997,4.3692946,4.4859004,4.722542,4.7671266,3.2512488,3.3987212,4.8288593,3.549623,3.5016088,2.750529,1.9994495,1.8108221,2.6167753,1.9582944,2.7813954,3.4398763,3.275256,2.609916,4.4104495,6.931196,6.8454566,4.3658648,3.2615378,3.0454736,3.7862647,4.7328305,4.852866,2.8225505,3.7553983,5.8371577,6.358455,4.695105,2.2909644,8.008087,9.9801,9.328478,7.1884155,4.698535,5.6142344,4.9488945,3.9646032,3.5393343,4.1429415,3.2443898,2.976882,3.0043187,3.4467354,4.8597255,6.23499,7.81603,7.671987,6.3207297,6.7459984,9.201583,11.355364,13.275933,15.172495,17.412016,10.367643,5.7239814,3.6765177,2.9700227,0.881404,0.9911508,1.3992717,1.5844694,1.7765263,2.959734,1.8554068,5.0449233,6.831738,5.48734,3.2272418,1.6907866,0.980862,1.1111864,1.7216529,2.0817597,2.7402403,3.0626216,3.3472774,3.7142432,4.1120753,3.3850029,3.4776018,3.8479972,4.2046742,4.4859004,5.267846,5.3330083,5.0414934,4.540774,3.7725463,3.5290456,3.3198407,3.4535947,3.8342788,3.9646032,2.9631636,2.8637056,2.7916842,2.4384367,2.0886188,1.3169615,0.8848336,0.7099246,0.6790583,0.64819205,1.1317638,1.4404267,1.920569,2.5070283,2.7368107,2.5893385,3.2512488,4.3624353,5.518206,6.2487082,6.1321025,6.2898636,6.111525,5.658819,5.6828265,4.6402316,4.431027,4.852866,5.675967,6.6568294,6.800872,5.48734,4.262977,3.532475,2.5310357,2.633923,2.9082901,3.1037767,3.0660512,2.7299516,2.1640697,2.5241764,3.059192,3.1072063,2.1057668,2.352697,2.3664153,2.7539587,3.3301294,3.1243541,2.194936,1.8965619,1.9102802,1.8245405,1.1489118,1.9891608,2.4487255,2.5996273,2.6613598,2.976882,2.9803114,3.4467354,3.5633414,3.1483612,2.6373527,2.0646117,2.1194851,2.3561265,2.5447538,2.7059445,3.2135234,2.959734,2.3218307,1.7422304,1.7319417,1.5330256,1.1592005,2.5996273,4.431027,1.8313997,6.7185616,4.4687524,2.5584722,3.2718265,3.6970954,4.616225,5.188966,4.863155,3.8479972,3.1312134,2.651071,2.318401,1.9239986,1.4953002,1.3238207,1.0425946,0.89169276,0.9259886,1.2106444,1.8245405,2.2600982,2.3046827,2.3252604,2.3972816,2.3286898,2.393852,2.8568463,3.2032347,3.7622573,5.7274113,6.910619,7.798882,8.22758,8.131552,7.582818,7.438775,6.8385973,6.0223556,5.4976287,6.060081,5.813151,5.206114,5.0277753,5.422178,5.885172,6.5710897,6.619104,6.1766872,5.422178,4.5784993,3.525616,3.0729103,2.6304936,2.177788,2.2395205,2.6785078,2.7299516,2.6373527,2.4555845,2.0646117,1.7490896,1.670209,1.6770682,1.6016173,1.2620882,0.9842916,0.84367853,0.84024894,0.922559,0.97057325,0.980862,1.0460242,1.1763484,1.3238207,1.3512574,1.2449403,1.3443983,1.5193073,1.7147937,1.9514352,2.054323,2.2360911,2.5241764,2.668219,2.1572106,2.534465,2.7985435,3.0900583,3.2478194,2.8294096,2.4075704,1.8416885,1.4369972,1.1797781,0.7613684,0.69963586,0.7510797,0.69963586,0.69963586,1.2620882,1.5330256,1.9445761,2.4007113,2.8911421,3.474172,2.9631636,3.3472774,3.8720043,3.9886103,3.3438478,3.309552,3.6970954,3.8274195,3.5461934,3.2135234,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.041155048,0.1097468,0.28122616,0.50757897,0.64133286,0.83681935,1.0871792,1.3684053,1.6599203,1.9514352,2.0749004,2.170929,2.1263442,1.978872,1.8931323,1.8416885,2.0886188,2.3424082,2.5550427,2.884283,2.8225505,2.935727,2.9494452,2.843128,2.867135,3.1380725,3.3232703,3.542764,3.841138,4.197815,4.537344,4.40359,4.434457,4.681387,4.6093655,4.547633,4.413879,4.1635194,3.6868064,2.8088322,2.7470996,3.0797696,3.2821152,3.083199,2.4727325,2.668219,2.3767042,2.1400626,2.1023371,2.0303159,2.6647894,3.316411,3.9165888,4.307562,4.273266,4.6402316,6.341307,7.963502,8.549961,7.599966,7.7097125,8.1487,8.793462,9.091836,8.042382,8.762596,10.388221,11.46854,11.71547,12.010415,11.849225,11.729189,12.1921835,12.9707,12.9707,11.235329,10.813489,11.269625,11.948683,11.948683,11.982979,11.516555,11.742908,12.826657,13.900118,12.55915,11.938394,11.375941,10.765475,10.5597,12.034423,13.999576,15.066177,15.2033615,15.717799,15.680074,15.158776,14.212211,13.46799,14.112752,13.419975,13.684054,14.898128,16.173935,15.748666,15.577187,15.388559,14.750656,13.989287,14.160767,15.3817,16.894148,18.348293,19.356592,19.514353,18.440891,17.504614,17.662374,19.21255,21.77445,21.626978,20.546658,18.965618,17.271402,15.806969,15.162207,15.155347,15.357693,15.481158,15.395418,15.604623,15.755525,15.6526375,15.46058,15.717799,15.412566,15.415996,15.501736,15.525743,15.443433,15.721229,16.177364,16.21509,15.868701,15.806969,15.7966795,15.693792,15.8138275,15.892709,15.076467,14.918706,15.79325,16.55119,16.671225,16.280252,15.597764,15.837835,16.362562,16.835844,17.226818,17.63151,18.005335,17.919594,17.470318,17.288551,16.578627,16.191082,16.228807,16.424294,16.143068,15.227368,14.5414505,14.085316,14.003006,14.603184,14.589465,14.815818,14.901558,14.918706,15.395418,14.7369375,14.095605,14.448852,16.101913,18.677534,20.361462,20.186552,19.459478,18.917604,18.722118,17.905876,17.29884,17.189093,17.391438,17.257685,17.28169,17.655516,18.307138,18.739265,18.022482,17.923023,17.367432,16.80498,16.63007,17.165085,17.984756,17.703531,17.271402,17.250826,17.837284,18.20425,17.809847,16.96274,15.844694,14.527733,14.733508,15.498305,15.927004,15.758954,15.3817,15.196502,15.134769,15.035312,14.867262,14.7095,15.477728,15.971589,16.362562,16.774113,17.271402,16.650646,16.300829,15.748666,14.973578,14.435134,13.581166,13.275933,13.227919,13.173045,12.895248,13.234778,13.248496,13.491997,13.697772,12.758065,12.792361,13.022143,12.418536,11.372512,11.705182,11.763485,12.723769,13.258785,12.991278,12.466551,13.749216,15.028452,13.279363,10.820349,15.350834,11.931535,11.619442,13.392539,15.361122,14.740367,14.363112,15.885849,17.065628,17.141079,16.859852,17.250826,15.4914465,17.4566,23.568125,28.791388,17.367432,12.689473,10.254466,8.186425,7.2467184,4.636802,6.042933,12.394529,16.317978,2.1194851,2.510458,9.740028,15.752095,16.976458,14.328816,4.0023284,6.9380555,6.992929,2.942586,8.484799,6.543653,5.271276,4.695105,5.703404,10.024684,10.477389,10.103564,8.186425,6.0806584,7.2158523,9.146709,10.103564,10.415657,10.443094,10.590566,12.493987,13.574307,11.506266,7.6616983,7.1266828,5.6485305,8.848335,8.855195,6.217842,9.901219,11.050131,12.106443,9.736599,5.761707,7.140401,5.9434752,6.468202,4.722542,1.3101025,1.4198492,3.0900583,3.216953,4.0537724,5.2506986,3.8445675,3.5873485,2.7573884,1.821111,1.1249046,0.8711152,0.48014224,0.26407823,0.12689474,0.041155048,0.030866288,0.041155048,0.1371835,0.31895164,0.65505123,1.2655178,1.1317638,0.9877212,0.8711152,0.7990939,0.7613684,0.48357183,0.3841138,0.41498008,0.4698535,0.39783216,0.5178677,0.6241849,0.7510797,0.89169276,0.9774324,1.1111864,0.9259886,0.864256,0.9774324,0.91569984,0.7442205,0.764798,0.8505377,0.90198153,0.84024894,0.9842916,1.1043272,1.1660597,1.1249046,0.9294182,0.96714365,1.2895249,1.3546871,1.2037852,1.4507155,1.8999915,2.0680413,2.0989075,2.0406046,1.845118,1.9925903,2.201795,2.287535,2.2566686,2.318401,2.4898806,2.5138876,2.7951138,3.2546785,3.340418,3.7931237,4.108646,4.3933015,4.5784993,4.3933015,3.4913201,2.9082901,3.525616,4.5510626,3.525616,2.9391565,2.9940298,2.651071,2.054323,2.5173173,2.1640697,2.4315774,2.651071,2.901431,4.012617,2.2669573,6.7391396,7.257007,3.0900583,2.9460156,3.7622573,5.4496145,5.627953,4.2389703,3.5564823,2.651071,5.658819,7.73372,6.492209,1.9994495,11.008976,12.490558,9.108984,4.3590055,2.5653315,3.333559,4.029765,4.338428,5.0586414,8.086967,6.3790326,5.0277753,3.391862,1.6839274,0.9774324,3.6627994,5.8337283,7.7885933,9.445084,10.360784,15.755525,27.916842,30.969175,23.27318,17.425734,12.775213,7.0443726,3.1072063,1.821111,2.0303159,0.91912943,4.3761535,4.5647807,1.6770682,3.9371665,4.0229063,5.4804807,9.057541,10.525404,0.6859175,0.6241849,0.7099246,0.9911508,1.4575747,2.0440342,2.3149714,2.7299516,3.093488,3.4535947,4.0880685,3.7108135,3.5976372,3.8548563,4.389872,4.914599,5.597087,5.703404,5.5147767,5.103226,4.3349986,3.9543142,3.6319332,4.0023284,5.0003386,5.844017,3.474172,3.350707,3.7108135,3.6387923,3.0523329,1.3924125,0.8745448,0.881404,0.9294182,0.67219913,0.84367853,1.5090185,2.2223728,2.7985435,3.309552,3.2512488,3.508468,3.974892,4.7602673,6.2247014,5.7377,5.1580997,4.822,4.523626,3.508468,2.8396983,2.9631636,3.3369887,3.9200184,5.2026844,6.375603,6.210983,5.562791,4.605936,2.8225505,3.2855449,3.5599117,3.5873485,3.4776018,3.4638834,3.059192,3.57363,4.170378,4.180667,3.083199,3.4844608,3.309552,2.9494452,3.1140654,4.822,3.0043187,2.037175,1.5638919,1.3169615,1.097468,1.8416885,2.386993,2.4727325,2.1812177,1.937717,2.3046827,2.3046827,2.352697,2.503599,2.4418662,2.0131679,1.8897027,2.037175,2.194936,1.8759843,1.961724,2.3595562,2.609916,2.5619018,2.3801336,1.5261664,0.864256,1.4678634,3.0146074,3.782835,6.6396813,4.0606318,2.270387,3.0386145,3.6627994,3.7108135,4.0434837,4.0674906,3.74168,3.5702004,3.0214665,2.8568463,2.3389788,1.5433143,1.371835,1.1900668,1.0631721,1.0631721,1.2998136,1.9239986,2.386993,2.301253,2.0989075,1.9239986,1.6324836,1.8656956,2.435007,2.9117198,3.4947495,5.020916,6.8763227,7.936065,8.134981,7.534804,6.3035817,6.5470824,6.368744,5.802862,5.2438393,5.4633327,5.2438393,5.1066556,5.06893,5.2026844,5.6313825,6.509357,7.0306544,6.7459984,5.7377,4.6402316,3.4776018,2.860276,2.4144297,2.1057668,2.2292318,2.3149714,2.5721905,2.9563043,3.1655092,2.6407824,2.369845,1.7559488,1.3752645,1.2998136,1.0666018,0.89855194,0.70649505,0.67219913,0.7613684,0.7613684,0.90884066,0.89169276,1.0425946,1.3752645,1.5707511,1.4267083,1.1489118,1.1214751,1.4267083,1.8931323,1.5638919,1.6084765,1.9925903,2.3664153,2.061182,1.9514352,1.99602,2.318401,2.7916842,3.0351849,2.877424,2.0886188,1.371835,0.9842916,0.70306545,0.6276145,0.64819205,0.66533995,0.7510797,1.1283343,1.8005334,2.253239,2.784825,3.3129816,3.3884325,2.935727,3.2889743,3.6970954,3.6387923,2.8088322,2.976882,3.707384,4.2389703,4.2526884,3.8617156,0.0,0.010288762,0.020577524,0.037725464,0.09602845,0.23664154,0.3566771,0.47328308,0.5761707,0.69963586,0.922559,1.155771,1.2620882,1.3684053,1.6736387,2.452155,2.136633,2.1572106,2.1674993,2.07833,2.0508933,2.0886188,2.2841053,2.4624438,2.5927682,2.784825,2.9288676,2.9254382,2.860276,2.8088322,2.843128,2.935727,3.1243541,3.3884325,3.6559403,3.806842,3.806842,3.9886103,4.190956,4.3624353,4.57164,4.108646,3.8617156,3.5873485,3.1037767,2.2841053,2.5447538,2.4967396,2.3835633,2.277246,2.0577524,1.8313997,1.7799559,1.7525192,1.7765263,2.054323,2.7162333,3.223812,3.6525106,3.8685746,3.5290456,4.0606318,5.5559316,7.6445503,9.414218,9.417647,8.913498,9.386781,9.870353,10.000677,10.041832,10.30591,10.206452,10.045261,9.945804,9.849775,10.48082,11.084427,11.866373,12.507706,12.164746,11.369082,10.834066,11.122152,12.092726,12.922686,12.854094,13.004995,13.272504,13.680624,14.363112,13.354814,12.079007,11.588576,11.931535,12.133881,11.979549,12.919256,14.421415,15.666355,15.54632,15.333686,14.54831,13.564018,12.902108,13.234778,13.917266,14.085316,15.268523,17.254255,18.115082,18.440891,18.070496,16.87357,15.645778,16.088194,17.53548,18.722118,19.70298,20.4472,20.872469,20.217419,18.893597,17.61779,17.247395,18.79757,20.310017,20.807306,20.100813,18.71183,17.87158,17.096493,16.187653,15.621771,15.443433,15.261664,15.323397,15.717799,16.002455,16.016174,15.861842,15.978448,15.9921665,16.12935,16.417435,16.722668,16.654078,16.938732,17.175373,17.069057,16.431154,16.331696,16.101913,16.21852,16.410576,15.662926,15.014734,16.002455,16.746675,16.616352,16.245956,15.542891,15.3817,15.662926,16.256245,17.007324,17.312557,17.449741,17.487467,17.439453,17.274832,16.29397,16.108772,16.287111,16.489456,16.47231,15.841265,15.54632,15.0456,14.452282,14.555169,15.323397,15.532601,15.193072,14.867262,15.666355,15.728088,15.450292,15.769243,16.942162,18.54378,20.412905,20.937632,20.656404,20.159115,20.100813,19.078794,18.478617,18.091074,17.802988,17.600643,18.053349,17.902447,17.751545,17.71382,17.436022,16.88729,16.489456,16.173935,16.11906,16.763824,16.935303,16.582056,16.232237,16.160215,16.386568,16.088194,15.659496,15.059319,14.407697,13.975569,14.359683,15.289101,15.700651,15.350834,14.79524,13.996146,13.4645605,13.423406,13.797231,14.184773,15.169065,15.29253,15.46744,15.837835,15.772673,15.676644,15.848124,15.728088,15.371411,15.46058,14.490007,14.006435,13.567448,13.059869,12.710052,13.121602,13.334236,13.564018,13.615462,12.891819,13.094165,12.682614,12.284782,12.5145645,13.985858,14.027013,14.256795,13.869251,13.317088,14.284232,12.538571,12.319078,12.30536,12.0138445,11.787492,11.97269,14.095605,14.997586,14.352823,14.668345,16.407146,17.079346,17.264544,17.610931,18.814716,20.104242,17.137648,16.918156,19.161106,16.317978,15.155347,13.958421,10.751757,6.2727156,3.9783216,2.6236343,4.2355404,5.7308407,5.7719955,4.756838,9.191295,14.839825,12.905538,6.3310184,9.774324,3.940596,5.658819,5.7377,3.4707425,6.6396813,5.020916,4.6436615,5.754848,7.3393173,7.1198235,9.211872,9.623423,9.297611,8.954653,9.084977,8.81747,9.863494,10.652299,10.741467,10.81006,11.091286,9.599416,8.786603,9.160428,9.297611,6.914048,7.06838,6.9380555,6.1904054,6.9963584,8.176137,8.086967,7.798882,7.5039372,6.5196457,6.1321025,5.7308407,4.629943,3.4124396,3.9200184,6.3653145,5.9812007,5.195825,4.5956473,2.9288676,3.4433057,3.1277838,2.2600982,1.255229,0.6379033,0.6859175,0.3806842,0.1097468,0.020577524,0.017147938,0.020577524,0.082310095,0.18519773,0.42526886,1.0357354,1.0460242,1.0288762,0.9328478,0.8128122,0.83681935,0.5658819,0.50757897,0.48014224,0.4081209,0.32238123,0.47328308,0.61389613,0.66876954,0.6790583,0.7922347,0.9294182,0.8505377,0.90198153,1.097468,1.1351935,1.0220171,0.90541106,0.7888051,0.72364295,0.77851635,0.83681935,0.77851635,0.7888051,0.88826317,0.96714365,1.1592005,1.3958421,1.4232788,1.2792361,1.2792361,1.4164196,1.5741806,1.6324836,1.5913286,1.5536032,1.4644338,1.5501735,1.6599203,1.6942163,1.5981878,1.7593783,2.1846473,2.5619018,2.7745364,2.8911421,3.3987212,3.7794054,3.8102717,3.4535947,2.8808534,2.4452958,2.3629858,2.7882545,3.7759757,5.271276,4.420738,4.197815,3.4467354,2.4007113,2.6887965,4.756838,5.219832,5.1580997,5.2987127,6.0395036,4.0777793,5.360445,5.953764,4.633373,2.8945718,2.201795,4.2869844,5.857735,5.6999745,4.6676683,4.4550343,4.756838,6.7391396,7.864044,1.8897027,3.9440255,3.5290456,2.9700227,3.234101,3.9303071,3.2443898,2.6750782,3.875434,6.451054,7.963502,4.3109913,2.877424,2.054323,2.3835633,6.56766,10.347065,12.0309925,11.423956,10.021255,10.995257,15.902997,22.096832,26.126596,25.564144,19.013634,9.410788,6.1321025,5.878313,5.3673043,1.3443983,1.0837497,1.4369972,1.9685832,3.0969174,6.0978065,4.465323,3.9783216,4.091498,3.649081,0.8711152,0.53501564,0.58988905,1.1249046,1.8382589,2.0337453,2.3218307,3.0626216,3.3987212,3.2821152,3.4673128,3.7931237,3.590778,3.6113555,4.016047,4.3761535,4.6779575,5.188966,5.346727,5.0414934,4.6127954,4.081209,3.923448,3.8925817,4.0434837,4.722542,4.091498,4.1943855,4.033195,3.5290456,3.5393343,3.0900583,2.3424082,1.6496316,1.2003556,1.0117283,0.84367853,1.2106444,1.7147937,2.1880767,2.702515,2.8156912,3.2512488,3.5290456,3.683377,4.249259,4.5030484,4.523626,4.5270553,4.530485,4.3761535,3.7519686,3.4295874,3.57363,4.0880685,4.616225,5.5833683,5.9914894,5.3913116,4.012617,2.7368107,3.1346428,3.7039545,4.0057583,3.957744,3.8171308,4.0023284,5.0346346,5.909179,6.108095,5.597087,4.2526884,3.3850029,3.0111778,3.234101,4.2595477,4.756838,4.0366244,3.000889,2.1572106,1.6221949,1.646202,1.8828435,2.085189,1.9685832,1.2175035,1.4850113,1.5776103,1.5364552,1.546744,1.9651536,2.153781,1.9411465,1.7353712,1.6256244,1.3752645,1.3924125,1.6324836,2.1126258,2.5756202,2.4898806,1.937717,2.1126258,1.9994495,2.1640697,4.7602673,3.2821152,2.633923,3.0283258,3.8514268,3.6627994,3.673088,4.1326528,4.383013,4.190956,3.765687,3.333559,3.0797696,2.568761,1.8108221,1.2895249,1.2895249,1.2243627,1.1317638,1.1866373,1.704505,1.8142518,1.8176813,1.7833855,1.704505,1.4987297,2.0337453,2.510458,2.7813954,3.1072063,4.15323,6.1766872,7.298162,7.56224,7.394191,7.596536,6.9037595,6.40304,5.919468,5.5422134,5.645101,5.5147767,5.501058,5.470192,5.353586,5.15467,5.456474,6.1492505,6.468202,6.0635104,5.003768,3.875434,2.9906003,2.3149714,1.8725548,1.7388009,2.0577524,2.3629858,2.760818,3.0969174,2.9322972,2.3629858,1.8313997,1.7113642,1.8348293,1.4953002,1.0494537,0.78537554,0.607037,0.5144381,0.59331864,0.7099246,0.6893471,0.7888051,0.99801,1.0460242,1.0666018,1.0082988,0.89169276,0.90198153,1.4164196,1.2826657,1.3409687,1.6907866,2.095478,1.9857311,1.7593783,1.6290541,1.9274281,2.49331,2.6716487,2.8739944,2.253239,1.4507155,0.85396725,0.59331864,0.45956472,0.53844523,0.6379033,0.7339317,0.94656616,1.5090185,2.0508933,2.5619018,3.000889,3.2889743,3.3747141,3.841138,4.1635194,4.256118,4.479041,4.5819287,4.4447455,4.0880685,3.8548563,4.420738,0.06516216,0.12003556,0.20234565,0.32581082,0.4698535,0.58302987,0.64819205,0.71678376,0.8265306,0.9534253,1.039165,1.2175035,1.2860953,1.4438564,1.8108221,2.452155,2.3149714,2.294394,2.2635276,2.2155135,2.2566686,2.4041407,2.5001693,2.5584722,2.5824795,2.5893385,2.8328393,2.9734523,3.0077481,3.0043187,3.07634,3.2786856,3.2889743,3.275256,3.3232703,3.450165,3.4981792,3.7382503,4.029765,4.197815,4.040054,3.4364467,3.0797696,2.7779658,2.4212887,2.0063086,2.2086544,2.1572106,2.0028791,1.8142518,1.5673214,1.4575747,1.5604624,1.7216529,1.8691251,2.0131679,2.4967396,3.0111778,3.3472774,3.4467354,3.3952916,4.5339146,5.754848,7.5725293,9.544542,10.2921915,9.801761,10.419086,10.851214,10.738038,10.652299,11.026124,10.326488,9.80862,9.671436,9.043822,9.321619,9.89436,10.460241,10.861504,11.05699,11.235329,11.279913,11.732618,12.566009,13.186764,13.433694,13.104454,12.686044,12.854094,14.479718,14.198492,13.413116,13.152468,13.272504,12.47341,12.576297,12.977559,13.886399,14.874121,14.88098,14.764374,14.057879,13.498857,13.354814,13.426835,13.858963,13.924125,14.428274,15.37827,15.9613,16.770683,17.899017,18.348293,18.149376,18.348293,19.555508,20.227707,20.45063,20.299728,19.836735,20.107672,19.997925,19.19197,18.094503,17.823566,18.331144,18.897026,18.996485,18.564358,17.974468,17.53548,17.031332,16.386568,15.512024,14.29452,14.421415,15.073037,15.553179,15.515453,14.973578,15.127911,15.3817,15.830976,16.424294,16.979887,17.662374,18.20082,18.142517,17.686382,17.665806,17.405157,17.408587,17.477179,17.353712,16.722668,15.9750185,16.146498,16.37971,16.317978,16.108772,15.676644,15.179354,14.956431,15.162207,15.772673,16.146498,16.45859,16.654078,16.746675,16.80498,16.37971,16.21166,16.167076,16.235666,16.54776,16.276823,15.721229,15.110763,14.678635,14.668345,15.042171,15.450292,15.443433,15.182784,15.440002,16.12249,16.448301,16.849564,17.590355,18.756414,20.35803,21.03709,21.071384,20.752434,20.392326,19.757853,18.938183,18.142517,17.645227,17.823566,18.362011,18.36544,18.097933,17.782412,17.62808,16.609491,16.20137,16.321407,16.698662,16.87357,16.643787,15.940722,15.391989,15.206791,15.179354,14.942713,14.79524,14.3974085,13.821238,13.557159,14.020154,14.55174,14.819247,14.726648,14.428274,13.680624,13.430264,13.430264,13.533153,13.670336,14.640909,14.808959,15.0250225,15.357693,15.083325,15.306249,15.861842,15.87899,15.518884,15.981877,15.374841,14.527733,13.906977,13.697772,13.807519,13.7526455,13.588025,13.642899,13.831526,13.618892,14.033872,13.437123,13.29994,14.037301,15.031882,15.083325,15.71437,17.315987,18.687822,17.055338,12.912396,11.821788,12.205902,12.257345,9.925226,10.909517,12.140739,12.672326,13.152468,15.810398,16.273392,16.832415,18.386019,20.056227,19.19197,19.11652,15.059319,15.453721,18.70154,13.162757,12.295071,10.89237,8.64256,5.686256,2.609916,1.4095604,1.9994495,2.1091962,2.9151495,9.040393,9.571979,12.116733,10.247607,6.293293,11.365653,6.3961806,6.4098988,6.4098988,5.130663,5.0277753,3.5461934,4.262977,6.3378778,8.052671,6.8145905,8.879202,9.39707,9.788043,10.233889,9.6817255,8.351046,10.034973,11.321068,10.607714,8.134981,7.473071,7.689135,7.9875093,8.436785,9.9869585,7.8503256,6.046363,5.761707,6.334448,5.2644167,6.5230756,5.8988905,5.9434752,6.9723516,7.058091,7.3427467,7.3358874,7.5416627,7.4284863,5.425607,5.2781353,4.664239,3.8274195,3.0969174,2.8945718,3.1552205,2.8637056,2.1297739,1.2380811,0.65162164,0.70306545,0.5007198,0.22292319,0.01371835,0.01371835,0.006859175,0.037725464,0.12003556,0.29494452,0.65505123,0.77851635,0.91912943,0.9774324,0.96371406,0.9911508,0.7373613,0.548734,0.45613512,0.41840968,0.34295875,0.4698535,0.5624523,0.61046654,0.6379033,0.70306545,0.70306545,0.8265306,0.9877212,1.138623,1.2346514,1.3203912,1.2483698,1.1146159,0.9568549,0.72707254,0.70306545,0.6756287,0.6927767,0.7579388,0.84024894,1.0185875,1.2655178,1.4164196,1.4129901,1.3101025,1.1592005,1.1694894,1.2620882,1.3889829,1.5364552,1.3512574,1.2723769,1.214074,1.1694894,1.1797781,1.3341095,1.6427724,2.0131679,2.3081124,2.3286898,2.6545007,3.0797696,3.199805,2.8396983,2.0440342,1.9171394,2.1297739,2.5447538,3.5221863,5.909179,5.2335505,4.5613513,3.625074,2.8739944,3.4913201,4.979761,4.822,5.0620713,5.802862,5.1821065,2.9048605,2.726522,4.3281393,5.9160385,4.2115335,3.0866287,4.2355404,5.796003,6.6568294,6.464772,7.085528,6.4098988,6.118384,6.025785,4.057202,4.1326528,3.8788633,3.6696587,4.4104495,7.5588107,6.258997,4.389872,4.8014226,6.4716315,4.5030484,3.40901,2.1880767,1.3546871,1.8279701,4.945465,6.2864337,8.512236,9.050681,8.004657,8.152129,10.357354,13.687484,17.312557,19.085653,15.54632,7.7748747,5.9880595,5.597087,4.139512,1.2586586,1.6770682,1.6942163,2.5619018,4.448175,6.416758,4.619654,2.7985435,1.7765263,1.4095604,0.59674823,0.4938606,0.5212973,1.0254467,1.786815,2.0028791,2.2429502,3.018037,3.316411,3.059192,3.0729103,3.6627994,3.4981792,3.4947495,3.8034124,3.8205605,3.9543142,4.413879,4.846007,5.0174866,4.8322887,4.2423997,4.214963,4.105216,3.9200184,4.32128,4.139512,4.081209,3.9474552,3.7348208,3.6079261,3.2478194,2.8054025,2.1194851,1.4198492,1.3443983,1.2860953,1.3752645,1.5947582,2.0646117,3.0523329,3.333559,3.532475,3.6285036,3.6147852,3.4878905,3.7382503,4.0057583,4.2595477,4.372724,4.125794,4.012617,3.6044965,3.6936657,4.2081037,4.2046742,4.822,5.2987127,4.9351764,3.9303071,3.4192986,2.877424,3.4707425,4.091498,4.32471,4.4550343,4.417309,5.07236,5.7651367,6.108095,5.970912,4.976331,4.3178506,3.940596,3.9165888,4.413879,4.57164,4.7019644,4.2835546,3.3678548,2.5893385,2.07833,1.8931323,1.8108221,1.6221949,1.138623,1.0666018,1.0494537,0.94999576,0.922559,1.4164196,1.7353712,1.611906,1.3375391,1.1249046,1.1146159,0.89512235,1.0837497,1.5364552,2.1091962,2.6647894,2.4658735,3.0866287,2.976882,2.3252604,3.0557625,2.0131679,2.1880767,3.0317552,3.7039545,3.0489032,3.3850029,3.957744,4.389872,4.4447455,4.0434837,3.765687,3.5153272,3.0866287,2.411,1.5604624,1.5124481,1.5913286,1.5776103,1.546744,1.8691251,1.8108221,1.937717,2.1297739,2.2395205,2.07833,2.534465,2.9185789,3.1346428,3.3198407,3.8445675,5.9228973,7.058091,7.377043,7.157549,6.848886,6.4990683,6.2247014,5.970912,5.7719955,5.7274113,5.113515,5.038064,5.171818,5.3432975,5.528495,6.090947,6.7940125,7.2535777,7.0923867,5.9469047,4.3281393,3.2409601,2.5961976,2.2669573,2.1023371,2.2669573,2.5173173,2.7402403,2.843128,2.7779658,2.07833,1.6942163,1.6976458,1.821111,1.4472859,1.0357354,0.8162418,0.6893471,0.61389613,0.58645946,0.6001778,0.70649505,0.7956643,0.8162418,0.77851635,0.8471081,0.8128122,0.72707254,0.70306545,0.91227025,1.0185875,1.0666018,1.2380811,1.5536032,1.8588364,1.6599203,1.529596,1.7388009,2.1229146,2.085189,2.3321195,2.0406046,1.5844694,1.1934965,0.9568549,0.6859175,0.7099246,0.9602845,1.3375391,1.7147937,1.8142518,2.2841053,2.7128036,3.0454736,3.5770597,3.8548563,4.32471,4.7499785,5.003768,5.0826488,5.3570156,5.456474,5.003768,4.431027,4.972902,0.33266997,0.3806842,0.45270553,0.5624523,0.7133542,0.88826317,0.9328478,0.97400284,1.08032,1.2106444,1.1900668,1.3203912,1.4987297,1.7525192,2.1091962,2.5893385,2.4418662,2.3492675,2.2909644,2.301253,2.49331,2.5447538,2.4624438,2.4041407,2.4007113,2.3561265,2.651071,2.942586,3.1552205,3.2615378,3.2649672,3.40901,3.3266997,3.1895163,3.1586502,3.40901,3.5187566,3.6113555,3.7348208,3.7485392,3.2958336,2.7985435,2.4761622,2.1880767,1.920569,1.7902447,1.9171394,1.8999915,1.7971039,1.6153357,1.3238207,1.3272504,1.4953002,1.821111,2.1434922,2.1194851,2.5756202,2.9700227,3.2135234,3.3678548,3.666229,5.164959,6.3138704,7.706283,9.146709,9.671436,9.716022,10.600855,11.177026,11.156448,11.111863,11.880091,11.38623,10.786053,10.275044,9.091836,8.971801,9.136421,9.3079,9.534253,10.203023,10.902658,11.441104,12.082437,12.734058,12.943263,13.077017,12.46998,11.96926,12.195613,13.560589,13.745787,13.306799,13.149038,13.341095,13.13189,13.677195,13.306799,13.011855,13.334236,14.366542,14.781522,14.819247,14.874121,14.994157,14.887839,14.5243025,14.160767,13.965281,13.965281,14.057879,14.507155,15.87213,17.525192,18.924463,19.61724,20.35803,20.76958,20.714708,20.20027,19.384027,19.569225,19.644676,19.288,18.519772,17.693241,17.29541,17.315987,17.370861,17.29541,17.134218,17.158226,17.391438,17.031332,15.80011,13.9481325,13.598314,14.359683,15.172495,15.357693,14.589465,14.685493,14.88441,15.429714,16.235666,16.88729,17.988186,18.838724,18.910746,18.478617,18.61923,18.187103,18.115082,18.115082,18.070496,18.02934,17.703531,17.161655,16.63007,16.194511,15.7966795,15.6697855,15.29939,14.819247,14.46943,14.599753,14.71636,15.001016,15.275383,15.4914465,15.738377,15.9750185,16.163645,16.20137,16.184223,16.393429,16.170506,15.755525,15.22051,14.7369375,14.589465,14.493437,14.898128,15.223939,15.309678,15.409137,15.999025,16.671225,17.233677,17.734396,18.437462,19.871029,20.659836,20.923914,20.773012,20.320305,20.152256,19.178253,18.12537,17.525192,17.71382,18.118511,18.190533,17.919594,17.61436,17.909306,16.986746,16.475739,16.558048,16.955881,16.928444,16.482597,15.570327,14.730078,14.260224,14.225929,14.284232,14.198492,13.749216,13.166186,13.104454,13.413116,13.780083,14.013294,14.037301,13.893259,13.588025,13.954991,14.174485,14.033872,13.924125,14.627191,14.699212,14.956431,15.429714,15.371411,15.556609,15.837835,15.738377,15.556609,16.37285,16.047039,15.364552,14.819247,14.706071,15.134769,14.500296,13.893259,13.780083,14.174485,14.658057,15.066177,14.747226,14.898128,15.563468,15.635489,15.704081,16.393429,18.231688,19.442331,15.944152,12.188754,11.852654,12.089295,11.382801,9.56512,10.549411,10.268185,10.88551,13.029003,15.786391,15.374841,17.384579,20.063087,21.067955,17.477179,15.069608,10.288762,10.796341,14.987297,12.003556,9.692014,8.018375,6.5299344,4.6779575,1.845118,0.83681935,1.3581166,2.5241764,5.857735,15.29253,11.4376745,9.301042,7.534804,7.2707253,12.147599,8.1212635,7.870903,7.7028537,6.2727156,4.5990767,5.096367,6.3138704,7.8983397,8.999237,8.285883,8.834618,9.040393,9.853205,10.8958,10.48082,9.081548,10.299051,10.539123,9.160428,8.488229,6.279575,6.9552035,7.31531,7.3187394,10.086417,8.100685,5.8371577,5.5730796,6.3961806,4.214963,6.5230756,6.0086374,5.9571934,7.0889573,7.548522,7.6033955,7.380472,8.025234,8.381912,4.979761,2.9460156,2.2806756,2.2498093,2.5173173,3.1449318,2.5996273,2.2395205,1.8691251,1.3684053,0.6962063,0.5590228,0.5693115,0.36353627,0.01371835,0.01371835,0.0034295875,0.030866288,0.09259886,0.20920484,0.42526886,0.70306545,1.0666018,1.155771,1.0254467,1.138623,0.8128122,0.53501564,0.40126175,0.39097297,0.36696586,0.42869842,0.4629943,0.52815646,0.607037,0.6173257,0.61389613,0.8128122,1.0357354,1.1866373,1.2415106,1.5227368,1.5638919,1.529596,1.3992717,0.96371406,0.805953,0.7510797,0.72707254,0.7099246,0.7339317,0.91569984,1.1214751,1.3306799,1.471293,1.430138,1.1420527,0.9945804,1.039165,1.2312219,1.430138,1.2483698,1.1008976,0.9259886,0.77851635,0.83338976,0.9294182,1.0666018,1.371835,1.7216529,1.7113642,1.7216529,2.1297739,2.3664153,2.1332035,1.3855534,1.4404267,1.7388009,2.2052248,3.0248961,4.6573796,4.3487167,4.2115335,4.1429415,4.07435,3.9851806,4.149801,4.341858,5.295283,6.6739774,7.0752387,4.839148,4.7979927,6.276145,7.4181976,5.212973,5.7582774,7.932636,9.414218,8.988949,6.550512,7.846896,7.8331776,6.0086374,4.1772375,6.4887795,5.0312047,5.346727,5.73427,6.543653,10.179015,9.009526,8.05953,8.049242,7.5039372,2.7368107,3.6044965,2.3595562,1.2929544,1.611906,3.4433057,2.5481834,4.928317,6.8454566,6.6568294,4.8082814,7.332458,8.903209,10.981539,12.614022,10.456812,5.871454,5.7239814,4.98662,2.6887965,1.9239986,2.5996273,2.2326615,2.4658735,3.5530527,4.355576,3.9268777,2.1229146,1.2106444,1.3821237,0.7407909,0.6241849,0.6927767,1.08032,1.6804979,2.16064,2.6716487,3.1415021,3.309552,3.1552205,2.8911421,3.2203827,3.1312134,3.2443898,3.4981792,3.1792276,3.457024,3.6970954,4.1429415,4.6882463,4.8905916,4.2938433,4.3521466,4.3761535,4.190956,4.1326528,4.1429415,3.974892,3.9611735,4.012617,3.625074,3.1826572,2.9631636,2.4555845,1.7696671,1.6187652,1.5364552,1.5741806,1.6599203,2.0920484,3.508468,3.7382503,3.7313912,3.7759757,3.8342788,3.5564823,3.3609958,3.5290456,3.8034124,3.9371665,3.7039545,4.0949273,3.957744,3.9200184,4.064061,3.9200184,4.383013,4.6608095,4.4756117,3.9783216,3.724532,2.9906003,3.3952916,4.0846386,4.623084,4.98662,4.866585,5.2575574,5.6210938,5.778855,5.9126086,5.206114,4.4756117,3.9303071,3.7142432,3.9063,3.9714622,4.6402316,4.7979927,4.2218223,3.5873485,2.976882,2.4247184,1.9137098,1.4610043,1.1214751,0.8676856,0.8093826,0.7407909,0.6859175,0.8848336,1.2483698,1.1866373,0.980862,0.88826317,1.1214751,0.7099246,0.78194594,1.0768905,1.5913286,2.5893385,2.9871707,3.6970954,3.8342788,3.2409601,2.4795918,2.1880767,2.2463799,2.767677,3.2512488,2.5721905,3.0626216,3.6970954,4.338428,4.722542,4.4516044,4.256118,3.957744,3.5393343,2.9494452,2.1263442,1.8348293,1.937717,2.0749004,2.1572106,2.3732746,2.2738166,2.4452958,2.7813954,3.0900583,3.1037767,3.350707,3.5118976,3.6936657,3.8891523,3.9851806,5.610805,6.351596,6.660259,6.636252,6.018926,6.1629686,6.042933,5.970912,5.994919,5.9160385,5.130663,4.8905916,4.931747,5.1169443,5.4324665,6.355026,7.006647,7.349606,7.2467184,6.447624,4.928317,3.8960114,3.2203827,2.784825,2.49331,2.6887965,2.7985435,2.860276,2.901431,2.942586,2.3458378,1.821111,1.5947582,1.5707511,1.3478279,1.1180456,0.8779744,0.75450927,0.7373613,0.6962063,0.6379033,0.7476501,0.8025235,0.75450927,0.7339317,0.72707254,0.6859175,0.66876954,0.6824879,0.7099246,0.84367853,0.8848336,0.9294182,1.0734608,1.430138,1.4644338,1.5021594,1.5707511,1.6324836,1.5776103,1.6153357,1.5433143,1.4987297,1.4610043,1.2586586,1.0871792,1.097468,1.4541451,2.0749004,2.6064866,2.5001693,2.9322972,3.175798,3.2272418,3.8102717,4.437886,4.8494368,5.3261495,5.7582774,5.6313825,5.90575,6.1904054,6.183546,5.90575,5.6828265,0.69963586,0.69963586,0.69963586,0.71678376,0.8162418,1.1180456,1.2072148,1.2277923,1.2963841,1.4061309,1.4267083,1.5536032,1.8759843,2.170929,2.435007,2.877424,2.4830213,2.301253,2.218943,2.2600982,2.6167753,2.4487255,2.2120838,2.1091962,2.16064,2.2395205,2.551613,2.8259802,3.1209247,3.3129816,3.100347,3.0248961,3.0111778,3.0214665,3.1312134,3.5016088,3.532475,3.3952916,3.2306714,3.0489032,2.7230926,2.4212887,2.218943,1.978872,1.7079345,1.5673214,1.7010754,1.6736387,1.6667795,1.6496316,1.3924125,1.3615463,1.546744,2.0028791,2.4795918,2.417859,2.901431,3.0969174,3.2718265,3.6079261,4.2046742,5.675967,6.8557453,7.9189177,8.601405,8.220721,8.954653,10.010965,10.768905,11.170166,11.739478,12.881531,12.922686,12.325937,11.317638,9.89093,9.568549,9.153569,8.992378,9.270175,10.0041065,10.587136,11.156448,11.907528,12.668896,12.898679,12.542002,12.103014,12.116733,12.439114,12.233338,12.394529,11.718901,11.393089,12.113303,14.068168,14.788382,13.790371,12.607163,12.439114,14.167625,14.96672,15.875561,16.496315,16.70895,16.657507,16.0539,15.196502,14.459141,14.023583,13.872682,13.615462,13.766364,15.206791,17.638369,19.572655,20.073376,20.69413,20.982216,20.845032,20.563807,20.011642,19.13024,18.557497,18.358582,18.019053,17.62808,17.29541,16.664366,15.978448,16.108772,16.506605,17.182234,17.20624,16.263103,14.627191,13.344524,13.900118,15.021593,15.638919,14.918706,14.994157,15.035312,15.481158,16.252815,16.732958,17.682953,18.650097,19.1954,19.250275,19.11995,18.684393,18.197392,17.974468,18.163095,18.739265,19.106232,18.523201,17.504614,16.424294,15.512024,15.450292,15.539461,15.182784,14.428274,13.978998,13.529722,13.371962,13.629181,14.143619,14.472859,14.96672,15.765814,16.276823,16.338554,16.21852,15.861842,15.920145,15.6252,14.928994,14.500296,14.208781,14.335675,14.699212,15.172495,15.707511,15.769243,16.37285,17.055338,17.55263,17.79613,18.972477,19.87446,20.37518,20.436913,20.141968,20.35803,19.490345,18.399736,17.62465,17.357141,17.432592,17.226818,16.767254,16.53747,17.470318,17.37772,17.021042,16.767254,16.695232,16.619781,16.012743,15.169065,14.157337,13.354814,13.426835,13.728639,13.509145,12.871242,12.274493,12.5145645,12.562579,13.094165,13.461131,13.4474125,13.282792,13.540011,14.352823,14.79524,14.754086,14.908417,15.103903,14.843254,14.997586,15.642348,16.04361,16.21509,15.752095,15.361122,15.532601,16.55119,16.53404,16.393429,15.923574,15.453721,15.824117,14.918706,14.243076,14.126471,14.682064,15.789821,16.143068,16.221949,16.510035,16.774113,16.081335,16.033321,15.906426,15.6869335,14.812388,12.175035,11.0981455,12.140739,11.845795,10.189304,10.563129,10.834066,9.712592,10.731179,13.526293,13.838386,15.357693,19.078794,20.803877,18.70154,13.330807,9.3764925,5.0895076,5.2747054,8.927217,9.218731,7.160979,6.23156,4.955754,3.018037,1.2792361,0.84024894,3.4947495,6.9517736,11.399949,19.500635,14.249936,9.14328,5.871454,5.7891436,9.932085,7.840037,8.927217,8.724871,6.5950966,5.7102633,8.752307,9.746887,10.055551,10.213311,9.935514,8.944365,8.669997,9.451943,10.768905,11.228469,10.583707,10.652299,9.156999,7.689135,11.718901,7.606825,6.5950966,6.3618846,6.800872,10.038403,9.129561,7.740579,7.14726,6.742569,4.0537724,7.706283,7.6959944,7.610255,8.213862,7.459353,6.478491,5.4667625,5.5422134,5.7308407,2.9871707,1.4507155,0.9259886,1.728512,3.1552205,3.4981792,2.2909644,1.903421,1.99602,1.937717,0.7956643,0.5144381,0.65162164,0.50757897,0.072021335,0.01371835,0.006859175,0.041155048,0.07888051,0.15090185,0.36696586,0.7339317,1.255229,1.2895249,0.9602845,1.1592005,0.7579388,0.51100856,0.37039545,0.31895164,0.34638834,0.34638834,0.34295875,0.4115505,0.5144381,0.51100856,0.64819205,0.7888051,1.0048691,1.196926,1.1214751,1.4747226,1.6290541,1.7388009,1.7490896,1.4095604,1.138623,0.9602845,0.881404,0.8745448,0.8745448,0.9945804,1.0460242,1.1694894,1.3752645,1.5536032,1.3203912,1.1008976,1.0185875,1.0940384,1.2312219,1.0940384,0.94999576,0.7579388,0.5658819,0.5212973,0.5212973,0.6036074,0.823101,1.0631721,1.0631721,0.83338976,1.1523414,1.4267083,1.3581166,0.922559,0.97400284,1.1660597,1.6187652,2.1743584,2.4041407,2.4007113,3.333559,4.4756117,5.0003386,3.99204,3.4364467,4.5201964,6.1972647,8.097256,10.545981,9.510246,10.209882,10.213311,8.453933,5.2438393,8.567109,12.939834,13.978998,10.573419,4.8597255,5.9434752,7.4936485,6.0326443,3.508468,7.281014,4.040054,4.3452873,6.258997,8.447074,10.172156,9.630281,11.547421,11.856084,9.033533,4.1326528,4.5201964,3.0317552,1.9651536,2.294394,3.6559403,2.369845,3.9783216,5.8988905,5.98463,2.510458,7.949784,9.002667,9.139851,9.006097,6.4304767,4.2286816,5.147811,4.671098,2.7642474,3.882293,3.799983,2.1091962,1.0357354,1.2072148,1.6359133,2.983741,2.0886188,1.5261664,1.7971039,1.3375391,0.922559,1.0494537,1.3409687,1.7490896,2.534465,3.4878905,3.5599117,3.6044965,3.6182148,2.7299516,2.7573884,2.7985435,2.9906003,3.1209247,2.6476414,3.0557625,3.216953,3.5050385,4.029765,4.6402316,4.149801,4.2252517,4.40359,4.3590055,3.8925817,4.201245,4.1360826,4.1292233,4.1360826,3.6525106,3.3541365,3.1517909,2.8088322,2.3046827,1.8656956,1.4747226,1.5913286,1.762808,2.1743584,3.649081,3.7313912,3.789694,4.0023284,4.2423997,4.0606318,3.175798,3.0454736,3.2272418,3.4295874,3.5050385,4.1292233,4.386442,4.197815,3.8171308,3.8479972,4.2389703,4.2526884,4.166949,3.998899,3.4844608,3.3884325,3.5393343,4.0434837,4.729401,5.164959,5.0586414,5.5593615,5.7719955,5.610805,5.8062916,4.835718,3.7348208,2.9734523,2.7333813,2.9220085,3.625074,4.2046742,4.434457,4.3487167,4.2252517,3.8925817,3.2306714,2.4384367,1.6736387,1.0700313,0.77508676,0.75450927,0.77851635,0.7099246,0.5178677,0.8676856,0.8196714,0.7373613,0.84367853,1.2243627,0.82996017,0.7339317,0.8265306,1.2106444,2.1743584,3.234101,3.882293,4.2526884,4.2526884,3.5942078,2.942586,2.527606,2.568761,2.8019729,2.4898806,2.8122618,3.3438478,4.170378,4.955754,4.955754,4.7945633,4.338428,3.7931237,3.2683969,2.7642474,2.2738166,2.2463799,2.469303,2.784825,3.059192,2.9700227,3.1106358,3.4913201,3.981751,4.2835546,4.3007026,4.1635194,4.256118,4.5099077,4.389872,5.188966,5.2026844,5.4599032,5.9812007,5.809721,6.186976,6.018926,6.0086374,6.2727156,6.334448,5.7822843,5.2987127,4.9351764,4.715683,4.6676683,5.6142344,6.1904054,6.447624,6.4990683,6.550512,5.8817425,5.0277753,4.0880685,3.2203827,2.6545007,3.1140654,3.1072063,3.0900583,3.2306714,3.4021509,3.0866287,2.301253,1.6770682,1.4438564,1.4267083,1.3443983,1.0048691,0.77165717,0.75450927,0.8025235,0.78194594,0.78537554,0.78194594,0.7888051,0.8848336,0.7442205,0.6756287,0.70649505,0.8025235,0.8711152,0.7956643,0.8162418,0.8471081,0.8711152,0.939707,1.2243627,1.5398848,1.5604624,1.3889829,1.5330256,1.1351935,1.0666018,1.255229,1.4850113,1.4129901,1.4507155,1.5158776,1.9342873,2.651071,3.2546785,3.4364467,3.7759757,3.649081,3.350707,4.0709205,5.0757895,5.4324665,5.7822843,6.2487082,6.39961,6.680836,6.677407,7.181556,7.7542973,6.742569,0.8093826,0.85739684,0.91569984,1.0254467,1.1900668,1.371835,1.4335675,1.3306799,1.3306799,1.4850113,1.6324836,1.7799559,2.0268862,2.287535,2.510458,2.6716487,2.5481834,2.335549,2.1091962,2.0303159,2.335549,2.2360911,2.1194851,2.1023371,2.2292318,2.4727325,2.7642474,2.7573884,2.784825,2.784825,2.2566686,2.270387,2.3664153,2.5790498,2.867135,3.0969174,2.9631636,2.719663,2.585909,2.6373527,2.8088322,2.4795918,2.2395205,2.0097382,1.728512,1.371835,1.4472859,1.529596,1.7593783,1.9514352,1.587899,1.6359133,1.8759843,2.3767042,2.8808534,2.8088322,2.7951138,3.0866287,3.3644254,3.789694,4.972902,6.4133286,7.2604365,7.997798,8.464222,7.8434668,8.769455,9.424506,10.0041065,10.751757,11.948683,13.118172,13.392539,13.114742,12.5145645,11.732618,10.80663,9.640571,9.373062,10.065839,10.710602,10.652299,10.81006,11.712041,13.169616,14.267084,13.999576,13.344524,13.125031,13.200482,12.466551,12.295071,11.190743,10.422516,10.991828,13.642899,15.093615,15.062748,14.726648,14.486577,13.96185,13.642899,14.150477,15.114192,16.108772,16.6335,17.473747,16.87014,15.501736,14.1299,13.581166,14.105893,14.13676,14.647768,16.191082,18.890167,20.073376,21.349182,22.117409,22.333473,22.491234,22.820475,22.20658,21.397196,20.53294,19.164536,18.578075,18.807858,18.03277,16.280252,15.426285,15.999025,16.520323,16.842705,16.702091,15.700651,13.920695,13.80409,14.517444,15.172495,14.832966,14.928994,15.604623,16.280252,16.599203,16.403717,17.63494,18.338005,18.61923,18.862732,19.730417,19.754423,19.109661,18.214539,17.494326,17.394867,18.115082,18.248835,17.840714,16.96617,15.731518,15.22051,15.440002,15.333686,14.627191,13.807519,13.029003,12.1921835,12.428825,13.533153,13.9481325,13.982429,14.990726,15.837835,16.167076,16.386568,16.414005,16.060759,15.885849,15.806969,15.138199,14.500296,14.363112,14.63062,15.193072,15.913286,16.184223,16.479168,17.034761,17.737827,18.1288,18.04306,18.653526,19.5315,20.104242,19.654966,20.347742,19.973917,18.900457,17.700102,17.151367,16.588915,16.026463,15.179354,14.5414505,15.395418,16.578627,17.278261,17.418875,16.96274,15.899568,14.959861,14.339106,13.540011,12.696333,12.572867,13.001566,13.025573,12.4802685,11.746337,11.732618,11.818358,12.243628,12.758065,13.13532,13.183334,13.841815,14.30138,14.445422,14.651197,15.762384,15.285671,14.819247,14.71636,15.079896,15.762384,16.811838,16.050468,15.309678,15.37827,15.9750185,17.12393,16.832415,15.88242,15.066177,15.21365,14.7369375,14.7197895,14.973578,15.580616,16.877,17.717249,17.62808,17.54234,17.398296,16.12935,15.604623,14.198492,13.169616,12.922686,13.032433,13.80066,13.845244,12.178465,10.429376,12.833516,9.853205,8.423067,9.925226,12.456262,10.834066,18.097933,20.361462,17.988186,12.500846,6.591667,4.1155047,2.9631636,5.844017,9.537683,4.897451,3.4467354,2.760818,2.3835633,1.9857311,1.3889829,1.4369972,8.755736,14.352823,15.021593,13.337666,9.15014,9.431366,7.7097125,4.5030484,7.3084507,6.2727156,8.666568,9.033533,7.160979,8.100685,9.688584,10.278474,10.593996,10.583707,9.400499,9.568549,8.889491,8.309891,8.519095,9.932085,10.679735,11.423956,10.751757,9.668007,11.595435,7.006647,5.90575,6.101236,7.0478024,9.8429165,14.249936,14.29795,11.784062,8.385342,5.675967,8.704293,9.067829,8.663138,8.155559,6.958633,5.079219,4.7088237,4.4413157,3.391862,1.2072148,1.8759843,1.7799559,2.4624438,3.8377085,4.180667,3.3747141,2.8808534,3.100347,3.2272418,1.2346514,1.0528834,0.9431366,0.6859175,0.29494452,0.01371835,0.01371835,0.01371835,0.058302987,0.14747226,0.24350071,0.31895164,0.66533995,0.8848336,0.89169276,0.91569984,0.70649505,0.5453044,0.41840968,0.31895164,0.26064864,0.31895164,0.28122616,0.29837412,0.39097297,0.42869842,0.61046654,0.764798,0.90541106,0.9602845,0.77851635,0.9842916,1.2209331,1.4472859,1.605047,1.6187652,1.4815818,1.2586586,1.3066728,1.5604624,1.5090185,1.1797781,0.9877212,0.939707,1.1008976,1.6016173,1.5638919,1.4369972,1.2483698,1.1214751,1.2826657,1.1729189,0.89855194,0.66533995,0.53501564,0.4115505,0.31552204,0.37382504,0.50757897,0.5727411,0.36696586,0.30523327,0.47328308,0.8265306,1.1763484,1.1900668,0.90884066,0.8676856,1.097468,1.4781522,1.7079345,1.6976458,2.177788,2.6064866,3.0283258,4.0880685,3.8445675,3.7211025,5.5319247,8.179566,7.630832,10.069269,10.233889,9.067829,7.14726,4.6676683,8.8929205,11.753197,10.048691,5.284994,3.6627994,2.503599,5.079219,5.3158607,3.1792276,4.671098,2.534465,1.9274281,4.90431,9.071259,7.582818,7.7542973,11.698323,11.739478,7.6342616,6.560801,5.4736214,4.0846386,3.566771,3.4124396,1.4335675,1.1523414,1.3958421,2.194936,2.74367,1.3889829,6.258997,10.278474,9.349055,5.209543,5.4153185,5.8817425,4.7431192,3.1860867,3.2958336,8.056101,5.2472687,2.3492675,0.89855194,1.1832076,2.2566686,3.5290456,2.819121,1.903421,1.5570327,1.5570327,1.2517995,1.2929544,1.5570327,2.061182,2.976882,3.8788633,3.9680326,4.1943855,4.180667,2.2292318,2.959734,3.316411,3.2683969,2.952875,2.6853669,2.4658735,3.0043187,3.3301294,3.3438478,3.8445675,3.7965534,3.7759757,3.841138,3.8788633,3.5873485,4.012617,4.1120753,4.0674906,3.8960114,3.433017,3.3472774,3.3644254,3.2958336,2.9631636,2.1812177,1.5090185,1.4541451,1.786815,2.4418662,3.4776018,3.782835,4.197815,4.8837323,5.381023,4.623084,2.877424,2.534465,2.9048605,3.3712845,3.3712845,3.8960114,4.2115335,4.187526,4.0194764,4.2252517,4.029765,3.9268777,4.0194764,4.0709205,3.508468,3.4124396,3.4981792,3.8377085,4.3692946,4.8837323,3.8685746,4.338428,4.914599,4.976331,4.6848164,4.122364,3.4707425,2.884283,2.651071,3.1895163,3.3472774,3.4981792,3.6010668,3.7382503,4.105216,4.091498,3.806842,3.1826572,2.3046827,1.3889829,0.7407909,0.58988905,0.65162164,0.6893471,0.5178677,0.45613512,0.53501564,0.58988905,0.6756287,1.0528834,0.9911508,0.8676856,0.78194594,0.91569984,1.5261664,2.7711067,3.5873485,4.1292233,4.290414,3.6936657,3.216953,2.9322972,2.5961976,2.318401,2.5619018,2.6613598,2.702515,3.4844608,4.7979927,5.4324665,5.4084597,4.715683,3.9714622,3.450165,3.083199,2.8739944,2.702515,2.8088322,3.192946,3.6319332,3.532475,3.6559403,4.1326528,4.822,5.3090014,5.0414934,4.7534084,4.6882463,4.804852,4.804852,5.0757895,4.557922,4.7808447,5.6999745,5.675967,6.334448,6.252138,6.2830043,6.6636887,7.0203657,6.3961806,5.5902276,4.8082814,4.266407,4.180667,4.6573796,5.1238036,5.6656785,6.3790326,7.3530354,7.490219,6.5059276,5.0414934,3.6696587,2.8980014,3.3884325,3.4810312,3.3781435,3.2683969,3.340418,3.3301294,2.8225505,2.2360911,1.8313997,1.7079345,1.5364552,1.1832076,0.8711152,0.71678376,0.71678376,0.90198153,0.9568549,0.9362774,0.9568549,1.1900668,1.0185875,0.7373613,0.7922347,1.1283343,1.1900668,0.86082643,0.7888051,0.89169276,1.0494537,1.097468,1.2586586,1.8108221,2.1400626,2.177788,2.411,1.3478279,1.138623,1.2483698,1.4507155,1.8142518,1.5604624,1.6770682,2.201795,2.9974594,3.7519686,4.57164,4.372724,3.5804894,3.2272418,4.972902,5.610805,5.9880595,6.018926,6.0566516,6.910619,7.9737906,7.5519514,7.9189177,9.002667,8.3922,0.9568549,1.2277923,1.4438564,1.488441,1.371835,1.2517995,1.2037852,1.1626302,1.2072148,1.3649758,1.6221949,1.7971039,2.1915064,2.4898806,2.6064866,2.6579304,2.527606,2.3389788,2.2566686,2.335549,2.5413244,2.4555845,2.3252604,2.2498093,2.2258022,2.1674993,2.253239,2.1194851,1.9274281,1.8039631,1.8554068,1.8176813,1.8725548,2.0063086,2.194936,2.3767042,2.4590142,2.3561265,2.3389788,2.428148,2.4041407,2.0165975,1.9239986,1.6873571,1.3066728,1.214074,1.2963841,1.4987297,1.8039631,2.095478,2.16064,2.1812177,2.2155135,2.3732746,2.551613,2.428148,2.4555845,3.3987212,4.297273,5.0003386,6.193835,7.888051,8.81404,8.995808,8.752307,8.683716,9.253027,9.325048,9.688584,10.669447,12.120162,12.576297,12.696333,12.531713,12.339656,12.562579,11.705182,10.525404,10.364213,11.249047,11.897239,11.921246,11.825217,11.921246,12.411677,13.365103,13.38911,13.708061,14.640909,15.512024,14.651197,13.035862,12.329367,12.041282,12.233338,13.543441,13.893259,13.951562,13.728639,13.594885,14.291091,15.028452,15.22051,16.009314,17.267973,17.607502,18.20768,18.684393,18.44432,17.446312,16.204802,15.909856,15.985307,16.506605,17.182234,17.339994,17.401728,17.919594,19.13024,20.78673,22.175713,21.849901,21.630407,21.599543,21.390337,20.179693,19.562366,19.147387,18.87645,18.667244,18.430603,18.77699,19.13024,18.674105,17.600643,17.117071,15.656067,14.757515,14.688923,15.22051,15.611482,15.6697855,15.031882,14.685493,14.856973,15.0250225,15.9921665,16.945591,17.532051,17.799559,18.180243,18.437462,18.327715,17.744686,16.925014,16.45516,16.636929,16.739817,16.732958,16.54776,16.084764,15.066177,14.760944,14.273943,13.38225,12.562579,12.260776,12.212761,12.452832,12.88839,13.262215,13.37882,13.817808,14.404267,14.932424,15.193072,15.909856,16.427725,16.362562,15.9921665,16.245956,16.160215,15.724659,15.700651,16.225378,16.818697,16.938732,16.393429,16.62321,17.806417,18.8593,18.910746,18.639809,18.595222,18.831865,18.907316,19.03764,18.900457,18.547209,17.95732,17.079346,16.729528,16.143068,15.275383,14.496866,14.589465,15.326826,16.352274,17.408587,17.751545,16.143068,14.959861,14.46257,14.023583,13.505715,13.255356,12.950122,12.624311,12.295071,11.96926,11.622872,11.924676,12.833516,13.224489,12.871242,12.452832,13.450842,14.177915,14.565458,14.757515,15.127911,14.867262,14.400838,14.225929,14.531162,15.21365,17.315987,17.065628,16.12935,15.549749,15.769243,15.978448,16.252815,16.067617,15.553179,15.494876,14.706071,14.959861,15.7795315,16.79126,17.741257,17.28512,16.811838,16.852993,16.952452,15.666355,15.227368,14.232788,13.354814,13.001566,13.337666,13.118172,12.764925,11.653738,10.281903,10.244178,9.328478,11.595435,12.404818,11.609154,13.567448,22.333473,17.182234,10.593996,7.949784,7.5210853,4.016047,2.0097382,4.0434837,7.840037,6.276145,3.3198407,2.8705647,2.5207467,1.646202,1.3889829,1.6324836,8.580828,11.777204,10.432805,13.433694,9.89093,9.541112,8.659708,7.6857057,11.214751,8.947794,9.482809,9.410788,8.416207,9.287323,10.326488,8.779744,8.385342,9.170717,7.459353,8.371623,8.073249,7.431916,7.431916,9.201583,11.177026,13.584596,13.083877,10.034973,8.508806,6.125243,6.2144127,5.8405876,4.5167665,4.1772375,7.970361,8.436785,8.9100685,9.074688,4.9694724,6.0703697,6.81802,6.48535,5.1238036,3.5770597,3.6696587,4.2115335,4.2286816,3.3129816,1.5947582,3.2443898,3.0454736,2.8945718,3.4947495,4.3624353,4.9351764,4.537344,4.0434837,3.6387923,2.8122618,1.9137098,1.1420527,0.69963586,0.490431,0.09945804,0.05144381,0.024007112,0.09259886,0.1920569,0.13375391,0.17833854,0.6276145,0.805953,0.6001778,0.48700142,0.58302987,0.65848076,0.53844523,0.29151493,0.20920484,0.24350071,0.22292319,0.25721905,0.32581082,0.29151493,0.4355576,0.58988905,0.6756287,0.70649505,0.77851635,0.8779744,1.0563129,1.3272504,1.5707511,1.5433143,1.6942163,1.7422304,1.845118,2.0234566,2.170929,2.1915064,1.9685832,1.7319417,1.6256244,1.7353712,1.7182233,1.3821237,1.0528834,0.9328478,1.1111864,1.0700313,0.90541106,0.6893471,0.5007198,0.44927597,0.4081209,0.39440256,0.39783216,0.41840968,0.4629943,0.5212973,0.5624523,0.72707254,0.94656616,0.9568549,1.0494537,1.1729189,1.6084765,2.1812177,2.2566686,2.527606,3.0248961,3.2718265,3.316411,3.724532,2.8259802,2.7779658,3.3850029,4.3692946,5.3707337,4.7362604,3.7622573,3.350707,4.3452873,7.548522,5.552502,5.885172,5.6793966,4.3590055,3.625074,6.975781,6.6465406,5.2472687,4.8185706,6.8043017,2.9494452,2.170929,6.824879,11.880091,4.9214582,4.791134,5.545643,5.7136927,5.5593615,7.0752387,6.046363,5.813151,5.086078,3.450165,1.3855534,0.9294182,0.7099246,0.8745448,1.155771,0.8745448,1.8416885,6.742569,9.493098,8.1041155,4.7088237,4.341858,4.887162,4.537344,5.377593,13.38911,4.8905916,1.6530612,0.89855194,1.3649758,3.309552,3.4844608,2.503599,1.7971039,1.8554068,2.2292318,1.3066728,1.371835,1.4644338,1.7559488,3.5599117,4.729401,4.187526,3.957744,4.108646,2.7539587,2.6647894,2.5310357,2.3321195,2.2738166,2.7951138,2.194936,2.5310357,3.0146074,3.2581081,3.2581081,3.707384,3.4673128,3.2958336,3.4433057,3.6593697,4.105216,4.4584637,4.4584637,4.139512,3.82399,3.649081,3.3952916,3.0900583,2.7573884,2.4144297,1.9171394,1.7730967,2.0680413,2.6819375,3.2581081,3.7211025,3.9097297,4.32471,4.856296,4.7808447,1.9720128,2.1434922,3.2203827,3.9474552,3.9097297,4.122364,4.307562,4.554492,4.5819287,3.7142432,4.064061,4.0194764,3.9200184,3.8205605,3.474172,3.210094,3.2443898,3.7108135,4.437886,4.979761,4.962613,4.7602673,4.5819287,4.5510626,4.7088237,4.2046742,3.457024,2.9117198,2.6853669,2.5653315,2.901431,3.3369887,3.4844608,3.4913201,4.0434837,3.3952916,3.2512488,3.0866287,2.627064,1.8416885,1.0357354,0.6344737,0.5178677,0.5521636,0.5555932,0.4938606,0.5041494,0.5212973,0.5796003,0.8196714,0.8779744,0.7510797,0.6310441,0.6893471,1.0871792,2.0886188,2.7470996,3.275256,3.6765177,3.7519686,3.532475,3.0900583,2.6716487,2.4624438,2.5893385,2.568761,2.8808534,3.5942078,4.5613513,5.4187484,6.0497923,5.6656785,4.852866,4.0194764,3.3987212,2.7333813,2.6304936,2.8911421,3.3472774,3.875434,3.532475,3.6593697,4.064061,4.496189,4.664239,4.773986,4.7671266,4.605936,4.4927597,4.8425775,5.267846,5.1340923,5.353586,6.1629686,7.116394,7.805741,7.9429245,7.822889,7.699424,7.798882,6.8763227,5.7891436,4.9934793,4.633373,4.557922,5.31929,5.7239814,5.8234396,5.7479887,5.720552,6.060081,5.675967,5.0449233,4.3624353,3.5461934,3.5770597,3.549623,3.40901,3.2443898,3.2683969,3.316411,2.9254382,2.3252604,1.8108221,1.7593783,1.6736387,1.5981878,1.4678634,1.2312219,0.8505377,0.9842916,1.0666018,1.0220171,0.9602845,1.1523414,1.1694894,1.0494537,1.0666018,1.2449403,1.371835,1.0631721,0.83338976,0.7579388,0.8505377,1.0871792,1.2175035,1.5707511,1.9239986,2.194936,2.4487255,2.2635276,1.9582944,1.7010754,1.6976458,2.170929,2.2635276,2.3904223,2.651071,3.1483612,3.974892,3.7382503,3.9851806,3.642222,3.07634,4.108646,6.2967224,7.3701835,7.1266828,6.1766872,5.9469047,6.667118,7.531374,8.80718,10.031544,10.014396,0.94656616,1.0768905,1.2175035,1.3203912,1.3341095,1.2209331,1.1489118,1.0597426,1.0871792,1.2655178,1.5158776,1.786815,2.0817597,2.3321195,2.4452958,2.2806756,2.335549,2.435007,2.4315774,2.386993,2.5481834,2.2738166,2.2429502,2.1743584,1.9823016,1.7525192,2.0440342,1.9994495,1.786815,1.6084765,1.7010754,1.6804979,1.8005334,1.9445761,1.9823016,1.786815,1.862266,1.8999915,2.0028791,2.1332035,2.1126258,2.0234566,1.8931323,1.6633499,1.4610043,1.605047,1.6976458,1.903421,2.1194851,2.2806756,2.386993,2.3561265,2.4830213,2.534465,2.452155,2.3629858,2.3904223,3.1689389,4.125794,5.1580997,6.619104,8.567109,9.030104,9.006097,8.961512,8.81404,9.098696,9.163857,9.438225,10.2236,11.694893,12.267634,12.397959,12.157887,11.941824,12.459691,12.065289,11.375941,11.008976,11.22161,11.89038,11.7257595,11.787492,12.144169,12.555719,12.46998,12.778643,13.533153,14.260224,14.428274,13.450842,12.679185,13.087306,13.481709,13.529722,13.738928,14.030442,14.027013,13.951562,14.013294,14.390549,16.19794,17.830425,19.161106,19.823015,19.215979,18.728977,18.62266,18.756414,18.674105,17.593784,16.287111,15.9750185,16.283682,16.911295,17.63151,17.71039,17.70696,17.929884,18.183672,17.7927,18.022482,19.017063,20.155685,20.827885,20.430052,19.243416,18.866161,19.03764,19.342873,19.236557,19.12681,19.408035,19.322296,18.660385,17.765263,16.774113,15.776102,15.289101,15.5085945,16.300829,16.235666,15.340545,14.472859,13.992717,13.783512,14.613472,15.391989,16.012743,16.45173,16.767254,16.45516,16.184223,15.964729,15.745236,15.395418,15.738377,16.256245,16.365992,16.098484,16.091625,15.851553,15.433144,14.445422,12.956982,11.465111,11.091286,11.372512,11.784062,12.154458,12.651748,12.55915,12.593445,13.029003,13.817808,14.599753,15.182784,15.54632,15.724659,15.865272,16.21509,16.818697,16.280252,15.680074,15.676644,16.486027,17.267973,16.969599,16.955881,17.600643,18.30028,18.739265,18.608942,18.197392,17.7927,17.717249,17.61436,17.648657,17.837284,17.933313,17.408587,17.017612,16.328266,15.529172,14.953001,15.076467,15.193072,15.597764,16.554619,17.439453,16.726099,15.597764,14.699212,14.099034,13.660047,13.042721,12.562579,12.466551,12.360233,12.05843,11.578287,12.13731,13.001566,13.395968,13.234778,13.090735,13.526293,13.985858,14.376831,14.620332,14.658057,15.100473,14.932424,14.651197,14.688923,15.422854,16.743246,16.832415,16.414005,15.964729,15.697222,15.285671,15.278812,15.141628,14.839825,14.832966,13.831526,14.393978,15.196502,15.830976,16.770683,16.558048,16.671225,16.736387,16.345413,15.035312,14.4317045,13.282792,12.538571,12.55229,13.073587,13.056439,13.13532,12.315649,10.8958,10.477389,10.432805,10.827208,11.070708,12.922686,20.505503,20.155685,11.612583,6.636252,6.9209075,4.0880685,2.6579304,1.4918705,6.90033,13.958421,6.495639,5.9228973,4.856296,3.4295874,2.0440342,1.3615463,8.025234,10.38479,8.961512,6.9723516,10.319629,9.462232,9.208443,9.105555,8.676856,7.421627,5.658819,8.224151,10.196163,10.203023,10.398509,9.184435,7.140401,6.4544835,6.917478,5.90232,7.449064,7.2535777,7.0375133,7.7440085,9.541112,11.214751,12.30193,11.921246,10.172156,8.131552,6.2830043,5.686256,5.2164025,4.3658648,3.2649672,4.4859004,4.1772375,4.804852,5.785714,3.4913201,3.6079261,4.331569,4.2835546,3.4878905,3.3438478,3.0146074,3.4192986,4.170378,4.2835546,2.177788,4.012617,3.765687,3.1037767,3.0146074,3.7862647,4.8185706,4.557922,4.2869844,4.386442,4.3041325,3.4055803,1.9720128,0.9328478,0.4938606,0.15776102,0.12003556,0.08573969,0.10288762,0.15090185,0.13375391,0.14061308,0.3806842,0.5555932,0.5453044,0.39097297,0.5761707,0.8848336,0.91912943,0.59674823,0.15090185,0.20577525,0.22978236,0.28465575,0.36010668,0.37039545,0.4081209,0.61389613,0.84024894,0.9877212,0.9877212,0.9602845,1.0048691,1.2346514,1.5536032,1.6633499,2.1229146,2.270387,2.3286898,2.4555845,2.7368107,2.884283,2.5207467,2.0920484,1.8691251,1.9514352,2.1160555,1.8485477,1.5570327,1.4198492,1.3992717,1.3306799,1.1283343,0.84024894,0.5590228,0.44927597,0.45956472,0.4081209,0.40126175,0.4698535,0.5796003,0.5555932,0.5555932,0.7442205,0.9842916,0.8265306,1.0528834,1.2998136,1.7147937,2.1846473,2.3218307,2.8122618,3.2718265,3.3026927,3.1655092,3.806842,3.4673128,3.4673128,3.4535947,3.4776018,3.99204,3.234101,2.9151495,2.7916842,2.9288676,3.7039545,4.698535,6.8626046,8.508806,8.536243,6.427047,9.184435,7.4284863,4.979761,5.0414934,10.179015,5.284994,4.650521,9.338767,13.481709,4.2835546,5.360445,6.5985265,6.1046658,4.8940215,6.910619,4.605936,5.3432975,5.4187484,3.765687,1.9514352,0.89855194,0.5796003,1.0700313,2.510458,5.1066556,2.6407824,6.111525,9.619993,9.39707,3.8274195,6.725421,7.1061053,6.0978065,5.504488,7.8126,3.1312134,1.5604624,1.5844694,2.4247184,4.0366244,3.4913201,2.7539587,2.1091962,1.8588364,2.3218307,2.0028791,1.9685832,1.978872,2.1915064,3.175798,4.6436615,4.4447455,4.098357,3.923448,3.0214665,2.6990852,2.3904223,2.0337453,1.8348293,2.2841053,2.0474637,2.1469216,2.6304936,3.192946,3.1689389,3.6765177,3.357566,3.0283258,3.07634,3.4844608,3.841138,4.57164,5.0483527,4.955754,4.32471,4.149801,3.8891523,3.4913201,3.07634,2.9117198,2.4658735,2.1126258,2.2223728,2.6716487,2.867135,3.2992632,3.4295874,3.6182148,3.9954693,4.437886,2.1812177,2.170929,2.9631636,3.6525106,3.8960114,4.3178506,4.266407,4.2218223,4.091498,3.2203827,3.7382503,4.0194764,3.9268777,3.5359046,3.1243541,3.0317552,3.2512488,3.6319332,4.0091877,4.2081037,4.3590055,4.3624353,4.214963,4.081209,4.2835546,3.9131594,3.3232703,2.7402403,2.2738166,1.9239986,2.3321195,3.3301294,3.7931237,3.5599117,3.4227283,3.1380725,3.0111778,2.877424,2.603057,2.0817597,1.3786942,0.8471081,0.548734,0.48357183,0.59331864,0.65505123,0.5658819,0.51100856,0.5693115,0.6790583,0.8093826,0.7133542,0.65505123,0.7922347,1.1763484,1.7388009,2.3286898,2.74367,3.0214665,3.457024,3.4535947,3.1723683,2.9117198,2.7642474,2.620205,3.07634,3.5873485,4.214963,4.9831905,5.8474464,6.077229,6.1149545,5.693115,4.9077396,4.201245,3.5153272,3.0420442,2.9494452,3.2889743,3.99204,3.8960114,3.875434,4.046913,4.32471,4.4104495,4.273266,4.4721823,4.413879,4.184097,4.557922,4.804852,5.1992545,5.6828265,6.279575,7.1026754,8.045813,8.217292,8.169277,8.086967,7.795452,6.9689217,5.857735,5.130663,4.911169,4.773986,5.3981705,5.7308407,5.7891436,5.6313825,5.3741636,5.435896,5.24041,5.1238036,5.003768,4.3933015,3.8171308,4.0434837,4.3487167,4.4721823,4.633373,4.773986,3.6044965,2.4315774,1.862266,1.786815,1.9239986,1.9857311,1.8519772,1.5193073,1.0940384,1.0288762,1.0220171,0.9842916,0.9328478,0.99801,1.08032,1.1077567,1.2037852,1.4267083,1.7936742,1.5330256,1.3238207,1.155771,1.0494537,1.0734608,1.138623,1.4815818,1.8828435,2.1915064,2.3458378,2.287535,2.2360911,2.1229146,2.085189,2.469303,2.7093742,2.935727,3.210094,3.5770597,4.046913,3.82399,4.1120753,4.187526,4.0880685,4.6127954,6.2384195,7.4181976,7.534804,6.8385973,6.447624,6.8626046,7.963502,9.119273,9.836057,9.770895,0.8471081,0.85739684,0.922559,1.0357354,1.1489118,1.1351935,1.08032,0.9945804,1.0357354,1.2175035,1.3992717,1.7147937,1.8828435,2.0920484,2.270387,2.07833,2.1572106,2.386993,2.4555845,2.3561265,2.3904223,2.054323,1.9685832,1.9171394,1.7799559,1.5433143,1.7971039,1.8039631,1.6290541,1.4164196,1.4061309,1.4164196,1.4815818,1.5638919,1.5707511,1.3649758,1.5673214,1.728512,1.8519772,1.9480057,2.0440342,2.201795,2.201795,2.0714707,1.9651536,2.1674993,2.2052248,2.3595562,2.527606,2.651071,2.702515,2.5790498,2.5378947,2.4658735,2.4315774,2.6716487,2.8499873,3.223812,3.923448,5.120374,7.010077,8.460793,8.477941,8.573969,9.023245,8.868914,8.440215,8.539673,8.985519,9.788043,11.163307,12.092726,12.449403,12.312219,12.068718,12.418536,12.233338,11.674315,11.115293,10.950673,11.595435,11.125582,11.166737,11.509696,11.664027,10.858074,11.838936,12.4802685,12.634601,12.394529,12.089295,12.3533745,13.279363,14.009865,14.321958,14.616901,15.076467,14.671775,14.291091,14.147048,13.783512,15.806969,18.276272,20.052797,20.61525,20.045938,19.387459,18.687822,18.420315,18.389448,17.744686,16.904436,16.87357,17.051908,17.312557,18.025911,18.838724,18.492336,17.734396,16.729528,15.062748,15.868701,16.877,18.03277,19.219408,20.248285,19.60695,19.46291,19.757853,20.251715,20.512363,20.234566,20.19341,20.011642,19.480057,18.574646,17.682953,16.558048,15.858413,15.79325,16.108772,16.033321,15.326826,14.555169,13.924125,13.282792,13.910407,14.582606,15.22051,15.721229,15.940722,15.512024,15.193072,14.96672,14.743796,14.369971,14.781522,15.885849,16.362562,16.04018,15.913286,15.875561,15.649208,14.805529,13.227919,11.087856,10.511685,10.5597,10.97468,11.574858,12.250486,12.068718,11.838936,12.0309925,12.788932,13.917266,14.167625,14.359683,14.644339,15.073037,15.590904,16.434584,16.245956,15.6697855,15.405707,16.187653,17.364002,17.761833,17.833855,17.861292,17.940172,18.338005,18.217968,17.71382,17.04505,16.53747,16.45173,16.352274,16.654078,17.182234,17.182234,16.993607,16.321407,15.573756,15.103903,15.193072,15.302819,15.230798,15.539461,16.064188,15.927004,14.939283,13.80066,13.128461,12.908967,12.476839,12.034423,12.21619,12.404818,12.274493,11.790922,12.336226,12.895248,13.320518,13.63604,14.057879,14.177915,14.428274,14.616901,14.634049,14.448852,15.4742985,15.62863,15.5085945,15.614912,16.328266,16.582056,16.763824,16.760393,16.486027,15.892709,15.121051,14.637479,14.102464,13.642899,13.862392,13.491997,14.147048,14.606613,14.788382,15.738377,15.748666,16.033321,15.782962,14.990726,14.46257,14.009865,13.104454,12.713481,12.891819,12.775213,12.542002,12.459691,11.880091,11.019264,10.940384,10.192734,9.671436,11.393089,15.776102,21.633839,14.13333,7.6445503,5.48734,6.090947,2.9974594,2.6990852,5.8234396,11.818358,15.484588,6.992929,8.1384115,5.689686,4.6127954,5.8371577,6.279575,10.583707,11.14273,9.3079,7.164408,7.5279446,8.162418,7.9943686,7.716572,7.1369715,5.144381,4.5990767,9.283894,12.202472,11.4754,10.319629,7.870903,6.276145,5.5079174,5.178677,4.557922,6.4373355,6.23156,6.5333643,8.045813,9.589127,10.607714,10.268185,9.897789,9.846346,9.458802,6.4579134,4.887162,4.1429415,3.6010668,2.620205,3.6765177,2.5481834,2.3595562,3.3815732,3.0454736,2.5378947,2.9734523,3.0489032,2.8465576,3.8342788,3.210094,3.649081,4.4996185,4.698535,2.7573884,3.923448,3.9131594,3.5461934,3.3987212,3.806842,4.7259717,4.4756117,4.431027,4.8597255,4.914599,4.3624353,3.0214665,1.6530612,0.6962063,0.274367,0.17147937,0.13375391,0.12689474,0.1371835,0.15090185,0.15433143,0.20920484,0.33952916,0.47671264,0.4389872,0.4938606,0.980862,1.1729189,0.82996017,0.20234565,0.25378948,0.2503599,0.28122616,0.3566771,0.4115505,0.42526886,0.7442205,1.097468,1.2998136,1.2312219,1.2037852,1.2346514,1.430138,1.7490896,1.9994495,2.627064,2.8396983,2.8396983,2.8294096,3.0043187,3.1346428,2.7745364,2.3835633,2.2258022,2.3492675,2.551613,2.3424082,2.095478,1.9411465,1.7765263,1.6770682,1.4164196,1.0528834,0.69963586,0.5212973,0.5144381,0.51100856,0.5555932,0.64476246,0.7442205,0.6379033,0.61389613,0.85739684,1.2037852,1.1489118,1.3203912,1.4850113,1.7113642,1.9720128,2.1503513,2.702515,3.1963756,3.2375305,3.0660512,3.542764,3.899441,4.262977,4.2698364,3.9680326,3.8342788,3.3369887,3.4638834,3.4021509,2.7951138,1.7353712,3.7485392,7.2124224,10.415657,11.214751,7.051232,8.659708,8.110974,5.65539,4.1772375,9.177576,7.9120584,8.080108,10.281903,11.492548,5.0826488,7.1266828,8.207003,7.1541195,5.521636,7.5931067,4.0057583,4.331569,4.756838,3.7862647,2.2600982,1.2312219,1.0700313,1.7456601,3.6113555,7.407909,4.197815,5.871454,9.901219,11.434244,3.2889743,8.100685,7.239859,5.6039457,4.746549,2.8877127,2.5961976,1.8108221,1.6770682,2.6167753,4.3007026,3.457024,2.9391565,2.49331,2.1640697,2.2669573,2.3629858,2.3561265,2.49331,2.726522,2.726522,3.8205605,4.122364,3.882293,3.3712845,2.8808534,2.568761,2.2052248,1.8176813,1.5433143,1.6290541,2.0303159,2.1057668,2.4830213,3.0797696,3.100347,3.40901,3.2409601,3.0386145,3.0351849,3.2546785,3.6285036,4.6916757,5.6793966,6.0669403,5.579939,4.9934793,4.448175,3.9131594,3.4604537,3.2581081,2.9460156,2.3595562,2.1983654,2.5824795,3.0489032,3.1620796,3.2683969,3.3369887,3.4878905,3.998899,2.8945718,2.6133456,2.884283,3.391862,3.7862647,4.383013,4.1155047,3.7451096,3.5359046,3.2683969,3.789694,4.033195,3.940596,3.5804894,3.1380725,3.0043187,3.3301294,3.7142432,3.8960114,3.7519686,3.666229,3.858286,3.9646032,3.923448,3.9611735,3.7553983,3.4878905,2.9254382,2.218943,1.8691251,1.9514352,2.9460156,3.7862647,3.8960114,3.216953,2.9151495,2.74367,2.5996273,2.4007113,2.0646117,1.5021594,1.0666018,0.75450927,0.5796003,0.6036074,0.7613684,0.66191036,0.5761707,0.59674823,0.6241849,0.7442205,0.70306545,0.66876954,0.7613684,1.08032,1.4164196,2.1400626,2.568761,2.668219,3.0420442,3.4673128,3.316411,3.1243541,3.0454736,2.8396983,3.4535947,4.2218223,4.9694724,5.641671,6.293293,6.200694,6.5024977,6.509357,6.025785,5.3330083,4.5956473,3.8925817,3.5050385,3.5530527,3.974892,4.2355404,4.173808,4.1360826,4.2252517,4.3007026,4.105216,4.417309,4.3624353,3.9886103,4.2835546,4.5099077,5.312431,5.826869,6.0326443,6.776865,7.805741,7.9772205,8.018375,8.032094,7.500508,6.9071894,6.1972647,5.7411294,5.535354,5.212973,5.470192,5.768566,5.8817425,5.744559,5.442755,5.6142344,5.425607,5.346727,5.3913116,5.1340923,4.465323,4.629943,4.962613,5.2266912,5.645101,6.0326443,4.3281393,2.644212,1.8931323,1.8313997,2.0131679,2.1229146,2.020027,1.7147937,1.3512574,1.2346514,1.1146159,1.0048691,0.939707,0.9602845,1.0117283,1.1180456,1.3272504,1.6427724,2.037175,2.0474637,1.7902447,1.5090185,1.3546871,1.4027013,1.3101025,1.4953002,1.9171394,2.3595562,2.4452958,2.1812177,2.0474637,2.0063086,2.0714707,2.3218307,2.7951138,3.234101,3.5290456,3.6799474,3.7965534,4.033195,4.2252517,4.280125,4.448175,5.3330083,6.012067,6.931196,7.39762,7.4113383,7.682276,7.3393173,7.9257765,8.766026,9.537683,10.285333,0.7099246,0.78537554,0.8676856,0.9294182,0.97400284,1.0425946,1.0220171,0.9945804,1.08032,1.255229,1.3478279,1.6084765,1.7079345,1.903421,2.153781,2.1229146,1.99602,2.1057668,2.201795,2.1846473,2.0989075,1.8176813,1.611906,1.5776103,1.6324836,1.5227368,1.430138,1.3375391,1.1626302,0.96371406,0.9259886,0.9431366,0.881404,0.8711152,0.9602845,1.1146159,1.5055889,1.7388009,1.8176813,1.8656956,2.085189,2.311542,2.5927682,2.6853669,2.609916,2.668219,2.6304936,2.7985435,3.0214665,3.1826572,3.1860867,2.9700227,2.551613,2.352697,2.603057,3.333559,3.690236,3.9371665,4.355576,5.336438,7.3701835,7.805741,7.699424,8.107545,8.944365,8.98209,7.936065,8.097256,8.7283,9.510246,10.515115,11.55771,12.236768,12.507706,12.483699,12.415107,12.380811,11.732618,11.1393,10.981539,11.358793,10.600855,10.336777,10.206452,9.908078,9.239308,10.600855,10.803201,10.679735,10.820349,11.5645685,12.274493,13.035862,13.831526,14.760944,16.026463,16.2974,15.529172,14.7026415,14.088745,13.258785,14.832966,16.732958,18.307138,19.19197,19.28457,19.339443,18.852442,18.149376,17.562918,17.422304,18.001905,18.770132,19.11652,18.900457,18.437462,19.562366,18.921034,17.861292,16.846134,15.446862,16.20137,16.101913,16.20137,17.161655,19.250275,20.443771,20.78673,20.937632,21.273731,21.894485,21.921923,21.606401,20.827885,19.853882,19.318867,18.348293,16.997036,16.149927,15.834405,15.21365,15.282242,14.778092,14.263655,13.845244,13.173045,13.526293,14.116182,14.791811,15.343974,15.5085945,15.522313,15.45715,15.004445,14.21564,13.505715,13.622321,14.88098,15.865272,16.029892,15.704081,15.049029,15.018164,14.784951,13.783512,11.684605,10.909517,10.347065,10.405369,11.026124,11.705182,11.64345,11.413667,11.379372,11.828648,12.956982,13.049581,13.399398,13.660047,13.924125,14.7369375,15.46058,16.009314,16.156786,16.091625,16.410576,17.312557,18.190533,18.451181,18.118511,17.826996,17.916164,17.532051,17.021042,16.438013,15.584045,15.560039,15.1862135,15.261664,15.803539,16.050468,16.2974,15.861842,15.217079,14.664916,14.363112,14.922135,14.898128,14.579176,14.174485,13.838386,12.878101,11.869802,11.369082,11.430815,11.612583,11.393089,11.691463,12.109874,12.325937,12.082437,12.346515,12.596875,13.039291,13.732068,14.616901,15.114192,15.522313,15.577187,15.258235,14.808959,15.851553,16.204802,16.46888,16.928444,17.573206,17.37772,17.470318,17.432592,17.089634,16.520323,15.789821,15.049029,14.099034,13.289652,13.522863,14.243076,14.634049,14.743796,14.887839,15.638919,15.37827,15.158776,14.441993,13.673765,14.29795,13.920695,13.601744,13.591455,13.443983,12.024134,11.622872,10.81006,10.456812,10.64201,10.676306,8.759167,9.767465,13.272504,16.588915,14.774663,8.186425,6.6568294,5.878313,4.629943,4.7499785,5.703404,14.503725,16.523752,10.377932,7.8777623,12.624311,8.498518,7.0478024,10.834066,13.419975,8.193284,11.55771,12.744347,9.218731,6.694555,7.208993,6.6293926,5.6656785,5.353586,7.034084,8.05953,12.164746,13.605173,11.314209,8.889491,6.7700057,5.9571934,5.3707337,4.5853586,3.8205605,5.5387836,5.3913116,6.0737996,7.9086285,8.858624,9.774324,9.386781,8.738589,8.937505,11.159878,6.3447366,4.6848164,3.690236,2.4727325,1.7593783,3.8720043,3.0248961,2.719663,3.6627994,3.799983,2.8705647,3.1655092,3.2272418,3.0660512,4.184097,3.8342788,4.5990767,4.931747,4.2766957,3.0729103,3.316411,3.6936657,4.108646,4.386442,4.2869844,4.914599,4.629943,4.4927597,4.65395,4.355576,4.180667,3.799983,2.7813954,1.3581166,0.4389872,0.216064,0.16119061,0.17147937,0.17490897,0.14747226,0.18176813,0.20234565,0.2469303,0.34981793,0.53844523,0.36353627,0.9362774,1.196926,0.86082643,0.41498008,0.36696586,0.29151493,0.274367,0.32238123,0.36696586,0.47328308,0.8676856,1.2037852,1.3752645,1.4987297,1.605047,1.821111,2.07833,2.3492675,2.644212,3.1963756,3.4673128,3.4192986,3.2032347,3.1312134,3.175798,2.9220085,2.7230926,2.7162333,2.836269,2.9322972,2.7093742,2.4624438,2.311542,2.177788,2.0577524,1.7799559,1.3821237,0.980862,0.78194594,0.64819205,0.72364295,0.84024894,0.9259886,1.0220171,0.8848336,0.7956643,1.0117283,1.4610043,1.7593783,1.7799559,1.7319417,1.7353712,1.845118,2.037175,2.568761,3.1449318,3.3952916,3.309552,3.216953,3.8137012,4.616225,4.976331,4.7842746,4.496189,3.5976372,3.4124396,3.3472774,3.216953,3.2375305,2.5207467,4.623084,8.045813,9.729739,5.0620713,6.3653145,8.460793,7.425057,4.355576,5.3570156,9.400499,10.089847,9.537683,8.327039,5.5250654,8.580828,8.676856,7.2535777,6.341307,8.539673,4.7774153,4.2218223,4.1189346,3.2718265,2.054323,1.879414,1.8416885,2.1983654,3.5290456,6.7459984,4.7534084,5.778855,10.295622,13.272504,4.149801,7.846896,5.439326,3.8788633,4.338428,2.2120838,2.9734523,2.0474637,1.4232788,2.1263442,4.2115335,3.5221863,3.0214665,2.7985435,2.6853669,2.2600982,2.1332035,2.3835633,2.877424,3.1895163,2.6064866,2.836269,3.2443898,3.1860867,2.6785078,2.411,2.2292318,1.9102802,1.6736387,1.5021594,1.1317638,1.8656956,2.2738166,2.7539587,3.2032347,3.000889,3.0729103,3.1689389,3.2512488,3.2649672,3.1277838,3.5702004,4.804852,6.0703697,6.869464,6.9517736,5.744559,4.8254294,4.1635194,3.7005248,3.3232703,3.3541365,2.603057,2.1469216,2.5001693,3.6044965,3.4364467,3.590778,3.625074,3.5290456,3.7005248,3.642222,3.2683969,3.1792276,3.457024,3.6936657,4.32471,3.9954693,3.4947495,3.309552,3.625074,3.9611735,3.923448,3.858286,3.7862647,3.4124396,3.1380725,3.340418,3.7313912,3.9783216,3.7039545,3.3644254,3.4295874,3.6970954,3.9165888,3.806842,3.8479972,3.8685746,3.4467354,2.7230926,2.3904223,2.0577524,2.369845,3.3061223,4.187526,3.666229,2.843128,2.510458,2.335549,2.1332035,1.8588364,1.3821237,1.196926,1.0288762,0.7888051,0.59674823,0.7476501,0.72021335,0.64819205,0.61389613,0.6207553,0.66876954,0.6893471,0.6241849,0.5555932,0.7099246,1.0220171,1.8519772,2.4658735,2.6922262,2.9460156,3.7965534,3.6696587,3.316411,3.1517909,3.2546785,3.5770597,4.413879,5.2987127,5.9914894,6.492209,6.550512,6.8866115,7.1987042,7.208993,6.660259,5.7479887,5.0483527,4.6127954,4.3692946,4.125794,4.4413157,4.461893,4.355576,4.262977,4.280125,4.372724,4.6779575,4.4927597,3.9543142,4.029765,4.437886,5.5387836,5.9469047,5.796003,6.759717,7.589677,7.7885933,7.8126,7.706283,7.1198235,6.835168,6.725421,6.591667,6.3001523,5.7822843,5.761707,6.0978065,6.217842,6.001778,5.7479887,6.48535,6.451054,6.101236,5.7994323,5.8062916,5.5422134,5.2781353,5.113515,5.2266912,5.8988905,6.3961806,4.770556,2.9151495,1.879414,1.8485477,1.9239986,2.1126258,2.1640697,1.9823016,1.6187652,1.5981878,1.4129901,1.2277923,1.138623,1.1729189,1.1214751,1.2243627,1.4850113,1.8176813,2.037175,2.3801336,2.0646117,1.7079345,1.6564908,1.9651536,1.7799559,1.6736387,2.0063086,2.6133456,2.8156912,2.3081124,1.7799559,1.5981878,1.7422304,1.8416885,2.6064866,3.2443898,3.4638834,3.3712845,3.4604537,3.9440255,4.232111,3.9886103,3.8514268,5.4084597,5.9331865,6.5779486,7.1369715,7.723431,8.766026,7.8194594,7.5210853,7.9600725,9.2153015,11.348505,0.5658819,0.83338976,1.0117283,1.0768905,1.0940384,1.1900668,1.1763484,1.1489118,1.2312219,1.3992717,1.4335675,1.5570327,1.587899,1.7593783,2.0131679,2.0131679,1.6599203,1.6256244,1.6256244,1.5981878,1.7079345,1.2346514,1.2792361,1.3443983,1.2895249,1.3272504,1.1077567,0.77851635,0.5453044,0.48357183,0.53501564,0.5212973,0.6001778,0.69963586,0.8093826,0.9911508,1.1489118,1.3375391,1.5021594,1.6564908,1.8759843,2.1812177,2.5070283,2.9082901,3.216953,3.0214665,3.0317552,3.474172,3.7382503,3.6627994,3.5393343,3.333559,3.0043187,2.9460156,3.3438478,4.2115335,4.383013,5.219832,5.686256,5.857735,6.941485,7.0786686,7.2295704,7.9017696,8.786603,8.772884,8.772884,9.523964,9.764035,9.345626,9.246168,9.770895,10.597425,11.47197,11.952112,11.413667,12.511135,12.6586075,12.157887,11.4205265,10.957532,10.041832,9.56512,9.458802,9.592556,9.750318,9.493098,9.355915,9.571979,10.096705,10.635151,11.760056,12.788932,14.109323,15.721229,17.271402,16.660936,16.482597,16.20137,15.62863,14.908417,16.578627,17.264544,17.69667,17.806417,16.70895,16.53747,17.034761,17.384579,17.521763,18.142517,18.410025,19.054789,20.008213,20.76958,20.416334,19.586374,18.499195,17.724108,17.182234,16.143068,16.095055,15.971589,15.642348,15.477728,16.359133,19.349733,21.047379,21.11597,20.207129,19.987637,20.62554,21.03023,20.735287,19.757853,18.584934,18.279701,17.168514,16.108772,15.395418,14.784951,14.980438,14.479718,13.375391,12.247057,12.161317,12.308789,12.288212,12.840376,13.896688,14.616901,14.582606,14.637479,14.496866,13.954991,12.895248,12.614022,12.679185,13.570878,14.935853,15.594335,14.898128,14.55174,14.30138,13.920695,13.197053,12.05157,10.995257,10.275044,10.007536,10.179015,10.22703,10.504827,10.679735,10.957532,12.055,12.274493,12.785502,13.176475,13.406258,13.810948,14.846684,16.13278,17.017612,17.226818,16.859852,17.079346,17.53891,17.38115,16.70552,16.571766,17.058767,17.024471,16.482597,15.618341,14.802099,14.592895,14.339106,14.30481,14.4145565,14.267084,14.668345,14.71636,14.435134,13.872682,13.090735,13.4474125,13.670336,13.440554,12.836946,12.360233,11.1393,10.38479,9.97667,9.853205,10.024684,10.501397,10.868362,11.105004,11.348505,11.8869505,11.934964,12.113303,12.600305,13.409687,14.373401,15.63206,16.606062,17.117071,17.031332,16.249386,16.46888,16.88386,17.322845,17.802988,18.523201,18.718689,18.749556,18.38259,17.837284,17.775553,17.851004,17.226818,16.427725,15.707511,15.059319,15.830976,15.536031,15.700651,16.482597,16.678083,16.300829,15.728088,15.014734,14.5414505,15.028452,13.282792,12.840376,12.614022,11.718901,9.462232,11.461681,10.854645,10.542552,11.015835,10.347065,9.403929,10.854645,11.050131,8.841476,5.56965,7.596536,7.39762,5.885172,4.187526,3.6627994,12.157887,22.100262,19.078794,6.9620624,7.888051,27.820814,22.570116,13.22106,10.014396,12.343085,8.669997,16.064188,15.721229,7.023795,7.5382333,8.745448,7.034084,6.619104,8.241299,9.170717,12.442543,11.482259,9.952662,8.927217,6.914048,5.055212,4.7842746,5.003768,5.0414934,4.6402316,5.518206,5.7102633,6.5710897,7.857185,7.7371492,9.72631,10.799771,9.263316,7.4113383,11.550851,6.3618846,6.2727156,6.0532217,4.4584637,4.2252517,1.8348293,3.532475,5.2918534,5.360445,4.2869844,3.40901,4.3624353,4.7019644,4.256118,5.1100855,3.9508848,4.331569,4.623084,4.07435,2.7916842,3.1346428,3.5221863,4.1017866,4.4584637,3.6147852,4.214963,4.170378,3.9200184,3.5599117,2.8534167,2.8054025,3.7519686,3.882293,2.5996273,0.548734,0.30523327,0.22635277,0.22635277,0.2194936,0.12346515,0.19548649,0.24007112,0.2469303,0.31895164,0.6859175,0.42869842,0.97057325,1.1523414,0.8162418,0.7922347,0.4629943,0.39097297,0.39783216,0.39097297,0.36696586,0.61046654,0.85396725,0.9774324,1.1694894,1.937717,2.170929,2.750529,3.2546785,3.549623,3.7691166,3.9886103,4.190956,4.057202,3.6936657,3.6319332,3.6182148,3.2306714,2.9631636,2.9803114,3.1277838,3.275256,3.1277838,2.9254382,2.8122618,2.8396983,2.6167753,2.3904223,1.9857311,1.5124481,1.3443983,0.96371406,0.9877212,1.1763484,1.3752645,1.5090185,1.3032433,1.0597426,1.1317638,1.5364552,1.9514352,1.9171394,1.8142518,1.7662375,1.8897027,2.3046827,2.976882,3.5461934,3.875434,4.0091877,4.180667,4.4721823,4.9694724,5.346727,5.360445,4.835718,3.3232703,3.000889,2.9700227,2.8465576,2.760818,3.2272418,1.9411465,2.819121,5.3570156,4.623084,4.695105,7.332458,9.458802,9.510246,7.4456344,8.508806,7.208993,9.040393,11.201033,2.5927682,9.040393,11.262765,8.944365,5.2918534,7.051232,5.1340923,6.217842,5.3570156,2.335549,1.6633499,2.5893385,2.1743584,2.0749004,3.6079261,7.720001,5.2438393,7.874333,10.566559,10.679735,7.9943686,9.630281,6.159539,4.852866,5.703404,1.4198492,1.0288762,1.8279701,2.5893385,3.100347,4.149801,4.0777793,3.590778,3.0557625,2.627064,2.2738166,1.786815,2.4795918,3.4776018,3.875434,2.7162333,2.644212,2.4795918,2.503599,2.534465,1.9239986,2.0817597,2.0749004,2.1469216,2.0234566,0.90198153,1.0117283,2.1091962,3.4947495,4.245829,3.2203827,3.292404,3.4398763,3.4878905,3.3952916,3.2512488,3.457024,4.664239,5.8234396,6.427047,6.4990683,5.3878818,4.9180284,4.479041,3.8617156,3.2512488,3.8960114,3.1517909,2.4144297,2.4452958,3.3712845,3.7622573,4.2081037,4.214963,3.82399,3.6147852,4.105216,3.7519686,3.4878905,3.532475,3.3884325,4.2526884,4.149801,3.649081,3.234101,3.2958336,2.9665933,3.3061223,3.566771,3.450165,3.083199,3.3266997,3.2032347,3.1552205,3.2272418,3.083199,2.8019729,2.750529,3.0077481,3.3781435,3.4021509,3.9165888,3.9063,3.7039545,3.4021509,2.8534167,2.9494452,2.4898806,2.784825,3.82399,4.2869844,3.5564823,2.767677,2.1812177,1.8588364,1.6633499,1.2346514,1.2037852,1.1592005,0.9362774,0.59674823,0.6790583,0.65505123,0.59674823,0.5590228,0.59674823,0.59674823,0.64133286,0.61046654,0.5418748,0.6241849,0.66191036,1.0014396,1.8142518,2.9220085,3.799983,4.396731,4.383013,3.6868064,2.983741,3.6936657,3.9371665,4.0057583,4.4516044,5.3570156,6.3310184,6.6876955,6.9380555,7.5245147,8.210432,8.086967,7.14726,6.307011,5.857735,5.638242,5.0655007,4.6882463,4.6676683,4.7019644,4.6436615,4.4859004,4.705394,4.852866,4.6402316,4.081209,3.4947495,3.8720043,5.442755,6.3001523,6.3207297,7.1266828,7.6616983,7.9086285,7.747438,7.2295704,6.5470824,6.8283086,6.8591747,6.684266,6.3447366,5.90575,6.135532,6.615674,6.7185616,6.526505,6.8214493,7.8331776,8.525954,8.100685,6.9792104,6.8214493,6.759717,6.276145,5.7651367,5.641671,6.3618846,6.166398,4.791134,3.0866287,1.8382589,1.7388009,1.9239986,2.3801336,2.6613598,2.534465,1.9994495,1.8897027,1.7593783,1.7353712,1.7696671,1.646202,1.488441,1.5124481,1.6530612,1.8554068,2.0749004,2.318401,2.2806756,2.1160555,2.0131679,2.1983654,2.3424082,2.1880767,2.2120838,2.609916,3.2821152,2.633923,2.1332035,1.8965619,1.8279701,1.6324836,2.4384367,2.959734,3.083199,3.093488,3.6936657,3.5221863,4.4584637,4.396731,3.5153272,4.273266,6.0669403,6.8900414,7.4456344,8.05953,8.683716,8.961512,7.888051,7.2364297,7.9086285,9.932085,0.6241849,0.8848336,0.91912943,0.9328478,0.9877212,1.0082988,1.3649758,1.3409687,1.2483698,1.2243627,1.2037852,1.1489118,1.1146159,1.255229,1.4541451,1.3169615,1.2277923,1.2003556,1.2106444,1.2517995,1.3443983,1.2175035,1.2860953,1.1249046,0.7888051,0.8265306,0.6276145,0.52815646,0.4938606,0.48700142,0.4972902,0.44584638,0.42183927,0.4355576,0.5144381,0.69963586,0.88826317,1.0734608,1.2758065,1.5021594,1.7319417,2.2292318,2.9974594,3.4055803,3.4021509,3.508468,3.6696587,4.190956,4.386442,4.1155047,3.8102717,3.4535947,3.3198407,3.5359046,4.3178506,5.9571934,4.7019644,4.722542,5.0895076,5.6039457,6.807731,6.5813785,6.5710897,6.708273,6.9346256,7.174697,8.200144,9.2153015,9.846346,9.702303,8.344186,8.086967,8.573969,9.788043,11.255906,12.034423,12.363663,12.483699,12.349944,11.965831,11.396519,11.2593355,10.48082,9.788043,9.496528,9.517105,9.39021,9.194724,10.415657,12.315649,11.952112,13.066729,13.941273,14.568888,15.05246,15.6252,16.029892,16.506605,16.767254,16.647217,16.091625,15.858413,15.7966795,16.53404,17.38115,16.331696,15.340545,15.776102,16.417435,16.928444,17.861292,17.700102,17.658945,18.238546,19.188541,19.486916,18.36544,17.28512,16.657507,16.492886,16.414005,16.938732,18.410025,18.979338,18.176813,16.907866,18.70497,18.862732,19.246845,20.141968,20.244854,20.176264,19.881319,18.893597,17.600643,17.230247,18.241976,17.477179,15.4914465,13.54687,13.601744,13.697772,13.004995,12.744347,13.121602,13.320518,12.627741,12.157887,12.092726,12.432255,13.004995,13.7526455,14.500296,14.661487,14.05102,12.881531,11.808069,11.540562,12.127021,13.351384,14.7026415,14.994157,14.328816,13.786942,13.615462,13.234778,12.411677,11.640019,11.043272,10.621432,10.275044,10.285333,9.791472,9.884071,10.88894,12.360233,12.041282,11.821788,12.147599,12.922686,13.491997,14.568888,15.738377,16.715809,17.271402,17.226818,17.309128,17.12736,16.736387,16.208231,15.608052,15.830976,15.755525,15.402277,14.894698,14.445422,13.917266,13.745787,13.670336,13.437123,12.80265,13.430264,13.759505,13.937843,13.917266,13.457702,13.022143,12.764925,12.418536,11.996697,11.773774,11.012405,10.196163,9.616563,9.3079,9.047252,9.650859,10.285333,10.772334,11.194174,11.897239,11.938394,12.075578,12.5145645,13.162757,13.629181,15.05246,16.221949,17.027903,17.38115,17.21653,16.6335,17.37429,18.11165,18.427174,18.804428,18.910746,18.694681,18.145947,17.662374,18.019053,18.560926,18.694681,18.588364,18.12537,16.904436,17.312557,16.904436,16.88386,17.470318,17.909306,16.71238,16.311117,16.067617,15.71437,15.323397,13.478279,13.917266,13.999576,12.80265,11.122152,11.873232,9.928656,9.6988735,11.070708,9.3936405,8.433355,6.6636887,5.2918534,4.979761,5.8371577,5.521636,5.3227196,9.054111,12.758065,4.722542,15.347404,10.823778,10.261326,18.3723,25.502413,12.46998,13.05301,14.695783,13.872682,16.067617,10.302481,8.920357,6.7185616,4.180667,7.4765005,9.14328,8.762596,8.580828,9.016385,8.64599,9.623423,8.340756,7.363324,6.9963584,5.2781353,4.8288593,4.8322887,4.9420357,5.055212,5.346727,5.90232,6.0223556,6.6293926,7.630832,7.9189177,9.949233,10.827208,10.278474,9.3936405,10.611144,6.368744,5.288424,4.705394,3.5564823,2.3458378,2.0131679,3.7313912,5.439326,5.936616,4.8734436,3.4981792,2.9700227,3.532475,5.0757895,7.15069,8.587687,6.166398,3.9097297,2.9151495,1.3409687,3.9165888,4.6093655,5.103226,5.658819,5.06893,4.7499785,3.6044965,3.1243541,3.4638834,3.4398763,3.9268777,3.765687,3.3129816,2.5447538,1.0494537,0.39440256,0.1920569,0.19548649,0.23664154,0.20920484,0.4081209,0.4046913,0.33266997,0.32238123,0.5041494,0.45270553,0.91227025,0.9877212,1.0117283,2.551613,0.9534253,0.67219913,0.65162164,0.4664239,0.30523327,0.59674823,0.8093826,1.1043272,1.4610043,1.6942163,2.3149714,3.2066643,4.1017866,4.7808447,5.038064,5.103226,4.90431,4.40359,3.8960114,4.0229063,3.8342788,3.6799474,3.5599117,3.549623,3.8102717,3.9783216,3.5359046,3.1689389,3.117495,3.1792276,3.192946,3.1792276,2.7985435,2.1400626,1.6839274,1.5398848,1.3615463,1.3443983,1.4850113,1.5707511,1.6770682,1.6187652,1.7730967,2.1160555,2.2566686,2.386993,2.270387,2.1469216,2.2052248,2.5619018,3.018037,3.0660512,3.2958336,3.7176728,3.74168,4.249259,5.425607,6.2075534,6.217842,5.7891436,4.996909,4.197815,3.4124396,2.8225505,2.7368107,3.6010668,2.901431,2.5241764,3.3301294,5.137522,5.1409516,5.8474464,7.363324,9.280463,10.693454,12.682614,14.815818,12.826657,8.515666,9.73317,7.3118806,13.612033,12.812939,5.1512403,6.9380555,7.034084,6.8214493,5.4187484,3.450165,3.0420442,3.532475,3.2066643,2.9254382,4.383013,10.13786,6.3790326,7.798882,11.489118,13.22106,7.4113383,6.5059276,5.381023,5.346727,5.5730796,3.0557625,2.527606,2.0028791,1.6976458,2.1812177,4.3933015,4.173808,4.588788,3.974892,2.6613598,2.9803114,2.16064,2.2086544,2.7916842,3.2821152,2.7299516,2.627064,2.3081124,2.218943,2.3218307,2.0920484,2.5927682,2.5207467,2.386993,2.3081124,1.9754424,1.7422304,2.1126258,2.5310357,3.000889,4.07435,3.2306714,3.0729103,3.5359046,4.2595477,4.5819287,4.681387,4.8117113,5.4941993,6.3035817,5.888602,5.5422134,5.2815647,5.130663,4.9934793,4.6676683,4.2766957,3.765687,3.3644254,3.3369887,3.9714622,4.029765,4.420738,4.3109913,3.8205605,4.0434837,4.852866,4.396731,4.0606318,4.166949,3.974892,4.4413157,4.4996185,4.046913,3.4192986,3.3815732,3.433017,3.4844608,3.5564823,3.6147852,3.5702004,3.8925817,3.9131594,3.57363,3.0489032,2.7642474,2.7951138,2.7333813,2.633923,2.568761,2.620205,3.5942078,3.8102717,3.9131594,3.6868064,2.0234566,3.3609958,2.3595562,1.99602,2.9631636,3.7005248,4.1017866,4.125794,3.6182148,2.8019729,2.2841053,1.7525192,1.4267083,1.3992717,1.4267083,0.94999576,0.82996017,0.805953,0.7133542,0.5796003,0.59674823,0.6927767,0.78537554,0.6962063,0.5144381,0.58988905,0.84024894,0.881404,1.2449403,2.1023371,3.275256,4.420738,4.972902,4.57164,3.7622573,4.0229063,4.314421,4.3178506,4.396731,4.8014226,5.662249,6.0840883,6.697984,7.5382333,8.289313,8.296172,8.186425,7.5245147,6.8866115,6.5024977,6.262427,5.425607,4.8425775,4.629943,4.7979927,5.254128,5.5250654,5.336438,4.870014,4.3281393,3.9474552,4.0709205,5.254128,6.5127864,7.3393173,7.675417,7.2364297,6.5196457,5.826869,5.6210938,6.509357,7.267296,7.4010496,7.2364297,7.016936,6.883182,6.5779486,6.7974424,6.9826403,7.15069,7.881192,9.472521,11.012405,10.847785,9.352485,8.920357,8.31332,8.40249,7.8674736,6.708273,6.2658563,6.090947,5.192395,3.998899,2.8396983,1.9582944,2.0440342,2.668219,3.0866287,2.9494452,2.3046827,2.1743584,2.4967396,2.726522,2.7093742,2.6853669,2.633923,2.4452958,2.2292318,2.0989075,2.1743584,2.1332035,2.2052248,2.153781,1.978872,1.9274281,2.037175,2.3767042,2.4795918,2.5447538,3.450165,2.8534167,2.4315774,2.2806756,2.3252604,2.3149714,2.8877127,2.9906003,3.2992632,3.957744,4.5853586,3.7485392,4.2252517,4.664239,4.547633,4.2115335,4.8837323,5.360445,6.2384195,7.205563,7.0478024,8.05953,7.366754,6.7185616,6.9792104,8.128122,0.72364295,0.8128122,0.77508676,0.823101,0.9602845,0.9877212,1.4095604,1.5055889,1.3615463,1.1043272,0.91569984,0.9294182,1.0528834,1.1832076,1.2106444,1.0151579,1.0151579,0.922559,0.8848336,0.90198153,0.84024894,0.7888051,0.7682276,0.64476246,0.45613512,0.42869842,0.34981793,0.37039545,0.40126175,0.41840968,0.4698535,0.34295875,0.31209245,0.3806842,0.51100856,0.6344737,0.8162418,0.9431366,1.0906088,1.3169615,1.6564908,2.2566686,2.8465576,3.1723683,3.2821152,3.532475,3.8514268,4.15666,4.40702,4.400161,3.7759757,3.8308492,3.789694,4.256118,5.147811,5.6965446,4.73969,4.6127954,4.7088237,4.9351764,5.7136927,5.953764,6.1766872,6.3035817,6.2418494,5.895461,6.6053853,7.582818,8.39563,8.652849,7.997798,7.7885933,7.9737906,9.033533,10.525404,11.094715,10.796341,10.912948,11.046701,10.820349,9.884071,10.55284,10.816919,10.693454,10.388221,10.31277,11.050131,12.133881,13.838386,15.05246,13.282792,14.003006,14.400838,14.452282,14.400838,14.774663,15.71094,16.071047,16.108772,16.13621,16.516893,16.722668,16.647217,16.732958,16.719238,15.63206,15.028452,15.940722,17.058767,17.63151,17.470318,17.408587,17.734396,18.831865,20.03908,19.668684,17.878439,17.274832,17.449741,17.943602,18.217968,17.909306,18.650097,19.147387,18.670673,17.051908,17.566347,17.20624,17.514904,18.70154,19.6241,19.853882,19.342873,18.993055,18.934752,18.492336,18.656956,17.929884,16.283682,14.428274,13.790371,13.279363,12.830087,13.186764,14.085316,14.243076,13.337666,12.466551,11.945253,11.869802,12.099585,13.231348,13.852104,13.982429,13.656617,12.950122,11.427385,10.55284,10.834066,12.161317,13.80409,14.839825,13.975569,13.2862215,13.317088,13.097594,12.373952,11.996697,11.605724,11.177026,10.995257,11.382801,10.834066,10.388221,10.666017,11.842365,12.041282,11.777204,11.787492,12.154458,12.30536,13.368532,14.730078,16.016174,16.931873,17.243965,17.497755,16.78783,16.208231,15.988737,15.501736,15.772673,15.518884,15.323397,15.237658,14.788382,14.054449,13.519434,12.895248,12.130451,11.399949,12.13731,12.476839,12.833516,13.186764,13.101024,12.504276,12.140739,11.808069,11.547421,11.646879,11.249047,10.690024,10.124143,9.589127,8.995808,9.441654,9.89436,10.233889,10.600855,11.38966,11.924676,12.490558,13.056439,13.488567,13.55373,14.586036,15.707511,16.45859,16.767254,16.96274,16.890718,17.703531,18.341434,18.554068,18.883308,18.427174,18.012194,17.679523,17.576635,17.943602,18.567787,19.092514,19.154245,18.722118,18.077356,18.725548,18.231688,17.940172,18.180243,18.265984,17.250826,17.528622,17.29541,16.307688,15.909856,13.982429,14.006435,13.38911,11.756626,10.950673,11.602294,10.823778,11.314209,11.595435,6.0326443,8.114404,5.284994,3.7279615,4.636802,4.2286816,3.3850029,3.4810312,6.6225333,10.72775,9.530824,10.55284,6.742569,10.789482,22.851341,30.547335,9.829198,15.391989,16.636929,8.567109,11.790922,6.7631464,5.6142344,5.5662203,6.262427,9.788043,8.999237,9.006097,9.177576,9.0369625,8.2310095,8.522525,7.3118806,6.3961806,5.895461,4.2526884,4.880303,4.650521,4.3624353,4.537344,5.394741,5.6073756,6.2864337,6.077229,5.6656785,7.764586,8.865483,7.9463544,7.2638664,7.3598948,7.0443726,4.40359,5.8234396,5.9400454,3.7622573,2.6922262,8.032094,11.050131,10.72775,7.870903,5.137522,3.5050385,2.527606,3.0660512,4.8014226,6.2212715,8.1212635,6.0978065,3.3644254,1.7559488,1.728512,4.170378,5.127233,5.535354,5.693115,5.2781353,5.020916,4.4859004,4.0366244,3.8514268,3.9337368,4.32128,4.4104495,4.1772375,3.5564823,2.4555845,0.8196714,0.34295875,0.28808534,0.25721905,0.20234565,0.32924038,0.4389872,0.48014224,0.48357183,0.5693115,0.66191036,0.8128122,0.8093826,0.91227025,1.8382589,1.0048691,0.8711152,0.83338976,0.66876954,0.5555932,0.764798,0.8676856,1.0117283,1.2689474,1.6496316,2.218943,3.3644254,4.4584637,5.1512403,5.3741636,5.353586,4.0057583,3.8514268,4.8288593,4.2766957,4.314421,4.3658648,4.197815,3.9611735,4.173808,4.0674906,3.7725463,3.5633414,3.590778,3.9063,3.7519686,3.7965534,3.5187566,2.9391565,2.6407824,2.7162333,2.277246,1.9411465,1.8897027,1.862266,1.9068506,2.0577524,2.2155135,2.277246,2.16064,2.6545007,2.836269,2.860276,2.8739944,3.018037,3.333559,3.4638834,3.7553983,4.2046742,4.4550343,4.722542,5.3570156,5.857735,6.0532217,6.0806584,5.669108,5.2266912,4.40702,3.391862,2.8945718,3.683377,3.5461934,2.7951138,2.860276,6.2898636,8.028665,9.537683,10.028113,10.175586,12.127021,16.839275,14.102464,8.7283,5.5730796,9.523964,6.725421,10.381361,9.767465,4.90431,6.5813785,7.4970784,5.802862,3.9028704,2.843128,2.287535,2.3595562,2.6579304,3.590778,6.4407654,13.38911,5.919468,5.785714,9.071259,12.22648,12.041282,12.421966,10.666017,8.525954,6.550512,4.0503426,2.8054025,1.8519772,1.3101025,1.4678634,2.7985435,4.1017866,4.6127954,4.372724,3.6696587,3.0214665,2.2120838,2.218943,2.486451,2.5653315,2.1194851,2.2052248,2.2292318,2.3904223,2.5893385,2.4212887,2.6407824,2.5550427,2.4795918,2.5070283,2.527606,1.7696671,2.411,2.8980014,3.069481,4.1772375,3.7931237,3.6010668,4.0949273,4.979761,5.178677,5.552502,5.610805,6.0703697,6.6876955,6.2692857,5.9914894,5.521636,5.284994,5.305572,5.2026844,4.4687524,3.8205605,3.5016088,3.6387923,4.266407,4.2115335,4.5784993,4.3933015,3.7451096,3.765687,4.6436615,4.7602673,4.681387,4.6436615,4.557922,4.1943855,3.9851806,3.7176728,3.4810312,3.6696587,3.974892,3.8720043,3.7348208,3.707384,3.6936657,4.1017866,4.417309,4.201245,3.5359046,3.0043187,3.234101,3.199805,3.0626216,2.9151495,2.7573884,3.3952916,3.6147852,3.566771,3.2718265,2.6133456,3.5359046,2.9700227,2.5756202,2.9665933,3.7211025,4.372724,4.547633,4.4413157,4.1463714,3.6593697,3.1106358,2.7093742,2.4247184,2.1846473,1.862266,1.5227368,1.2483698,1.0185875,0.85739684,0.823101,0.91569984,0.9259886,0.805953,0.6310441,0.5796003,0.7613684,0.8505377,0.96371406,1.3546871,2.4007113,3.625074,4.4275975,4.5956473,4.431027,4.746549,5.1752477,5.305572,5.07236,4.698535,4.722542,5.127233,5.970912,6.9071894,7.6788464,8.117833,8.2310095,8.100685,7.781734,7.366754,6.9826403,6.3447366,5.4770513,4.928317,5.0655007,6.0326443,6.159539,5.7754254,5.130663,4.5339146,4.341858,4.746549,5.888602,7.291303,8.429926,8.700864,8.076678,6.7631464,5.7582774,5.689686,6.848886,7.390761,7.48336,7.442205,7.4936485,7.7748747,7.407909,7.1987042,7.3564653,7.9086285,8.707723,10.14129,11.4205265,11.729189,11.2593355,11.211322,10.065839,9.451943,8.625413,7.5039372,6.660259,6.15268,5.4907694,4.65395,3.666229,2.5996273,2.3389788,2.4418662,2.702515,2.860276,2.5893385,2.603057,2.819121,3.0283258,3.2135234,3.5599117,3.5118976,3.1243541,2.7642474,2.585909,2.534465,2.3972816,2.335549,2.2395205,2.0474637,1.7696671,1.7730967,2.2498093,2.5584722,2.867135,4.15323,3.2375305,2.5996273,2.3492675,2.4075704,2.4967396,3.3987212,3.4878905,3.7108135,4.2218223,4.40359,4.2218223,4.7808447,5.302142,5.4804807,5.48734,5.7891436,5.8405876,6.0395036,6.355026,6.3173003,7.2192817,7.4044795,7.2947326,7.346176,8.069819,0.7305021,0.70649505,0.6927767,0.7476501,0.8505377,0.90198153,1.1729189,1.2723769,1.1660597,0.9362774,0.77508676,0.8128122,1.0014396,1.1077567,1.039165,0.84367853,0.7956643,0.70649505,0.67219913,0.66533995,0.5418748,0.40126175,0.33609957,0.29494452,0.26064864,0.22635277,0.24007112,0.26750782,0.26750782,0.26407823,0.35324752,0.25721905,0.29837412,0.44584638,0.6207553,0.6962063,0.91227025,0.980862,1.0666018,1.2860953,1.704505,2.170929,2.469303,2.6990852,2.9220085,3.175798,3.532475,3.7279615,4.0263357,4.2526884,3.7931237,4.4413157,4.7979927,5.435896,5.9640527,5.0140567,4.7671266,4.8014226,4.770556,4.712253,5.0586414,5.744559,6.0840883,6.111525,5.871454,5.4153185,5.284994,6.018926,6.694555,7.0135064,7.298162,7.394191,7.682276,8.443645,9.445084,9.945804,9.740028,9.801761,9.89093,9.767465,9.194724,10.062409,11.063849,11.612583,11.770344,12.240198,13.725209,15.385129,16.163645,15.700651,14.373401,14.476289,14.339106,14.160767,14.260224,15.073037,15.848124,15.851553,15.4742985,15.261664,15.923574,16.561478,16.441442,15.920145,15.371411,15.179354,15.158776,15.96816,16.846134,17.113642,16.177364,15.9613,16.70895,18.307138,19.895037,19.847023,18.602083,17.936743,17.71382,17.912735,18.62266,18.341434,18.262554,18.591793,18.746124,17.364002,16.074476,15.313108,15.854982,17.525192,19.164536,19.222837,18.557497,18.62266,19.438902,19.61038,19.301718,18.28999,17.12736,16.13621,15.402277,14.13333,13.491997,13.742357,14.483148,14.644339,14.123041,13.2862215,12.63117,12.377381,12.452832,13.155897,13.471419,13.516005,13.272504,12.617453,11.101575,10.268185,10.261326,11.039842,12.397959,13.80066,13.5503,13.094165,13.015285,13.018714,12.109874,11.756626,11.530273,11.303921,11.2593355,11.821788,11.739478,11.46854,11.372512,11.732618,12.63803,12.607163,12.229909,11.876661,11.688034,12.88839,14.342535,15.604623,16.516893,17.226818,17.765263,17.36057,16.822126,16.335125,15.470869,15.676644,15.676644,15.8138275,15.988737,15.662926,14.308239,13.22106,12.291641,11.489118,10.864933,11.1393,11.327928,11.626302,12.048141,12.411677,11.924676,11.578287,11.279913,11.122152,11.38966,11.55771,11.406808,10.967821,10.360784,9.80862,9.736599,9.839486,9.9801,10.295622,11.211322,12.082437,12.812939,13.402828,13.783512,13.821238,14.435134,15.319967,15.985307,16.335125,16.681513,17.055338,17.768692,18.279701,18.468328,18.6158,17.744686,17.343424,17.271402,17.425734,17.748116,18.547209,18.999914,18.9519,18.691252,18.927893,19.768143,19.558937,19.363451,19.346302,18.766703,18.193962,18.95876,18.79414,17.446312,16.684942,14.249936,13.71492,13.039291,12.017275,12.253916,11.866373,11.509696,11.756626,11.019264,5.552502,8.584257,5.2644167,4.5030484,6.842027,4.437886,4.256118,3.1380725,5.7582774,10.487679,9.403929,6.4716315,9.55826,16.311117,22.573545,22.381487,9.760606,14.836395,13.371962,4.064061,8.536243,4.7259717,5.6313825,7.1232533,8.182996,10.916377,8.457363,8.567109,8.899779,8.357904,7.082098,7.0478024,6.1561093,5.4496145,5.0174866,3.9851806,5.1340923,4.7431192,4.341858,4.6848164,5.7308407,5.73427,6.334448,5.950334,5.3432975,7.6171136,7.8606143,6.228131,5.23698,5.1752477,4.1189346,3.1963756,7.2295704,8.14527,5.0106273,4.040054,11.187314,15.134769,13.049581,7.222711,5.096367,2.983741,2.2429502,3.0043187,4.437886,4.7774153,6.5642304,5.675967,3.433017,1.6153357,2.435007,4.822,5.717122,5.7822843,5.4736214,5.06893,5.2609873,5.295283,4.928317,4.5442033,5.1409516,5.305572,5.422178,5.2575574,4.7259717,3.8960114,1.920569,0.90541106,0.4664239,0.30523327,0.23664154,0.29494452,0.4698535,0.607037,0.6756287,0.7888051,0.90541106,0.83338976,0.78194594,0.83681935,0.9534253,0.97400284,0.9842916,0.89169276,0.7442205,0.72707254,0.84367853,0.9328478,1.0254467,1.255229,1.8588364,2.1572106,3.3026927,4.3658648,5.020916,5.562791,5.0174866,3.5599117,3.3472774,4.386442,4.5270553,4.7362604,4.996909,4.955754,4.715683,4.846007,4.3933015,4.280125,4.1772375,4.1292233,4.554492,4.149801,4.15666,4.0366244,3.7142432,3.5599117,3.6970954,3.1243541,2.5756202,2.318401,2.1674993,2.16064,2.3458378,2.4555845,2.3458378,2.020027,2.627064,2.9906003,3.2032347,3.3266997,3.3952916,3.5599117,3.940596,4.5442033,5.2335505,5.720552,5.6313825,5.6519604,5.809721,6.090947,6.4133286,5.8543057,5.501058,5.003768,4.2081037,3.175798,3.316411,3.6765177,3.433017,3.2683969,5.3570156,8.169277,10.487679,11.677745,12.298501,14.099034,15.690363,11.31078,6.591667,5.1169443,8.419638,6.0737996,5.802862,4.8117113,3.57363,5.830299,6.4133286,4.5201964,3.2821152,3.2546785,2.3972816,1.8485477,2.2052248,3.7211025,6.584808,10.916377,6.001778,4.7259717,7.4696417,12.740917,17.158226,21.723007,17.53548,10.9541025,5.888602,3.7862647,3.292404,2.4830213,1.9514352,1.9068506,2.1880767,3.0969174,3.882293,4.389872,4.297273,3.117495,2.16064,2.318401,2.4898806,2.270387,1.9651536,2.170929,2.1640697,2.294394,2.5447538,2.5310357,2.6133456,2.5173173,2.503599,2.627064,2.7333813,1.7490896,2.4418662,3.07634,3.3061223,4.197815,4.290414,4.180667,4.629943,5.3707337,5.1169443,5.8474464,5.9400454,6.1766872,6.5470824,6.2487082,6.217842,5.960623,5.65539,5.4496145,5.4599032,4.90431,4.417309,4.0503426,3.9886103,4.547633,4.7191124,5.0757895,4.7431192,3.8925817,3.7519686,4.5167665,5.0929375,5.15467,4.839148,4.712253,4.0674906,3.7279615,3.6044965,3.6456516,3.8342788,4.091498,4.091498,4.0366244,4.0194764,4.029765,4.434457,4.835718,4.705394,4.0674906,3.4947495,3.532475,3.4535947,3.3541365,3.2478194,3.059192,3.357566,3.4673128,3.3266997,3.0386145,2.8945718,3.357566,3.1312134,2.884283,3.000889,3.5976372,4.3349986,4.513337,4.7945633,5.1409516,4.787704,4.396731,4.057202,3.5393343,2.959734,2.7882545,2.5756202,2.1057668,1.6290541,1.2792361,1.0871792,1.0563129,0.99801,0.881404,0.7339317,0.64819205,0.66533995,0.78537554,0.82996017,0.9328478,1.546744,2.760818,3.7485392,4.4859004,5.0140567,5.422178,5.6656785,6.018926,5.686256,4.763697,4.2355404,4.5201964,5.3501563,6.385892,7.3564653,8.049242,8.193284,8.169277,8.069819,7.8674736,7.4284863,6.9037595,6.0978065,5.5490727,5.675967,6.773435,6.6465406,6.1286726,5.429037,4.9180284,5.1238036,5.6793966,6.5710897,7.864044,9.081548,9.225591,8.556821,7.2604365,6.385892,6.4236174,7.2947326,7.795452,7.98065,7.9909387,8.06639,8.525954,8.179566,7.956643,8.196714,8.769455,9.084977,10.278474,11.005547,11.30049,11.396519,11.732618,10.827208,10.199594,9.575408,8.755736,7.6274023,6.776865,5.919468,5.0620713,4.187526,3.2649672,2.6785078,2.417859,2.4452958,2.651071,2.8705647,3.1312134,3.0454736,3.0729103,3.4604537,4.2355404,4.0777793,3.6079261,3.216953,3.0077481,2.7813954,2.6545007,2.568761,2.3561265,2.0303159,1.8073926,1.6736387,1.99602,2.4041407,3.000889,4.355576,3.683377,3.093488,2.7985435,2.819121,2.9906003,3.8342788,4.029765,4.125794,4.386442,4.8014226,5.24041,5.446185,5.6519604,5.9160385,6.138962,5.953764,5.802862,5.6656785,5.703404,6.245279,6.684266,7.3358874,7.6685576,7.6788464,7.881192,0.6859175,0.6344737,0.6893471,0.70306545,0.66533995,0.6962063,0.78194594,0.764798,0.72707254,0.71678376,0.7579388,0.72021335,0.7922347,0.8265306,0.764798,0.6344737,0.53501564,0.5178677,0.5178677,0.4972902,0.4424168,0.22635277,0.17833854,0.16804978,0.15433143,0.17490897,0.20920484,0.1920569,0.14061308,0.12003556,0.216064,0.25378948,0.40126175,0.607037,0.7888051,0.85739684,1.1008976,1.1351935,1.2072148,1.4335675,1.7936742,1.9480057,2.1091962,2.2498093,2.386993,2.5790498,2.959734,3.2512488,3.5804894,3.9268777,4.125794,5.120374,5.950334,6.591667,6.492209,4.5990767,4.8905916,5.219832,5.3158607,5.23698,5.3741636,6.0532217,6.1732574,5.90232,5.518206,5.4084597,4.852866,5.394741,5.919468,6.183546,6.81802,7.058091,7.534804,7.9600725,8.4264965,9.400499,9.849775,9.853205,9.709162,9.640571,9.798331,10.220171,11.156448,11.965831,12.648318,13.845244,15.46401,16.585485,16.005884,14.5414505,15.031882,14.589465,14.171056,14.164196,14.733508,15.830976,15.930434,15.758954,15.268523,14.740367,14.760944,14.88441,14.490007,13.87954,13.646329,14.682064,14.863832,14.973578,15.13134,15.0078745,13.831526,13.070158,14.092175,15.930434,17.809847,19.157675,19.233126,17.960749,16.417435,15.649208,16.654078,17.820137,17.998474,18.265984,18.478617,17.250826,14.863832,13.862392,14.860402,17.243965,19.1954,18.653526,17.782412,17.525192,18.183672,19.401176,19.744135,18.389448,17.333136,17.117071,16.808409,15.364552,14.29795,13.944703,14.191633,14.496866,14.582606,14.119612,13.63604,13.437123,13.615462,13.512574,13.6086035,13.543441,13.077017,12.092726,10.916377,10.583707,10.374502,10.251037,10.871792,12.21619,12.860953,12.908967,12.668896,12.662037,11.664027,11.187314,11.0981455,11.166737,11.06042,11.489118,11.928105,12.339656,12.542002,12.21619,13.457702,13.663476,13.114742,12.325937,12.072148,13.251926,14.555169,15.539461,16.273392,17.346853,18.025911,18.434032,18.180243,17.175373,15.635489,15.337115,15.707511,16.239098,16.602633,16.6335,14.726648,13.166186,12.22648,11.777204,11.266195,10.854645,10.72775,10.714031,10.871792,11.482259,11.314209,11.05699,10.772334,10.618003,10.816919,11.543991,11.732618,11.506266,11.094715,10.813489,10.275044,10.158438,10.247607,10.590566,11.509696,12.404818,12.953552,13.38225,13.735497,13.876111,14.369971,15.059319,15.755525,16.324837,16.70552,16.921585,17.436022,17.940172,18.193962,18.025911,17.075916,16.849564,16.904436,17.072487,17.446312,18.636377,18.728977,18.584934,18.825006,19.809298,20.433481,20.721567,20.930773,20.872469,19.901896,19.726988,20.508932,20.443771,19.157675,17.682953,14.925565,14.387119,14.081886,13.618892,14.2190695,12.425395,11.084427,9.966381,9.156999,9.040393,9.438225,5.977771,6.1972647,9.290752,6.121814,6.8111606,3.649081,6.23156,11.537132,3.9165888,6.975781,13.622321,19.085653,18.70497,7.9429245,8.988949,9.3593445,6.9346256,4.3487167,8.992378,6.427047,7.6925645,8.484799,8.182996,9.863494,7.682276,7.888051,8.008087,7.0718093,5.597087,5.1580997,4.6573796,4.629943,4.9008803,4.554492,5.8337283,5.3707337,5.219832,5.936616,6.5882373,6.711703,6.420188,6.368744,6.776865,7.4113383,7.4524937,6.5985265,5.446185,4.249259,2.9391565,3.0900583,8.272165,9.547972,5.9914894,4.681387,9.719451,12.164746,9.338767,4.0194764,4.4516044,2.153781,1.9582944,3.3026927,4.98662,5.164959,7.0889573,6.121814,4.0366244,2.4384367,2.7711067,5.627953,6.276145,5.8474464,5.1992545,4.931747,5.188966,5.2472687,5.137522,5.2438393,6.3035817,6.416758,5.9812007,5.5662203,5.2438393,4.57507,3.2478194,1.7696671,0.77165717,0.4046913,0.33266997,0.38754338,0.5796003,0.75450927,0.8848336,1.0528834,1.1146159,1.0597426,0.9945804,0.9259886,0.764798,0.96371406,0.9945804,0.8676856,0.7133542,0.77165717,0.8471081,1.039165,1.2792361,1.6256244,2.2566686,2.2806756,3.210094,4.1120753,4.729401,5.4633327,4.90431,3.9714622,3.0626216,2.9391565,4.73969,5.192395,5.7102633,6.018926,6.0395036,5.878313,5.0586414,4.9660425,4.863155,4.6779575,5.003768,4.448175,4.3933015,4.434457,4.372724,4.201245,4.2835546,3.7553983,3.1895163,2.8568463,2.7162333,2.8396983,2.8396983,2.8328393,2.7573884,2.3664153,2.750529,3.0317552,3.2992632,3.5187566,3.5393343,3.5530527,4.064061,4.9523244,5.9160385,6.4579134,6.334448,6.279575,6.358455,6.5882373,6.9380555,6.0703697,5.48734,5.3330083,5.130663,3.806842,3.0317552,3.4638834,3.9954693,3.9303071,3.0077481,4.8151407,7.2535777,10.655728,14.037301,15.114192,10.161868,9.4862385,8.450503,6.5882373,7.579388,4.9008803,2.9048605,2.1126258,2.8739944,5.3570156,5.6828265,4.6436615,4.420738,4.8425775,3.3952916,2.5173173,2.335549,3.2649672,4.6848164,4.9488945,7.490219,6.2487082,8.7145815,15.498305,20.340883,27.676771,21.002794,11.170166,4.6402316,3.5016088,4.1017866,3.4055803,3.0900583,3.3712845,3.018037,1.7250825,2.9288676,4.0229063,4.0229063,3.5461934,2.294394,2.4041407,2.5961976,2.417859,2.2326615,2.4384367,2.1160555,1.9514352,2.1194851,2.2978237,2.5070283,2.4452958,2.5070283,2.7059445,2.6990852,1.9823016,2.3321195,2.9563043,3.6216443,4.671098,4.671098,4.506478,4.9180284,5.521636,4.8151407,5.638242,5.5902276,5.6313825,5.888602,5.6348124,6.0669403,6.420188,6.210983,5.662249,5.689686,5.576509,5.641671,5.271276,4.671098,4.8905916,5.2644167,5.717122,5.425607,4.530485,4.1155047,4.7431192,5.394741,5.3432975,4.6779575,4.290414,4.1120753,3.998899,3.9543142,3.9680326,4.0229063,4.07435,4.341858,4.5099077,4.5167665,4.5682106,4.914599,5.209543,5.0003386,4.389872,4.012617,3.6868064,3.5290456,3.4364467,3.357566,3.2546785,3.508468,3.5118976,3.4776018,3.316411,2.6407824,2.9288676,2.6545007,2.4967396,2.7059445,3.0900583,4.15323,4.4584637,4.9077396,5.5250654,5.470192,5.435896,5.171818,4.465323,3.6182148,3.4398763,3.5359046,3.1312134,2.503599,1.879414,1.4129901,1.1523414,1.0494537,0.939707,0.7990939,0.7579388,0.67219913,0.70306545,0.764798,0.83338976,0.9602845,2.0714707,3.2718265,4.479041,5.446185,5.7651367,5.641671,6.125243,5.919468,4.938606,4.331569,4.448175,5.0826488,6.2144127,7.4765005,8.1384115,8.416207,8.152129,7.9943686,8.025234,7.764586,7.1129646,6.64997,6.416758,6.584808,7.4284863,7.1849856,6.6739774,5.970912,5.521636,6.1321025,6.560801,6.999788,7.9943686,9.078118,8.779744,8.354475,7.6616983,7.2604365,7.3598948,7.822889,8.601405,9.170717,9.331907,9.1810055,9.129561,8.529384,8.573969,8.971801,9.287323,8.958082,10.007536,10.422516,10.436234,10.381361,10.696883,10.576848,10.789482,10.683165,9.9698105,8.700864,7.857185,6.6876955,5.5662203,4.647091,3.8514268,3.0969174,2.7745364,2.5447538,2.4590142,2.9494452,3.4535947,3.234101,3.1209247,3.5153272,4.420738,4.197815,3.8479972,3.5221863,3.2478194,2.9391565,2.8568463,2.8705647,2.5619018,2.0406046,1.9274281,1.7490896,1.7833855,2.037175,2.5824795,3.5564823,3.7348208,3.690236,3.5564823,3.4810312,3.6319332,4.0537724,4.2595477,4.2355404,4.4275975,5.720552,6.608815,6.279575,6.0052075,6.077229,5.826869,5.3090014,5.099797,5.161529,5.5490727,6.420188,6.3653145,6.790583,7.2604365,7.438775,7.1095347,0.8093826,0.65162164,0.6824879,0.6790583,0.5727411,0.48700142,0.6241849,0.6207553,0.5693115,0.548734,0.61046654,0.5727411,0.490431,0.37039545,0.26750782,0.30523327,0.39097297,0.37382504,0.28465575,0.18519773,0.19891608,0.1371835,0.08573969,0.06859175,0.07545093,0.07545093,0.11317638,0.13032432,0.15090185,0.1920569,0.29151493,0.42526886,0.64133286,0.8779744,1.0768905,1.1763484,1.2586586,1.2620882,1.3855534,1.611906,1.7079345,1.6496316,1.8348293,1.8588364,1.7353712,1.9068506,2.6887965,3.059192,3.508468,4.197815,4.945465,5.579939,6.077229,6.385892,6.0635104,4.256118,5.0277753,5.813151,6.2212715,6.252138,6.3001523,6.5230756,6.1904054,5.7891436,5.4084597,4.7602673,5.2609873,6.0806584,7.143831,8.158989,8.635701,8.56368,8.323608,8.241299,8.604835,9.705732,10.497967,10.621432,10.508256,10.299051,9.873782,9.72631,10.477389,11.159878,11.537132,12.099585,13.114742,13.7697935,14.287662,14.750656,15.107333,14.640909,14.572317,15.001016,15.536031,15.306249,14.791811,14.911846,15.05246,14.846684,14.174485,13.334236,12.785502,12.55915,12.644889,12.984418,12.874671,12.764925,13.083877,13.097594,10.926665,9.716022,11.482259,13.680624,15.323397,16.983316,16.678083,15.237658,13.900118,13.272504,13.320518,16.177364,17.778982,17.63151,16.21509,14.970149,15.042171,14.987297,15.769243,17.473747,19.318867,19.342873,18.37916,17.638369,17.655516,18.265984,19.349733,18.132229,16.88386,16.149927,14.7095,14.757515,14.332246,13.831526,13.615462,14.006435,14.2533655,13.900118,13.694343,13.858963,14.112752,14.140189,13.989287,13.560589,12.922686,12.312219,11.399949,10.738038,10.542552,10.64201,10.484249,11.38623,11.4754,11.835506,12.233338,11.122152,10.978109,11.105004,11.317638,11.4754,11.4754,11.866373,12.120162,12.168177,12.154458,12.435684,13.375391,13.711491,13.588025,13.22106,12.878101,13.059869,14.078457,15.261664,16.383139,17.638369,18.005335,18.334574,18.434032,18.073925,17.014183,15.536031,15.21365,15.776102,16.660936,17.014183,16.12249,14.424845,13.125031,12.511135,11.962401,11.756626,11.070708,10.401938,10.041832,10.100135,10.686595,10.734609,10.494537,10.220171,10.1481495,10.696883,10.871792,10.991828,11.05699,10.72775,10.679735,10.792912,11.039842,11.362224,11.705182,12.668896,13.248496,13.461131,13.337666,12.922686,13.728639,14.644339,15.45715,16.071047,16.510035,16.276823,16.530611,17.075916,17.525192,17.319416,16.37971,16.191082,16.245956,16.396858,16.859852,18.410025,18.324286,18.44432,19.504065,21.102251,21.006224,21.345753,21.712719,21.843042,21.62012,21.925352,22.422644,21.887627,20.344313,19.071936,17.840714,18.108221,16.496315,13.179905,11.8869505,11.55771,9.798331,7.466212,7.1952744,13.395968,9.72288,7.641121,7.805741,8.354475,4.914599,5.329579,2.4555845,0.4355576,0.48700142,0.90198153,11.080997,7.915488,7.970361,11.362224,1.7559488,11.080997,9.678296,7.0718093,7.4181976,9.506817,9.6645775,9.760606,8.97866,7.8366075,8.179566,6.848886,7.0375133,6.543653,5.305572,5.4016004,4.863155,4.6402316,5.761707,7.226141,5.9812007,7.5450926,6.550512,6.601956,7.9429245,7.4936485,8.296172,7.2158523,6.550512,6.800872,6.667118,7.301592,6.8111606,5.363875,3.5599117,2.4247184,2.0097382,7.116394,8.196714,4.170378,2.411,8.796892,4.870014,1.5741806,2.2429502,2.609916,1.8999915,2.1194851,4.187526,7.449064,9.657719,11.989838,8.344186,4.5819287,3.1140654,2.867135,5.1409516,5.970912,5.3570156,4.3349986,5.003768,3.99204,4.297273,5.0655007,5.5490727,5.096367,5.4153185,4.705394,4.32128,4.3795834,3.7691166,3.5873485,2.4967396,1.3375391,0.58988905,0.3806842,0.4664239,0.7888051,1.0837497,1.2243627,1.2346514,1.2963841,1.5227368,1.4850113,1.1214751,0.71678376,0.8265306,0.864256,0.8711152,0.89512235,0.9911508,1.0768905,1.371835,1.7216529,2.1126258,2.6853669,2.5996273,3.3850029,4.245829,4.5853586,3.998899,6.3790326,3.9714622,2.369845,3.3232703,4.715683,6.2041235,7.0615206,7.7028537,7.891481,6.7459984,5.425607,5.223262,5.2506986,5.223262,5.4941993,4.9077396,4.887162,4.979761,4.9351764,4.715683,4.8734436,4.482471,4.07435,3.9474552,4.180667,4.557922,4.2698364,4.0366244,4.040054,3.9063,4.0023284,4.0846386,4.1017866,3.9440255,3.4192986,3.3815732,3.782835,4.280125,4.712253,5.127233,5.8234396,6.279575,6.584808,6.8626046,7.2775846,6.852316,6.715132,6.5950966,6.210983,5.295283,4.0606318,3.4776018,3.782835,4.280125,3.3266997,1.6530612,4.852866,9.410788,12.072148,9.825768,7.39762,8.484799,8.532814,6.1046658,2.8705647,3.4913201,3.5187566,5.007198,7.222711,6.636252,9.201583,8.155559,6.5710897,5.164959,2.335549,2.627064,2.3424082,2.4487255,3.6696587,6.4990683,9.9801,10.731179,12.699762,16.921585,21.500084,22.487804,15.577187,9.692014,7.675417,6.2727156,4.0503426,2.5241764,3.117495,4.65395,3.3712845,1.8965619,2.551613,3.093488,3.1312134,4.1189346,2.9974594,2.4795918,2.4658735,2.503599,1.7696671,2.0646117,2.1743584,2.1229146,1.9823016,1.845118,1.9068506,2.095478,2.49331,2.819121,2.4418662,2.428148,2.9117198,3.8274195,4.976331,6.025785,5.5387836,4.8117113,5.055212,5.830299,5.0346346,5.2918534,5.254128,5.442755,5.744559,5.4016004,5.754848,6.228131,6.1904054,5.761707,5.7994323,6.018926,6.584808,6.4579134,5.6348124,5.171818,4.8905916,5.693115,6.2967224,5.885172,4.105216,4.787704,5.425607,5.1512403,4.108646,3.450165,3.875434,4.2218223,4.3109913,4.338428,4.852866,5.0106273,5.381023,5.312431,4.8494368,4.715683,5.0826488,5.4736214,5.267846,4.6127954,4.4413157,4.280125,4.1772375,4.1155047,3.974892,3.525616,3.865145,3.8960114,3.940596,3.8720043,3.1277838,2.5790498,2.3424082,2.2120838,2.1880767,2.4555845,4.201245,4.804852,5.0895076,5.545643,6.3001523,6.8145905,6.4304767,5.336438,4.122364,3.7691166,3.6593697,3.6868064,3.4433057,2.8294096,2.061182,1.4850113,1.2312219,1.097468,0.96371406,0.7922347,0.7579388,0.7579388,0.7682276,0.77851635,0.77851635,1.3032433,2.6785078,4.314421,5.545643,5.6313825,5.641671,5.919468,5.909179,5.40503,4.5613513,4.5613513,5.0655007,6.1149545,7.346176,7.98065,8.687145,8.766026,8.532814,8.251588,8.117833,7.5450926,7.473071,7.442205,7.4524937,7.963502,8.172707,8.021805,7.1678376,6.1904054,6.6053853,6.9963584,7.332458,8.004657,8.498518,7.4010496,8.450503,8.676856,8.621983,8.591117,8.652849,9.421077,10.7586155,11.653738,11.413667,9.644,8.189855,7.936065,8.268735,8.601405,8.4093485,9.115844,9.73317,10.336777,10.744898,10.511685,10.4533825,10.731179,10.381361,9.431366,8.89635,8.786603,7.98065,6.869464,5.693115,4.547633,3.8034124,3.1312134,2.527606,2.1674993,2.411,2.983741,3.199805,3.2546785,3.3232703,3.5564823,3.6525106,3.7142432,3.5976372,3.4021509,3.4638834,3.3541365,3.2615378,2.9940298,2.4898806,1.8313997,1.9171394,1.7730967,1.546744,1.4541451,1.786815,2.5927682,3.4776018,3.7794054,3.4844608,3.2649672,3.9131594,3.8720043,3.6147852,3.8308492,5.4153185,7.6514096,8.06296,7.610255,6.8283086,5.813151,6.5470824,5.967482,5.809721,6.324159,6.2864337,5.857735,5.7239814,6.1904054,6.8797526,6.7459984,0.4664239,0.5144381,0.6859175,0.7956643,0.7476501,0.52472687,0.64819205,0.6790583,0.6379033,0.58645946,0.64819205,0.3566771,0.2469303,0.20234565,0.17490897,0.17147937,0.20920484,0.18862732,0.14404267,0.10288762,0.07545093,0.0548734,0.048014224,0.0548734,0.06516216,0.07545093,0.13375391,0.17147937,0.2469303,0.34638834,0.37382504,0.5590228,0.8676856,1.1694894,1.3512574,1.3203912,1.2998136,1.4164196,1.5707511,1.6393428,1.4644338,1.4918705,1.5398848,1.5158776,1.5604624,2.054323,2.9117198,3.2375305,3.858286,4.7362604,4.945465,5.130663,5.0895076,5.06893,5.0243454,4.623084,5.3158607,6.6533995,7.6857057,8.097256,8.207003,7.3530354,6.81802,6.293293,5.610805,4.7499785,5.2575574,6.4990683,7.829748,8.752307,8.916927,8.347616,8.152129,8.179566,8.543102,9.630281,10.463672,10.655728,10.696883,11.043272,12.116733,11.074138,10.741467,10.714031,10.381361,8.951223,10.912948,11.314209,12.175035,13.498857,13.275933,12.000127,13.245067,14.819247,15.642348,15.745236,15.4742985,14.805529,14.054449,13.241637,12.099585,11.423956,11.105004,10.679735,10.055551,9.517105,9.97667,10.710602,11.211322,11.043272,9.825768,9.3593445,9.884071,10.573419,11.046701,11.379372,12.3533745,12.493987,12.5145645,12.562579,12.2093315,14.157337,15.789821,16.249386,15.951012,16.578627,17.278261,17.343424,17.082775,17.240536,18.975908,19.185112,17.748116,16.691803,16.592344,16.568336,17.772121,17.487467,15.9750185,14.284232,14.270514,14.534592,14.599753,14.479718,14.496866,15.289101,15.63206,14.836395,13.807519,13.094165,12.881531,13.073587,12.891819,12.6586075,12.55229,12.593445,11.941824,11.2250395,10.830637,10.875222,11.214751,11.862943,11.331357,11.043272,11.279913,11.183885,10.597425,10.528833,10.792912,11.214751,11.633161,12.63803,12.987847,12.88496,12.535142,12.130451,12.456262,13.128461,13.567448,13.63604,13.63604,14.177915,14.743796,15.014734,15.076467,15.405707,16.55119,17.37772,17.484037,17.051908,16.818697,16.228807,15.536031,15.340545,15.724659,16.245956,16.184223,15.79325,15.0250225,14.033872,13.183334,12.730629,12.315649,11.777204,11.159878,10.710602,10.768905,10.251037,9.729739,9.462232,9.3764925,9.427936,9.918367,10.251037,10.371073,10.762046,11.094715,10.940384,11.087856,11.489118,11.262765,11.543991,12.30536,12.908967,13.114742,13.070158,13.145609,13.906977,15.055889,16.047039,16.095055,16.067617,16.475739,16.798119,16.88043,16.914726,16.660936,16.115631,15.827546,15.985307,16.420864,17.580065,18.097933,18.811287,19.771572,20.248285,21.489796,22.926792,23.550978,23.406935,23.585274,22.817045,22.69358,21.85676,20.313446,19.46291,17.88873,15.772673,13.810948,13.200482,15.645778,12.288212,11.533703,9.870353,7.116394,6.40304,7.034084,7.208993,5.9160385,3.8891523,3.6182148,2.726522,1.3272504,0.97400284,2.1263442,4.170378,11.413667,7.8263187,10.432805,16.678083,4.417309,9.678296,7.9429245,6.5813785,7.267296,5.967482,7.442205,9.119273,9.270175,8.47451,9.606275,6.351596,6.543653,6.560801,5.4496145,4.914599,5.178677,6.1046658,7.579388,8.433355,6.4579134,8.14527,7.2295704,6.9517736,7.8434668,7.723431,9.057541,8.268735,9.167287,10.655728,6.742569,5.411889,6.1972647,5.219832,2.7128036,3.0111778,1.7765263,5.813151,6.1458206,2.1915064,1.7525192,5.0106273,4.1155047,2.7951138,2.7230926,3.4878905,2.8294096,3.210094,3.7279615,5.960623,13.978998,14.339106,10.065839,6.591667,5.5113473,4.6127954,4.5510626,3.899441,3.6353626,3.9028704,4.029765,3.649081,4.4275975,5.329579,5.6210938,4.8768735,5.0174866,4.839148,4.4516044,3.9303071,3.2821152,3.0489032,2.386993,1.529596,0.7888051,0.5521636,0.64819205,0.84024894,1.0528834,1.2346514,1.3958421,1.3581166,1.5227368,1.7147937,1.7147937,1.255229,1.0117283,1.0117283,1.0048691,1.0597426,1.5776103,1.7319417,2.5070283,3.0797696,3.1552205,2.9665933,3.2409601,3.9028704,4.4927597,5.0243454,5.9983487,3.8685746,2.3252604,2.702515,4.8254294,6.9963584,7.596536,7.9189177,8.134981,8.107545,7.380472,6.451054,5.7239814,5.919468,6.773435,7.0306544,6.0737996,5.7274113,5.909179,6.310441,6.4133286,6.2075534,5.5662203,4.914599,4.588788,4.839148,5.627953,5.73427,5.796003,5.977771,5.967482,5.5490727,5.271276,5.137522,4.98662,4.479041,4.091498,4.1120753,4.016047,3.923448,4.602506,5.0346346,5.2644167,5.3501563,5.4976287,6.0703697,6.5299344,6.759717,6.5813785,6.042933,5.381023,5.768566,5.0620713,4.2938433,4.012617,4.290414,2.7539587,2.3252604,4.396731,7.425057,6.944915,9.184435,9.578837,8.762596,8.628842,12.329367,10.247607,7.671987,7.5553813,8.961512,7.0786686,16.067617,11.283342,6.526505,5.5319247,1.9548649,3.4810312,3.6216443,4.5784993,6.9723516,9.832627,6.9826403,6.848886,9.523964,13.166186,14.006435,16.029892,15.601193,12.984418,9.246168,6.2727156,9.126132,10.124143,7.4353456,2.9871707,2.4555845,2.0920484,2.3321195,2.6990852,3.059192,3.6182148,3.1517909,2.750529,2.486451,2.2738166,1.8931323,2.1263442,2.2223728,2.3732746,2.5550427,2.5310357,2.4555845,2.603057,2.6853669,2.6167753,2.503599,2.8019729,3.5016088,4.2115335,4.928317,6.025785,6.0086374,6.0635104,5.8543057,5.439326,5.2918534,5.4599032,5.4976287,5.5730796,5.778855,6.121814,5.9880595,6.40304,6.1766872,5.4804807,5.857735,6.012067,6.7357097,7.3564653,7.380472,6.5162163,5.669108,5.535354,6.3001523,6.944915,5.24041,5.1512403,5.7377,5.435896,4.2183924,3.5599117,4.3281393,4.90431,5.192395,5.254128,5.3158607,5.3673043,5.717122,5.90232,5.7994323,5.6073756,5.6210938,5.778855,5.703404,5.394741,5.2335505,4.7431192,4.461893,4.3795834,4.331569,3.9886103,4.0846386,4.290414,4.2835546,3.9783216,3.5050385,2.6853669,2.253239,2.0508933,1.9994495,2.1023371,3.2615378,4.712253,5.579939,5.861165,6.4236174,7.0718093,7.0306544,6.310441,5.206114,4.307562,3.7965534,3.8857226,3.9131594,3.5359046,2.719663,1.9308578,1.4095604,1.2380811,1.2415106,1.0014396,1.0425946,0.9877212,0.91227025,0.91569984,1.1317638,1.4335675,2.3218307,3.7039545,4.976331,5.0312047,4.8597255,5.3673043,5.857735,6.0052075,5.857735,5.31929,5.2987127,5.977771,7.034084,7.6376915,8.06296,7.9737906,8.052671,8.388771,8.460793,8.011517,7.8434668,7.6171136,7.5416627,8.368194,8.711152,8.340756,7.363324,6.23156,5.7274113,6.608815,7.298162,7.9943686,8.3922,7.6925645,8.587687,9.3079,9.242738,8.484799,7.8331776,8.330468,8.858624,9.578837,10.100135,9.472521,8.371623,7.4010496,7.455923,8.213862,8.114404,8.433355,9.081548,10.371073,11.862943,12.394529,11.80464,11.135871,10.089847,8.951223,8.577398,8.752307,8.471081,7.7371492,6.7528577,5.9400454,4.804852,3.8308492,2.8294096,2.1640697,2.7402403,2.8054025,2.8019729,2.867135,2.9494452,2.8122618,2.8980014,3.0900583,3.1483612,3.1895163,3.6696587,3.3369887,2.9906003,2.7711067,2.633923,2.3561265,2.1297739,1.6942163,1.3066728,1.1866373,1.5158776,1.920569,2.877424,3.7211025,3.940596,3.2032347,4.057202,4.413879,4.2286816,3.923448,4.3795834,7.747438,9.561689,9.846346,8.958082,7.582818,6.842027,5.7274113,5.305572,5.597087,5.5902276,4.8322887,4.996909,5.892031,6.869464,6.7940125,0.490431,0.45613512,0.48357183,0.5555932,0.5590228,0.29494452,0.33609957,0.35324752,0.34638834,0.32581082,0.29151493,0.14061308,0.10288762,0.106317215,0.10288762,0.082310095,0.08573969,0.06859175,0.05144381,0.044584636,0.037725464,0.030866288,0.05144381,0.07545093,0.11317638,0.20577525,0.274367,0.31895164,0.3841138,0.490431,0.6241849,0.939707,1.1729189,1.3615463,1.471293,1.3958421,1.3238207,1.3341095,1.4232788,1.5055889,1.4232788,1.6256244,1.7147937,1.7765263,1.9480057,2.411,3.333559,3.426158,3.8171308,4.647091,5.07236,5.0003386,4.695105,4.4859004,4.523626,4.787704,5.7377,6.7528577,7.548522,7.966932,7.949784,7.2947326,7.082098,6.7185616,6.0978065,5.6073756,6.090947,6.90033,7.891481,8.680285,8.64942,7.8126,7.421627,7.390761,7.654839,8.1384115,9.009526,9.914937,10.432805,10.899229,12.38767,12.545431,12.586586,11.567999,9.904649,9.39021,10.6488695,10.840926,11.465111,12.363663,11.729189,12.103014,12.847235,13.526293,13.96871,14.270514,14.232788,13.588025,12.922686,12.151029,10.528833,9.314759,8.879202,8.745448,8.611694,8.330468,8.093826,8.47451,8.460793,8.117833,8.591117,8.611694,8.570539,8.954653,9.417647,8.790032,9.554831,9.760606,10.566559,11.976119,12.830087,13.738928,14.743796,15.577187,16.112202,16.369421,17.62122,17.775553,16.87357,15.772673,16.13621,15.614912,15.54632,15.611482,15.450292,14.651197,15.494876,15.645778,15.234227,14.79867,15.29596,14.706071,14.490007,14.603184,14.949572,15.409137,15.004445,14.006435,13.118172,12.768354,13.114742,12.665466,11.948683,11.441104,11.290202,11.30049,11.616013,11.30735,11.197603,11.399949,11.317638,11.550851,11.238758,10.9198065,10.950673,11.4754,10.39165,10.069269,10.155008,10.477389,11.06042,11.852654,12.21619,12.644889,13.018714,12.620882,12.46998,13.371962,14.260224,14.634049,14.565458,15.018164,15.323397,15.395418,15.247946,15.001016,15.326826,16.187653,16.328266,15.71437,15.515453,15.529172,15.563468,15.662926,15.71094,15.440002,15.481158,15.388559,15.148488,14.815818,14.496866,13.677195,13.046151,12.363663,11.612583,11.002116,10.563129,10.007536,9.530824,9.301042,9.47938,9.15014,9.019815,9.126132,9.527394,10.316199,10.604284,10.854645,11.4033785,11.976119,11.701753,11.931535,12.418536,12.878101,13.231348,13.601744,13.762935,14.2362175,15.0078745,15.755525,15.854982,15.762384,16.112202,16.37628,16.414005,16.475739,16.516893,15.841265,15.580616,15.999025,16.486027,17.336565,17.820137,18.722118,20.066517,21.095392,22.868488,23.427511,23.832203,24.401514,24.710178,23.520111,23.142857,21.915064,19.9602,19.178253,17.53891,16.695232,16.527182,15.560039,10.9369545,11.276484,9.026674,7.205563,7.438775,9.952662,9.187865,8.1487,7.5245147,7.346176,6.975781,2.8911421,1.5638919,2.085189,6.1766872,18.20768,17.610931,13.697772,15.1862135,18.269413,6.608815,10.710602,7.623973,6.852316,9.496528,8.2481575,9.256456,9.002667,7.963502,7.1712675,8.224151,5.120374,6.7700057,7.507367,6.0806584,5.6793966,5.336438,6.7940125,8.450503,8.80718,6.495639,8.477941,7.582818,7.4456344,8.416207,7.5450926,8.40249,7.517656,8.279024,9.455373,5.2026844,4.139512,4.3487167,3.6147852,2.085189,2.2600982,6.461343,6.893471,4.4756117,1.6393428,2.3286898,2.6887965,4.8151407,5.171818,3.5153272,2.9117198,3.6353626,3.74168,4.0709205,6.427047,13.588025,11.701753,9.054111,6.8900414,5.3741636,3.5942078,3.1620796,3.1209247,3.1140654,3.117495,3.426158,4.2183924,4.400161,4.5270553,4.537344,3.7794054,4.184097,4.338428,4.184097,3.758828,3.1860867,2.5893385,1.978872,1.2929544,0.7339317,0.7682276,0.8162418,0.94656616,1.0768905,1.214074,1.4610043,1.5090185,1.5776103,1.8965619,2.2566686,1.9925903,1.2689474,1.1283343,1.1866373,1.4164196,2.1263442,2.5893385,3.2821152,3.5804894,3.2649672,2.5413244,2.9665933,3.5599117,3.998899,4.331569,4.9523244,3.789694,3.3678548,4.07435,5.5422134,6.680836,7.3598948,7.8674736,8.303031,8.275595,6.8969,6.3447366,5.9640527,6.1458206,6.7528577,7.1061053,6.917478,6.6739774,6.8043017,7.3290286,7.870903,7.407909,6.759717,6.2487082,6.0326443,6.121814,6.625963,6.7219915,6.9037595,7.1781263,7.0718093,6.691125,6.3001523,5.98463,5.693115,5.219832,5.5422134,5.669108,5.271276,4.705394,5.0003386,5.535354,5.9160385,6.001778,5.857735,5.7479887,6.0978065,6.526505,6.725421,6.4887795,5.7308407,6.4133286,6.2247014,5.4633327,4.756838,5.0346346,4.2938433,3.457024,3.433017,4.2286816,4.9523244,9.705732,12.233338,12.562579,12.30536,14.685493,9.685155,7.3118806,6.975781,8.285883,11.050131,14.116182,9.877212,6.3001523,5.3158607,2.8225505,3.3712845,3.1620796,3.5770597,5.7411294,10.528833,8.110974,7.3290286,10.47396,14.147048,9.273604,14.990726,13.495427,10.587136,8.597976,6.39961,9.098696,9.547972,6.807731,3.1655092,4.149801,3.223812,3.4192986,3.3609958,2.6647894,1.9754424,2.7162333,2.3561265,1.8759843,1.7559488,1.9685832,2.452155,2.2360911,1.8725548,1.8039631,2.3629858,2.0406046,2.3389788,2.620205,2.7470996,3.0866287,3.74168,4.2286816,4.763697,5.3261495,5.6519604,5.9914894,6.392751,6.4064693,6.0086374,5.610805,5.926327,5.919468,6.101236,6.5470824,6.9071894,6.56766,6.831738,6.7219915,6.121814,5.7754254,5.586798,6.492209,7.250148,7.233,6.420188,6.451054,6.108095,6.4304767,7.040943,6.1561093,5.874883,6.138962,5.926327,5.103226,4.400161,4.7191124,5.288424,5.895461,6.4373355,6.914048,6.574519,6.5024977,6.444195,6.307011,6.159539,6.4373355,6.910619,6.8214493,6.1458206,5.6073756,5.7068334,5.675967,5.6039457,5.4976287,5.267846,5.0757895,5.086078,5.0174866,4.7808447,4.48933,3.6936657,2.9082901,2.3218307,1.9891608,1.821111,2.6304936,4.245829,5.6348124,6.4304767,6.948344,7.8434668,8.604835,7.466212,4.911169,3.6627994,3.673088,4.214963,4.5819287,4.482471,4.0091877,3.0351849,2.0886188,1.529596,1.3924125,1.3649758,1.4404267,1.4918705,1.3786942,1.2483698,1.5227368,1.670209,2.1023371,2.9665933,3.9646032,4.341858,3.940596,4.3795834,5.0895076,5.693115,5.9983487,5.970912,6.0532217,6.416758,7.016936,7.606825,7.7920227,7.740579,7.8331776,8.114404,8.289313,8.179566,7.874333,7.4936485,7.4524937,8.450503,8.632272,7.939495,7.2158523,6.697984,6.0395036,6.7631464,7.0615206,7.6445503,8.47451,8.783174,8.985519,8.985519,8.97866,8.766026,7.7680154,8.333898,8.320179,8.515666,9.102125,9.668007,9.424506,8.268735,7.64798,8.056101,9.030104,9.654288,10.573419,11.835506,13.073587,13.485138,12.435684,11.396519,10.14129,8.923786,8.453933,8.471081,8.292743,7.98408,7.658269,7.4765005,6.1046658,4.619654,3.333559,2.5310357,2.4658735,2.5447538,2.6545007,2.6167753,2.428148,2.2841053,2.2978237,2.386993,2.6064866,2.9391565,3.2821152,3.333559,2.9631636,2.7745364,2.884283,2.935727,2.5138876,1.9171394,1.3924125,1.1317638,1.2860953,1.471293,2.0920484,3.0489032,3.724532,2.9974594,3.9063,4.880303,5.288424,4.955754,4.173808,6.5127864,8.083538,8.923786,9.167287,9.043822,7.160979,5.6348124,4.852866,4.705394,4.57507,4.280125,4.4584637,5.1238036,6.0052075,6.56766,0.4424168,0.32924038,0.26064864,0.26750782,0.2777966,0.106317215,0.09602845,0.08916927,0.10288762,0.1097468,0.041155048,0.0274367,0.037725464,0.0548734,0.058302987,0.041155048,0.037725464,0.030866288,0.0274367,0.0274367,0.030866288,0.044584636,0.08573969,0.14061308,0.2194936,0.3806842,0.4389872,0.47328308,0.53501564,0.64819205,0.84024894,1.1523414,1.3581166,1.4918705,1.546744,1.4610043,1.371835,1.2792361,1.2929544,1.3924125,1.4541451,1.7490896,1.920569,2.1194851,2.411,2.784825,3.7451096,3.8342788,4.0091877,4.5030484,4.835718,4.722542,4.3624353,4.262977,4.5613513,5.0620713,6.077229,6.5367937,6.8969,7.157549,6.8866115,6.8454566,6.742569,6.4304767,6.0635104,6.1321025,6.691125,7.2124224,8.080108,8.999237,8.988949,8.193284,7.4181976,7.023795,7.0615206,7.284444,8.186425,9.263316,9.849775,10.127572,11.122152,12.253916,12.80608,11.934964,10.5597,11.348505,10.823778,10.909517,11.7086115,12.47341,11.588576,12.487128,12.298501,12.075578,12.233338,12.566009,12.329367,11.880091,11.375941,10.63858,9.167287,7.8777623,7.2021337,7.010077,7.023795,6.835168,6.1732574,6.0703697,5.950334,5.9743414,7.06495,7.2295704,7.267296,7.870903,8.56025,7.6651278,8.207003,8.694004,9.908078,11.742908,13.190193,13.320518,13.4474125,14.037301,14.726648,14.318527,15.8138275,16.269962,15.676644,14.490007,13.642899,12.905538,13.46799,13.906977,13.697772,13.210771,14.764374,15.563468,15.374841,14.836395,15.446862,15.326826,14.668345,14.400838,14.616901,14.572317,14.325387,13.776653,13.313659,13.118172,13.149038,12.504276,11.910957,11.478829,11.14273,10.690024,11.273054,11.204462,11.345076,11.739478,11.609154,11.214751,11.146159,10.947243,10.799771,11.523414,10.978109,10.583707,10.4533825,10.604284,10.991828,11.211322,11.465111,12.109874,12.895248,12.9707,13.049581,13.858963,14.603184,14.977009,15.189643,15.529172,15.621771,15.566897,15.391989,15.031882,14.88441,15.580616,15.618341,14.856973,14.514014,14.568888,14.956431,15.350834,15.450292,14.973578,14.832966,14.712931,14.627191,14.644339,14.887839,14.188204,13.395968,12.586586,11.790922,10.988399,10.052121,9.692014,9.421077,9.277034,9.825768,9.496528,8.862054,8.594546,8.913498,9.599416,9.788043,10.343636,11.14273,11.897239,12.175035,12.734058,13.035862,13.262215,13.54687,13.978998,14.400838,14.870691,15.316538,15.731518,16.163645,16.112202,16.167076,16.235666,16.300829,16.434584,16.462019,15.834405,15.587475,16.005884,16.61292,17.730967,18.21111,19.106232,20.683842,22.456938,23.897366,24.0174,24.43581,25.20061,24.789059,24.17859,23.544119,21.85333,19.589804,18.766703,17.20967,16.300829,15.014734,12.8197975,9.6988735,12.493987,8.64599,5.9812007,7.267296,10.216741,8.495089,6.694555,6.680836,7.8983397,7.366754,4.650521,3.1860867,3.8445675,9.156999,23.300617,17.508043,16.486027,16.47231,14.544881,8.635701,12.425395,7.2192817,5.9160385,9.637141,7.73029,8.073249,6.8591747,5.90232,5.8645945,6.276145,4.5442033,6.8797526,7.490219,5.960623,7.2432885,5.658819,6.8969,8.285883,8.347616,6.773435,8.224151,7.414768,7.8674736,9.225591,7.257007,7.7611566,7.332458,7.4936485,7.610255,4.8905916,3.8308492,3.1895163,2.6236343,2.1400626,2.095478,9.362774,7.301592,3.5702004,2.1091962,3.1517909,2.2978237,4.5682106,5.147811,3.5942078,3.8342788,4.32128,3.5702004,3.9131594,6.451054,11.06042,8.124693,7.466212,6.81802,5.096367,2.4041407,2.0097382,2.633923,2.8499873,2.5721905,3.0489032,4.1463714,3.9543142,3.6079261,3.5187566,3.3747141,3.765687,4.184097,4.2286816,3.8857226,3.532475,2.7230926,1.9274281,1.2689474,0.91569984,1.0940384,1.0082988,1.1283343,1.2209331,1.2380811,1.3409687,1.4953002,1.5193073,1.8759843,2.4418662,2.510458,1.6839274,1.4644338,1.4747226,1.7353712,2.6990852,3.0386145,3.3609958,3.316411,2.9322972,2.609916,3.357566,3.82399,4.0674906,4.170378,4.2389703,4.461893,4.5270553,4.729401,5.329579,6.5710897,7.0546613,8.056101,8.841476,8.663138,6.7631464,6.3961806,6.183546,6.200694,6.351596,6.3721733,6.866034,6.9963584,7.257007,7.829748,8.567109,8.289313,7.73372,7.3598948,7.2604365,7.14726,7.5862474,7.582818,7.548522,7.599966,7.56567,7.2638664,6.948344,6.6568294,6.2864337,5.5833683,5.8371577,6.2555676,6.094377,5.4941993,5.4907694,5.8062916,6.166398,6.334448,6.2075534,5.8234396,5.857735,6.1561093,6.5539417,6.783724,6.464772,6.4579134,6.6465406,6.39961,5.7891436,5.6039457,5.5113473,4.7842746,3.789694,3.223812,4.1120753,8.7145815,12.583157,13.327377,11.609154,11.170166,9.510246,8.779744,8.762596,9.644,11.996697,9.949233,7.514226,5.7994323,4.911169,3.9474552,3.2615378,2.411,2.2258022,3.7348208,8.186425,9.493098,8.721441,11.492548,14.918706,7.589677,12.782072,10.7757635,8.076678,7.7577267,9.455373,9.661148,8.64256,7.058091,5.9914894,6.944915,3.9714622,3.4707425,3.0386145,1.920569,1.039165,1.7422304,1.4575747,2.620205,4.1155047,1.2655178,1.9891608,2.0406046,1.5776103,1.2106444,2.0028791,1.6496316,2.0097382,2.3904223,2.603057,2.976882,3.8479972,4.1943855,4.7534084,5.48734,5.579939,5.892031,6.2384195,6.468202,6.4133286,5.8680243,5.9914894,5.953764,6.3378778,7.0923867,7.5107965,7.0272245,7.0032177,7.160979,7.0615206,6.1046658,5.3398676,5.9640527,6.543653,6.495639,6.090947,7.130112,7.2432885,7.1712675,7.085528,6.5882373,6.15268,6.125243,6.159539,5.9160385,5.0895076,4.698535,5.1409516,6.077229,7.1232533,7.8606143,7.233,6.7391396,6.5024977,6.495639,6.5539417,6.807731,7.3393173,7.257007,6.543653,6.0532217,6.56766,6.81802,6.8763227,6.790583,6.5779486,6.0703697,5.751418,5.518206,5.2472687,4.7945633,4.0846386,3.309552,2.651071,2.2223728,2.0406046,2.503599,3.6285036,5.096367,6.4716315,7.2124224,8.488229,8.357904,6.375603,3.673088,2.9665933,3.4467354,4.0537724,4.5784993,4.9591837,5.2747054,4.636802,3.525616,2.4967396,1.8554068,1.6770682,1.7353712,2.0028791,2.1091962,2.0131679,2.0097382,1.9925903,2.0440342,2.2841053,2.8054025,3.683377,3.3747141,3.566771,4.2389703,5.147811,5.830299,6.3378778,6.9071894,7.1987042,7.346176,7.963502,8.014946,7.9463544,7.932636,8.080108,8.4093485,8.258447,7.8331776,7.548522,7.764586,8.766026,8.844906,8.258447,7.5759587,7.016936,6.4373355,6.783724,7.0889573,7.654839,8.512236,9.386781,9.537683,9.006097,8.930646,9.122703,8.097256,8.275595,8.152129,8.182996,8.611694,9.472521,9.56512,8.848335,8.464222,9.050681,10.7586155,11.8869505,12.775213,13.395968,13.670336,13.46799,12.6757555,11.677745,10.467101,9.31133,8.735159,8.639131,8.3922,8.169277,8.141841,8.477941,7.2707253,5.363875,3.7142432,2.7470996,2.3424082,2.5721905,2.6167753,2.3904223,2.0474637,1.9857311,1.9582944,2.0440342,2.2978237,2.6716487,2.9974594,3.3541365,3.1483612,3.0866287,3.3472774,3.5839188,3.059192,2.4967396,1.8897027,1.3992717,1.3649758,1.4850113,1.8073926,2.568761,3.309552,2.9048605,3.7176728,4.897451,5.7651367,5.861165,4.938606,5.5319247,5.9812007,6.560801,7.500508,8.98209,8.001227,6.4133286,5.1066556,4.3692946,3.9097297,3.9028704,4.2355404,4.7808447,5.470192,6.2864337,0.22292319,0.14061308,0.11317638,0.09945804,0.07545093,0.0548734,0.058302987,0.041155048,0.037725464,0.044584636,0.0274367,0.017147938,0.0274367,0.041155048,0.041155048,0.030866288,0.041155048,0.048014224,0.05144381,0.058302987,0.06859175,0.12689474,0.1920569,0.2709374,0.37725464,0.52472687,0.5624523,0.59331864,0.6824879,0.83338976,0.99801,1.2312219,1.4850113,1.6256244,1.6153357,1.5227368,1.4369972,1.3203912,1.2826657,1.3752645,1.5638919,1.903421,2.085189,2.3732746,2.784825,3.07634,3.9646032,4.2938433,4.461893,4.5339146,4.232111,4.214963,4.057202,4.3521466,5.0757895,5.5593615,6.090947,6.1972647,6.210983,6.159539,5.73427,6.2384195,6.0566516,5.754848,5.7308407,6.186976,6.9037595,7.599966,8.594546,9.585697,9.661148,9.283894,8.261876,7.366754,7.0546613,7.4456344,8.080108,8.488229,8.676856,8.80718,9.187865,10.329918,10.947243,11.22161,11.585147,12.71691,10.964391,10.899229,12.024134,13.121602,12.267634,12.257345,11.561139,11.026124,10.88551,10.772334,10.175586,9.952662,9.427936,8.498518,7.6205435,6.9209075,6.121814,5.5079174,5.099797,4.650521,4.290414,4.173808,4.4927597,5.120374,5.6073756,5.645101,6.046363,6.835168,7.5759587,7.349606,7.81603,8.796892,10.038403,11.255906,12.106443,11.595435,11.187314,11.581717,12.38767,12.123591,13.203912,13.745787,13.924125,13.701202,12.836946,12.593445,12.6586075,12.507706,12.284782,12.782072,15.446862,16.973028,16.115631,14.064738,14.424845,15.909856,15.134769,14.212211,13.954991,13.862392,14.4145565,14.479718,14.273943,13.80066,12.840376,12.408247,12.535142,12.545431,12.140739,11.396519,11.509696,11.286773,11.4033785,11.907528,12.21619,11.458252,11.297061,11.032983,10.738038,11.252477,11.89038,11.701753,11.461681,11.427385,11.355364,11.029553,11.201033,11.732618,12.401388,12.902108,13.536582,14.006435,14.174485,14.315098,15.127911,15.488017,15.450292,15.2033615,14.932424,14.79524,15.028452,15.518884,15.278812,14.4145565,14.123041,13.978998,14.088745,14.38026,14.675205,14.682064,14.5585985,14.476289,14.246507,14.023583,14.308239,13.9481325,13.183334,12.47341,11.869802,10.998687,9.832627,9.678296,9.537683,9.345626,9.993818,9.983529,9.294182,8.772884,8.745448,9.023245,9.266746,9.81205,10.47396,11.211322,12.092726,13.008426,13.505715,13.790371,14.006435,14.225929,14.685493,15.29253,15.635489,15.865272,16.719238,16.87357,16.671225,16.516893,16.595774,16.859852,16.767254,16.287111,15.9613,16.115631,16.849564,18.362011,19.061647,19.991066,21.496655,23.225166,24.216316,25.02227,25.649885,25.701328,24.36036,24.672453,23.725885,21.880768,19.826445,18.584934,16.71238,13.790371,10.508256,9.342196,14.54831,14.79867,10.563129,7.905199,7.6514096,5.4016004,4.355576,3.1517909,2.942586,3.5942078,3.6799474,5.8645945,4.822,5.3570156,9.496528,16.486027,11.149589,14.572317,14.068168,8.930646,10.419086,11.629731,5.7102633,4.355576,7.5931067,3.7691166,4.5613513,4.1463714,4.32471,5.161529,4.9660425,4.8494368,6.560801,6.464772,5.453044,8.968371,6.159539,6.9037595,7.6925645,7.421627,7.363324,7.750868,7.0443726,8.032094,9.688584,7.1712675,7.2604365,7.582818,7.4456344,6.6122446,5.3158607,3.899441,3.1449318,2.9082901,2.9460156,2.9048605,9.002667,6.3961806,3.5187566,3.3884325,3.5839188,3.093488,3.2306714,3.1792276,3.3815732,5.521636,4.972902,3.292404,3.1106358,5.144381,8.193284,5.8165803,7.0135064,7.500508,5.5490727,1.9925903,1.3992717,1.9720128,2.411,2.4555845,2.9048605,3.350707,3.5016088,3.3472774,3.2272418,3.8377085,3.8960114,4.479041,4.547633,4.081209,4.081209,3.3438478,2.5138876,1.862266,1.546744,1.6016173,1.3409687,1.430138,1.5124481,1.4404267,1.2860953,1.4575747,1.471293,1.762808,2.3218307,2.6750782,2.1503513,1.9514352,1.8142518,1.978872,3.2066643,3.0214665,2.959734,2.9220085,2.9940298,3.4638834,4.4721823,4.7362604,4.7431192,4.7499785,4.7842746,5.007198,4.976331,4.712253,4.9248877,7.010077,7.2878733,8.498518,9.31133,8.995808,7.4044795,6.9654922,6.447624,6.210983,6.1458206,5.6656785,6.23156,6.7185616,7.239859,7.8503256,8.543102,8.769455,8.31675,7.9600725,7.8606143,7.5725293,8.193284,8.193284,7.8503256,7.5279446,7.671987,7.459353,7.3255987,7.281014,7.058091,6.108095,5.453044,5.892031,6.0978065,5.7925735,5.761707,5.521636,5.6793966,5.9160385,6.018926,5.888602,5.885172,5.8062916,5.9812007,6.4544835,6.9963584,6.245279,6.3790326,6.6705475,6.632822,6.025785,6.1561093,5.3158607,4.437886,4.125794,4.6436615,6.4064693,9.832627,10.1481495,7.363324,6.2898636,11.828648,12.356804,12.555719,12.905538,9.695444,8.056101,6.725421,5.826869,5.2266912,4.530485,3.4364467,2.1229146,2.0817597,3.4055803,4.8151407,10.659158,9.139851,9.9869585,12.874671,7.4113383,7.781734,7.750868,6.944915,7.284444,12.9809885,12.322508,10.734609,9.757176,9.942374,10.847785,4.9660425,2.8637056,2.1332035,1.5776103,1.2312219,0.9774324,0.69963586,3.6216443,6.6225333,0.22978236,0.89169276,1.5536032,1.5570327,1.2277923,1.8588364,1.6221949,1.8999915,2.2155135,2.3835633,2.503599,3.0729103,3.4947495,4.3452873,5.4770513,6.0052075,5.9228973,5.9160385,6.0566516,6.1629686,5.785714,5.5250654,5.5833683,6.111525,6.927767,7.5416627,7.1541195,7.016936,7.373613,7.723431,6.8454566,5.6656785,5.576509,5.8062916,5.9331865,5.885172,7.2295704,7.9909387,7.936065,7.257007,6.601956,5.9160385,5.7582774,6.0326443,6.200694,5.305572,4.602506,4.9488945,5.970912,7.133542,7.750868,7.239859,6.632822,6.427047,6.6431108,6.8283086,6.6636887,6.924337,6.9346256,6.6396813,6.615674,7.0375133,7.4044795,7.6445503,7.6857057,7.442205,6.8591747,6.351596,5.878313,5.3261495,4.537344,3.8102717,3.3301294,2.9220085,2.5893385,2.5070283,2.6956558,3.1792276,4.331569,5.874883,6.8591747,8.405919,6.56766,3.9131594,2.301253,2.867135,3.4192986,3.6456516,4.07435,4.870014,5.8165803,6.1046658,5.411889,4.232111,3.0386145,2.2635276,2.16064,2.469303,2.843128,2.9460156,2.4452958,2.2841053,2.0989075,1.8485477,1.879414,2.9254382,3.1380725,3.2135234,3.724532,4.7019644,5.6313825,6.2418494,7.2775846,7.7131424,7.654839,8.337327,8.505377,8.381912,8.268735,8.381912,8.841476,8.488229,8.107545,8.14527,8.707723,9.561689,9.921797,9.849775,8.838047,7.31531,6.636252,6.540223,7.3427467,8.107545,8.580828,9.194724,9.911508,9.592556,9.328478,9.225591,8.4264965,8.080108,8.100685,8.375052,8.738589,8.98209,8.766026,8.7283,9.270175,10.443094,11.952112,13.443983,13.776653,13.509145,13.066729,12.744347,12.651748,11.849225,10.844356,10.000677,9.527394,9.414218,9.006097,8.498518,8.213862,8.615124,7.7920227,5.7274113,3.7382503,2.6167753,2.620205,2.8911421,2.6785078,2.3218307,2.0406046,1.920569,1.8965619,2.07833,2.294394,2.5447538,3.0214665,3.3061223,3.3712845,3.532475,3.8479972,4.1120753,3.6044965,3.223812,2.6407824,1.961724,1.7079345,1.903421,2.07833,2.510458,3.0420442,3.083199,3.649081,4.554492,5.4770513,6.0978065,6.118384,5.5902276,4.8768735,4.5099077,5.07236,7.2295704,8.443645,7.291303,5.6965446,4.530485,3.6079261,3.4604537,4.108646,4.8254294,5.3501563,5.8817425,0.07545093,0.05144381,0.0548734,0.0548734,0.041155048,0.030866288,0.09259886,0.061732575,0.017147938,0.0034295875,0.01371835,0.01371835,0.041155048,0.0548734,0.041155048,0.030866288,0.041155048,0.06516216,0.082310095,0.12003556,0.22978236,0.36353627,0.432128,0.48700142,0.53844523,0.548734,0.59674823,0.6756287,0.8196714,1.0357354,1.2655178,1.646202,1.8759843,1.845118,1.6324836,1.5090185,1.4747226,1.3443983,1.2655178,1.3958421,1.9068506,2.4795918,2.5138876,2.7402403,3.210094,3.2958336,3.8342788,4.2526884,4.605936,4.636802,3.7691166,3.782835,4.214963,5.0449233,5.926327,6.193835,5.535354,5.6656785,5.377593,4.636802,4.5613513,5.4770513,5.7719955,5.977771,6.3207297,6.697984,7.455923,8.467651,9.091836,9.15014,8.940934,9.441654,8.879202,7.8606143,7.0786686,7.3255987,6.824879,6.3035817,6.2487082,6.8214493,7.857185,8.934075,9.321619,10.010965,11.008976,11.338216,11.653738,11.046701,11.094715,11.780633,11.4754,12.109874,11.653738,10.556271,9.112414,7.4765005,7.3290286,7.723431,7.4010496,6.2658563,5.3878818,5.2026844,4.6093655,4.0606318,3.7485392,3.6010668,3.649081,4.1189346,4.5956473,4.897451,5.0826488,4.9351764,5.3090014,5.8234396,6.5539417,8.056101,7.4696417,7.414768,8.110974,9.091836,9.201583,7.5279446,7.7611566,9.73317,12.271064,13.200482,12.734058,12.041282,11.955542,12.627741,13.519434,13.481709,13.694343,13.7526455,13.646329,13.732068,15.05246,16.37971,16.177364,14.695783,13.96185,15.426285,15.217079,14.490007,14.225929,15.227368,14.973578,14.421415,14.057879,13.900118,13.533153,12.397959,12.562579,12.644889,12.336226,12.421966,12.651748,12.068718,11.941824,12.421966,12.55915,12.7272,12.212761,11.530273,11.043272,10.971251,11.567999,11.818358,11.684605,11.2593355,10.7586155,10.244178,10.693454,11.736049,12.744347,12.816368,13.011855,13.227919,13.176475,13.173045,14.112752,14.503725,14.647768,14.496866,14.232788,14.280802,14.819247,15.090185,14.500296,13.488567,13.5503,13.903547,14.064738,14.109323,14.04759,13.838386,14.500296,14.582606,14.428274,14.160767,13.670336,12.706621,11.907528,11.664027,11.814929,11.657167,11.094715,11.029553,10.607714,9.873782,9.750318,9.993818,9.331907,8.940934,9.098696,9.170717,9.709162,10.271614,10.590566,10.734609,11.1393,11.96926,13.073587,14.037301,14.654627,14.922135,15.055889,15.227368,15.247946,15.415996,16.523752,16.79469,16.942162,17.082775,17.264544,17.470318,17.446312,17.130789,16.87357,16.983316,17.71382,18.351723,19.1954,20.526081,21.942501,22.36777,24.36036,25.917393,26.157463,25.300066,24.6896,24.60386,23.557837,22.645567,21.599543,18.766703,15.265094,12.109874,15.138199,21.321745,18.78385,11.924676,8.752307,9.89436,11.602294,5.768566,3.2649672,1.8897027,1.3889829,1.371835,1.313532,3.4364467,3.7211025,4.73969,7.5245147,11.567999,10.820349,13.756075,13.2862215,9.870353,11.506266,3.6936657,2.5653315,5.3158607,7.6376915,3.707384,7.0889573,6.324159,4.8837323,4.355576,4.4413157,5.0757895,6.0395036,6.210983,6.540223,10.055551,6.550512,7.6342616,7.9772205,6.7665763,7.706283,8.131552,7.2878733,7.7577267,9.050681,7.599966,5.693115,5.6210938,5.785714,5.0346346,2.6545007,2.8019729,3.1312134,3.7348208,4.187526,3.5393343,9.119273,5.936616,4.1360826,5.4736214,3.3266997,3.1312134,2.9460156,3.7451096,4.7774153,3.5564823,5.751418,4.214963,2.6716487,3.1517909,5.9983487,5.1409516,8.985519,9.873782,6.0566516,1.6633499,0.89512235,1.196926,1.8691251,2.5378947,3.1723683,3.210094,4.1429415,4.3452873,3.7622573,3.9200184,3.981751,4.4447455,4.3487167,3.8617156,4.2869844,3.724532,3.6593697,3.2615378,2.5550427,2.3972816,2.0165975,1.9308578,1.9754424,2.0063086,1.9068506,1.9445761,1.8348293,1.9308578,2.2841053,2.6407824,2.3458378,2.1743584,2.0680413,2.2909644,3.4021509,3.059192,2.867135,3.549623,4.647091,4.4996185,4.856296,4.897451,4.835718,4.846007,5.0655007,5.346727,5.638242,5.857735,5.9469047,5.874883,7.706283,8.080108,8.220721,8.453933,8.210432,7.4765005,6.6431108,6.1732574,6.090947,5.9812007,6.2247014,6.625963,7.0889573,7.6376915,8.405919,8.858624,8.515666,8.189855,8.045813,7.582818,7.7680154,7.949784,7.870903,7.5862474,7.4765005,7.829748,7.874333,8.093826,8.364764,7.949784,7.267296,6.8111606,6.444195,6.15268,6.042933,5.579939,5.857735,6.0806584,5.950334,5.645101,6.012067,5.6828265,5.3090014,5.3501563,6.0566516,6.0086374,5.813151,6.3138704,7.06495,6.3310184,6.492209,6.5230756,6.0395036,5.6073756,6.742569,3.4364467,6.262427,7.8126,6.7528577,7.8263187,13.162757,12.260776,12.127021,13.38225,10.268185,10.816919,9.016385,8.086967,7.706283,3.981751,3.532475,2.3664153,3.4707425,5.9126086,4.852866,14.544881,8.279024,4.8254294,7.7440085,5.3878818,3.3712845,3.5359046,4.5853586,6.245279,9.246168,14.3974085,14.651197,12.233338,11.190743,17.37772,8.759167,4.7019644,3.4810312,3.1483612,1.5261664,1.8691251,1.2037852,0.70306545,0.65505123,0.47328308,0.51100856,0.764798,0.9842916,1.2723769,2.0920484,1.6393428,1.8554068,2.4418662,3.100347,3.5393343,2.7333813,3.2272418,4.6093655,6.1149545,6.6533995,6.090947,5.610805,5.442755,5.4084597,4.945465,4.955754,5.360445,5.7479887,6.025785,6.4544835,7.0032177,7.5725293,7.7611566,7.5759587,7.431916,6.759717,6.0532217,5.7582774,5.751418,5.3261495,5.888602,6.6225333,7.06838,7.0272245,6.5779486,5.830299,5.65539,5.8200097,5.90575,5.295283,5.4770513,5.9160385,6.385892,6.8728933,7.5690994,7.798882,7.582818,7.3564653,7.205563,6.852316,6.5710897,6.910619,7.058091,6.8728933,6.8969,7.1541195,7.455923,7.7131424,7.822889,7.675417,7.7851634,7.548522,6.8763227,5.953764,5.2335505,4.280125,3.724532,3.2786856,2.7985435,2.2738166,2.6407824,3.3369887,4.245829,5.1752477,5.861165,7.0443726,6.5779486,4.273266,1.9651536,3.5393343,4.040054,4.1017866,4.3041325,4.7191124,4.914599,6.355026,6.842027,6.420188,5.329579,3.998899,3.3747141,3.0351849,3.1277838,3.2512488,2.4555845,2.3458378,2.136633,1.8554068,1.6324836,1.6942163,2.7059445,3.2889743,3.765687,4.3349986,5.0826488,5.5079174,6.392751,6.9380555,7.164408,7.936065,8.680285,8.766026,8.618553,8.56025,8.803751,9.132992,9.225591,9.541112,10.158438,10.7586155,12.075578,12.404818,10.933525,8.419638,7.1884155,6.4544835,7.298162,8.436785,9.071259,8.865483,9.561689,9.89093,9.517105,8.707723,8.31675,8.7317295,8.64256,8.934075,9.482809,9.139851,8.748878,8.762596,9.177576,9.815479,10.316199,11.814929,11.156448,10.432805,10.789482,12.452832,12.281353,11.451392,10.875222,10.81006,10.834066,10.405369,9.657719,8.827758,8.162418,7.9189177,7.0786686,5.1821065,3.2718265,2.2806756,3.0351849,3.1106358,2.9734523,2.8122618,2.603057,2.0920484,2.0165975,2.1091962,2.4247184,2.8499873,3.083199,2.9974594,3.3061223,3.6696587,3.9440255,4.149801,3.8445675,3.6044965,3.2135234,2.6236343,1.9514352,2.3801336,2.3218307,2.534465,3.1312134,3.5702004,3.765687,4.420738,5.0655007,5.641671,6.48535,6.667118,5.6519604,4.540774,4.081209,4.65395,6.1801167,5.994919,5.2506986,4.3624353,3.0214665,2.7779658,3.5393343,4.273266,4.636802,4.99005,0.041155048,0.034295876,0.06516216,0.08573969,0.07888051,0.06859175,0.041155048,0.030866288,0.048014224,0.06859175,0.05144381,0.024007112,0.0274367,0.041155048,0.05144381,0.07888051,0.12003556,0.16462019,0.22635277,0.33266997,0.51100856,0.5453044,0.6207553,0.6756287,0.6893471,0.67219913,0.72021335,0.8128122,0.99801,1.2655178,1.5364552,2.1091962,2.3252604,2.2292318,1.99602,1.9137098,1.5947582,1.4678634,1.5364552,1.8279701,2.4075704,3.0111778,3.1243541,3.1895163,3.4295874,3.858286,4.2286816,5.051782,5.5079174,5.284994,4.57507,4.0194764,4.290414,4.7671266,5.212973,5.754848,6.228131,6.6053853,6.574519,6.2418494,6.101236,5.8817425,5.562791,5.521636,5.7719955,5.953764,7.414768,8.742019,9.22216,9.0369625,9.259886,9.829198,8.711152,7.2638664,6.5024977,7.130112,6.7459984,6.4407654,6.1904054,6.2384195,7.1026754,8.450503,9.050681,9.551401,10.134431,10.532263,10.525404,9.866923,9.146709,8.786603,9.057541,9.078118,8.755736,7.6514096,6.2555676,5.9743414,5.4976287,5.3330083,4.99005,4.4927597,4.386442,3.7725463,3.7382503,3.5599117,3.2615378,3.6147852,3.673088,3.8960114,4.0777793,4.1429415,4.1292233,4.4996185,4.57164,4.7328305,4.98662,4.945465,4.4859004,4.4687524,4.7259717,5.130663,5.6005163,6.1732574,7.2295704,8.40249,9.482809,10.439664,10.240748,9.541112,9.551401,10.374502,10.991828,10.779194,11.561139,12.926115,14.112752,14.013294,14.757515,15.018164,14.781522,14.424845,14.706071,15.028452,15.453721,15.536031,15.608052,16.815268,15.611482,14.658057,14.335675,14.407697,14.009865,13.87954,13.104454,12.1921835,11.509696,11.273054,11.670886,11.856084,11.859513,12.048141,13.118172,13.728639,13.104454,12.161317,11.399949,10.88551,10.9369545,11.2250395,11.616013,11.770344,11.173596,11.578287,11.451392,11.595435,12.089295,12.281353,12.229909,12.106443,11.931535,11.842365,12.089295,13.13189,13.704632,13.937843,14.027013,14.232788,14.116182,14.064738,13.7526455,13.179905,12.634601,12.782072,13.282792,13.533153,13.437123,13.375391,13.858963,13.831526,13.519434,12.953552,11.986408,10.621432,10.213311,10.168727,10.110424,9.863494,10.39508,10.909517,11.029553,10.765475,10.508256,10.14472,9.932085,9.760606,9.6645775,9.818909,10.511685,10.347065,9.863494,9.626852,10.2236,10.64201,11.485688,12.569438,13.735497,14.826107,15.282242,15.138199,15.062748,15.29939,15.659496,16.20137,16.80498,17.326277,17.826996,18.581505,18.235117,18.437462,18.451181,18.231688,18.44775,18.612371,19.377169,20.556948,21.747015,22.319756,25.18003,25.951689,25.824793,25.725336,26.325514,24.343212,22.69358,21.211998,19.387459,16.352274,12.202472,18.142517,21.28402,17.806417,12.97413,11.122152,12.30193,13.869251,12.696333,5.1821065,2.952875,2.0337453,1.7388009,1.6770682,1.762808,7.949784,5.874883,6.824879,12.034423,12.6757555,12.010415,13.96185,14.205351,11.317638,6.7802944,4.955754,6.5299344,7.2878733,5.8988905,3.9508848,8.203573,5.552502,4.2389703,5.98463,5.9914894,6.324159,6.7631464,7.058091,7.4970784,8.934075,7.3427467,8.838047,8.573969,6.5470824,7.596536,7.349606,7.623973,8.176137,8.64256,8.525954,7.414768,7.0923867,6.468202,4.90431,2.1915064,3.4398763,3.2992632,2.9460156,3.4295874,5.662249,6.9552035,4.3281393,4.746549,7.2021337,2.6785078,2.170929,3.093488,3.8548563,3.6970954,2.702515,6.012067,5.0312047,3.4021509,3.8205605,8.021805,5.7925735,6.660259,7.449064,5.9914894,1.138623,0.64133286,1.0494537,1.6496316,2.1846473,2.867135,3.0111778,4.170378,4.554492,4.0091877,4.029765,4.2766957,4.040054,3.6147852,3.391862,3.8479972,3.9303071,4.0263357,3.9646032,3.7176728,3.3850029,2.5961976,2.0714707,1.8656956,1.9102802,2.0165975,2.3286898,2.4315774,2.651071,2.8877127,2.6167753,2.4487255,2.277246,2.2360911,2.5824795,3.683377,3.625074,3.9337368,4.32471,4.5613513,4.4516044,4.4241676,4.695105,5.0106273,5.096367,4.650521,4.8734436,5.0312047,5.4153185,6.018926,6.5230756,7.2878733,7.5862474,7.7097125,7.9189177,8.464222,8.457363,7.870903,7.2878733,6.9346256,6.677407,6.667118,6.667118,6.8969,7.3598948,7.846896,8.30646,7.98065,7.606825,7.5588107,7.8263187,7.239859,6.81802,6.790583,7.06838,7.2707253,8.296172,8.587687,8.663138,8.738589,8.742019,8.498518,8.220721,8.1041155,8.093826,7.8846216,7.3839016,6.632822,6.135532,5.90575,5.4633327,5.4976287,5.5387836,5.5319247,5.470192,5.3878818,5.9331865,5.9228973,6.2144127,6.7357097,6.492209,6.169828,6.632822,6.475061,5.346727,3.9131594,3.0454736,3.6182148,7.610255,13.251926,15.028452,13.275933,9.283894,7.3393173,8.320179,9.719451,10.065839,8.525954,7.7542973,7.438775,4.3109913,3.6456516,2.3664153,3.3712845,5.796003,5.0483527,7.2878733,6.2075534,5.442755,5.813151,5.312431,3.2992632,3.333559,3.8445675,4.1600895,4.4996185,9.798331,8.261876,7.2947326,9.002667,10.189304,5.9743414,4.5201964,3.5976372,2.935727,4.2115335,7.298162,4.3007026,1.3375391,0.64476246,0.5590228,0.7133542,0.84367853,1.4335675,2.2258022,2.2258022,2.085189,2.218943,2.5653315,3.0111778,3.3815732,3.806842,3.4810312,4.091498,5.528495,5.857735,5.552502,5.377593,5.2609873,5.099797,4.773986,4.9008803,5.5559316,6.3035817,6.697984,6.2967224,6.697984,7.1266828,7.1541195,6.9689217,7.3701835,6.8043017,6.118384,5.7719955,5.7377,5.4976287,5.7274113,6.0326443,6.0875177,5.9743414,6.1972647,5.754848,5.3707337,5.3673043,5.658819,5.720552,6.667118,6.526505,6.3138704,6.4990683,7.0203657,7.466212,7.4936485,7.2707253,6.9792104,6.790583,6.5299344,6.4887795,6.608815,6.807731,6.9689217,7.0032177,7.3427467,7.7028537,7.8983397,7.857185,7.6651278,7.431916,6.8866115,6.0737996,5.3432975,4.537344,3.7142432,3.0900583,2.7059445,2.4452958,2.750529,3.2443898,3.8308492,4.48933,5.2609873,5.977771,5.9297566,4.681387,3.391862,4.8082814,3.3952916,3.9680326,4.770556,4.962613,4.619654,5.4667625,6.375603,6.5539417,5.9228973,5.120374,3.9611735,3.2478194,2.9974594,2.9460156,2.5413244,2.4727325,2.301253,2.1503513,2.0028791,1.6942163,2.0234566,2.7642474,3.5290456,4.098357,4.434457,4.8905916,5.2335505,5.689686,6.427047,7.5690994,8.2653055,8.292743,8.004657,7.720001,7.73029,8.64599,9.410788,9.928656,10.278474,10.72089,11.38623,11.763485,10.902658,9.054111,7.675417,7.0203657,7.099246,8.080108,9.277034,9.146709,9.489669,9.403929,9.095266,8.81061,8.827758,8.707723,9.208443,10.103564,10.755186,10.127572,9.729739,9.297611,9.054111,9.146709,9.668007,10.281903,9.832627,9.5205345,9.791472,10.326488,10.899229,10.686595,10.624862,11.303921,12.956982,11.4754,10.81006,9.6645775,8.011517,7.06495,5.686256,4.2046742,3.0317552,2.4658735,2.6956558,3.1209247,3.2032347,3.1415021,2.952875,2.469303,2.2669573,2.270387,2.4075704,2.6785078,3.1552205,3.100347,3.333559,3.7142432,4.122364,4.4687524,3.9783216,3.6593697,3.3541365,2.9117198,2.2086544,2.4315774,2.767677,2.9940298,3.210094,3.865145,4.262977,4.822,5.3090014,5.693115,6.1561093,6.708273,6.468202,5.645101,4.705394,4.3624353,4.8322887,5.0414934,4.897451,4.3452873,3.3747141,3.1792276,3.6627994,4.122364,4.4687524,5.2335505,0.11317638,0.14061308,0.08573969,0.044584636,0.05144381,0.06859175,0.09259886,0.06859175,0.061732575,0.07888051,0.061732575,0.037725464,0.037725464,0.08573969,0.17833854,0.26407823,0.26407823,0.28122616,0.33952916,0.45270553,0.6241849,0.6379033,0.77508676,0.83338976,0.77508676,0.7305021,0.7407909,0.84367853,1.0666018,1.4061309,1.8142518,2.4727325,2.6476414,2.5481834,2.3321195,2.095478,1.7559488,1.7490896,1.9514352,2.2978237,2.7711067,3.0386145,3.2992632,3.5187566,3.7108135,3.9508848,4.5613513,5.223262,5.4839106,5.1992545,4.5647807,4.2423997,4.712253,5.2609873,5.672538,6.23156,6.8214493,6.869464,6.756287,6.6431108,6.48535,6.0223556,5.662249,5.4976287,5.693115,6.4716315,8.042382,8.752307,8.597976,8.213862,8.879202,9.1810055,8.601405,7.599966,6.800872,7.016936,6.341307,6.0566516,6.0086374,6.39961,7.7714453,8.347616,8.549961,9.074688,10.021255,10.899229,9.633711,8.721441,7.6857057,6.636252,6.2830043,6.324159,6.293293,5.785714,4.962613,4.557922,4.091498,3.6216443,3.192946,2.9460156,3.1277838,3.1106358,3.391862,3.1072063,2.4830213,2.819121,3.234101,3.6079261,3.8137012,3.806842,3.642222,3.858286,3.7348208,3.8720043,4.1292233,3.642222,3.0489032,2.9220085,2.8088322,2.7299516,3.1792276,4.0434837,5.195825,6.036074,6.6705475,7.9292064,8.021805,7.2295704,6.756287,7.2021337,8.546532,8.694004,9.606275,10.827208,11.866373,12.178465,12.456262,12.740917,12.939834,13.001566,12.922686,13.320518,14.29795,14.682064,14.63062,15.645778,14.843254,14.692352,14.479718,14.003006,13.560589,13.612033,12.524854,11.71547,11.461681,10.902658,11.05699,11.698323,12.130451,12.511135,13.845244,13.985858,13.540011,12.572867,11.670886,11.924676,11.746337,11.526843,11.667457,12.000127,11.780633,11.732618,11.194174,11.026124,11.286773,11.211322,10.926665,10.854645,11.05699,11.629731,12.699762,12.404818,12.641459,13.179905,13.7526455,14.04759,13.649758,13.509145,13.313659,12.80608,11.773774,11.821788,11.880091,11.825217,11.650309,11.454823,12.260776,12.507706,12.281353,11.664027,10.734609,9.3936405,9.3936405,9.695444,9.674867,9.112414,9.595985,10.076128,10.381361,10.525404,10.714031,10.326488,10.425946,10.460241,10.31277,10.299051,10.518545,10.38479,9.887501,9.349055,9.407358,9.602845,10.278474,11.351934,12.600305,13.666906,14.599753,14.819247,14.826107,14.863832,14.946142,15.697222,16.688372,17.549198,18.20082,18.842154,18.605513,18.924463,19.181683,19.13024,18.87645,19.404606,19.881319,20.474638,21.45893,23.232025,25.6053,25.787067,26.256922,27.073164,25.883097,23.986534,23.122278,20.666695,17.243965,16.715809,20.045938,22.889067,20.4472,14.620332,13.999576,13.989287,13.848674,12.6757555,9.740028,4.4756117,2.3732746,2.0337453,2.0577524,1.9651536,2.1880767,13.440554,9.746887,8.351046,12.38424,10.858074,10.47396,14.438563,15.223939,11.177026,6.4887795,5.8200097,6.697984,6.293293,4.880303,5.844017,6.941485,4.938606,6.1286726,9.345626,5.9571934,5.8680243,6.944915,7.881192,8.258447,8.549961,8.282454,9.736599,9.242738,7.3050213,8.584257,6.279575,7.373613,8.570539,8.663138,8.539673,7.98065,7.455923,7.06495,5.9434752,2.277246,4.166949,3.0900583,2.2463799,3.1072063,5.381023,5.576509,4.1600895,5.802862,8.64256,4.2766957,4.0263357,3.1723683,3.3438478,4.4721823,4.7842746,6.7185616,5.7822843,4.166949,4.417309,9.434795,4.3349986,4.9420357,6.118384,5.003768,1.0254467,0.5178677,1.3443983,2.1640697,2.6613598,3.532475,3.799983,4.170378,4.1360826,3.9543142,4.65395,4.389872,4.355576,4.245829,4.040054,4.012617,4.307562,4.3281393,4.2286816,4.057202,3.758828,3.2478194,2.7813954,2.369845,2.1023371,2.1469216,2.5310357,2.6579304,2.9631636,3.2958336,2.9117198,2.6887965,2.3595562,2.3904223,3.0077481,4.1943855,4.1600895,4.32471,4.400161,4.3521466,4.386442,4.197815,4.5030484,5.0826488,5.4599032,4.887162,5.086078,5.1100855,5.3432975,5.8165803,6.2075534,6.2898636,6.6053853,6.924337,7.2021337,7.5588107,8.05953,8.2653055,8.189855,7.846896,7.2535777,6.917478,7.0203657,7.205563,7.284444,7.2295704,7.3187394,7.380472,7.3221693,7.250148,7.459353,7.233,6.852316,6.711703,6.914048,7.2535777,8.038953,8.467651,8.635701,8.700864,8.879202,8.669997,8.56025,8.673427,8.865483,8.711152,8.018375,7.0786686,6.324159,5.950334,5.919468,5.871454,5.813151,5.7102633,5.4839106,5.0346346,5.6519604,6.025785,6.368744,6.7219915,6.9517736,6.125243,6.1732574,6.042933,5.305572,4.1463714,3.1586502,2.5824795,4.0537724,7.239859,9.836057,11.207891,11.036412,10.124143,8.999237,7.915488,8.004657,8.176137,10.017825,11.619442,7.5725293,5.0414934,2.976882,3.765687,5.8371577,3.649081,3.6696587,3.8034124,4.0777793,4.588788,5.504488,4.3487167,3.5633414,3.7382503,4.297273,3.4776018,8.951223,7.81603,5.7582774,5.147811,5.0414934,5.2815647,4.016047,2.8225505,3.0900583,5.9983487,5.65539,4.266407,2.5824795,1.3649758,1.3855534,1.1008976,1.155771,1.5570327,2.0165975,1.9548649,2.4007113,2.9185789,3.2066643,3.1655092,2.9220085,3.2135234,3.340418,3.9714622,4.9008803,5.055212,4.2869844,4.4516044,4.65395,4.6436615,4.8117113,5.5730796,5.658819,6.0875177,6.7665763,6.48535,6.3310184,6.6225333,6.7665763,6.7219915,6.989499,6.7940125,6.1801167,5.6656785,5.5147767,5.7582774,5.926327,6.1561093,6.025785,5.675967,5.809721,5.809721,5.2609873,4.9180284,5.0346346,5.360445,6.1972647,6.39961,6.475061,6.591667,6.560801,6.601956,6.728851,6.917478,7.023795,6.7665763,6.6122446,6.5059276,6.5230756,6.708273,7.0786686,7.281014,7.4113383,7.599966,7.874333,8.141841,8.028665,7.7851634,7.2947326,6.5985265,5.9126086,5.1580997,4.32128,3.5530527,2.9734523,2.6990852,2.9974594,3.192946,3.6044965,4.2046742,4.616225,4.7259717,5.0449233,4.7945633,4.2389703,4.6882463,3.0969174,3.4810312,4.307562,4.8837323,5.3432975,5.8474464,6.461343,6.835168,6.728851,6.0052075,4.9694724,4.2389703,3.6627994,3.1689389,2.784825,2.510458,2.503599,2.4898806,2.3286898,2.0063086,2.1263442,2.4830213,3.0900583,3.7725463,4.1360826,4.3487167,4.461893,4.7774153,5.48734,6.6636887,6.8043017,6.931196,7.1712675,7.582818,8.158989,8.275595,9.163857,10.106995,10.72089,10.978109,10.693454,10.840926,10.350495,9.067829,7.723431,7.1987042,7.06838,7.623973,8.683716,9.599416,9.914937,9.73317,9.338767,9.095266,9.458802,9.877212,11.255906,12.308789,12.394529,11.537132,11.201033,10.251037,9.386781,9.246168,10.39508,11.238758,10.816919,10.179015,9.863494,9.914937,10.196163,10.179015,10.549411,11.543991,12.950122,11.694893,10.669447,9.191295,7.239859,5.4496145,4.3452873,3.5290456,3.0969174,3.0043187,3.059192,4.105216,4.057202,3.7691166,3.525616,3.059192,2.767677,2.5927682,2.527606,2.6133456,2.952875,2.9700227,3.117495,3.5118976,4.0777793,4.537344,4.1326528,3.8479972,3.625074,3.3198407,2.6853669,2.651071,3.1723683,3.5187566,3.590778,3.9097297,4.763697,5.2164025,5.5250654,5.7822843,5.936616,6.6568294,6.848886,6.48535,5.785714,5.2472687,4.8254294,4.8734436,4.647091,4.0606318,3.666229,3.8342788,4.420738,4.7842746,5.055212,6.1561093,0.12003556,0.15776102,0.09259886,0.061732575,0.09259886,0.07888051,0.10288762,0.07545093,0.061732575,0.072021335,0.07888051,0.072021335,0.09602845,0.17490897,0.28122616,0.34638834,0.35324752,0.33266997,0.37382504,0.4938606,0.64476246,0.6859175,0.7922347,0.805953,0.72021335,0.66876954,0.6756287,0.8162418,1.1249046,1.5673214,2.0577524,2.6167753,2.6750782,2.5378947,2.3458378,2.0646117,2.0131679,2.1263442,2.3664153,2.6476414,2.8396983,2.8294096,3.1723683,3.4981792,3.7005248,3.9028704,4.8425775,5.329579,5.435896,5.2335505,4.8082814,4.3692946,5.1238036,5.7068334,5.796003,6.090947,6.691125,6.4887795,6.166398,6.025785,5.9914894,5.936616,5.8474464,5.830299,6.15268,7.2467184,8.4264965,8.56025,8.131552,7.7542973,8.1487,8.141841,8.141841,7.747438,7.0306544,6.5230756,5.878313,5.8817425,5.9812007,6.1561093,6.924337,6.975781,7.486789,8.268735,9.019815,9.335337,7.9429245,7.2432885,6.2967224,5.113515,4.6402316,4.5613513,4.5099077,4.32471,3.9165888,3.2683969,2.8054025,2.633923,2.452155,2.2566686,2.3286898,2.5173173,2.719663,2.551613,2.1160555,2.0097382,2.435007,2.702515,2.8465576,2.8465576,2.6304936,2.8225505,2.8328393,3.0523329,3.3232703,2.952875,2.1915064,1.9651536,1.7696671,1.587899,1.8691251,2.469303,3.6593697,4.40702,4.6916757,5.518206,5.6073756,5.3673043,4.791134,4.557922,6.0566516,6.8454566,7.5279446,8.237869,8.934075,9.421077,10.13786,10.185875,10.175586,10.367643,10.683165,11.012405,12.349944,12.939834,12.751206,13.474849,13.371962,13.38911,13.234778,12.881531,12.548861,12.041282,11.293632,11.2250395,11.585147,10.971251,11.2421875,12.339656,13.025573,13.248496,14.140189,14.363112,14.150477,13.560589,13.169616,14.057879,13.54687,12.809509,12.439114,12.428825,12.151029,11.578287,11.039842,10.72775,10.55284,10.168727,9.829198,9.935514,10.326488,11.022695,12.22305,11.7257595,11.952112,12.343085,12.614022,12.785502,12.576297,12.871242,12.809509,12.130451,11.149589,11.080997,10.72089,10.381361,10.082987,9.589127,10.110424,10.799771,10.950673,10.484249,9.932085,9.112414,9.342196,9.770895,9.791472,9.0644,8.985519,9.345626,9.791472,10.1652975,10.508256,10.515115,10.940384,11.122152,10.81006,10.179015,10.093276,10.182446,10.079557,9.702303,9.249598,9.541112,10.007536,10.834066,11.945253,13.035862,14.291091,14.802099,14.832966,14.7369375,14.96672,15.6526375,16.62664,17.545769,18.214539,18.598652,18.643238,19.071936,19.394318,19.353163,18.914175,19.987637,20.556948,21.03709,22.007662,24.240324,25.704758,25.996273,26.76107,27.368109,24.891945,24.391226,23.393215,21.325174,20.53294,26.256922,22.463799,19.092514,15.079896,11.495977,11.543991,12.21962,11.640019,11.303921,10.161868,4.623084,2.020027,1.903421,2.3424082,3.7553983,8.923786,13.046151,11.351934,11.129011,12.367092,7.7714453,10.847785,12.792361,12.751206,10.89237,8.399059,7.414768,6.166398,4.976331,4.839148,7.4181976,5.518206,5.206114,7.380472,9.47938,5.4736214,7.0375133,7.9292064,8.299602,8.47451,8.964942,8.824328,9.901219,9.445084,7.9120584,8.988949,6.042933,7.4524937,8.786603,8.628842,8.587687,7.599966,8.272165,8.491658,6.8763227,2.7642474,5.254128,3.2409601,1.9137098,2.7951138,3.7519686,6.0978065,5.689686,7.034084,9.386781,6.776865,5.3330083,3.3301294,2.6407824,3.6387923,5.1992545,5.7068334,5.0174866,4.1292233,4.8151407,9.637141,4.5682106,4.6402316,4.962613,3.4878905,1.0117283,0.4081209,1.1866373,2.0989075,2.8054025,3.8891523,4.2286816,3.99204,3.724532,3.899441,4.928317,4.479041,4.722542,4.972902,5.0106273,5.0757895,5.096367,4.8082814,4.465323,4.2081037,4.0537724,3.9097297,3.5221863,3.0351849,2.6716487,2.7128036,3.100347,3.1689389,3.4707425,3.8479972,3.4364467,3.0969174,2.726522,2.8054025,3.5050385,4.681387,4.2938433,4.262977,4.2698364,4.297273,4.636802,4.461893,4.7945633,5.336438,5.669108,5.2781353,5.6656785,5.5319247,5.4324665,5.597087,5.885172,5.8680243,6.0497923,6.307011,6.56766,6.800872,7.4456344,8.021805,8.22758,8.025234,7.6616983,7.2432885,7.3358874,7.56224,7.579388,7.0718093,6.927767,6.869464,6.8900414,6.9620624,7.0443726,7.3358874,7.281014,7.2124224,7.3118806,7.6033955,8.289313,8.724871,8.947794,9.026674,9.054111,8.632272,8.549961,8.748878,8.951223,8.639131,7.8983397,7.390761,7.010077,6.7940125,6.9209075,6.5127864,6.1629686,5.9331865,5.7925735,5.6210938,5.8645945,6.23156,6.6122446,6.992929,7.4284863,6.7528577,6.4236174,5.9880595,5.312431,4.5922174,3.4776018,2.7779658,2.1229146,1.9685832,3.6044965,6.3721733,8.423067,9.362774,8.858624,6.615674,7.7783046,9.424506,13.361672,16.688372,11.794352,6.941485,4.2286816,4.2526884,5.0757895,2.2292318,2.3732746,2.3389788,2.6613598,3.525616,4.7499785,4.465323,4.108646,4.99005,6.1766872,4.4756117,7.936065,8.165848,6.4236174,4.931747,6.866034,6.0086374,4.8768735,3.5118976,3.1517909,6.2212715,3.6970954,3.549623,3.3301294,2.5619018,2.7573884,2.2978237,2.1434922,2.4007113,2.726522,2.335549,2.6373527,3.0248961,3.2683969,3.2615378,3.018037,2.719663,3.1963756,3.8308492,4.173808,3.940596,3.525616,3.6147852,3.8308492,4.0606318,4.465323,5.528495,5.6313825,6.0052075,6.667118,6.4373355,6.3207297,6.6465406,6.924337,7.0032177,7.0786686,7.1026754,6.684266,6.0840883,5.703404,6.0875177,5.8508763,5.950334,6.001778,5.895461,5.785714,5.994919,5.6999745,5.2164025,4.8734436,5.0003386,5.6039457,6.0978065,6.475061,6.574519,6.0840883,6.159539,6.186976,6.468202,6.8557453,6.7665763,6.5813785,6.375603,6.3721733,6.608815,6.927767,7.473071,7.682276,7.8983397,8.275595,8.769455,8.64942,8.368194,7.9463544,7.431916,6.869464,6.2075534,5.4633327,4.57164,3.7176728,3.3198407,3.5770597,3.566771,3.6593697,3.9268777,4.122364,4.1189346,4.420738,4.57507,4.5201964,4.588788,3.6525106,3.7553983,4.290414,4.9934793,5.953764,6.3035817,6.667118,7.0272245,7.1129646,6.3893213,5.8165803,5.360445,4.8837323,4.2286816,3.2272418,2.7402403,2.7711067,2.8019729,2.6785078,2.633923,2.5756202,2.5619018,3.0146074,3.8857226,4.6608095,4.73969,4.6916757,4.7671266,5.1752477,6.101236,6.2418494,6.636252,7.3221693,8.172707,8.913498,8.81747,9.613133,10.456812,10.916377,10.971251,10.429376,10.415657,10.106995,9.201583,7.9017696,7.723431,7.582818,7.6925645,8.361334,9.9801,10.703742,10.97468,10.803201,10.590566,11.115293,11.537132,12.932974,13.540011,13.094165,12.80265,12.956982,11.372512,9.650859,9.012956,10.271614,11.7257595,11.441104,10.816919,10.600855,10.88551,10.696883,10.515115,10.755186,11.499407,12.507706,11.89038,10.333347,8.484799,6.4373355,3.758828,3.5290456,3.192946,3.1106358,3.3678548,3.782835,4.5099077,4.3692946,4.1292233,4.0366244,3.8274195,3.5564823,3.175798,2.8054025,2.5927682,2.6990852,2.8945718,3.0214665,3.3541365,3.882293,4.2938433,4.3178506,4.1429415,3.981751,3.799983,3.2958336,3.0557625,3.3609958,3.74168,4.016047,4.256118,5.219832,5.717122,5.90575,5.8817425,5.6793966,6.0154963,6.1561093,6.252138,6.2898636,6.090947,5.5559316,5.2815647,4.8768735,4.396731,4.341858,4.7259717,5.346727,5.8234396,6.2212715,7.040943,0.048014224,0.082310095,0.082310095,0.12346515,0.17490897,0.09602845,0.058302987,0.0548734,0.061732575,0.07888051,0.12003556,0.12689474,0.17833854,0.2469303,0.28808534,0.26064864,0.33609957,0.29837412,0.33266997,0.47328308,0.6036074,0.6790583,0.6790583,0.6344737,0.5727411,0.5418748,0.6173257,0.8128122,1.1866373,1.6736387,2.1057668,2.4590142,2.3972816,2.2395205,2.1332035,2.0508933,2.4075704,2.5070283,2.6304936,2.7711067,2.620205,2.603057,2.9665933,3.2889743,3.532475,4.0194764,5.0895076,5.5387836,5.6313825,5.56965,5.4976287,4.7842746,5.579939,5.967482,5.535354,5.3913116,6.0840883,5.8645945,5.394741,5.086078,5.1066556,5.6039457,5.926327,6.3173003,6.8900414,7.630832,8.05953,8.090397,7.8983397,7.6033955,7.284444,7.205563,7.3221693,7.2878733,6.842027,5.830299,5.4907694,5.8234396,5.826869,5.24041,4.523626,4.605936,5.9126086,6.8454566,6.7459984,5.8817425,5.6348124,5.5387836,4.955754,4.1120753,4.098357,3.666229,3.2821152,2.983741,2.6887965,2.218943,1.7525192,2.0920484,2.3046827,2.136633,2.0268862,1.8554068,1.7353712,1.8554068,1.978872,1.4541451,1.5741806,1.4918705,1.4267083,1.4061309,1.2620882,1.6324836,1.9102802,2.177788,2.3767042,2.3046827,1.5913286,1.3512574,1.2758065,1.2963841,1.587899,1.9480057,3.0283258,3.6387923,3.549623,3.5050385,3.2272418,3.9440255,3.8342788,3.0969174,3.9303071,5.171818,5.5730796,6.018926,6.6431108,6.8283086,8.303031,7.888051,7.239859,7.4044795,8.80718,8.591117,9.97667,10.940384,11.091286,11.650309,11.862943,11.132441,10.789482,11.019264,10.875222,9.884071,9.89436,10.679735,11.537132,11.303921,12.205902,13.540011,14.164196,14.04759,14.2533655,14.959861,14.874121,14.7369375,15.011304,15.906426,15.138199,14.174485,13.5503,13.248496,12.686044,11.825217,11.351934,10.834066,10.179015,9.623423,9.314759,9.544542,9.801761,9.949233,10.22703,10.710602,11.348505,11.451392,11.070708,10.991828,11.211322,12.020704,12.133881,11.434244,10.950673,10.738038,10.257896,9.801761,9.379922,8.683716,8.412778,9.314759,9.887501,9.764035,9.692014,9.571979,9.839486,10.158438,10.175586,9.513676,8.834618,9.084977,9.613133,10.007536,10.065839,10.55284,11.156448,11.417097,11.039842,9.904649,9.774324,9.959522,10.172156,10.168727,9.774324,10.381361,10.738038,11.303921,12.22648,13.341095,14.490007,15.038741,15.127911,15.134769,15.690363,16.184223,16.825556,17.477179,17.95046,18.019053,18.272842,18.886738,19.198832,19.082224,18.948471,20.186552,21.098822,21.959648,23.02968,24.569565,25.67732,26.620459,26.970276,26.407824,24.710178,25.317215,22.638706,22.563255,27.11089,34.450207,16.29397,9.784613,9.167287,9.205012,5.1580997,6.159539,7.1541195,9.942374,12.140739,7.191845,4.4516044,3.6799474,4.033195,7.1198235,16.96617,7.905199,10.799771,13.937843,11.900668,5.56965,12.6586075,9.517105,8.038953,10.419086,9.153569,8.611694,6.1321025,4.887162,5.7102633,7.0923867,4.9180284,6.3138704,7.267296,6.6465406,6.200694,9.877212,9.167287,7.9600725,8.05953,9.177576,8.669997,9.56512,9.201583,7.822889,8.597976,7.0203657,8.169277,8.958082,8.484799,8.025234,6.684266,9.047252,9.938945,7.4970784,3.1860867,6.018926,3.7313912,1.9925903,2.2909644,1.9411465,7.881192,7.2295704,7.0615206,8.769455,8.076678,4.5613513,3.5461934,2.4658735,1.4198492,3.1620796,3.1449318,2.9288676,3.0660512,4.633373,9.235879,7.531374,5.9400454,3.940596,1.8519772,0.8162418,0.34295875,0.77851635,1.6976458,2.7985435,3.9028704,4.1772375,3.899441,3.7794054,4.1292233,4.846007,4.7259717,4.9008803,5.2026844,5.6210938,6.3001523,5.874883,5.284994,4.695105,4.273266,4.2218223,4.307562,3.9783216,3.6319332,3.5187566,3.7313912,4.0606318,3.9646032,4.0777793,4.314421,3.8548563,3.5153272,3.40901,3.6319332,4.187526,4.996909,4.139512,4.1292233,4.3007026,4.5167665,5.1752477,5.15467,5.562791,5.9228973,6.025785,5.9228973,6.478491,6.217842,5.8508763,5.7411294,5.919468,6.1629686,6.1972647,6.1561093,6.2144127,6.6122446,7.06838,7.4627824,7.6274023,7.6857057,8.06296,7.7920227,7.699424,7.891481,8.05953,7.4936485,7.298162,6.715132,6.5162163,6.773435,6.852316,7.3358874,7.613684,7.798882,7.956643,8.131552,9.016385,9.448513,9.661148,9.709162,9.5033865,8.937505,8.7317295,8.80718,8.841476,8.289313,7.6376915,7.6857057,7.9017696,7.9909387,7.874333,7.040943,6.509357,6.3138704,6.4304767,6.756287,6.5950966,6.632822,6.958633,7.48336,7.932636,7.9086285,7.5416627,6.701414,5.5662203,4.5956473,3.8034124,3.6285036,3.100347,2.1332035,1.5055889,1.4164196,1.9342873,4.108646,6.6053853,5.720552,8.656279,10.281903,13.937843,17.693241,14.342535,9.218731,6.327589,4.770556,3.5564823,1.5673214,2.054323,1.903421,1.9445761,2.4075704,2.935727,3.100347,3.9851806,5.9469047,7.4765005,5.212973,5.844017,7.0786686,7.4181976,7.7748747,11.492548,6.6293926,6.742569,5.874883,3.7039545,5.521636,4.1635194,3.4021509,3.3061223,3.690236,4.1155047,3.7553983,3.292404,3.542764,4.07435,3.2135234,2.8945718,2.7128036,2.819121,3.1826572,3.5804894,2.9974594,3.3129816,3.7382503,3.7519686,3.083199,3.542764,3.3026927,3.3061223,3.74168,4.029765,4.763697,5.4324665,6.142391,6.608815,6.183546,6.636252,7.208993,7.579388,7.675417,7.682276,7.675417,7.4044795,6.852316,6.327589,6.468202,5.6793966,5.5662203,5.9126086,6.310441,6.159539,6.4407654,6.5196457,6.125243,5.4324665,5.0655007,5.5147767,5.970912,6.310441,6.358455,5.857735,6.341307,6.15268,6.135532,6.5162163,6.8797526,6.742569,6.355026,6.3653145,6.7631464,6.852316,7.589677,8.165848,8.580828,8.951223,9.517105,9.325048,8.961512,8.577398,8.203573,7.7714453,7.3118806,6.7048435,5.7994323,4.7808447,4.1943855,4.314421,4.187526,3.8514268,3.5461934,3.7211025,4.040054,4.1600895,4.256118,4.465323,4.866585,4.8940215,4.9934793,5.1992545,5.5902276,6.293293,6.478491,6.7802944,6.9723516,6.869464,6.3207297,6.138962,6.0395036,6.046363,5.73427,4.214963,3.4364467,3.2306714,3.1449318,3.1106358,3.3987212,3.210094,3.0489032,3.3781435,4.341858,5.7754254,6.094377,5.9571934,5.7994323,5.919468,6.4819202,7.016936,7.6651278,8.457363,9.242738,9.685155,9.952662,10.6317215,11.022695,10.981539,10.912948,10.978109,11.163307,10.882081,10.021255,8.9100685,9.019815,8.707723,8.419638,8.704293,10.216741,11.55428,12.614022,12.987847,12.922686,13.2862215,12.816368,13.392539,13.402828,12.953552,13.869251,14.30138,12.370522,10.045261,8.738589,9.297611,11.118723,11.358793,11.303921,11.619442,12.339656,11.773774,11.321068,11.094715,11.290202,12.171606,12.020704,10.388221,8.320179,5.9914894,2.7093742,3.210094,3.1037767,3.0557625,3.4535947,4.420738,4.1600895,4.214963,4.400161,4.57164,4.65395,4.461893,3.9611735,3.3369887,2.8225505,2.702515,3.0248961,3.1826572,3.4638834,3.858286,4.064061,4.482471,4.417309,4.262977,4.15323,3.974892,3.7519686,3.6285036,3.9200184,4.5167665,4.8768735,5.4839106,6.118384,6.375603,6.1458206,5.6039457,5.2335505,5.0346346,5.4153185,6.1732574,6.495639,6.324159,5.892031,5.48734,5.271276,5.2918534,5.627953,6.0669403,6.677407,7.239859,7.2158523,0.061732575,0.13375391,0.106317215,0.09602845,0.106317215,0.044584636,0.058302987,0.08916927,0.106317215,0.12003556,0.16804978,0.20577525,0.21263443,0.20920484,0.18519773,0.1371835,0.22292319,0.216064,0.26407823,0.39783216,0.5178677,0.5418748,0.5418748,0.53501564,0.52815646,0.5041494,0.7339317,0.9568549,1.2072148,1.471293,1.6770682,1.9342873,1.9720128,2.0131679,2.1846473,2.503599,2.9665933,2.760818,2.603057,2.609916,2.3046827,2.510458,3.0043187,3.4227283,3.8102717,4.5922174,5.302142,5.6245236,5.6965446,5.717122,5.936616,6.327589,6.5710897,6.5779486,6.307011,5.7822843,6.111525,5.7822843,5.360445,5.020916,4.530485,4.9214582,5.717122,6.6431108,7.3393173,7.3393173,6.8385973,7.143831,7.1026754,6.5642304,6.392751,6.7219915,6.550512,6.495639,6.492209,5.7822843,5.147811,4.9523244,4.73969,4.2526884,3.450165,3.4227283,4.2423997,4.540774,4.07435,3.707384,4.0880685,4.197815,4.040054,3.6456516,3.0969174,2.6956558,2.136633,1.8245405,1.7662375,1.5707511,1.4369972,1.4232788,1.4027013,1.4027013,1.587899,1.5638919,1.3169615,1.1111864,1.0117283,0.91569984,1.1351935,1.1729189,1.0117283,0.8128122,0.8848336,0.97057325,1.0014396,1.2209331,1.5844694,1.7559488,1.5604624,1.4267083,1.2689474,1.3443983,2.2566686,2.16064,2.1091962,2.201795,2.417859,2.6236343,1.8313997,2.6579304,3.0248961,2.6613598,3.1140654,3.9440255,4.4996185,5.096367,5.597087,5.4016004,5.9743414,6.3035817,6.142391,5.950334,6.866034,6.3173003,7.298162,8.927217,10.429376,11.1393,10.9198065,9.849775,8.786603,8.162418,7.98065,8.114404,8.81747,9.993818,11.255906,11.900668,13.488567,14.078457,14.517444,15.049029,15.302819,15.121051,14.973578,14.5243025,14.112752,14.771234,14.55174,13.735497,13.642899,14.335675,14.603184,13.039291,11.71547,10.909517,10.501397,9.962952,9.403929,9.592556,9.829198,9.798331,9.568549,9.201583,9.760606,10.449953,10.81006,10.710602,11.029553,11.245617,11.427385,11.523414,11.351934,11.084427,10.511685,9.901219,9.403929,9.0644,8.783174,9.078118,9.585697,10.021255,10.192734,10.278474,10.539123,10.868362,10.978109,10.39165,9.403929,9.191295,9.400499,9.661148,9.613133,10.151579,10.31277,10.604284,10.981539,10.834066,10.271614,10.350495,10.206452,9.908078,10.484249,11.262765,12.044711,12.898679,13.63604,13.7938,14.160767,14.911846,15.498305,15.87213,16.496315,17.165085,17.645227,17.87158,17.737827,17.089634,17.247395,17.909306,18.516342,19.010202,19.850452,20.37518,21.03709,21.918493,22.87192,23.544119,25.862518,27.165762,26.826233,25.77335,26.503853,25.392666,20.594673,22.820475,27.320093,13.855534,11.561139,8.268735,8.217292,9.551401,4.3041325,4.8151407,5.1169443,3.9886103,4.5682106,14.359683,14.332246,11.423956,10.028113,10.652299,9.935514,7.160979,12.308789,12.542002,7.023795,6.910619,10.329918,7.9909387,7.1884155,8.200144,4.256118,6.0532217,5.90575,6.492209,7.1026754,3.6627994,4.8940215,7.473071,7.5279446,6.334448,10.316199,11.170166,8.207003,6.5470824,7.2124224,7.1266828,7.7611566,9.595985,9.088407,7.058091,8.683716,8.865483,9.211872,9.493098,8.611694,4.6093655,5.8543057,7.2535777,8.851766,8.680285,2.7470996,4.8597255,3.765687,2.294394,1.611906,1.2209331,8.556821,5.137522,3.391862,5.878313,5.2781353,2.020027,3.6319332,3.8445675,1.7319417,1.7079345,1.5261664,1.3443983,1.3684053,3.2409601,10.041832,11.478829,8.399059,3.899441,0.5144381,0.18176813,0.5007198,1.4027013,2.7711067,4.1600895,4.804852,4.756838,4.554492,4.5956473,4.931747,5.2506986,5.3330083,5.055212,4.979761,5.3227196,5.919468,5.552502,5.178677,4.537344,3.8171308,3.6456516,3.974892,4.0674906,4.1463714,4.3658648,4.804852,4.928317,4.400161,3.998899,3.8788633,3.5873485,3.5976372,4.149801,4.870014,5.336438,5.0826488,4.3109913,4.4859004,4.7534084,4.955754,5.6142344,5.857735,6.2967224,6.8763227,7.4010496,7.5210853,7.5588107,7.377043,7.1198235,6.7631464,6.1046658,6.2864337,6.6876955,6.6396813,6.2727156,6.5162163,6.6876955,7.040943,7.4970784,8.06296,8.820899,8.587687,8.621983,8.48137,8.186425,8.224151,7.747438,7.298162,7.0615206,6.9963584,6.852316,7.2158523,7.630832,7.9086285,8.069819,8.299602,8.923786,9.592556,9.959522,9.990388,9.9801,9.832627,9.47595,9.187865,9.019815,8.790032,8.018375,8.001227,8.069819,7.936065,7.689135,7.3358874,7.0546613,6.989499,7.0752387,7.051232,7.1712675,7.2947326,7.579388,8.090397,8.772884,8.906639,8.556821,7.73372,6.6465406,5.7068334,4.046913,4.355576,4.5819287,3.8617156,2.5173173,2.2258022,1.6667795,3.5942078,6.23156,3.2649672,6.036074,5.329579,5.5902276,8.289313,11.900668,12.401388,9.633711,5.6245236,2.3389788,1.6770682,1.3238207,1.4198492,1.4987297,1.3615463,1.0666018,1.2037852,1.3649758,2.5961976,4.016047,2.8088322,4.7842746,5.2609873,6.193835,7.2192817,5.645101,4.7671266,7.191845,7.966932,6.3618846,5.874883,5.7754254,3.865145,3.0660512,3.9097297,4.530485,3.7519686,3.1243541,3.083199,3.40901,3.2512488,3.309552,3.2546785,3.0900583,3.0420442,3.5564823,3.6147852,3.8514268,4.2526884,4.4996185,3.9371665,3.6559403,3.6044965,3.9165888,4.434457,4.715683,4.715683,5.0277753,5.7822843,6.560801,6.3790326,6.7940125,7.720001,8.299602,8.292743,8.073249,8.035523,7.449064,6.9620624,6.8214493,6.883182,6.4064693,6.341307,6.4133286,6.4990683,6.6225333,7.390761,7.016936,6.6053853,6.3721733,5.6142344,5.6656785,6.142391,6.385892,6.334448,6.5299344,6.6053853,6.2727156,6.169828,6.550512,7.2947326,7.939495,7.56224,7.3530354,7.630832,7.8263187,8.207003,8.858624,9.122703,9.102125,9.688584,9.846346,9.3764925,8.790032,8.296172,7.781734,7.6342616,7.2707253,6.615674,5.7308407,4.791134,4.6676683,4.3281393,3.789694,3.2546785,3.0969174,3.426158,3.9680326,4.3349986,4.5030484,4.804852,5.967482,6.468202,6.6122446,6.7322803,7.1712675,6.8797526,6.8043017,6.574519,6.210983,6.1492505,5.7822843,5.7822843,6.1629686,6.5813785,6.3618846,4.8734436,4.098357,3.7313912,3.6559403,3.9371665,4.15666,3.899441,3.765687,4.40702,6.5299344,7.654839,7.7131424,7.6033955,7.750868,8.117833,8.056101,8.56368,9.3764925,10.261326,11.015835,10.247607,10.851214,11.516555,11.729189,11.780633,12.696333,13.646329,13.279363,11.924676,11.595435,11.218181,10.22703,9.462232,9.458802,10.436234,12.000127,13.516005,14.321958,14.335675,14.068168,12.689473,12.8197975,13.114742,13.502286,15.21365,14.054449,12.902108,11.485688,10.117283,9.688584,11.118723,12.562579,12.977559,12.569438,12.80265,11.64345,11.252477,11.177026,11.194174,11.290202,11.180455,10.906088,9.1810055,6.0806584,3.0523329,2.867135,3.0248961,3.2375305,3.566771,4.4104495,4.2766957,4.9180284,5.4941993,5.6073756,5.3261495,5.0929375,4.7499785,4.2869844,3.7794054,3.3884325,3.3747141,3.508468,3.9851806,4.5647807,4.5784993,4.5167665,4.4275975,4.184097,4.0503426,4.6848164,4.928317,4.7602673,4.955754,5.4153185,5.1580997,5.3158607,5.895461,6.5779486,6.910619,6.2864337,5.7136927,5.442755,5.7102633,6.3721733,6.8969,6.3481665,6.1629686,5.909179,5.6210938,5.830299,6.0978065,6.3207297,6.64997,6.800872,6.0566516,0.13375391,0.13032432,0.09602845,0.07888051,0.09602845,0.13032432,0.17147937,0.14404267,0.12346515,0.14061308,0.17833854,0.22635277,0.2469303,0.22978236,0.1920569,0.17490897,0.18176813,0.1920569,0.274367,0.4081209,0.4698535,0.4938606,0.47671264,0.53501564,0.6379033,0.61389613,0.805953,0.90198153,0.9911508,1.155771,1.471293,1.7765263,1.9274281,2.1469216,2.49331,2.867135,2.959734,2.942586,2.8465576,2.6819375,2.4247184,2.534465,3.1140654,3.6696587,4.0434837,4.386442,4.9180284,5.0655007,5.288424,5.7754254,6.4373355,6.3961806,6.540223,6.8454566,6.835168,5.586798,5.926327,6.0840883,5.861165,5.3741636,5.0312047,5.5113473,6.831738,7.6376915,7.363324,6.2418494,6.5813785,7.2124224,7.082098,6.2727156,6.001778,6.018926,5.885172,5.638242,5.2918534,4.8185706,4.7019644,4.9077396,4.629943,3.6936657,2.5584722,2.503599,2.627064,2.5893385,2.3904223,2.3767042,2.5413244,2.6133456,2.5824795,2.4418662,2.194936,1.8691251,1.5947582,1.4678634,1.3821237,1.0117283,1.0117283,1.0837497,1.1900668,1.2860953,1.2929544,1.3101025,1.0528834,0.89855194,0.91227025,0.84367853,0.8471081,0.94656616,0.9294182,0.84024894,0.97057325,0.89855194,0.8162418,0.8676856,0.9945804,0.9602845,0.90198153,1.0460242,0.980862,0.78537554,1.0254467,0.9945804,1.0425946,1.0563129,1.0528834,1.1729189,1.0425946,1.3341095,1.605047,1.786815,2.16064,2.843128,3.3541365,3.6799474,3.7176728,3.2786856,3.7142432,4.0880685,4.232111,4.190956,4.2183924,4.5167665,5.7102633,7.267296,8.697433,9.551401,8.796892,8.110974,7.8194594,7.781734,7.394191,7.051232,7.140401,7.997798,9.273604,9.959522,10.336777,11.180455,12.367092,13.471419,13.766364,12.703192,12.984418,13.454271,13.766364,14.366542,14.225929,14.088745,13.958421,14.054449,14.808959,14.205351,13.039291,12.041282,11.375941,10.621432,9.856634,9.908078,10.189304,10.261326,9.836057,9.849775,9.846346,10.216741,10.820349,10.9541025,11.156448,11.029553,11.338216,12.006986,12.109874,11.790922,11.38623,10.422516,9.242738,8.97866,9.067829,9.39021,9.89436,10.333347,10.278474,9.640571,9.692014,10.288762,11.070708,11.454823,10.923236,10.2921915,9.650859,9.194724,9.22216,9.709162,9.846346,10.041832,10.261326,10.028113,10.628291,10.662587,10.662587,10.964391,11.701753,12.144169,12.531713,13.066729,13.680624,14.013294,14.400838,14.819247,15.158776,15.529172,16.249386,17.487467,18.533491,19.154245,19.095943,18.077356,17.926455,18.03963,18.180243,18.403166,19.071936,19.809298,20.649546,21.767591,22.769032,22.690151,25.26234,26.256922,26.119738,25.886526,27.17605,22.967947,21.527521,22.210009,21.53095,13.13532,8.261876,4.389872,2.7779658,3.2992632,4.4241676,3.981751,5.120374,9.794902,13.704632,6.279575,5.521636,6.0395036,7.425057,8.968371,9.6645775,11.063849,9.863494,7.5725293,7.905199,16.798119,8.783174,6.842027,6.5196457,5.8337283,5.2575574,6.6533995,6.2658563,6.2384195,6.6705475,5.638242,7.623973,6.4887795,5.4667625,6.3618846,9.5205345,7.8366075,6.7871537,7.2364297,8.333898,7.517656,7.915488,9.671436,9.945804,9.006097,10.220171,9.084977,9.263316,9.441654,8.663138,6.327589,9.849775,7.966932,6.7871537,7.14726,4.6127954,3.2683969,3.216953,2.7162333,1.7147937,1.8313997,6.8626046,4.139512,2.2052248,4.1635194,7.6959944,5.9297566,6.495639,5.545643,2.7573884,1.3169615,2.9700227,2.1126258,2.170929,5.312431,12.445972,12.744347,8.4093485,3.4398763,0.36353627,0.2194936,1.1317638,2.2052248,3.4364467,4.523626,4.866585,5.1100855,4.8494368,4.681387,4.7774153,4.870014,4.5956473,4.4275975,4.647091,5.223262,5.809721,5.425607,5.271276,4.8597255,4.105216,3.3301294,3.1792276,3.5633414,4.1017866,4.5442033,4.770556,3.974892,3.5393343,3.3712845,3.292404,3.0489032,3.3541365,4.266407,5.56965,6.680836,6.619104,5.761707,5.130663,5.0003386,5.31929,5.7239814,6.183546,6.6876955,7.0478024,7.438775,8.388771,8.573969,8.471081,8.100685,7.534804,6.883182,6.7940125,6.5299344,6.3035817,6.2384195,6.3447366,6.2041235,6.619104,7.1884155,7.870903,8.97866,9.009526,9.205012,9.088407,8.718011,8.676856,8.453933,7.8194594,7.363324,7.140401,6.680836,6.8626046,7.298162,7.459353,7.394191,7.750868,8.285883,8.89635,9.451943,9.89093,10.209882,9.997248,9.56512,8.940934,8.340756,8.179566,8.532814,8.443645,8.100685,7.723431,7.5553813,7.5039372,7.4456344,7.4524937,7.4799304,7.366754,7.6342616,7.2295704,7.349606,8.193284,8.944365,9.273604,8.995808,8.169277,7.2364297,6.989499,5.6313825,4.880303,4.4996185,4.098357,3.117495,2.74367,2.0577524,1.8725548,2.3252604,2.8739944,3.974892,3.9783216,4.040054,4.6745276,5.7377,4.7259717,4.5167665,3.8102717,2.5447538,1.8862731,1.6393428,1.4678634,1.2243627,0.9294182,0.7613684,0.9842916,1.3821237,2.510458,3.6319332,2.6853669,5.113515,6.931196,7.6788464,7.257007,5.926327,4.461893,5.672538,5.528495,4.081209,5.446185,6.7357097,5.861165,4.846007,4.6127954,4.972902,7.1678376,4.012617,3.7622573,6.1286726,2.2978237,2.8294096,2.8877127,2.884283,2.9254382,2.8225505,3.333559,3.093488,5.5593615,8.64942,4.7671266,4.633373,4.091498,3.99204,4.3281393,4.2252517,4.763697,4.7191124,5.271276,6.478491,7.281014,7.5588107,8.107545,8.258447,8.086967,8.412778,8.385342,7.750868,7.116394,6.776865,6.711703,6.5779486,7.226141,7.534804,7.3050213,7.281014,8.2653055,8.200144,7.750868,7.0718093,5.7994323,5.7891436,6.4887795,7.0546613,7.3255987,7.8263187,6.8728933,6.5367937,6.8728933,7.490219,7.548522,8.303031,8.303031,8.213862,8.457363,9.218731,9.537683,9.729739,9.753747,9.602845,9.297611,9.105555,8.916927,8.738589,8.522525,8.196714,8.032094,7.8503256,7.5107965,6.81802,5.535354,4.681387,4.1360826,3.8034124,3.525616,3.0729103,3.0797696,3.4021509,3.9611735,4.623084,5.171818,5.346727,6.492209,7.442205,7.7440085,7.6959944,7.2192817,6.8214493,6.451054,6.142391,6.001778,5.7719955,5.662249,5.7479887,6.046363,6.509357,5.7411294,4.979761,4.4687524,4.256118,4.2046742,4.4721823,4.6848164,5.1066556,6.077229,7.9943686,9.362774,9.088407,8.460793,8.621983,10.569988,10.950673,10.964391,11.063849,11.180455,10.734609,10.532263,11.002116,11.592006,11.958971,11.938394,13.138749,14.277372,14.874121,14.771234,14.160767,13.584596,12.435684,11.180455,10.449953,11.046701,12.171606,13.54687,14.616901,15.13134,15.165636,14.081886,13.612033,13.797231,14.613472,15.981877,13.951562,11.684605,10.240748,9.822338,9.774324,10.882081,12.034423,12.415107,11.917816,11.153018,10.6488695,10.319629,10.6317215,11.050131,10.034973,9.788043,9.668007,8.796892,6.773435,3.6868064,2.935727,2.9734523,3.3678548,3.974892,4.9351764,5.161529,5.40503,5.9434752,6.6053853,6.7528577,6.090947,5.422178,4.955754,4.7259717,4.6093655,4.4687524,4.650521,5.0826488,5.552502,5.6999745,4.8494368,4.5339146,4.4104495,4.4550343,4.9523244,5.528495,5.686256,5.6999745,5.703404,5.669108,5.3707337,5.579939,6.2144127,6.941485,7.1781263,6.574519,6.2727156,6.375603,6.7528577,7.0443726,6.444195,6.2212715,6.0806584,6.0086374,6.2555676,6.3893213,6.4887795,6.5299344,6.5299344,6.5470824,0.17147937,0.12346515,0.09259886,0.07888051,0.10288762,0.17833854,0.16462019,0.1371835,0.12003556,0.12689474,0.15433143,0.20577525,0.22978236,0.2469303,0.24350071,0.20234565,0.19548649,0.2194936,0.2709374,0.32581082,0.33952916,0.41498008,0.4664239,0.59674823,0.7442205,0.66876954,0.8162418,0.91227025,1.1077567,1.4232788,1.7593783,2.0303159,2.270387,2.4727325,2.6647894,2.9220085,2.9734523,3.0660512,3.0351849,2.8705647,2.6853669,2.7711067,3.1552205,3.4981792,3.7759757,4.2869844,4.386442,4.4275975,4.8597255,5.6176643,6.121814,6.0840883,6.279575,6.608815,6.5710897,5.2747054,5.909179,6.276145,6.108095,5.521636,5.0106273,5.5422134,7.346176,8.110974,7.346176,6.3961806,6.433906,6.783724,6.742569,6.193835,5.593657,5.079219,4.856296,4.547633,4.064061,3.5976372,3.875434,3.9303071,3.433017,2.534465,1.8862731,1.8828435,1.605047,1.4644338,1.4918705,1.3409687,1.4644338,1.6530612,1.786815,1.7971039,1.6496316,1.4369972,1.313532,1.2998136,1.2312219,0.7510797,0.7442205,0.90541106,1.0425946,1.0563129,0.94656616,0.9568549,0.84024894,0.7476501,0.71678376,0.6790583,0.6962063,0.77851635,0.83338976,0.86082643,0.96371406,0.83338976,0.70649505,0.6859175,0.7305021,0.65162164,0.5624523,0.5796003,0.5555932,0.47328308,0.4424168,0.45270553,0.44584638,0.41840968,0.39440256,0.432128,0.4629943,0.5658819,0.8162418,1.1866373,1.546744,1.9171394,2.527606,3.0077481,3.1380725,2.867135,2.5961976,2.6579304,2.819121,2.983741,3.199805,3.9680326,4.698535,5.7239814,6.914048,7.671987,7.140401,6.9689217,7.226141,7.531374,7.0546613,6.6431108,6.8043017,7.6205435,8.7283,9.328478,8.971801,9.602845,10.686595,11.842365,12.850664,12.857523,13.313659,13.745787,13.906977,13.745787,13.858963,14.596324,15.066177,15.073037,15.155347,15.0456,14.445422,13.255356,11.780633,10.741467,10.254466,10.39165,10.436234,10.367643,10.827208,11.111863,10.830637,10.779194,11.015835,10.861504,11.523414,11.4033785,11.543991,12.154458,12.610593,12.449403,11.746337,10.563129,9.331907,8.838047,9.249598,9.770895,10.39508,10.827208,10.491108,10.010965,9.932085,10.106995,10.429376,10.840926,11.05356,10.714031,10.05898,9.438225,9.280463,9.493098,9.626852,9.609704,9.441654,9.177576,9.839486,10.113853,10.569988,11.348505,12.13731,12.006986,12.21962,12.548861,12.926115,13.437123,14.143619,14.898128,15.21022,15.2033615,15.604623,16.647217,18.231688,19.716698,20.560377,20.313446,19.8676,19.689262,19.53836,19.349733,19.233126,20.025362,21.153696,22.43979,23.52354,23.849352,25.300066,25.9414,26.19176,26.36324,26.647894,23.60242,21.45893,19.404606,15.608052,7.2432885,3.8548563,3.5976372,8.711152,13.200482,2.843128,3.758828,3.1655092,4.729401,6.8454566,2.6373527,2.7059445,3.5633414,4.636802,5.586798,6.293293,6.5950966,5.5833683,5.096367,6.3138704,9.73317,5.5559316,5.6656785,6.0806584,5.6793966,6.2041235,6.869464,5.6348124,5.579939,6.728851,6.0532217,6.869464,5.717122,5.857735,7.7268605,8.930646,6.5882373,7.5279446,8.128122,7.514226,7.5690994,8.752307,9.719451,10.155008,10.14472,10.155008,9.043822,9.949233,10.72775,10.05898,7.455923,12.291641,8.028665,4.434457,4.619654,5.0346346,2.627064,3.0557625,3.0489032,2.2120838,3.0351849,4.064061,3.6868064,3.99204,5.2609873,5.9743414,8.831187,8.519095,5.909179,2.942586,2.6579304,3.3781435,4.7979927,7.56224,11.351934,14.867262,9.849775,4.9420357,1.6839274,0.4698535,0.58645946,1.6633499,3.1826572,4.256118,4.7088237,5.0929375,5.284994,4.7259717,4.65395,5.1100855,4.914599,4.722542,4.7602673,4.773986,4.835718,5.360445,5.754848,5.672538,5.271276,4.7671266,4.4413157,3.6147852,3.6765177,4.1120753,4.4275975,4.173808,3.5359046,3.1689389,3.117495,3.2512488,3.2546785,3.6010668,4.513337,5.950334,7.349606,7.606825,6.8763227,6.121814,5.7925735,6.001778,6.540223,6.999788,7.4456344,7.654839,7.8091707,8.488229,8.742019,8.357904,8.042382,7.9429245,7.64798,7.160979,6.324159,5.970912,6.1321025,6.036074,6.4990683,7.2467184,7.874333,8.47451,9.640571,9.671436,9.633711,9.544542,9.469091,9.513676,8.971801,8.1212635,7.5450926,7.2364297,6.5813785,6.5196457,6.6293926,6.790583,6.8900414,6.81802,7.160979,7.846896,8.762596,9.695444,10.323058,9.873782,9.321619,8.889491,8.64942,8.546532,9.012956,8.886061,8.505377,8.124693,7.9257765,7.7097125,7.7748747,8.052671,8.333898,8.279024,8.114404,7.582818,7.589677,8.323608,9.263316,9.400499,9.493098,9.019815,8.097256,7.473071,6.6739774,5.970912,5.5079174,5.144381,4.4721823,3.782835,3.0797696,2.277246,1.786815,2.5207467,2.8019729,3.2889743,4.0880685,5.353586,7.281014,4.2355404,3.340418,4.547633,6.461343,6.324159,2.6613598,1.3855534,1.0494537,0.85739684,0.6790583,0.7373613,1.2037852,2.0097382,2.976882,3.789694,4.6608095,5.2918534,7.332458,10.206452,11.14273,10.415657,10.528833,9.674867,7.8503256,6.831738,6.5779486,6.447624,6.186976,5.65539,4.7979927,4.979761,3.841138,3.690236,4.588788,4.3590055,4.0229063,2.719663,2.0234566,2.2429502,2.411,2.585909,2.5138876,3.8685746,6.7357097,9.589127,5.8645945,5.518206,5.717122,5.206114,4.314421,4.955754,4.6745276,5.099797,6.3961806,7.233,7.4181976,8.117833,8.279024,7.949784,8.251588,8.337327,7.870903,7.5245147,7.449064,7.2707253,7.1712675,7.8366075,8.2481575,8.100685,7.7851634,8.697433,8.666568,8.244728,7.623973,6.667118,5.90232,6.279575,7.006647,7.723431,8.488229,7.514226,7.0032177,7.082098,7.500508,7.623973,8.844906,8.81747,8.501947,8.460793,8.879202,9.06097,9.3936405,9.692014,9.657719,8.851766,8.580828,8.31332,7.963502,7.517656,6.999788,7.1095347,7.3358874,7.226141,6.550512,5.2918534,4.5099077,4.0194764,3.625074,3.2581081,2.976882,3.100347,3.426158,3.7931237,4.214963,4.863155,4.955754,5.892031,7.0752387,7.8434668,7.4627824,7.1061053,6.90033,6.7494283,6.5127864,6.001778,5.5079174,5.3090014,5.3981705,5.7719955,6.4373355,6.0840883,5.586798,5.3570156,5.5079174,5.8645945,5.778855,6.0978065,6.9071894,8.073249,9.22216,9.184435,8.724871,8.608265,9.434795,11.670886,12.751206,13.166186,12.593445,11.362224,10.456812,10.4533825,11.022695,11.732618,12.178465,11.986408,12.932974,13.601744,14.164196,14.538021,14.390549,13.55373,12.332796,11.249047,10.786053,11.382801,12.97413,14.38026,15.594335,16.362562,16.163645,14.095605,12.977559,13.361672,14.88441,16.273392,14.373401,11.900668,10.398509,10.233889,10.573419,11.790922,12.490558,12.30536,11.506266,10.988399,10.031544,9.9698105,10.580277,11.050131,9.97667,9.006097,8.3922,7.7680154,6.701414,4.705394,3.6765177,3.2992632,3.625074,4.420738,5.164959,5.3878818,5.5593615,6.0497923,6.7494283,7.0546613,6.48535,5.7102633,5.3330083,5.3878818,5.360445,5.3227196,5.2987127,5.3878818,5.6210938,5.9812007,5.171818,5.055212,5.0483527,5.120374,5.761707,6.310441,6.8385973,6.866034,6.464772,6.2830043,5.6039457,5.562791,6.108095,6.8763227,7.181556,6.3961806,6.1904054,6.677407,7.6171136,8.433355,7.6205435,7.2295704,6.9654922,6.8043017,7.0032177,6.8728933,6.6568294,6.5642304,6.64997,6.8145905,0.16462019,0.10288762,0.08916927,0.106317215,0.14747226,0.20577525,0.13032432,0.1097468,0.11317638,0.13032432,0.17833854,0.20577525,0.20920484,0.2194936,0.22978236,0.20920484,0.23321195,0.23664154,0.2469303,0.274367,0.29494452,0.36696586,0.48357183,0.65162164,0.8162418,0.8505377,0.99801,1.1832076,1.4953002,1.8725548,2.1229146,2.3835633,2.5996273,2.7333813,2.8156912,2.9665933,2.9871707,3.2478194,3.3678548,3.292404,3.2821152,3.3198407,3.433017,3.5118976,3.7005248,4.386442,4.166949,4.029765,4.32471,5.003768,5.5902276,5.9640527,5.9297566,6.0703697,6.1801167,5.254128,5.8817425,6.3207297,6.307011,5.8508763,5.2472687,5.909179,7.164408,7.582818,6.9792104,6.4133286,5.9743414,5.892031,5.8508763,5.552502,4.7328305,4.0229063,3.8102717,3.5770597,3.1689389,2.7813954,2.8259802,2.585909,2.0680413,1.4747226,1.1900668,1.2209331,0.9294182,0.8025235,0.8676856,0.69963586,0.8471081,1.0631721,1.2826657,1.4095604,1.3238207,1.2895249,1.155771,1.0666018,0.97057325,0.6344737,0.5624523,0.67219913,0.764798,0.75450927,0.6276145,0.61046654,0.7476501,0.7407909,0.5761707,0.53844523,0.6173257,0.7407909,0.83338976,0.864256,0.8471081,0.7613684,0.66876954,0.6310441,0.6207553,0.5178677,0.51100856,0.36010668,0.26750782,0.26064864,0.1920569,0.20577525,0.16804978,0.14061308,0.1371835,0.12689474,0.14747226,0.19548649,0.35324752,0.6173257,0.881404,1.08032,1.6084765,2.1640697,2.5653315,2.7573884,2.170929,2.037175,2.1434922,2.352697,2.5824795,3.2375305,3.7759757,4.448175,5.2301207,5.7994323,5.6656785,5.672538,6.1629686,6.8111606,6.6225333,6.2864337,6.492209,7.222711,8.255017,9.177576,9.129561,9.349055,9.925226,10.827208,11.893809,12.339656,13.035862,13.591455,13.786942,13.557159,14.013294,15.076467,15.738377,15.707511,15.415996,15.247946,14.54831,13.392539,12.024134,10.844356,10.81006,10.799771,10.88551,11.231899,12.109874,12.199042,11.924676,11.694893,11.598865,11.4033785,12.22648,12.267634,12.247057,12.500846,12.977559,12.795791,11.965831,10.88551,9.884071,9.235879,9.956093,10.556271,11.108434,11.427385,11.046701,10.576848,10.439664,10.38479,10.388221,10.6317215,10.964391,11.05356,10.748327,10.209882,9.921797,9.582268,9.451943,9.294182,9.040393,8.803751,9.328478,9.6988735,10.350495,11.317638,12.257345,12.133881,12.432255,12.566009,12.620882,13.344524,13.7938,14.452282,14.781522,14.856973,15.385129,16.019604,17.840714,19.925903,21.500084,21.911634,21.527521,21.229147,20.827885,20.306587,19.847023,20.484926,21.596113,22.789608,23.931662,25.132017,26.033998,26.483274,26.69248,26.68219,26.301506,24.572994,19.692692,14.256795,8.930646,2.4555845,1.2860953,2.860276,8.786603,12.953552,1.5193073,2.4247184,1.1797781,1.1180456,2.784825,3.9680326,3.2649672,2.8054025,2.568761,2.5619018,2.784825,2.270387,2.6853669,3.7553983,4.506478,3.2615378,4.214963,5.5387836,6.101236,5.9469047,6.3138704,6.5882373,5.717122,6.1046658,7.2295704,5.6485305,6.310441,6.2075534,6.5470824,7.31531,7.2638664,6.15268,7.7748747,8.162418,7.181556,8.508806,9.266746,9.434795,10.374502,11.382801,9.692014,9.441654,10.182446,10.700313,9.918367,6.8626046,13.320518,8.093826,3.1620796,3.2718265,5.9126086,2.7882545,3.0283258,3.3266997,2.7745364,2.8911421,3.093488,3.3644254,5.07236,6.866034,4.664239,8.056101,7.675417,5.3981705,3.2546785,3.4021509,3.450165,7.0203657,12.127021,15.6526375,13.368532,5.662249,2.2120838,1.1214751,1.0460242,1.1832076,2.352697,3.7108135,4.465323,4.6402316,5.0826488,4.931747,4.413879,4.557922,5.219832,5.07236,5.1100855,5.161529,5.113515,5.1169443,5.593657,6.48535,6.4304767,6.036074,5.7136927,5.686256,4.314421,3.9371665,4.166949,4.3521466,3.5702004,3.1483612,2.952875,3.0660512,3.40901,3.758828,3.8857226,4.513337,5.6313825,6.759717,6.931196,6.790583,6.468202,6.310441,6.4544835,6.8557453,7.1541195,7.4627824,7.579388,7.548522,7.6616983,8.134981,7.857185,7.6376915,7.6033955,7.1884155,6.6122446,6.0326443,5.892031,6.0497923,5.7754254,7.051232,7.8606143,8.3922,8.968371,10.038403,10.2236,10.436234,10.467101,10.30591,10.14129,9.352485,8.457363,7.747438,7.2192817,6.5710897,6.2967224,6.262427,6.420188,6.601956,6.5230756,6.7940125,7.534804,8.512236,9.513676,10.347065,9.719451,9.084977,8.848335,9.002667,9.132992,9.5033865,9.386781,9.050681,8.683716,8.405919,8.2481575,8.251588,8.375052,8.433355,8.090397,7.720001,7.5725293,7.284444,7.0786686,7.747438,8.052671,8.724871,8.958082,8.628842,8.323608,7.870903,7.4284863,6.924337,6.3790326,5.9331865,5.2026844,4.530485,3.5564823,2.5550427,2.4487255,2.534465,3.192946,4.722542,6.715132,8.06296,4.914599,6.2658563,10.611144,13.941273,9.760606,3.309552,1.2586586,1.0323058,1.0906088,0.89855194,0.72707254,1.2072148,3.1072063,5.144381,3.9851806,3.683377,3.3644254,7.2467184,14.483148,19.137098,19.69955,18.643238,16.016174,12.370522,8.748878,7.133542,7.534804,7.81603,6.975781,5.164959,3.7142432,6.0497923,6.23156,3.858286,4.0777793,4.9694724,3.0489032,1.8965619,2.3835633,2.6853669,2.3492675,2.4830213,2.6133456,3.8720043,9.023245,6.142391,6.7871537,7.0478024,5.720552,4.290414,4.9214582,4.8151407,5.1169443,6.029215,6.7871537,6.924337,7.8366075,8.2481575,8.049242,8.31332,8.443645,8.001227,7.7440085,7.7783046,7.596536,8.320179,8.7317295,8.923786,8.851766,8.327039,8.587687,8.601405,8.519095,8.357904,8.011517,6.7048435,6.5196457,7.0478024,7.881192,8.621983,8.090397,7.723431,7.7714453,8.217292,8.769455,9.294182,8.848335,8.587687,8.865483,9.22902,9.3079,9.537683,9.654288,9.441654,8.738589,8.519095,8.330468,7.9875093,7.507367,7.1095347,7.133542,7.1884155,6.9071894,6.1458206,4.955754,4.0880685,3.6456516,3.316411,3.0214665,2.9151495,3.2135234,3.4604537,3.6936657,3.9371665,4.201245,4.4550343,4.856296,5.895461,7.1129646,7.0889573,7.040943,7.0546613,7.1266828,7.099246,6.667118,5.8645945,5.5730796,5.6793966,6.0497923,6.550512,6.694555,6.5059276,6.39961,6.601956,7.160979,7.284444,7.6205435,8.296172,9.023245,9.126132,8.399059,8.255017,8.913498,10.4533825,12.79922,13.392539,13.72178,13.505715,12.445972,10.240748,10.120712,10.563129,11.413667,12.168177,11.955542,12.80608,12.994707,12.88839,12.737488,12.679185,11.705182,10.768905,10.367643,10.72432,11.80464,14.030442,15.618341,17.031332,17.998474,17.53891,14.479718,12.847235,13.035862,14.4145565,15.354263,14.033872,12.421966,11.156448,10.669447,11.204462,12.127021,12.644889,12.397959,11.626302,11.190743,9.619993,9.105555,9.6988735,10.556271,9.945804,8.419638,7.5519514,7.040943,6.560801,5.768566,4.65395,3.981751,4.0537724,4.698535,5.2644167,5.1992545,5.254128,5.4633327,5.7891436,6.1458206,6.169828,5.7479887,5.4976287,5.535354,5.4667625,5.4770513,5.4667625,5.48734,5.6656785,6.2144127,5.909179,5.888602,5.8817425,5.9434752,6.451054,6.835168,7.143831,7.034084,6.6122446,6.4304767,5.6142344,5.3673043,5.693115,6.2898636,6.5710897,6.2384195,6.276145,6.8797526,7.8537555,8.625413,7.48336,7.181556,7.1678376,7.1987042,7.3564653,6.944915,6.5230756,6.2898636,6.3618846,6.7665763,0.14061308,0.09259886,0.09945804,0.14747226,0.19891608,0.19891608,0.12689474,0.13032432,0.15090185,0.17490897,0.23321195,0.23321195,0.21263443,0.18862732,0.18519773,0.22635277,0.2709374,0.24007112,0.23664154,0.29151493,0.37725464,0.4355576,0.5521636,0.7099246,0.91227025,1.1763484,1.3958421,1.6839274,1.9857311,2.2463799,2.4007113,2.6956558,2.877424,2.983741,3.0454736,3.0969174,3.0866287,3.4810312,3.7691166,3.8479972,4.033195,3.9886103,3.882293,3.82399,3.974892,4.557922,4.3041325,4.0229063,4.012617,4.448175,5.4016004,6.1149545,5.6656785,5.4976287,5.7754254,5.3844523,5.8508763,6.186976,6.2144127,5.970912,5.675967,6.375603,6.4236174,6.310441,6.159539,5.7136927,5.079219,4.7431192,4.523626,4.190956,3.457024,2.9734523,2.942586,2.884283,2.668219,2.4967396,1.879414,1.4095604,1.097468,0.86082643,0.548734,0.5624523,0.4972902,0.42869842,0.40126175,0.45270553,0.58645946,0.69963586,0.8848336,1.0940384,1.1111864,1.196926,1.0048691,0.77851635,0.6379033,0.5761707,0.44927597,0.42526886,0.45956472,0.48357183,0.4081209,0.40126175,0.6927767,0.7442205,0.52472687,0.490431,0.61389613,0.8128122,0.881404,0.7888051,0.66533995,0.66191036,0.64819205,0.61389613,0.53501564,0.3806842,0.51100856,0.34295875,0.16804978,0.10288762,0.07888051,0.082310095,0.072021335,0.06859175,0.06516216,0.041155048,0.0548734,0.06516216,0.08573969,0.13375391,0.22292319,0.4115505,0.67219913,1.0734608,1.6016173,2.1880767,1.9514352,1.8656956,1.937717,2.0508933,1.9720128,2.1812177,2.8259802,3.3952916,3.7691166,4.2115335,4.4550343,4.386442,4.804852,5.645101,5.9640527,5.861165,5.90575,6.341307,7.250148,8.573969,9.47938,9.551401,9.788043,10.429376,10.957532,10.717461,11.677745,12.593445,13.077017,13.6086035,14.452282,15.258235,15.498305,15.275383,15.29253,14.685493,13.481709,12.603734,12.096155,11.146159,11.358793,11.077567,11.430815,12.449403,13.056439,12.785502,12.744347,12.672326,12.562579,12.627741,13.063298,13.1593275,13.087306,13.018714,13.121602,12.785502,12.22648,11.55771,10.89237,10.353925,11.070708,11.492548,11.818358,12.0309925,11.9040985,11.231899,11.122152,11.22161,11.30735,11.286773,11.1393,11.417097,11.379372,10.930096,10.624862,9.966381,9.523964,9.314759,9.22216,8.988949,9.506817,9.788043,10.326488,11.255906,12.377381,12.586586,13.107883,13.248496,13.214201,14.13676,13.886399,13.906977,14.147048,14.658057,15.570327,16.160215,17.823566,19.836735,21.421204,21.740154,21.688711,21.541239,21.187992,20.738716,20.519222,20.755863,21.640697,22.751883,24.02426,25.759632,27.217207,27.807095,27.649334,27.086882,26.702768,24.912523,17.058767,8.707723,3.0660512,0.94999576,1.0768905,1.6564908,2.0577524,1.8862731,0.9842916,0.432128,0.59331864,2.369845,5.020916,6.186976,4.1635194,3.1380725,2.177788,1.214074,1.0254467,1.6153357,2.4967396,3.1483612,3.3747141,3.309552,4.98662,5.8062916,6.0326443,5.857735,5.4153185,5.9160385,6.557371,7.3050213,7.377043,5.2266912,6.8763227,7.2604365,6.550512,5.518206,5.5079174,6.1046658,7.2467184,7.73372,7.915488,9.709162,8.615124,8.772884,10.607714,12.202472,9.301042,10.528833,9.89436,9.506817,8.937505,5.2301207,12.456262,8.224151,3.415869,3.1963756,7.040943,3.0557625,2.7299516,3.4638834,3.450165,1.646202,3.758828,3.0626216,5.23698,8.81404,5.192395,5.1821065,5.0277753,4.8254294,4.479041,3.7211025,4.081209,8.06296,13.1421795,15.230798,8.687145,2.5893385,1.7525192,2.177788,2.1023371,1.9994495,3.07634,3.74168,3.9851806,4.0709205,4.530485,4.214963,4.170378,4.537344,5.1169443,5.3432975,5.5422134,5.521636,5.717122,6.1904054,6.6053853,7.5039372,7.3873315,6.9517736,6.550512,6.210983,4.705394,4.1463714,4.2526884,4.3178506,3.2512488,2.8019729,2.8911421,3.223812,3.6353626,4.0777793,3.899441,4.187526,4.839148,5.446185,5.2781353,5.895461,6.166398,6.327589,6.447624,6.4236174,6.5299344,6.608815,6.619104,6.550512,6.4304767,7.130112,7.421627,7.346176,6.866034,5.8680243,5.6485305,5.8234396,6.029215,6.0532217,5.830299,7.4765005,8.086967,8.549961,9.22216,9.956093,10.38479,11.146159,11.38966,10.995257,10.573419,9.767465,9.006097,8.210432,7.431916,6.869464,6.56766,6.680836,6.776865,6.824879,7.1884155,7.407909,8.004657,8.707723,9.414218,10.189304,9.582268,9.057541,8.9100685,9.153569,9.513676,9.832627,9.784613,9.554831,9.266746,8.961512,9.318189,9.136421,8.738589,8.131552,7.010077,6.574519,6.9689217,6.5642304,5.4839106,5.5833683,6.2041235,7.1129646,7.8606143,8.416207,9.184435,8.947794,8.7283,8.155559,7.39762,7.160979,6.948344,6.341307,5.120374,3.6353626,2.784825,2.9563043,3.5702004,5.267846,7.2638664,7.3221693,6.186976,10.957532,18.073925,20.903336,9.740028,3.1723683,1.2003556,1.255229,1.6942163,1.8142518,1.2277923,2.2292318,5.8234396,9.081548,5.144381,4.938606,3.9543142,7.5690994,15.731518,22.95423,25.907104,23.715597,19.19197,14.363112,10.4533825,8.577398,8.820899,8.988949,8.052671,6.125243,4.705394,8.724871,9.355915,5.127233,1.9239986,4.6779575,3.6319332,2.7951138,3.316411,3.4981792,2.8465576,2.9974594,3.0043187,2.8911421,3.6353626,5.188966,6.5196457,6.4819202,5.195825,4.064061,4.65395,5.0895076,5.2575574,5.4153185,6.193835,6.3378778,7.250148,7.9600725,8.217292,8.508806,8.56368,8.117833,7.747438,7.599966,7.414768,9.22902,9.56512,9.506817,9.383351,8.772884,8.237869,8.471081,8.81747,8.999237,9.119273,7.9017696,7.250148,7.3118806,7.81603,8.093826,8.004657,8.258447,8.793462,9.506817,10.254466,9.451943,8.793462,8.995808,9.89093,10.432805,10.340206,10.079557,9.616563,9.098696,8.879202,8.522525,8.591117,8.539673,8.200144,7.8023114,7.5210853,7.1129646,6.495639,5.6828265,4.8117113,3.5599117,3.018037,2.8637056,2.8534167,2.7916842,3.1517909,3.2512488,3.508468,3.8308492,3.6010668,3.8891523,3.8891523,4.588788,5.8988905,6.6533995,6.948344,7.1129646,7.301592,7.514226,7.599966,6.931196,6.6225333,6.694555,6.975781,7.130112,7.6376915,7.5588107,7.250148,7.0752387,7.421627,8.2310095,8.690575,8.868914,8.80718,8.536243,8.176137,8.258447,9.249598,11.214751,13.797231,13.368532,12.857523,13.313659,13.536582,10.117283,9.654288,9.777754,10.63858,11.688034,11.667457,12.524854,12.548861,11.80464,10.779194,10.38479,9.541112,9.050681,9.414218,10.600855,12.065289,14.46943,16.252815,17.840714,18.969048,18.70154,15.772673,13.790371,13.190193,13.591455,13.821238,13.022143,12.648318,11.859513,10.943813,11.331357,11.2250395,11.677745,12.05843,11.921246,10.984968,9.314759,8.207003,8.652849,9.928656,9.599416,8.1384115,7.500508,7.1678376,6.8900414,6.684266,5.6313825,4.8905916,4.6127954,4.773986,5.1992545,4.7774153,4.4756117,4.2869844,4.2938433,4.65395,5.3261495,5.5662203,5.4839106,5.2506986,5.1066556,5.055212,5.24041,5.501058,5.8817425,6.608815,6.81802,6.759717,6.800872,6.941485,6.8454566,7.0786686,6.7459984,6.351596,6.159539,6.169828,5.645101,5.305572,5.3844523,5.8165803,6.228131,6.684266,6.8763227,7.099246,7.3393173,7.281014,5.977771,5.926327,6.307011,6.6636887,6.8900414,6.5299344,6.101236,5.720552,5.6348124,6.2212715,0.15090185,0.16462019,0.15090185,0.16119061,0.18519773,0.1371835,0.17490897,0.28465575,0.30866286,0.23321195,0.18176813,0.23321195,0.25378948,0.26407823,0.28808534,0.33609957,0.31209245,0.28808534,0.28808534,0.34295875,0.48700142,0.72021335,0.7407909,0.8745448,1.1866373,1.4815818,1.8588364,2.153781,2.3252604,2.4384367,2.6716487,3.0111778,3.4192986,3.5839188,3.450165,3.2203827,3.450165,3.6387923,3.899441,4.2046742,4.3624353,4.280125,4.0846386,4.057202,4.2526884,4.4859004,4.4241676,4.389872,4.629943,5.219832,6.0737996,6.121814,5.7136927,5.212973,4.8940215,4.945465,6.018926,5.830299,5.127233,4.698535,5.3707337,5.5559316,5.5079174,5.312431,4.9934793,4.5167665,3.9303071,3.7005248,3.2512488,2.5790498,2.2738166,2.054323,2.2909644,2.4247184,2.3389788,2.3492675,1.5090185,0.939707,0.7373613,0.70649505,0.36696586,0.32924038,0.34638834,0.36696586,0.39097297,0.48700142,0.47671264,0.5007198,0.61046654,0.78194594,0.91569984,0.805953,0.7407909,0.7099246,0.6756287,0.5658819,0.41840968,0.490431,0.5144381,0.42183927,0.33609957,0.4938606,0.45956472,0.42869842,0.48014224,0.5658819,0.7339317,0.8505377,0.7613684,0.5418748,0.5178677,0.50757897,0.5418748,0.51100856,0.3806842,0.19891608,0.11317638,0.072021335,0.0548734,0.041155048,0.030866288,0.041155048,0.037725464,0.037725464,0.041155048,0.030866288,0.041155048,0.044584636,0.05144381,0.06516216,0.07545093,0.1371835,0.28122616,0.4938606,0.7613684,1.0528834,1.3821237,1.4095604,1.4232788,1.5570327,1.8005334,1.9239986,2.1263442,2.3424082,2.6236343,3.1723683,3.9543142,4.187526,4.3521466,4.681387,5.1580997,5.720552,5.7411294,5.686256,5.878313,6.4990683,7.599966,8.495089,9.270175,10.014396,10.834066,10.381361,11.22161,11.763485,11.873232,12.864383,14.109323,14.784951,14.634049,14.109323,14.390549,13.413116,12.88496,12.315649,11.705182,11.537132,11.341646,11.327928,11.561139,12.065289,12.847235,13.018714,13.289652,13.55373,13.701202,13.642899,13.519434,13.2862215,13.173045,13.111313,12.758065,12.586586,12.5145645,12.363663,12.123591,11.979549,11.7086115,11.753197,12.082437,12.528283,12.771784,12.576297,12.644889,12.754636,12.569438,11.64345,11.38623,11.396519,11.156448,10.624862,10.206452,10.539123,10.436234,10.151579,9.794902,9.369633,9.80862,10.127572,10.734609,11.670886,12.634601,12.21962,12.812939,13.622321,14.38026,15.319967,15.100473,14.79867,14.7369375,14.973578,15.289101,16.777542,18.02934,19.20912,19.9602,19.408035,19.483486,20.004784,20.663265,21.10568,20.934202,20.508932,21.565247,23.328054,25.063425,26.078583,28.287237,29.49788,29.480734,28.558174,27.618467,25.409813,15.902997,6.776865,1.7902447,0.77851635,1.3169615,1.9514352,3.8377085,4.996909,0.33609957,0.4081209,2.3389788,2.9803114,1.7422304,0.59674823,1.961724,4.4996185,4.465323,2.136633,1.8313997,3.1620796,4.4275975,3.8308492,2.4315774,4.166949,4.7774153,4.0880685,4.557922,5.672538,3.9508848,5.171818,6.5230756,6.5813785,5.6313825,5.6313825,6.7528577,6.4407654,6.0497923,6.228131,6.910619,6.8626046,8.049242,8.673427,8.460793,8.683716,6.094377,7.936065,10.203023,10.6317215,8.7283,12.085866,10.048691,10.079557,11.406808,5.0346346,8.601405,7.8983397,4.6916757,2.4007113,6.0875177,2.1812177,1.5810398,3.2581081,4.671098,1.7559488,2.7573884,2.959734,7.720001,13.104454,5.888602,6.025785,4.756838,5.3261495,7.2364297,6.2727156,6.368744,8.865483,10.597425,9.832627,6.2555676,2.5824795,2.4315774,3.1895163,3.4638834,3.0969174,3.3061223,3.7965534,3.4055803,2.551613,3.234101,3.8205605,4.2698364,4.8425775,5.5250654,6.025785,6.1972647,6.495639,6.917478,7.3530354,7.582818,8.64599,8.158989,7.3255987,6.5779486,5.6005163,4.6127954,4.417309,4.3521466,4.0057583,3.2512488,2.9563043,3.3061223,3.7794054,3.99204,3.6627994,3.5050385,3.7759757,4.40359,5.055212,5.1409516,5.8371577,6.2041235,6.228131,6.046363,5.936616,6.0703697,5.7102633,5.4667625,5.586798,5.967482,6.4407654,7.1369715,7.3701835,6.831738,5.6005163,6.0154963,6.090947,6.0669403,6.1629686,6.5779486,7.5279446,8.251588,9.112414,9.880642,9.736599,9.932085,10.2921915,10.772334,11.231899,11.427385,10.511685,9.880642,9.294182,8.639131,7.9189177,7.966932,8.189855,8.213862,8.117833,8.423067,8.203573,8.2481575,8.738589,9.421077,9.626852,9.273604,9.304471,9.451943,9.56512,9.613133,9.637141,9.6988735,9.873782,10.045261,9.887501,10.998687,10.762046,10.213311,9.352485,7.157549,5.813151,6.0806584,6.680836,6.999788,7.1095347,7.0375133,6.835168,6.8283086,7.2432885,8.210432,8.673427,9.016385,8.700864,8.025234,8.1487,9.050681,8.580828,7.0752387,5.113515,3.5393343,3.625074,4.2252517,5.3707337,7.613684,12.006986,12.936404,12.572867,16.314548,19.336014,6.591667,2.503599,1.3786942,1.7936742,2.8396983,4.1189346,2.5070283,5.5490727,8.182996,9.589127,13.152468,13.690913,9.668007,6.475061,6.8385973,10.820349,19.143957,16.235666,12.867812,12.590015,11.732618,9.438225,7.7748747,7.500508,7.870903,6.636252,4.07435,4.5784993,5.638242,5.7102633,4.1943855,3.1106358,3.6627994,3.8925817,3.5702004,4.180667,3.5702004,3.666229,4.0674906,4.331569,3.9508848,3.6593697,3.0729103,3.0489032,3.649081,4.149801,4.5030484,5.453044,5.5319247,4.914599,5.4016004,5.6210938,6.217842,7.1266828,7.9463544,7.936065,7.8606143,7.98065,7.956643,7.658269,7.1712675,8.172707,9.054111,9.517105,9.39707,8.652849,8.357904,9.026674,9.174147,8.680285,8.790032,8.213862,7.5588107,7.2775846,7.2021337,6.5299344,6.468202,7.654839,8.868914,9.458802,9.338767,9.191295,9.72288,10.388221,10.738038,10.422516,9.750318,9.14328,8.800322,8.735159,8.759167,7.548522,7.5690994,7.5759587,6.7528577,4.715683,4.8117113,5.0655007,4.729401,4.105216,4.530485,3.2992632,2.4967396,2.201795,2.2669573,2.3046827,2.633923,2.8705647,3.0900583,3.3198407,3.5393343,3.7108135,3.789694,4.139512,4.835718,5.675967,6.1766872,6.7219915,7.051232,7.1952744,7.4765005,7.9909387,7.936065,8.093826,8.471081,8.299602,8.251588,7.8091707,7.2124224,6.8111606,7.0786686,7.8983397,8.707723,8.711152,8.536243,10.206452,9.585697,8.268735,8.467651,10.539123,12.953552,13.735497,12.476839,11.492548,11.190743,10.055551,9.163857,9.325048,9.918367,10.484249,10.72775,10.909517,11.074138,10.696883,9.9698105,9.81205,9.493098,8.937505,9.458802,10.830637,11.30735,12.943263,14.640909,16.077906,17.151367,18.005335,17.322845,15.018164,13.327377,13.063298,13.625751,12.809509,12.504276,12.020704,11.355364,11.183885,9.4862385,9.211872,10.264755,11.348505,9.932085,9.102125,9.335337,10.096705,10.525404,9.414218,8.803751,8.460793,8.289313,8.06296,7.414768,6.550512,5.8200097,5.195825,4.773986,4.7602673,4.2595477,3.292404,3.0660512,3.642222,3.9200184,4.396731,5.103226,5.2781353,4.9351764,4.835718,4.7774153,4.7602673,5.07236,5.7925735,6.8043017,7.0135064,7.2192817,7.798882,8.261876,7.2467184,7.442205,7.034084,6.5333643,6.23156,6.193835,6.5985265,6.461343,6.5882373,7.143831,7.6445503,7.8263187,7.606825,7.298162,6.914048,6.193835,5.3878818,5.1683884,5.0277753,4.962613,5.4633327,6.0978065,5.73427,5.3501563,5.219832,4.914599,0.17833854,0.17833854,0.16119061,0.16804978,0.1920569,0.17490897,0.24007112,0.29837412,0.29837412,0.26064864,0.28122616,0.30866286,0.29837412,0.28122616,0.28465575,0.32238123,0.32924038,0.37039545,0.4664239,0.58988905,0.64819205,0.77165717,0.8745448,1.0048691,1.2243627,1.6153357,1.9137098,2.177788,2.352697,2.5310357,2.9391565,3.5633414,3.6147852,3.508468,3.4433057,3.415869,3.5873485,3.7965534,3.9371665,4.091498,4.523626,4.32128,4.32128,4.420738,4.4447455,4.170378,4.0503426,4.3658648,4.8494368,5.3090014,5.645101,5.4324665,5.1821065,4.8494368,4.722542,5.442755,5.7479887,5.5490727,5.3158607,5.1512403,4.7979927,5.1855364,5.212973,5.0655007,4.7774153,4.2252517,3.5118976,3.2272418,2.7951138,2.1846473,1.9068506,1.8348293,2.1160555,2.2841053,2.1640697,1.8725548,1.196926,0.83338976,0.6962063,0.6344737,0.4389872,0.37382504,0.33952916,0.31895164,0.32581082,0.40126175,0.41840968,0.4355576,0.4972902,0.5693115,0.53844523,0.53501564,0.548734,0.5761707,0.5761707,0.4664239,0.7613684,0.6276145,0.4424168,0.37039545,0.37382504,0.39440256,0.3566771,0.35324752,0.4355576,0.58988905,0.7510797,0.7888051,0.7510797,0.6859175,0.65162164,0.4355576,0.29494452,0.19891608,0.13375391,0.07545093,0.030866288,0.01371835,0.010288762,0.006859175,0.006859175,0.006859175,0.030866288,0.030866288,0.006859175,0.006859175,0.006859175,0.010288762,0.010288762,0.020577524,0.05144381,0.0548734,0.1097468,0.216064,0.36353627,0.5418748,0.89855194,1.1180456,1.2449403,1.3238207,1.371835,1.6016173,1.99602,2.2738166,2.4007113,2.5893385,2.9700227,3.3198407,3.690236,4.125794,4.681387,5.2438393,5.5730796,5.9434752,6.444195,6.989499,7.548522,8.069819,9.084977,10.422516,11.211322,11.30735,11.317638,11.321068,11.4205265,11.71547,12.912396,13.900118,13.7526455,12.9638405,13.450842,13.13532,13.491997,13.55373,12.946692,11.876661,12.188754,11.873232,11.660598,12.05843,13.337666,13.536582,14.373401,14.760944,14.490007,14.21564,14.191633,14.13676,14.212211,14.38369,14.428274,14.373401,14.267084,14.061309,13.941273,14.321958,13.622321,13.032433,12.830087,13.001566,13.234778,12.7272,13.070158,13.2690735,12.908967,12.168177,12.017275,11.835506,11.773774,11.64345,10.916377,11.509696,11.365653,10.984968,10.659158,10.456812,10.357354,11.026124,12.085866,13.145609,13.817808,13.491997,13.642899,14.222499,15.114192,16.163645,15.913286,15.638919,15.350834,15.405707,16.523752,17.87501,18.11165,18.317427,18.427174,17.223389,17.532051,18.492336,19.147387,19.349733,19.764713,19.637817,20.601532,22.419212,24.645016,26.627317,28.35583,29.809975,30.629646,30.430729,28.777668,25.951689,18.331144,9.496528,2.7368107,1.0117283,0.805953,0.77508676,1.3958421,1.8999915,0.26407823,0.83338976,1.3581166,1.471293,1.8485477,4.1943855,5.113515,4.098357,2.9151495,2.4384367,2.6613598,3.0043187,3.4535947,3.192946,2.8259802,4.372724,3.8205605,3.7553983,5.086078,6.6568294,5.2575574,6.077229,6.6533995,7.0752387,7.5588107,8.436785,7.257007,7.3050213,7.425057,7.3221693,7.548522,6.756287,7.5245147,7.9463544,7.888051,8.988949,8.7145815,9.156999,9.712592,10.120712,10.460241,13.917266,12.123591,9.925226,8.567109,5.720552,6.5779486,7.970361,6.615674,3.3644254,3.1826572,1.8142518,2.5893385,3.4810312,3.340418,1.8759843,2.2223728,3.4295874,5.3090014,6.893471,6.427047,8.80718,6.1972647,5.768566,8.525954,9.297611,9.630281,9.088407,6.927767,4.647091,5.9640527,3.4021509,3.5530527,4.0057583,3.8137012,3.4776018,3.683377,4.232111,4.15666,3.3815732,2.7470996,3.3815732,4.149801,4.962613,5.8234396,6.831738,5.950334,6.6053853,7.349606,7.6651278,7.9875093,8.385342,7.610255,6.684266,5.98463,5.223262,4.65395,4.8151407,4.996909,4.722542,3.7519686,3.3198407,3.4947495,3.6593697,3.6696587,3.858286,3.7965534,3.7039545,3.858286,4.2183924,4.420738,4.746549,4.996909,5.038064,4.99005,5.24041,5.305572,5.2506986,5.2301207,5.3981705,5.892031,6.447624,6.9346256,7.0752387,6.694555,5.7479887,5.8405876,5.8337283,5.9126086,6.135532,6.4544835,7.699424,8.31332,8.89635,9.547972,9.870353,9.527394,9.72288,10.124143,10.607714,11.283342,11.080997,10.47396,9.863494,9.366203,8.820899,8.872343,8.755736,8.570539,8.368194,8.155559,7.8949103,7.6959944,7.840037,8.255017,8.529384,8.488229,8.862054,8.738589,8.14527,8.038953,8.279024,8.707723,9.3079,9.97667,10.521975,11.290202,11.111863,11.05356,11.129011,10.268185,8.759167,8.107545,8.30646,8.930646,9.136421,9.424506,9.102125,8.141841,7.298162,8.086967,8.512236,9.287323,9.794902,9.863494,9.760606,9.911508,9.80862,9.194724,7.822889,5.470192,4.479041,5.425607,6.636252,7.5416627,8.663138,8.488229,6.6705475,7.459353,9.513676,5.909179,2.9220085,2.1469216,2.0508933,2.5413244,4.98662,4.2252517,12.010415,14.308239,11.183885,16.79126,13.869251,14.63062,13.039291,8.597976,6.3378778,15.923574,15.145059,10.81006,7.8194594,9.170717,7.997798,9.194724,10.467101,10.2236,7.56567,6.8866115,4.184097,3.1243541,4.2389703,4.9420357,3.7553983,3.882293,3.9028704,3.782835,4.852866,4.770556,4.928317,5.411889,5.6348124,4.3795834,4.506478,3.5359046,3.1895163,3.7348208,3.99204,4.2766957,5.23698,5.693115,5.5833683,5.9743414,5.5422134,5.48734,5.8988905,6.4373355,6.334448,6.6053853,6.5950966,6.893471,7.473071,7.6959944,8.131552,8.447074,8.796892,8.97866,8.419638,8.23444,8.745448,8.937505,8.601405,8.351046,8.213862,8.093826,8.158989,8.22758,7.750868,7.8846216,8.429926,9.253027,10.14129,10.789482,11.4754,12.133881,12.247057,11.917816,11.873232,10.676306,9.561689,8.834618,8.4093485,7.8194594,7.3427467,8.268735,8.759167,7.514226,3.7862647,2.7916842,2.952875,3.0729103,2.8225505,2.760818,2.486451,1.8554068,1.471293,1.4335675,1.3649758,1.8108221,2.3424082,2.8637056,3.357566,3.8685746,4.0194764,4.0503426,4.2183924,4.605936,5.113515,5.3330083,6.416758,7.116394,7.1849856,7.380472,7.226141,7.0375133,7.274155,7.829748,8.018375,7.8434668,7.7885933,7.73029,7.822889,8.484799,8.803751,8.851766,8.690575,8.796892,10.048691,8.742019,7.5039372,7.963502,10.131001,12.394529,13.536582,12.205902,10.899229,10.593996,10.72775,10.422516,10.714031,10.823778,10.618003,10.618003,10.264755,9.877212,9.321619,8.7317295,8.505377,8.412778,8.292743,8.721441,9.743458,10.89237,12.4974165,13.869251,15.155347,16.208231,16.564907,17.082775,15.079896,12.96727,12.082437,12.662037,12.929544,13.004995,12.706621,12.1921835,11.952112,11.934964,11.749766,11.537132,10.960961,9.211872,8.587687,9.098696,9.798331,10.196163,10.257896,9.019815,8.505377,8.399059,8.337327,7.915488,7.1781263,5.7891436,4.6848164,4.0880685,3.5290456,3.3987212,2.7299516,2.5173173,2.976882,3.532475,4.046913,4.5647807,4.5647807,4.1155047,3.8617156,4.297273,4.523626,4.822,5.422178,6.5230756,6.948344,7.706283,8.40249,8.519095,7.4181976,7.8674736,7.6033955,7.205563,7.06495,7.390761,7.15069,6.7631464,6.773435,7.2604365,7.840037,7.7885933,7.8537555,7.822889,7.5210853,6.8283086,6.433906,6.1492505,5.7102633,5.288424,5.4736214,5.9160385,5.501058,4.98662,4.722542,4.681387,0.2194936,0.18176813,0.14404267,0.13032432,0.14061308,0.17490897,0.23321195,0.26407823,0.28808534,0.32238123,0.39783216,0.32581082,0.39440256,0.47328308,0.48357183,0.4115505,0.4081209,0.4355576,0.5555932,0.72364295,0.7956643,0.88826317,0.9568549,0.9911508,1.0666018,1.3272504,1.8073926,2.1674993,2.469303,2.767677,3.117495,3.474172,3.6182148,3.683377,3.7279615,3.7279615,3.9680326,4.091498,4.139512,4.2423997,4.616225,4.523626,4.479041,4.4687524,4.434457,4.273266,4.081209,4.180667,4.6265135,5.192395,5.3570156,5.2438393,5.079219,4.914599,4.8288593,4.928317,5.2438393,5.164959,5.161529,5.1821065,4.65395,5.0929375,5.15467,4.863155,4.338428,3.8034124,3.1312134,2.6956558,2.352697,2.0886188,2.0268862,1.9754424,2.1160555,2.170929,2.0063086,1.6187652,1.1660597,0.89169276,0.71678376,0.5796003,0.42183927,0.34638834,0.33609957,0.31895164,0.29837412,0.32581082,0.37382504,0.42183927,0.44927597,0.432128,0.34981793,0.3841138,0.39783216,0.45956472,0.548734,0.53501564,0.6379033,0.47328308,0.34638834,0.36696586,0.42869842,0.3566771,0.3566771,0.50757897,0.7682276,0.9877212,0.91227025,0.8745448,0.77508676,0.58988905,0.3841138,0.2194936,0.12003556,0.058302987,0.0274367,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.01371835,0.044584636,0.09945804,0.17490897,0.25721905,0.490431,0.7407909,1.0323058,1.2758065,1.2380811,1.5330256,1.8828435,2.0577524,2.095478,2.3046827,2.7299516,3.2718265,3.6525106,3.9440255,4.554492,5.086078,5.669108,6.217842,6.694555,7.1369715,7.874333,8.529384,9.331907,10.329918,11.434244,12.034423,11.760056,11.592006,11.698323,11.4376745,12.181894,13.059869,13.330807,13.066729,13.1421795,13.529722,13.910407,13.759505,12.9809885,11.897239,11.958971,11.660598,11.705182,12.295071,13.166186,13.841815,15.199932,15.820687,15.477728,15.127911,14.688923,14.438563,14.743796,15.409137,15.680074,15.734947,15.145059,14.452282,14.061309,14.222499,14.088745,13.560589,13.313659,13.37882,13.149038,12.528283,12.665466,12.665466,12.329367,12.161317,12.308789,12.394529,12.55229,12.562579,11.852654,12.517994,12.590015,12.22305,11.595435,10.899229,10.72775,11.849225,13.193623,14.119612,14.424845,14.195063,14.582606,15.062748,15.614912,16.746675,17.04162,16.691803,16.427725,16.691803,17.645227,18.523201,18.362011,18.248835,18.248835,17.401728,17.833855,18.36544,18.506054,18.348293,18.564358,18.931322,20.052797,21.733295,23.76361,25.913963,27.971716,29.412142,30.718815,31.216105,29.076042,26.099161,21.136547,13.937843,6.368744,2.4144297,1.0700313,0.4424168,0.41840968,0.7133542,0.8676856,2.2155135,2.3321195,2.3252604,3.2409601,6.077229,5.007198,3.8925817,3.875434,4.870014,5.5593615,4.6848164,4.2766957,4.547633,5.2472687,5.6793966,3.8548563,5.377593,6.3618846,5.7822843,5.4667625,6.420188,6.7391396,7.332458,8.388771,9.3764925,8.375052,8.81747,8.711152,7.6959944,7.0375133,7.517656,9.026674,9.678296,9.225591,9.071259,9.517105,9.355915,9.746887,10.823778,11.691463,13.083877,13.275933,11.115293,7.5210853,5.4599032,6.433906,6.6225333,5.8680243,4.149801,1.5947582,1.2380811,2.037175,3.1209247,3.6696587,2.9151495,2.4761622,4.5647807,6.2212715,6.8866115,8.436785,7.870903,7.0478024,8.069819,10.6488695,12.116733,7.781734,6.433906,5.4941993,4.6848164,6.046363,4.266407,4.6573796,4.6882463,3.9371665,4.091498,3.6627994,3.40901,3.1895163,3.0283258,3.1106358,4.173808,5.0346346,5.504488,5.6965446,6.018926,5.4941993,6.5882373,7.5725293,7.8606143,8.004657,7.5416627,6.677407,5.90232,5.3227196,4.650521,4.7362604,4.8940215,4.9214582,4.6848164,4.105216,3.6113555,3.4878905,3.4810312,3.525616,3.7313912,3.6868064,3.5873485,3.5564823,3.6387923,3.7759757,4.1463714,4.3692946,4.3795834,4.4413157,5.1580997,5.219832,5.0586414,5.020916,5.24041,5.6176643,5.950334,6.200694,6.1732574,5.844017,5.353586,5.56965,5.796003,6.046363,6.2727156,6.358455,7.4010496,8.131552,8.687145,9.167287,9.626852,9.585697,9.650859,9.9869585,10.590566,11.273054,11.05699,10.542552,9.9869585,9.510246,9.074688,9.153569,9.115844,8.999237,8.755736,8.261876,7.390761,7.181556,7.3393173,7.6171136,7.805741,7.599966,7.8606143,7.7920227,7.4696417,7.8263187,7.9875093,8.241299,8.580828,9.009526,9.554831,9.925226,9.942374,10.257896,10.7586155,10.569988,9.798331,8.7145815,8.309891,8.769455,9.469091,9.921797,10.017825,9.386781,8.515666,8.762596,8.508806,8.597976,8.882631,9.2153015,9.465661,9.626852,9.119273,8.64256,8.155559,6.8557453,6.464772,7.2295704,8.258447,8.868914,8.597976,7.9463544,6.1561093,4.8940215,4.98662,6.4133286,3.309552,2.6167753,2.4658735,2.3321195,3.0523329,2.6853669,8.742019,10.014396,6.9517736,11.677745,7.98065,10.854645,12.46998,9.911508,5.192395,15.37827,12.939834,8.484799,7.0718093,8.22758,7.0203657,9.626852,12.3533745,12.195613,6.8454566,5.4599032,3.7211025,2.9185789,3.6147852,5.638242,3.875434,3.8960114,4.1943855,4.3349986,4.945465,5.5387836,5.6519604,5.977771,6.1561093,4.7979927,5.219832,4.3795834,3.74168,3.8925817,4.5647807,4.8322887,5.4907694,6.0840883,6.540223,7.1712675,6.1492505,5.6142344,5.4667625,5.5079174,5.4599032,6.252138,6.2418494,6.5642304,7.366754,7.7920227,8.06296,8.076678,8.06639,8.114404,8.152129,8.98209,9.640571,9.784613,9.506817,9.349055,8.875772,8.772884,8.8929205,9.122703,9.338767,9.945804,10.072699,10.741467,11.756626,11.72233,11.859513,11.677745,11.55428,11.509696,11.211322,9.609704,8.299602,7.2947326,6.4579134,5.48734,5.40503,6.9654922,8.81404,8.584257,2.8877127,1.6530612,1.529596,1.7833855,1.9651536,1.8965619,1.7799559,1.4061309,1.1832076,1.2072148,1.2483698,1.5261664,1.961724,2.6133456,3.3884325,4.0263357,4.273266,4.32471,4.3933015,4.6608095,5.2575574,5.0449233,5.641671,6.3035817,6.64997,6.660259,6.4887795,6.355026,6.677407,7.3358874,7.675417,7.747438,8.004657,8.152129,8.340756,9.163857,9.469091,9.458802,9.112414,8.930646,9.918367,8.381912,7.8331776,8.553391,10.233889,11.979549,13.262215,12.932974,11.852654,11.187314,12.377381,12.020704,11.667457,11.38623,11.063849,10.388221,9.688584,9.31133,8.759167,8.114404,8.069819,8.368194,8.577398,9.266746,10.508256,11.849225,13.3033695,14.222499,15.090185,15.618341,14.767803,15.343974,14.435134,12.452832,10.655728,11.177026,11.989838,12.082437,12.041282,11.96926,11.478829,12.072148,12.161317,11.537132,10.528833,10.031544,9.441654,9.283894,9.321619,9.585697,10.347065,9.945804,9.095266,8.669997,8.7317295,8.525954,7.7748747,5.9331865,4.629943,4.15323,3.457024,3.3850029,2.983741,2.7059445,2.7368107,2.983741,3.532475,3.9303071,4.0263357,3.8479972,3.6079261,4.197815,4.804852,5.3432975,5.9571934,7.0203657,7.73372,8.368194,8.608265,8.292743,7.425057,7.682276,8.05953,8.083538,7.9429245,8.460793,8.107545,7.5519514,7.1781263,7.1884155,7.596536,7.7851634,8.268735,8.573969,8.375052,7.455923,7.0958166,6.5024977,5.830299,5.377593,5.6073756,5.761707,5.4599032,5.1409516,4.98662,4.9077396,0.18862732,0.17833854,0.15433143,0.12689474,0.12003556,0.18519773,0.2503599,0.28808534,0.34295875,0.4355576,0.59331864,0.5521636,0.5178677,0.5178677,0.52815646,0.48014224,0.48014224,0.52472687,0.64476246,0.7990939,0.8505377,0.91227025,0.91227025,0.88826317,0.9328478,1.1797781,1.786815,2.1743584,2.5447538,2.9494452,3.275256,3.3987212,3.6456516,3.8685746,4.016047,4.108646,4.4550343,4.6093655,4.715683,4.7808447,4.65395,4.5990767,4.355576,4.2286816,4.2252517,4.033195,3.9646032,4.040054,4.448175,4.9934793,5.099797,5.295283,5.425607,5.4770513,5.3330083,4.787704,4.979761,5.113515,5.2438393,5.23698,4.746549,4.9180284,4.763697,4.307562,3.673088,3.1140654,2.6716487,2.4624438,2.3046827,2.1503513,2.1057668,2.0989075,2.1194851,2.0268862,1.7936742,1.4781522,1.1317638,0.864256,0.67219913,0.52815646,0.36696586,0.30866286,0.29494452,0.29151493,0.28122616,0.2777966,0.34295875,0.4046913,0.4081209,0.34638834,0.2709374,0.28808534,0.31209245,0.37382504,0.44927597,0.45613512,0.4115505,0.31209245,0.29837412,0.37725464,0.40126175,0.33266997,0.4664239,0.7922347,1.1523414,1.2620882,1.0563129,0.89169276,0.66876954,0.38754338,0.15090185,0.08916927,0.041155048,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.041155048,0.08916927,0.18176813,0.24007112,0.4355576,0.77165717,1.0940384,1.0940384,1.3375391,1.5604624,1.6599203,1.7696671,2.2566686,3.093488,3.7622573,4.2355404,4.5853586,5.0106273,5.5147767,6.1492505,6.677407,6.9792104,7.051232,8.069819,8.882631,9.589127,10.343636,11.372512,12.123591,12.024134,12.003556,12.171606,11.828648,11.962401,12.517994,12.946692,12.847235,11.955542,12.994707,13.443983,13.313659,12.740917,11.979549,11.945253,11.427385,11.46854,12.229909,12.987847,14.188204,15.494876,16.03675,15.731518,15.316538,14.846684,14.764374,15.498305,16.571766,16.619781,16.04018,15.069608,14.263655,13.869251,13.810948,14.291091,14.027013,13.718349,13.560589,13.21763,12.583157,12.493987,12.253916,11.80121,11.71547,12.147599,12.679185,13.118172,13.231348,12.744347,13.073587,13.423406,13.231348,12.404818,11.321068,11.228469,12.281353,13.426835,14.174485,14.613472,14.534592,15.083325,15.481158,15.782962,16.877,17.36057,17.12736,17.113642,17.518333,17.809847,18.20082,18.344864,18.307138,18.094503,17.658945,17.909306,18.169954,18.169954,17.981327,18.025911,18.307138,19.411465,20.934202,22.61127,24.302057,26.68219,28.300955,29.734524,30.303835,28.10204,25.51613,21.959648,15.87899,8.7283,4.9351764,2.935727,1.471293,0.6276145,0.5041494,1.196926,2.2738166,2.9940298,3.5770597,4.3590055,5.802862,4.6848164,5.9571934,7.164408,7.4799304,7.73372,8.052671,7.5931067,7.1198235,6.776865,6.094377,4.9488945,6.608815,6.9071894,5.593657,6.307011,7.0032177,7.0306544,7.4456344,8.388771,9.078118,9.465661,10.024684,9.6988735,8.786603,8.954653,9.97324,10.556271,10.7757635,10.511685,9.47595,9.709162,9.650859,10.182446,11.321068,12.199042,12.411677,14.229359,12.435684,7.380472,4.9831905,7.0546613,6.3001523,5.48734,4.770556,1.6804979,1.1660597,1.5021594,2.620205,3.7176728,3.2615378,4.2286816,5.593657,6.0737996,6.2864337,8.755736,5.5730796,6.355026,9.362774,11.880091,10.206452,6.042933,5.857735,6.64997,6.948344,6.8454566,4.931747,5.689686,5.435896,3.9646032,4.5682106,3.7039545,3.1895163,2.8739944,2.9048605,3.6970954,4.8322887,5.504488,5.802862,5.802862,5.579939,5.6485305,6.5779486,7.346176,7.6171136,7.7371492,6.7219915,6.111525,5.5662203,5.0277753,4.7191124,4.99005,4.8768735,4.7328305,4.6402316,4.4275975,4.046913,3.841138,3.690236,3.549623,3.4707425,3.3815732,3.2855449,3.2615378,3.3198407,3.433017,3.8925817,4.173808,4.1772375,4.232111,5.103226,5.4599032,5.3844523,5.3330083,5.439326,5.5387836,5.5833683,5.6519604,5.552502,5.3227196,5.219832,5.6210938,5.9126086,6.245279,6.557371,6.5985265,6.8797526,7.5519514,8.2310095,8.745448,9.132992,9.523964,9.750318,10.055551,10.456812,10.755186,10.535692,10.106995,9.668007,9.349055,9.22902,9.287323,9.338767,9.349055,9.156999,8.47451,7.4456344,7.1952744,7.174697,7.1095347,7.0135064,6.866034,7.06495,7.1952744,7.2467184,7.6205435,7.630832,7.716572,7.8263187,8.038953,8.546532,8.388771,8.340756,8.80718,9.592556,9.880642,10.021255,9.006097,8.450503,8.903209,9.846346,10.172156,10.371073,10.069269,9.541112,9.695444,9.1810055,8.882631,8.735159,8.738589,8.940934,9.434795,9.054111,8.694004,8.529384,8.021805,8.718011,9.095266,9.637141,10.113853,9.585697,9.088407,7.846896,5.579939,3.8034124,5.830299,3.1106358,2.6579304,2.901431,2.7573884,1.611906,1.2449403,4.180667,6.4887795,7.2878733,8.776315,5.885172,9.89093,13.567448,12.524854,5.223262,14.757515,11.379372,8.484799,9.571979,8.241299,7.5279446,8.40249,10.179015,10.463672,5.192395,3.525616,3.7862647,3.8137012,3.8342788,6.451054,4.5099077,4.482471,4.7842746,4.8082814,4.90431,6.0669403,6.018926,6.118384,6.368744,5.4324665,6.036074,5.3707337,4.616225,4.4756117,5.1512403,5.377593,5.768566,6.392751,7.222711,8.131552,6.711703,5.8337283,5.360445,5.130663,4.9420357,6.018926,6.101236,6.475061,7.3084507,7.675417,8.141841,8.107545,7.7783046,7.5931067,8.207003,9.249598,10.096705,10.343636,10.254466,10.738038,9.770895,9.280463,9.280463,9.613133,9.97324,11.519984,11.746337,12.103014,12.651748,12.065289,12.055,11.279913,10.714031,10.377932,9.338767,7.9017696,6.7185616,5.4770513,4.314421,3.8274195,3.083199,4.870014,7.3084507,7.658269,2.318401,1.0460242,0.66876954,0.77851635,1.0082988,1.0323058,1.1008976,0.939707,0.922559,1.0940384,1.1763484,1.6599203,2.0028791,2.568761,3.309552,3.7759757,3.9851806,4.190956,4.232111,4.2526884,4.7019644,4.8082814,5.06893,5.65539,6.245279,6.036074,6.094377,6.0154963,6.3173003,6.8797526,6.924337,7.208993,7.720001,8.117833,8.412778,8.958082,9.23245,9.493098,9.22216,8.875772,9.856634,8.477941,8.519095,9.211872,10.110424,11.080997,11.88352,12.466551,12.291641,11.965831,13.245067,13.224489,12.542002,12.267634,12.439114,12.065289,10.902658,10.0041065,8.961512,7.9600725,7.8126,8.40249,8.964942,10.151579,11.928105,13.601744,15.083325,15.54632,15.717799,15.515453,14.04759,14.174485,13.718349,12.027563,10.048691,10.347065,11.125582,11.348505,11.362224,10.97468,9.458802,10.988399,11.821788,11.495977,10.624862,10.902658,10.213311,9.379922,8.803751,8.988949,10.539123,10.799771,9.410788,8.30646,8.213862,8.673427,8.515666,6.893471,5.3158607,4.4104495,3.9165888,3.8925817,3.7348208,3.433017,3.1106358,3.0523329,3.340418,3.6970954,3.9371665,4.0091877,3.9680326,4.6127954,5.3398676,5.8474464,6.258997,7.1198235,8.090397,8.56025,8.419638,7.8263187,7.2295704,7.5690994,8.172707,8.543102,8.64256,8.879202,8.659708,8.23444,7.8023114,7.5690994,7.7680154,8.1041155,8.923786,9.55826,9.496528,8.378482,7.64798,6.848886,6.1286726,5.686256,5.751418,5.6005163,5.178677,5.0140567,5.192395,5.363875,0.12689474,0.16804978,0.18519773,0.17490897,0.16119061,0.22635277,0.33952916,0.4424168,0.51100856,0.58302987,0.7476501,0.7990939,0.5624523,0.39097297,0.41498008,0.5144381,0.5178677,0.607037,0.7305021,0.8196714,0.7922347,0.823101,0.8162418,0.83338976,0.96371406,1.3101025,1.8828435,2.2052248,2.5653315,3.0214665,3.3815732,3.532475,3.799983,4.0709205,4.3178506,4.588788,4.880303,5.079219,5.2472687,5.219832,4.605936,4.496189,4.125794,3.9543142,3.9440255,3.5530527,3.673088,4.016047,4.4516044,4.8288593,4.9694724,5.394741,5.9640527,6.23499,5.994919,5.2506986,4.945465,5.24041,5.439326,5.2301207,4.722542,4.465323,4.091498,3.6525106,3.1655092,2.6373527,2.4624438,2.651071,2.6407824,2.3321195,2.0920484,2.0886188,2.0165975,1.8005334,1.5021594,1.3306799,1.0425946,0.7339317,0.5453044,0.4629943,0.30866286,0.2709374,0.22978236,0.22635277,0.2503599,0.23664154,0.29837412,0.33952916,0.34981793,0.32581082,0.25721905,0.22635277,0.26750782,0.29151493,0.26407823,0.20920484,0.25721905,0.24350071,0.28465575,0.3566771,0.31895164,0.38754338,0.7510797,1.2449403,1.6221949,1.5536032,1.2449403,0.86082643,0.490431,0.21263443,0.09945804,0.09259886,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.18176813,0.12346515,0.26064864,0.5041494,0.7510797,0.8711152,0.97057325,1.1180456,1.2312219,1.4507155,2.1194851,3.3026927,4.139512,4.9351764,5.6210938,5.73427,6.2075534,6.7459984,7.140401,7.2158523,6.8557453,7.720001,8.512236,9.3936405,10.2921915,10.899229,11.4376745,11.787492,12.120162,12.377381,12.274493,12.075578,12.154458,12.205902,11.746337,10.093276,11.262765,12.055,12.572867,12.734058,12.257345,12.22648,11.465111,11.399949,12.291641,13.241637,14.754086,15.584045,15.841265,15.604623,14.942713,14.829536,15.244516,16.314548,17.37429,16.976458,15.498305,14.400838,13.896688,13.927555,14.177915,14.771234,14.562028,14.009865,13.522863,13.4474125,12.874671,12.63117,12.267634,11.7257595,11.345076,11.938394,12.665466,13.203912,13.37882,13.155897,13.05301,13.443983,13.502286,12.939834,12.027563,12.178465,12.830087,13.471419,13.992717,14.661487,14.445422,14.726648,15.076467,15.481158,16.355703,16.715809,16.86671,17.158226,17.439453,17.058767,17.278261,17.885298,17.988186,17.556059,17.436022,17.302269,17.607502,17.820137,17.88873,18.241976,18.022482,18.670673,19.809298,21.109112,22.295748,24.538698,26.630747,28.023159,28.112328,26.246634,24.260902,20.663265,15.069608,9.3764925,7.7885933,5.909179,3.525616,1.670209,0.85739684,1.0837497,1.1111864,2.5070283,3.882293,4.7019644,5.271276,5.967482,9.095266,10.131001,8.738589,8.793462,11.756626,11.784062,9.863494,7.4765005,6.615674,7.596536,7.795452,7.3255987,6.931196,8.008087,7.699424,7.5553813,7.805741,8.347616,8.755736,10.295622,10.734609,10.604284,10.765475,12.415107,12.493987,11.187314,10.868362,11.478829,10.528833,10.22703,10.539123,10.837497,11.156448,12.181894,12.905538,14.987297,13.430264,8.4264965,5.3570156,7.3290286,7.380472,7.0375133,6.1458206,2.867135,1.6221949,1.5501735,2.369845,3.3541365,3.3301294,6.931196,6.1629686,4.715683,4.7019644,6.691125,4.7019644,6.2658563,9.990388,12.123591,6.557371,6.4716315,7.613684,8.64599,8.848335,8.114404,5.778855,6.5230756,6.001778,4.0674906,4.773986,3.9543142,3.8205605,3.549623,3.2546785,3.974892,4.712253,4.9694724,5.377593,5.874883,5.720552,6.210983,6.6705475,7.085528,7.394191,7.486789,6.307011,6.090947,5.768566,5.2609873,5.501058,5.3913116,4.911169,4.6848164,4.73969,4.5167665,4.3624353,4.2526884,3.974892,3.5564823,3.2375305,3.2032347,3.1106358,3.1312134,3.2821152,3.40901,3.8445675,4.2526884,4.355576,4.3658648,4.996909,5.6485305,5.9160385,5.953764,5.888602,5.8165803,5.610805,5.518206,5.4153185,5.3158607,5.377593,5.8474464,6.101236,6.451054,6.8728933,7.0135064,6.6636887,7.0786686,7.7783046,8.3922,8.669997,9.235879,9.760606,10.052121,10.052121,9.81205,9.695444,9.259886,8.889491,8.80718,9.067829,9.184435,9.301042,9.47595,9.496528,8.899779,8.303031,7.9257765,7.4765005,6.8900414,6.3310184,6.4716315,6.756287,7.023795,7.181556,7.1987042,7.0032177,7.140401,7.3084507,7.4799304,7.891481,7.466212,7.174697,7.5862474,8.553391,9.211872,9.908078,9.493098,9.301042,9.798331,10.566559,10.542552,10.491108,10.179015,9.870353,10.319629,10.158438,10.168727,9.935514,9.493098,9.318189,9.832627,9.997248,9.9801,9.80519,9.349055,10.549411,10.539123,10.484249,10.635151,10.347065,10.014396,9.455373,7.226141,4.3658648,4.40359,3.0523329,3.0043187,3.5187566,3.6353626,2.177788,1.2415106,2.7711067,6.543653,10.439664,10.443094,8.879202,14.030442,17.38115,14.565458,5.360445,14.256795,10.4705305,9.256456,12.373952,8.080108,8.656279,6.39961,5.4839106,5.9297566,3.5873485,2.7951138,4.5956473,5.130663,4.6127954,7.3393173,5.5490727,5.535354,5.6176643,5.2609873,5.0895076,6.6739774,6.5024977,6.4819202,6.9037595,6.447624,6.7357097,6.101236,5.456474,5.2609873,5.4976287,5.6005163,5.977771,6.495639,7.3290286,8.961512,7.0546613,5.809721,5.0346346,4.7259717,5.086078,5.826869,5.9812007,6.4133286,7.1266828,7.284444,8.131552,8.23444,7.949784,7.870903,8.80718,9.1810055,10.05898,10.429376,10.504827,11.732618,10.456812,9.719451,9.547972,9.712592,9.746887,12.199042,12.555719,12.30193,12.092726,11.763485,12.363663,11.417097,10.209882,9.084977,7.438775,6.478491,5.562791,4.256118,2.9906003,3.0557625,1.3546871,2.9322972,4.8905916,5.1066556,2.218943,0.805953,0.274367,0.13032432,0.10288762,0.13032432,0.4698535,0.432128,0.5796003,0.9431366,1.0151579,1.903421,2.411,2.8534167,3.2443898,3.3129816,3.2889743,3.6216443,3.673088,3.4433057,3.5564823,4.386442,4.7842746,5.3570156,5.953764,5.638242,5.885172,5.8543057,6.0326443,6.3138704,5.9914894,6.228131,6.800872,7.514226,8.114404,8.309891,8.309891,8.718011,8.735159,8.639131,9.788043,9.009526,9.170717,9.421077,9.554831,10.031544,10.017825,10.80663,11.688034,12.415107,13.193623,13.680624,13.21763,13.083877,13.584596,14.057879,13.111313,11.694893,10.038403,8.573969,7.9257765,8.48137,9.3764925,11.036412,13.248496,15.162207,16.674654,16.828985,16.365992,15.6697855,14.788382,14.733508,13.690913,11.958971,10.405369,10.467101,10.799771,11.423956,11.537132,10.439664,7.5450926,9.901219,11.413667,11.71547,11.266195,11.372512,10.573419,9.400499,8.570539,8.879202,11.218181,11.331357,9.3079,7.4524937,7.016936,8.200144,8.872343,8.100685,6.3035817,4.5442033,4.537344,4.705394,4.763697,4.5167665,4.081209,3.8788633,3.6559403,4.0023284,4.372724,4.5784993,4.7808447,5.3432975,5.813151,5.9880595,6.029215,6.4819202,7.490219,8.025234,7.881192,7.3118806,7.051232,7.675417,8.018375,8.450503,8.848335,8.56368,8.625413,8.580828,8.467651,8.354475,8.351046,8.64599,9.561689,10.463672,10.72775,9.743458,8.337327,7.442205,6.81802,6.3310184,5.9400454,5.5422134,4.8837323,4.7671266,5.336438,6.042933,0.21263443,0.16462019,0.16119061,0.19891608,0.2503599,0.274367,0.50757897,0.7476501,0.8196714,0.7099246,0.5658819,0.42869842,0.34981793,0.38754338,0.5144381,0.6241849,0.5418748,0.6001778,0.70649505,0.7579388,0.67219913,0.72021335,0.8779744,1.0494537,1.2106444,1.4198492,1.8965619,2.2429502,2.6407824,3.0626216,3.2958336,3.6147852,4.0674906,4.5201964,4.9180284,5.3090014,5.055212,4.8905916,4.681387,4.4584637,4.4104495,4.4104495,4.3349986,4.1120753,3.8342788,3.782835,3.6970954,4.033195,4.437886,4.7979927,5.2506986,5.4324665,6.135532,6.5162163,6.2144127,5.3707337,4.6265135,4.804852,4.911169,4.57507,4.07435,3.7211025,3.8137012,3.8102717,3.5873485,3.4776018,3.2821152,3.117495,2.9460156,2.726522,2.411,2.0920484,1.7765263,1.4472859,1.1592005,1.039165,1.0631721,0.7305021,0.44927597,0.34638834,0.26064864,0.22292319,0.20577525,0.18519773,0.16462019,0.15090185,0.16462019,0.17833854,0.28122616,0.40126175,0.30523327,0.20920484,0.17490897,0.14404267,0.09945804,0.07545093,0.16119061,0.17490897,0.19891608,0.25721905,0.30523327,0.70649505,1.3203912,2.0063086,2.5413244,2.6407824,1.7730967,1.0528834,0.5212973,0.19891608,0.07545093,0.07545093,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16462019,0.33609957,0.490431,0.7476501,0.7099246,0.94999576,1.1077567,1.1454822,1.3272504,2.0097382,3.3438478,4.7431192,5.7102633,5.844017,6.258997,6.8214493,7.0478024,6.883182,6.697984,6.478491,7.174697,8.237869,9.239308,9.873782,10.127572,10.943813,11.650309,11.921246,11.749766,12.127021,11.499407,10.765475,10.203023,9.445084,9.39707,10.374502,11.869802,13.025573,12.634601,11.657167,11.633161,12.596875,13.88983,14.143619,15.645778,16.386568,16.808409,16.736387,15.3817,15.110763,15.539461,16.12592,16.427725,16.098484,15.158776,13.951562,13.419975,13.9481325,15.350834,15.436573,14.760944,13.9309845,13.337666,13.169616,12.740917,12.168177,11.8869505,11.945253,11.993267,12.617453,12.689473,12.644889,12.63117,12.4974165,12.71691,12.5145645,12.672326,13.138749,13.015285,13.917266,14.832966,15.361122,15.367981,14.953001,13.588025,13.234778,13.704632,14.534592,15.001016,15.927004,16.571766,16.931873,16.911295,16.328266,17.034761,17.075916,16.969599,17.144508,17.912735,17.573206,17.54234,17.412016,17.473747,18.708399,18.670673,18.341434,18.272842,18.903887,20.539799,22.089973,24.710178,26.298077,26.10259,24.734184,22.758743,19.360022,15.21022,11.399949,9.458802,8.165848,5.4153185,3.0969174,1.8656956,1.1454822,1.1934965,1.4438564,2.510458,4.8425775,8.711152,9.469091,8.824328,7.641121,7.514226,10.772334,13.224489,12.915827,11.461681,10.412228,11.228469,12.72034,11.982979,10.281903,8.923786,9.277034,7.4456344,8.114404,9.091836,9.585697,10.206452,11.026124,11.495977,12.061859,12.535142,12.085866,11.022695,11.077567,12.315649,13.557159,12.360233,11.7257595,11.897239,11.46854,10.851214,12.267634,13.732068,14.812388,14.421415,12.096155,7.9943686,6.1286726,8.179566,10.590566,10.082987,3.6627994,1.9274281,1.7319417,2.702515,4.245829,5.5387836,8.748878,6.3481665,6.200694,8.155559,4.029765,8.495089,12.037852,13.498857,12.943263,11.670886,7.9737906,7.250148,7.630832,8.200144,9.016385,7.846896,6.9654922,5.6965446,4.4687524,4.822,4.249259,3.9474552,3.5221863,3.1312134,3.508468,3.8891523,3.642222,3.9200184,4.7088237,4.866585,5.9434752,6.914048,7.8674736,8.4264965,7.7680154,6.461343,6.245279,6.108095,5.90575,6.3310184,5.7719955,5.055212,4.681387,4.530485,3.8445675,3.8102717,3.542764,3.292404,3.175798,3.1895163,3.6044965,3.789694,3.7279615,3.542764,3.4947495,3.8617156,4.4275975,4.8425775,5.0449233,5.2644167,5.3981705,5.778855,5.994919,6.0497923,6.3790326,5.926327,5.5387836,5.271276,5.1340923,5.096367,5.535354,6.2212715,6.7459984,6.9654922,6.989499,7.5382333,7.8846216,8.1041155,8.31675,8.683716,9.071259,9.462232,9.764035,9.788043,9.263316,8.824328,8.14527,7.6205435,7.442205,7.613684,8.200144,8.676856,9.225591,9.777754,10.010965,9.716022,9.239308,8.556821,7.6616983,6.5779486,6.540223,6.7494283,6.8728933,6.9654922,7.4936485,6.8557453,7.1095347,7.390761,7.281014,6.8043017,7.2192817,7.0958166,7.3701835,8.162418,8.772884,9.321619,10.093276,10.261326,10.007536,10.484249,10.103564,10.264755,10.179015,9.846346,10.041832,10.199594,10.604284,10.861504,10.940384,11.183885,10.587136,10.172156,10.501397,11.266195,11.290202,11.427385,11.122152,10.816919,10.662587,10.528833,9.160428,9.599416,8.285883,5.4153185,4.928317,5.161529,5.2747054,4.7602673,4.046913,4.4859004,1.99602,4.9523244,4.5990767,2.4727325,10.405369,9.674867,16.283682,17.192522,10.535692,5.6142344,17.003895,8.471081,5.086078,10.340206,6.166398,7.6788464,6.042933,4.3521466,3.7211025,3.2821152,2.9391565,5.967482,6.7048435,5.3741636,8.073249,5.703404,6.090947,6.574519,6.2144127,5.7994323,7.8126,7.8503256,8.014946,8.570539,7.949784,6.6568294,6.012067,5.6348124,5.4736214,5.830299,5.693115,6.3653145,6.4407654,6.8283086,10.7586155,7.5588107,5.641671,3.8377085,3.1723683,6.883182,6.3310184,6.3035817,6.4579134,6.5162163,6.2727156,7.3839016,7.6959944,8.158989,9.0644,10.041832,10.39508,11.039842,11.029553,10.72089,11.794352,10.487679,10.600855,10.371073,9.6988735,10.161868,12.312219,11.574858,10.494537,10.275044,10.789482,11.691463,10.131001,8.611694,7.891481,6.989499,5.8405876,4.9214582,4.0846386,3.0797696,1.5398848,0.84367853,1.8245405,3.2786856,3.9508848,2.5481834,0.94999576,0.28465575,0.082310095,0.044584636,0.044584636,0.034295876,0.030866288,0.35324752,0.9294182,1.2963841,1.786815,2.784825,3.4707425,3.5461934,3.2649672,2.9494452,2.976882,3.0454736,3.117495,3.433017,3.8377085,4.2835546,4.7362604,5.055212,5.003768,5.212973,5.4187484,5.48734,5.4770513,5.662249,5.5250654,5.720552,6.4716315,7.5519514,8.285883,7.798882,7.6925645,7.8263187,8.309891,9.506817,9.9698105,9.774324,9.156999,8.858624,10.117283,9.945804,10.131001,11.05356,12.507706,13.718349,13.423406,13.104454,12.425395,11.55428,11.1393,13.008426,13.255356,12.271064,10.707172,9.47595,9.523964,10.4533825,12.2093315,14.171056,15.138199,16.016174,16.21852,15.844694,15.5085945,16.328266,17.267973,15.258235,12.535142,10.748327,10.9541025,10.81006,11.945253,12.9707,12.535142,9.338767,10.14472,10.930096,11.547421,11.907528,11.993267,11.321068,9.880642,9.14328,9.911508,12.329367,11.828648,9.314759,7.2158523,6.636252,7.3701835,7.6033955,7.7714453,6.420188,4.4756117,5.2335505,5.720552,5.936616,5.8062916,5.4153185,4.99005,4.3658648,4.6402316,5.2026844,5.662249,5.844017,5.8680243,5.874883,5.861165,5.7994323,5.6142344,6.166398,6.914048,7.0923867,6.866034,7.3530354,7.610255,7.966932,8.186425,8.1487,7.8434668,8.440215,8.700864,8.81747,8.800322,8.484799,8.934075,9.599416,10.690024,11.732618,11.550851,9.403929,8.186425,7.56567,7.1129646,6.3310184,5.857735,5.453044,5.545643,6.200694,7.140401,0.26407823,0.22292319,0.2503599,0.28465575,0.30866286,0.37382504,0.59331864,0.65162164,0.6344737,0.5727411,0.4046913,0.4389872,0.48700142,0.5693115,0.7099246,0.9568549,0.59674823,0.53158605,0.5693115,0.61389613,0.6344737,0.8196714,1.0494537,1.2792361,1.5433143,1.9548649,2.1503513,2.3252604,2.6064866,3.0557625,3.649081,3.957744,4.386442,5.1512403,5.9160385,5.7994323,4.887162,4.65395,4.4859004,4.2252517,4.166949,3.8925817,3.6696587,3.5359046,3.5050385,3.5530527,3.799983,4.2252517,4.715683,5.120374,5.2609873,5.3844523,5.658819,5.8474464,5.7411294,5.164959,4.3590055,3.9543142,3.6319332,3.3712845,3.426158,3.083199,2.702515,2.6750782,3.000889,3.3198407,3.5530527,3.1586502,2.7230926,2.4041407,1.9102802,1.4850113,1.2655178,1.0734608,0.84367853,0.6241849,0.5693115,0.4355576,0.33266997,0.2777966,0.20920484,0.1920569,0.15776102,0.13032432,0.12003556,0.12689474,0.14061308,0.17490897,0.2194936,0.22635277,0.1097468,0.1097468,0.08573969,0.0548734,0.034295876,0.041155048,0.116605975,0.2194936,0.26064864,0.31209245,0.6344737,1.4472859,2.6750782,3.8788633,4.3521466,3.1517909,2.1297739,1.0631721,0.3806842,0.1371835,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09945804,0.22635277,0.37039545,0.58988905,0.7373613,0.8025235,0.8162418,0.864256,1.0940384,1.4164196,2.1332035,3.340418,4.383013,3.8548563,4.180667,4.57507,4.897451,5.171818,5.576509,6.029215,6.680836,7.4799304,8.309891,8.992378,9.297611,9.671436,10.120712,10.477389,10.39508,10.185875,10.120712,10.240748,10.422516,10.398509,10.278474,10.611144,11.369082,12.257345,12.696333,12.130451,11.842365,12.566009,13.996146,14.778092,15.861842,16.204802,16.21166,15.951012,15.162207,15.333686,15.772673,16.0539,16.009314,15.755525,15.313108,14.160767,13.481709,13.663476,14.277372,14.723219,14.2190695,13.71492,13.564018,13.509145,12.603734,11.770344,11.290202,11.180455,11.201033,11.4205265,11.447963,11.4376745,11.543991,11.8869505,12.175035,11.976119,12.397959,13.564018,14.613472,14.699212,15.237658,15.656067,15.697222,15.415996,14.315098,13.759505,13.63261,13.848674,14.352823,15.083325,15.834405,16.400288,16.732958,16.94902,16.691803,16.328266,16.115631,16.146498,16.338554,16.523752,17.144508,17.53548,17.518333,17.412016,17.521763,17.422304,17.477179,17.895588,18.732407,19.901896,22.141417,24.226606,25.159454,24.171732,21.150267,18.636377,16.105343,13.358243,10.511685,8.98209,7.4936485,5.909179,4.2218223,2.5241764,1.371835,1.7833855,2.7882545,4.2389703,6.807731,6.2487082,7.5588107,9.314759,10.8958,12.504276,14.325387,14.901558,14.987297,14.781522,13.927555,13.649758,12.576297,11.482259,10.63858,9.801761,9.22216,9.06097,8.913498,8.944365,9.89093,10.124143,10.988399,12.116733,12.956982,12.768354,13.454271,14.1299,14.195063,13.63261,12.9809885,13.313659,13.505715,13.601744,13.910407,15.014734,15.103903,15.289101,13.965281,11.204462,8.752307,6.327589,6.680836,7.599966,7.2295704,4.040054,2.2669573,1.3958421,1.7182233,2.7745364,3.3541365,8.261876,8.416207,8.584257,10.257896,11.670886,13.001566,13.893259,13.821238,13.392539,14.359683,9.047252,7.4113383,7.7097125,8.577398,8.992378,7.723431,7.1198235,6.3824625,5.56965,5.5902276,4.664239,4.256118,3.9165888,3.566771,3.4844608,3.6113555,3.8377085,4.0537724,4.3933015,5.2472687,6.6122446,7.226141,7.7097125,8.021805,7.449064,6.444195,5.9743414,5.645101,5.4839106,5.9434752,5.7994323,5.442755,5.1683884,4.945465,4.40702,4.262977,3.9714622,3.7108135,3.5599117,3.4947495,3.841138,3.957744,3.9611735,3.9474552,4.0057583,4.2355404,4.4687524,4.6608095,4.856296,5.2026844,5.192395,5.353586,5.5113473,5.627953,5.778855,5.8165803,5.754848,5.7891436,5.9228973,5.9640527,5.953764,6.125243,6.4304767,6.7459984,6.8797526,7.4284863,7.73029,8.025234,8.450503,9.06097,9.139851,9.472521,9.743458,9.72631,9.297611,8.546532,7.8503256,7.6376915,7.8366075,7.870903,7.9600725,8.244728,8.573969,8.930646,9.434795,9.105555,8.618553,8.155559,7.7680154,7.394191,7.160979,6.759717,6.169828,5.7308407,6.135532,6.0395036,6.375603,6.81802,7.034084,6.684266,6.7357097,6.8454566,6.8728933,6.941485,7.394191,8.354475,9.050681,9.225591,9.297611,10.360784,10.676306,11.129011,11.077567,10.518545,10.089847,9.709162,10.39165,10.823778,10.703742,10.734609,10.88551,10.336777,10.30591,10.926665,11.255906,11.64345,11.585147,11.163307,10.628291,10.405369,8.920357,8.89635,8.56025,7.1712675,5.0003386,4.187526,7.394191,7.459353,4.07435,3.8034124,3.1483612,22.793037,23.02625,4.8425775,9.956093,6.245279,10.124143,13.361672,11.931535,6.0052075,11.125582,5.6176643,3.474172,6.7357097,5.4804807,7.2878733,7.205563,6.475061,5.9571934,6.125243,4.7671266,6.3618846,6.8763227,6.2212715,8.255017,6.5710897,6.725421,7.082098,6.831738,6.018926,7.8777623,8.532814,9.074688,9.547972,8.961512,8.001227,7.133542,6.1046658,5.353586,6.012067,5.4770513,5.8508763,5.446185,4.870014,7.023795,6.7631464,5.8817425,4.880303,4.636802,6.392751,6.927767,6.9380555,6.807731,6.8043017,7.0786686,8.296172,8.8929205,9.496528,10.13786,10.233889,10.14129,10.683165,10.9541025,11.146159,12.55229,11.852654,11.917816,11.640019,11.177026,11.931535,12.332796,10.960961,10.038403,9.952662,9.273604,9.602845,9.187865,9.626852,9.801761,5.90232,4.9008803,4.0263357,3.083199,3.5942078,8.803751,4.2115335,4.9214582,6.5985265,6.2692857,2.3149714,0.90198153,0.90541106,0.69963586,0.030866288,0.020577524,0.020577524,0.017147938,0.28808534,0.94656616,1.9685832,2.1640697,3.1346428,3.74168,3.8102717,4.1429415,3.690236,3.82399,3.923448,3.789694,3.6765177,3.7176728,3.9165888,4.4516044,4.9694724,4.588788,4.7979927,5.1512403,5.295283,5.2164025,5.2335505,5.1100855,5.593657,6.245279,7.016936,8.2481575,8.56025,8.14527,7.956643,8.549961,10.069269,10.532263,9.421077,8.539673,8.597976,9.201583,9.959522,10.185875,10.837497,12.236768,14.071597,13.9138365,13.101024,11.838936,10.566559,9.956093,10.8958,11.231899,11.187314,10.88551,10.367643,9.56512,10.251037,11.4376745,12.521424,13.282792,13.594885,14.109323,14.507155,14.939283,16.023033,16.005884,14.651197,12.953552,11.674315,11.334786,10.738038,10.998687,11.760056,12.175035,10.899229,10.995257,11.485688,11.797781,11.828648,11.931535,11.369082,10.628291,10.134431,10.347065,11.766914,10.192734,7.8331776,6.835168,7.486789,8.2481575,8.169277,7.3564653,6.375603,5.9880595,7.174697,7.6445503,7.7783046,7.56224,6.948344,5.8680243,5.206114,5.288424,5.6210938,5.967482,6.358455,6.0497923,6.0532217,6.166398,6.1801167,5.871454,5.90232,6.262427,6.550512,6.831738,7.623973,7.888051,8.1041155,8.008087,7.6171136,7.1952744,7.6959944,8.042382,8.2653055,8.39563,8.460793,8.899779,10.021255,10.542552,10.216741,9.829198,8.803751,8.110974,7.699424,7.4765005,7.3221693,7.1198235,7.1129646,7.010077,7.0958166,8.241299,0.31895164,0.2469303,0.33609957,0.44927597,0.53844523,0.6241849,0.72021335,0.6824879,0.6001778,0.5212973,0.42869842,0.58988905,0.7442205,0.7339317,0.6241849,0.70649505,0.66876954,0.6859175,0.7373613,0.7990939,0.8162418,1.0597426,1.3615463,1.646202,1.903421,2.1915064,2.2120838,2.294394,2.4761622,2.8980014,3.8034124,4.400161,5.161529,6.23156,6.999788,6.111525,4.636802,4.3452873,4.273266,3.9954693,3.6182148,3.4227283,3.2992632,3.2546785,3.2649672,3.2546785,3.426158,3.6799474,3.9508848,4.1943855,4.3933015,4.5613513,4.763697,4.9214582,4.931747,4.65395,3.8514268,3.2786856,2.9871707,2.901431,2.8156912,2.3732746,2.2395205,2.5447538,3.0351849,3.0900583,3.0729103,2.5996273,2.270387,2.1674993,1.8588364,1.3786942,1.0666018,0.83681935,0.64819205,0.490431,0.37382504,0.29837412,0.25378948,0.2194936,0.15090185,0.15433143,0.12346515,0.09602845,0.08916927,0.09602845,0.11317638,0.116605975,0.12003556,0.1097468,0.05144381,0.0548734,0.037725464,0.030866288,0.030866288,0.020577524,0.072021335,0.16119061,0.26750782,0.4972902,1.0940384,1.9137098,3.1277838,4.0606318,4.122364,2.8328393,1.5947582,0.72707254,0.26407823,0.11317638,0.06516216,0.020577524,0.020577524,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.12346515,0.25721905,0.3841138,0.6173257,0.6859175,0.6893471,0.7339317,0.9294182,0.99801,1.3992717,2.4555845,3.6044965,3.3850029,3.083199,3.4776018,3.9028704,4.170378,4.5819287,5.439326,6.121814,6.691125,7.3427467,8.399059,8.752307,8.865483,8.8929205,9.016385,9.424506,9.194724,9.702303,10.31277,10.799771,11.331357,11.753197,11.808069,11.955542,12.349944,12.830087,12.349944,12.257345,13.025573,14.407697,15.443433,15.6697855,15.683503,15.724659,15.662926,14.977009,14.791811,14.575747,14.712931,15.055889,14.911846,14.445422,13.817808,13.368532,13.265644,13.505715,13.9309845,13.4474125,12.80608,12.428825,12.397959,11.605724,10.981539,10.80663,11.032983,11.293632,11.101575,10.748327,10.63858,10.840926,11.094715,11.619442,11.96926,12.72034,13.954991,15.261664,15.556609,15.789821,15.940722,15.87899,15.350834,14.589465,13.982429,13.941273,14.387119,14.740367,15.2033615,15.659496,16.084764,16.407146,16.492886,16.2974,16.180794,15.88242,15.522313,15.608052,16.393429,17.559488,18.235117,18.159666,17.686382,17.069057,16.664366,16.564907,16.828985,17.466888,18.488907,19.922474,21.599543,22.885637,22.69701,19.740705,17.223389,15.29596,13.708061,11.797781,9.846346,8.584257,7.31531,5.7994323,4.2698364,2.9631636,2.7059445,2.8945718,3.5050385,5.06893,6.3310184,7.4181976,8.882631,10.511685,11.327928,13.207341,14.627191,15.121051,14.740367,14.071597,13.642899,13.766364,13.588025,12.867812,11.976119,12.154458,11.945253,11.677745,11.55771,11.650309,11.451392,12.024134,12.754636,13.279363,13.516005,14.565458,14.977009,14.839825,14.579176,14.959861,15.29939,15.752095,15.553179,15.0250225,15.580616,17.237106,16.486027,13.200482,8.97523,7.1198235,6.7528577,6.7185616,7.64798,7.888051,3.4844608,2.085189,1.2483698,1.5913286,2.6819375,3.0626216,6.4373355,7.085528,8.628842,10.984968,10.367643,9.599416,10.233889,10.182446,9.740028,11.595435,9.266746,8.39563,8.690575,9.22216,8.419638,7.857185,7.380472,6.6122446,5.761707,5.627953,4.9934793,4.3521466,3.882293,3.625074,3.4878905,3.7965534,4.122364,4.4275975,4.773986,5.3227196,6.48535,6.9517736,7.1987042,7.366754,7.250148,6.368744,5.645101,5.1409516,4.976331,5.360445,5.813151,6.0052075,5.9228973,5.658819,5.3981705,4.9934793,4.4104495,4.180667,4.2938433,4.1943855,4.4275975,4.417309,4.2355404,4.1017866,4.355576,4.506478,4.671098,4.6779575,4.647091,4.996909,4.756838,4.7602673,4.911169,5.0929375,5.1821065,5.5147767,5.6313825,5.6793966,5.802862,6.135532,6.0703697,6.166398,6.3653145,6.601956,6.8043017,7.034084,7.3427467,7.7131424,8.141841,8.659708,8.9100685,9.095266,9.167287,9.102125,8.89635,8.364764,7.795452,7.73029,8.1487,8.457363,8.237869,8.1384115,8.090397,8.080108,8.158989,7.8537555,7.5107965,7.3187394,7.274155,7.1952744,6.7974424,6.245279,5.761707,5.545643,5.761707,6.0703697,6.3138704,6.64997,6.807731,6.094377,6.327589,6.5127864,6.7494283,7.1026754,7.589677,8.745448,9.294182,9.56512,9.935514,10.816919,11.348505,11.790922,11.965831,11.859513,11.612583,10.645439,10.9541025,11.543991,11.72233,11.094715,11.290202,11.022695,10.9369545,11.14273,11.207891,11.96926,12.1921835,11.650309,10.600855,9.770895,9.355915,8.9100685,8.56368,7.9737906,6.293293,4.15666,5.470192,6.7219915,5.953764,2.7711067,2.6990852,12.977559,13.080446,4.331569,9.887501,6.324159,7.507367,10.010965,10.6317215,6.358455,10.299051,5.8371577,3.858286,5.9640527,4.496189,6.3035817,6.392751,6.3721733,6.7974424,7.174697,5.892031,6.8283086,7.517656,7.5279446,8.429926,6.9071894,7.332458,7.9086285,7.857185,7.407909,9.403929,9.626852,9.860064,10.278474,9.462232,8.738589,7.682276,6.5162163,5.7102633,5.9743414,5.5387836,5.6828265,5.305572,4.6436615,5.2815647,5.0620713,4.647091,4.0949273,3.8342788,4.650521,5.8817425,6.2418494,6.4887795,6.910619,7.3427467,8.244728,9.006097,9.757176,10.254466,9.89093,9.56512,9.788043,10.031544,10.611144,12.686044,12.706621,12.984418,12.826657,12.439114,12.88839,12.360233,10.998687,9.791472,9.14328,8.879202,7.997798,7.5279446,8.117833,8.330468,4.633373,3.4124396,2.9665933,3.457024,4.8288593,6.8043017,4.6265135,7.226141,7.9292064,5.1992545,2.6236343,1.0528834,3.6319332,3.4433057,0.17490897,0.13375391,1.0288762,1.08032,1.6187652,2.7642474,3.426158,2.9631636,3.3678548,3.8548563,4.180667,4.6402316,4.122364,4.3624353,4.5442033,4.3349986,3.9028704,3.6627994,3.625074,3.9337368,4.341858,4.1943855,4.314421,4.7842746,5.2026844,5.3741636,5.31929,5.336438,6.1286726,6.917478,7.5725293,8.632272,9.462232,9.132992,8.944365,9.445084,10.436234,10.88551,9.640571,9.088407,9.668007,9.897789,10.401938,10.655728,11.255906,12.291641,13.344524,13.677195,13.05301,11.653738,10.055551,9.218731,9.5033865,9.914937,10.412228,10.840926,10.9369545,10.196163,10.343636,11.235329,12.445972,13.282792,13.762935,14.486577,14.843254,14.894698,15.367981,14.928994,13.670336,12.476839,11.773774,11.547421,10.7586155,10.501397,10.875222,11.413667,11.091286,11.444533,11.561139,11.513125,11.46854,11.688034,11.581717,11.05356,10.494537,10.326488,11.012405,9.009526,7.7542973,7.7542973,8.529384,8.625413,8.244728,7.0752387,5.9743414,5.672538,6.7528577,7.4010496,7.891481,8.05953,7.8091707,7.1061053,6.4544835,6.262427,6.3173003,6.461343,6.584808,6.23156,5.936616,5.796003,5.809721,5.861165,5.7274113,6.042933,6.495639,7.0546613,7.963502,7.963502,8.056101,7.9086285,7.473071,6.9689217,7.3873315,7.630832,7.864044,8.1212635,8.279024,9.047252,9.47595,9.623423,9.575408,9.445084,8.855195,8.22758,7.8434668,7.7851634,7.9257765,8.114404,8.069819,7.8537555,7.997798,9.5033865,0.34981793,0.36010668,0.4972902,0.6173257,0.66876954,0.69963586,0.7442205,0.7682276,0.7133542,0.607037,0.5658819,0.64819205,0.7510797,0.72364295,0.6036074,0.6241849,0.7579388,0.805953,0.91227025,1.0940384,1.2277923,1.2346514,1.4850113,1.7730967,1.9754424,2.037175,2.1023371,2.2669573,2.5241764,2.9082901,3.4844608,4.5613513,5.826869,6.992929,7.377043,5.892031,4.187526,3.789694,3.7176728,3.4913201,3.1552205,3.117495,3.1037767,3.0900583,3.0317552,2.877424,2.9871707,3.1277838,3.1826572,3.2375305,3.5839188,3.765687,3.9474552,4.1600895,4.190956,3.6113555,3.1689389,2.8328393,2.6785078,2.6133456,2.3767042,2.0406046,2.2498093,2.6373527,2.8637056,2.5996273,2.4452958,2.0886188,1.9171394,1.9480057,1.821111,1.2517995,0.90198153,0.66876954,0.4972902,0.3806842,0.274367,0.21263443,0.18176813,0.15090185,0.10288762,0.106317215,0.09259886,0.07545093,0.06516216,0.06516216,0.07545093,0.058302987,0.048014224,0.048014224,0.041155048,0.0274367,0.020577524,0.020577524,0.024007112,0.01371835,0.072021335,0.15090185,0.29151493,0.6379033,1.4575747,2.5584722,3.6799474,4.2355404,4.1017866,3.625074,1.6324836,0.6344737,0.2194936,0.08916927,0.06516216,0.020577524,0.020577524,0.0274367,0.05144381,0.14061308,0.082310095,0.06516216,0.037725464,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.15090185,0.21263443,0.45613512,0.548734,0.5658819,0.58645946,0.70306545,0.6893471,0.90198153,1.6153357,2.5584722,2.9220085,2.4795918,3.0043187,3.4776018,3.5770597,3.683377,4.756838,5.4324665,5.885172,6.447624,7.630832,8.189855,8.453933,8.457363,8.488229,9.105555,8.961512,9.788043,10.64201,11.146159,11.509696,12.257345,12.548861,12.699762,12.922686,13.323947,13.022143,12.915827,13.351384,14.335675,15.532601,15.5085945,15.165636,15.093615,15.237658,14.88098,14.229359,13.536582,13.55373,14.071597,13.917266,13.992717,13.896688,13.7938,13.666906,13.289652,13.018714,12.593445,11.952112,11.372512,11.46854,11.183885,10.923236,11.101575,11.674315,12.123591,11.876661,11.180455,10.744898,10.81006,11.129011,11.917816,12.5145645,13.104454,13.920695,15.230798,15.854982,16.03675,16.023033,15.758954,14.898128,14.589465,14.088745,14.208781,14.922135,15.361122,15.7966795,15.841265,15.820687,15.789821,15.5085945,15.659496,15.649208,15.343974,15.004445,15.29596,16.554619,17.933313,18.732407,18.725548,18.166525,17.117071,16.479168,16.191082,16.283682,16.849564,17.700102,18.684393,19.713268,20.502073,20.553518,18.814716,16.70552,14.802099,13.3033695,12.0309925,10.501397,9.551401,8.567109,7.3530354,6.1321025,4.8940215,3.9063,3.4398763,3.549623,4.098357,5.717122,6.8728933,8.186425,9.695444,10.875222,12.212761,13.560589,14.270514,14.325387,14.335675,14.092175,14.661487,14.774663,14.260224,14.030442,14.400838,14.239647,14.188204,14.13676,13.22106,12.782072,13.080446,13.443983,13.817808,14.750656,15.46058,16.012743,16.37285,16.647217,17.04848,17.576635,18.883308,16.434584,12.260776,14.942713,18.169954,16.29054,11.80121,7.531374,6.6568294,6.2418494,5.754848,6.0875177,6.029215,2.277246,1.611906,1.4198492,2.1332035,3.2683969,3.4227283,4.619654,6.420188,7.7783046,7.874333,6.142391,5.2472687,5.809721,6.385892,6.7322803,7.8126,8.200144,8.196714,8.769455,9.5205345,8.711152,8.423067,7.6274023,6.632822,5.796003,5.528495,4.7808447,4.122364,3.7965534,3.7931237,3.8479972,4.1772375,4.4996185,4.7328305,4.8494368,4.8768735,5.970912,6.48535,6.608815,6.5985265,6.773435,6.2144127,5.518206,5.0655007,4.938606,4.938606,5.470192,5.8234396,5.7411294,5.363875,5.2472687,4.8597255,4.417309,4.307562,4.4721823,4.400161,4.698535,4.7808447,4.5784993,4.2938433,4.396731,4.523626,4.6745276,4.623084,4.5167665,4.866585,4.588788,4.431027,4.3933015,4.4516044,4.530485,4.945465,5.2438393,5.394741,5.5662203,6.135532,6.334448,6.56766,6.715132,6.8111606,7.06838,7.0752387,7.2467184,7.438775,7.64798,8.018375,8.4264965,8.553391,8.484799,8.327039,8.224151,8.042382,7.8434668,7.8983397,8.258447,8.766026,8.591117,8.292743,7.98408,7.6514096,7.1266828,6.7185616,6.4133286,6.341307,6.4407654,6.444195,6.0669403,5.744559,5.6073756,5.6519604,5.7377,6.121814,6.142391,6.334448,6.550512,5.9297566,6.2212715,6.293293,6.711703,7.5382333,8.309891,9.417647,9.921797,10.189304,10.443094,10.762046,11.125582,11.547421,11.952112,12.370522,12.905538,12.394529,12.349944,12.830087,13.306799,12.6586075,12.05157,11.646879,11.430815,11.4376745,11.732618,12.356804,12.600305,12.199042,11.194174,9.925226,9.709162,9.290752,8.793462,8.207003,7.366754,5.381023,3.899441,5.051782,6.680836,2.3252604,2.4315774,2.7573884,2.5790498,3.0969174,7.4456344,6.101236,7.6514096,10.573419,12.624311,10.851214,13.536582,7.517656,4.6848164,6.550512,4.232111,5.6965446,5.302142,5.4667625,6.893471,8.584257,6.64997,7.7131424,8.879202,9.259886,9.959522,8.107545,8.347616,8.927217,9.084977,9.033533,10.734609,10.484249,10.281903,10.39165,9.31133,8.81404,7.98065,7.14726,6.5642304,6.4098988,6.1286726,6.060081,5.7308407,5.2644167,5.3673043,4.557922,4.1189346,3.6559403,3.4192986,4.32128,5.4839106,5.9640527,6.711703,7.7028537,7.9292064,8.025234,7.9943686,8.488229,9.249598,9.108984,9.174147,9.39021,9.647429,10.340206,12.349944,12.655178,13.234778,13.279363,12.812939,12.703192,11.664027,10.497967,9.338767,8.556821,8.772884,6.077229,5.020916,4.90431,4.7088237,3.093488,2.1674993,5.4907694,6.334448,3.865145,3.1449318,3.3198407,7.675417,7.6651278,3.210094,2.7333813,1.5090185,3.5393343,3.2581081,0.8025235,1.99602,4.1326528,4.557922,4.8768735,5.2781353,4.506478,3.2958336,3.5702004,4.122364,4.4927597,4.955754,4.2835546,4.2526884,4.431027,4.4756117,4.1463714,3.9165888,3.8205605,3.8617156,3.9714622,4.0229063,4.125794,4.5922174,5.0586414,5.381023,5.638242,5.672538,6.560801,7.407909,7.9943686,8.748878,9.880642,9.829198,9.6645775,9.884071,10.401938,10.820349,10.072699,10.131001,11.0981455,11.207891,11.375941,11.55428,11.948683,12.504276,12.919256,13.474849,13.083877,11.838936,10.251037,9.256456,9.095266,9.510246,10.069269,10.539123,10.906088,10.271614,10.257896,10.97468,12.130451,13.035862,13.972139,14.640909,14.757515,14.520873,14.616901,13.725209,12.343085,11.519984,11.399949,11.211322,10.744898,10.419086,10.738038,11.444533,11.509696,11.739478,11.31078,11.05356,11.327928,12.006986,12.096155,11.338216,10.436234,9.901219,10.041832,8.800322,8.776315,9.23245,9.47938,8.855195,8.378482,7.4970784,6.4819202,5.909179,6.6431108,7.2364297,7.939495,8.412778,8.515666,8.299602,8.155559,7.740579,7.208993,6.677407,6.2247014,5.768566,5.3878818,5.188966,5.2918534,5.8371577,5.9297566,6.4407654,7.0546613,7.6959944,8.519095,8.080108,7.874333,7.6857057,7.486789,7.4456344,7.64798,7.56567,7.6857057,8.035523,8.162418,8.786603,8.669997,8.683716,9.383351,10.995257,9.873782,8.920357,8.515666,8.621983,8.779744,8.992378,8.752307,8.704293,9.270175,10.655728,0.36010668,0.5521636,0.7133542,0.764798,0.7339317,0.7373613,0.78194594,0.8676856,0.85396725,0.7510797,0.71678376,0.6241849,0.58302987,0.6173257,0.7099246,0.83338976,0.8848336,0.90198153,1.0357354,1.313532,1.6564908,1.3958421,1.4781522,1.6496316,1.7490896,1.704505,1.9342873,2.318401,2.7470996,3.069481,3.0729103,4.5819287,6.1149545,6.9654922,6.697984,5.130663,3.758828,3.2855449,3.093488,2.9391565,2.9494452,2.9700227,2.976882,2.8911421,2.719663,2.534465,2.7402403,2.877424,2.8396983,2.784825,3.1655092,3.3712845,3.4604537,3.6387923,3.6044965,2.510458,2.6373527,2.644212,2.5310357,2.3424082,2.153781,2.0680413,2.3389788,2.4967396,2.369845,2.0749004,2.0131679,1.8073926,1.6667795,1.6221949,1.5227368,0.97400284,0.71678376,0.5521636,0.38754338,0.24007112,0.1920569,0.15090185,0.116605975,0.08573969,0.06859175,0.061732575,0.06516216,0.058302987,0.041155048,0.041155048,0.041155048,0.037725464,0.034295876,0.030866288,0.0274367,0.01371835,0.01371835,0.006859175,0.0034295875,0.01371835,0.106317215,0.19548649,0.31895164,0.7305021,1.8897027,3.2855449,4.4275975,5.0929375,5.3741636,5.686256,2.668219,1.0082988,0.2709374,0.061732575,0.0034295875,0.0,0.010288762,0.10288762,0.32581082,0.70649505,0.30866286,0.17147937,0.09945804,0.020577524,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.061732575,0.11317638,0.29494452,0.36696586,0.38754338,0.4046913,0.45613512,0.48357183,0.5624523,0.8162418,1.2929544,1.9685832,1.9823016,2.5927682,3.018037,3.0317552,2.9563043,3.998899,4.681387,5.195825,5.802862,6.848886,7.5588107,8.196714,8.553391,8.738589,9.187865,9.0369625,9.73317,10.6317215,11.190743,10.978109,11.489118,12.116733,12.737488,13.289652,13.780083,13.7526455,13.440554,13.37882,13.87954,15.028452,15.340545,14.664916,14.256795,14.400838,14.411126,13.601744,13.193623,13.21763,13.371962,13.029003,14.006435,14.256795,14.46257,14.5243025,13.522863,12.271064,11.928105,11.547421,11.063849,11.314209,11.694893,11.773774,12.195613,12.96727,13.4474125,13.406258,12.607163,11.773774,11.423956,11.893809,12.943263,13.347955,13.457702,13.7697935,14.953001,15.728088,16.143068,16.187653,15.776102,14.757515,14.815818,14.476289,14.510585,15.117621,15.923574,16.328266,15.9921665,15.436573,14.911846,14.393978,14.582606,14.466,14.339106,14.483148,15.193072,16.506605,17.730967,18.519772,18.62266,17.878439,17.134218,16.592344,16.269962,16.29054,16.863281,17.477179,18.434032,18.999914,18.910746,18.351723,17.960749,16.911295,15.165636,13.118172,11.588576,10.844356,10.405369,9.839486,8.934075,7.6959944,6.392751,5.212973,4.705394,4.746549,4.5339146,4.355576,5.8988905,7.720001,9.349055,11.2593355,11.842365,12.566009,13.5503,14.613472,15.268523,15.014734,15.0078745,14.757515,14.417986,14.784951,14.953001,14.860402,15.090185,15.234227,13.896688,13.567448,13.88983,14.352823,15.049029,16.671225,16.897577,18.025911,18.842154,18.945042,18.742695,19.963629,21.640697,16.859852,9.716022,15.282242,19.092514,15.148488,10.1652975,7.5519514,7.39762,4.8185706,3.5770597,2.6476414,1.6770682,0.97057325,1.0528834,1.5947582,2.585909,3.549623,3.5461934,4.835718,7.997798,7.3427467,3.5221863,3.5290456,4.108646,3.9543142,4.887162,6.3824625,5.562791,6.9037595,7.239859,8.028665,9.3079,9.702303,9.160428,7.9875093,6.8866115,6.1492505,5.6656785,4.5819287,4.1463714,4.0434837,4.098357,4.2766957,4.173808,4.479041,4.5784993,4.32471,4.0366244,5.120374,5.826869,6.060081,5.9812007,6.0223556,5.926327,5.6656785,5.518206,5.4153185,4.9248877,4.976331,5.0483527,4.7979927,4.297273,4.057202,3.9165888,4.0057583,4.0709205,4.0503426,4.0880685,4.448175,4.756838,4.7602673,4.479041,4.187526,4.32471,4.448175,4.431027,4.420738,4.839148,4.671098,4.4104495,4.1155047,3.9063,3.9646032,4.3590055,4.8254294,5.212973,5.597087,6.2692857,6.708273,7.116394,7.267296,7.2638664,7.517656,7.500508,7.4284863,7.298162,7.226141,7.449064,7.7748747,7.891481,7.7920227,7.582818,7.455923,7.4970784,7.6925645,7.857185,8.042382,8.549961,8.697433,8.436785,8.06296,7.5862474,6.728851,6.101236,5.7136927,5.6142344,5.6999745,5.7308407,5.627953,5.6965446,5.778855,5.796003,5.7754254,6.0052075,5.8165803,5.874883,6.1766872,6.036074,6.228131,6.159539,6.574519,7.56224,8.56368,9.362774,10.082987,10.350495,10.233889,10.257896,10.233889,10.63858,11.105004,11.7086115,12.97413,13.982429,14.020154,14.126471,14.472859,14.349394,13.087306,12.277924,11.729189,11.612583,12.449403,12.830087,13.004995,12.816368,12.181894,11.067279,10.05898,9.897789,9.451943,8.512236,7.7680154,7.222711,4.461893,3.9371665,5.267846,3.2375305,2.9391565,1.762808,1.3752645,2.2806756,3.8171308,5.7719955,9.73317,14.205351,17.388008,17.178804,16.403717,8.570539,5.127233,7.040943,4.791134,5.535354,4.57507,4.715683,6.7871537,9.633711,6.924337,8.697433,10.30591,10.714031,12.504276,10.497967,10.024684,10.168727,10.367643,10.439664,11.331357,10.9198065,10.494537,10.182446,8.964942,8.762596,8.2481575,7.8194594,7.6274023,7.5759587,7.0272245,6.8385973,6.451054,5.977771,6.200694,5.2987127,4.8082814,4.3452873,4.214963,5.4084597,6.0875177,6.6533995,7.764586,9.119273,9.445084,8.508806,6.636252,6.355026,7.747438,8.460793,8.930646,9.3593445,9.81205,10.477389,11.657167,12.061859,12.843805,12.9707,12.380811,11.982979,10.72432,9.849775,9.294182,8.906639,8.433355,4.3007026,2.7573884,1.8759843,1.2072148,1.7593783,2.3801336,8.988949,8.913498,2.2326615,1.8073926,1.978872,7.016936,7.346176,2.7059445,2.153781,1.8519772,0.7682276,0.432128,1.5501735,4.0057583,6.9654922,8.584257,8.423067,6.8385973,4.972902,3.3369887,3.899441,4.5167665,4.554492,4.8494368,4.1463714,3.707384,3.858286,4.3349986,4.297273,4.3761535,4.372724,4.3041325,4.232111,4.2835546,4.2869844,4.705394,5.0174866,5.2335505,5.90232,5.857735,6.5882373,7.349606,7.888051,8.464222,9.794902,10.062409,9.945804,9.9698105,10.501397,10.782623,10.844356,11.478829,12.459691,12.528283,12.572867,12.572867,12.562579,12.624311,12.874671,13.22106,13.049581,12.298501,11.166737,10.110424,9.469091,9.462232,9.623423,9.846346,10.381361,9.925226,10.155008,10.72432,11.485688,12.500846,13.478279,13.910407,13.954991,13.841815,13.858963,12.439114,11.074138,10.628291,10.902658,10.6317215,10.748327,10.556271,11.036412,12.061859,12.397959,12.075578,11.002116,10.655728,11.393089,12.445972,12.456262,11.410237,10.124143,9.208443,9.06097,9.352485,10.264755,10.693454,10.213311,9.067829,8.772884,8.573969,8.021805,7.380472,7.6342616,7.966932,8.656279,9.225591,9.458802,9.383351,9.956093,9.287323,8.004657,6.6568294,5.6999745,5.020916,4.787704,4.822,5.1409516,5.960623,6.5470824,7.284444,7.8983397,8.347616,8.831187,8.217292,7.6445503,7.4284863,7.6514096,8.172707,8.141841,7.7440085,7.6959944,8.056101,8.213862,8.289313,8.220721,8.2653055,9.208443,12.370522,10.72775,9.702303,9.414218,9.674867,9.993818,10.093276,9.716022,9.911508,10.80663,11.602294,0.39783216,0.66533995,0.823101,0.922559,1.0563129,1.371835,1.2037852,0.9842916,0.8196714,0.75450927,0.77851635,0.8025235,0.7613684,0.72707254,0.7476501,0.8711152,1.0768905,1.2655178,1.2895249,1.2895249,1.6942163,1.8519772,1.7833855,1.6187652,1.5227368,1.6942163,1.9137098,2.4898806,2.8568463,3.0248961,3.5873485,5.1238036,6.0497923,5.9640527,5.06893,4.166949,3.8960114,3.590778,3.292404,3.059192,2.976882,2.877424,2.8156912,2.5481834,2.2395205,2.4727325,2.7779658,2.8088322,2.7299516,2.702515,2.884283,3.3369887,3.292404,3.1209247,2.9254382,2.5481834,2.8396983,2.7128036,2.49331,2.311542,2.1057668,1.9720128,1.8931323,1.9720128,2.136633,2.136633,1.8313997,1.4610043,1.1934965,1.0357354,0.84024894,0.77851635,0.6790583,0.53844523,0.37382504,0.22978236,0.18176813,0.14061308,0.10288762,0.06859175,0.044584636,0.044584636,0.044584636,0.034295876,0.017147938,0.030866288,0.06859175,0.06859175,0.048014224,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.13375391,0.15776102,0.26750782,0.9362774,2.9151495,3.450165,4.557922,6.3138704,7.857185,7.3701835,4.098357,1.6770682,0.39783216,0.06516216,0.01371835,0.0034295875,0.044584636,0.38754338,1.1111864,2.136633,0.72021335,0.22978236,0.12346515,0.09602845,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.044584636,0.01371835,0.07545093,0.09945804,0.13375391,0.21263443,0.32238123,0.39783216,0.42183927,0.47328308,0.5453044,0.69963586,1.0528834,1.2723769,1.6496316,1.9239986,2.1263442,2.5790498,3.1517909,4.046913,4.8768735,5.6656785,6.835168,7.06838,7.6651278,8.179566,8.505377,8.89635,8.724871,8.683716,9.438225,10.573419,10.573419,10.401938,10.508256,11.290202,12.47341,13.107883,13.070158,13.032433,13.38911,14.05102,14.466,14.661487,13.876111,13.351384,13.238208,12.603734,12.079007,13.001566,13.533153,13.101024,12.404818,13.149038,13.646329,14.057879,14.229359,13.718349,12.288212,11.869802,11.64345,11.38623,11.458252,12.38767,12.764925,13.461131,14.472859,14.939283,14.767803,14.201921,13.275933,12.356804,12.161317,13.55373,13.927555,14.123041,14.514014,15.014734,16.101913,16.904436,17.21996,16.96617,16.173935,16.112202,15.769243,15.426285,15.522313,16.6335,16.21852,15.573756,14.774663,13.96871,13.38225,12.905538,13.107883,13.461131,13.999576,15.306249,15.865272,16.702091,17.350283,17.339994,16.204802,16.252815,16.047039,15.978448,16.352274,17.364002,17.840714,18.574646,19.017063,18.667244,17.04505,16.081335,15.913286,15.46058,14.273943,12.528283,10.916377,10.302481,10.206452,9.89436,8.3922,6.999788,6.550512,6.6568294,6.9380555,7.0478024,6.159539,5.953764,6.64997,7.949784,9.047252,10.7586155,11.897239,12.764925,13.742357,15.306249,15.059319,15.22051,14.79867,13.88297,13.625751,13.625751,14.174485,14.88441,15.227368,14.555169,14.959861,15.470869,16.321407,17.600643,19.270851,19.28457,20.21056,20.19341,19.45262,20.29287,22.19972,21.246294,18.938183,17.528622,20.018501,24.377508,16.064188,9.434795,8.289313,5.861165,3.7108135,2.3046827,1.4438564,0.89855194,0.39783216,0.5693115,1.0220171,1.6256244,2.277246,2.8980014,9.794902,10.871792,8.495089,5.579939,5.56965,7.534804,6.560801,6.7871537,7.98065,5.5387836,7.9429245,8.361334,8.423067,8.882631,9.626852,9.3593445,8.834618,8.018375,7.0306544,6.1629686,5.9812007,5.6965446,4.9831905,4.091498,3.8617156,2.9082901,3.083199,3.4776018,3.5873485,3.2821152,3.6216443,4.5682106,5.501058,5.9126086,5.3878818,5.3981705,5.977771,6.2212715,5.90232,5.4633327,5.0826488,4.8905916,4.650521,4.2423997,3.6319332,3.4124396,3.649081,3.8205605,3.8445675,4.0880685,3.9303071,4.139512,4.307562,4.249259,3.9680326,4.125794,4.3109913,4.245829,4.1429415,4.729401,4.4721823,4.383013,4.173808,3.8788633,3.8308492,4.341858,4.763697,5.24041,5.8543057,6.6225333,6.6705475,7.15069,7.449064,7.455923,7.5519514,7.466212,7.3255987,7.2124224,7.133542,7.034084,7.1061053,6.9620624,6.8385973,6.807731,6.759717,6.8214493,6.8900414,7.051232,7.366754,7.905199,8.344186,8.097256,7.716572,7.363324,6.790583,6.046363,5.693115,5.6039457,5.658819,5.768566,6.183546,6.468202,6.475061,6.228131,5.936616,6.1561093,6.036074,5.8165803,5.5730796,5.219832,5.744559,5.874883,6.23499,6.9037595,7.414768,7.6616983,9.002667,9.668007,9.609704,10.511685,10.096705,10.268185,10.477389,10.714031,11.519984,14.085316,14.778092,14.479718,13.910407,13.642899,13.972139,13.63261,12.679185,11.739478,12.010415,13.485138,14.1299,13.612033,12.507706,12.312219,11.324498,10.792912,10.4533825,9.781183,8.011517,8.073249,6.3207297,3.841138,2.7368107,6.118384,3.642222,1.9857311,1.371835,2.0097382,4.1360826,9.568549,12.864383,15.789821,17.899017,16.554619,11.012405,6.444195,5.051782,5.9880595,5.3398676,4.962613,3.7794054,4.6093655,6.90033,6.728851,6.166398,8.793462,10.237319,10.515115,14.006435,13.334236,12.445972,11.814929,11.612583,11.674315,11.784062,11.2421875,10.88894,10.63858,9.489669,9.6988735,8.597976,7.9189177,8.30646,9.3079,7.548522,7.548522,7.2021337,6.15268,5.7994323,5.2987127,5.521636,5.545643,5.23698,5.2506986,6.1149545,7.6857057,9.016385,10.179015,12.253916,10.64201,6.557371,5.15467,7.1781263,8.971801,8.251588,8.4093485,9.160428,10.096705,10.679735,12.072148,12.703192,12.507706,11.996697,12.253916,11.228469,11.026124,11.331357,10.909517,7.613684,4.389872,3.0351849,2.0063086,1.1351935,1.6496316,5.689686,4.5099077,4.461893,5.885172,3.1140654,2.7573884,7.795452,9.6817255,6.036074,0.64133286,1.1283343,0.52815646,0.58302987,1.3821237,1.3581166,3.7005248,8.086967,8.433355,5.2266912,5.5079174,4.32471,4.5853586,4.6848164,4.1429415,3.6147852,3.6147852,3.5050385,3.865145,4.431027,4.0880685,4.5784993,4.5990767,4.7328305,5.0655007,5.188966,4.5167665,5.127233,5.535354,5.4633327,5.830299,5.90232,6.4064693,7.051232,7.671987,8.210432,9.770895,10.326488,10.576848,11.036412,12.037852,11.893809,12.569438,13.399398,13.869251,13.625751,13.272504,13.083877,12.764925,12.312219,12.010415,11.982979,12.517994,12.860953,12.576297,11.550851,9.962952,8.460793,7.8983397,8.501947,9.856634,10.55284,10.827208,11.231899,12.133881,13.732068,13.354814,13.670336,13.9481325,13.759505,13.015285,11.489118,10.669447,10.467101,10.645439,10.803201,10.998687,10.55284,10.707172,11.667457,12.617453,12.617453,11.015835,10.405369,11.149589,11.382801,11.640019,10.960961,9.654288,8.450503,8.498518,9.719451,11.252477,11.71547,10.7757635,9.139851,9.287323,9.644,9.589127,9.074688,8.635701,8.97866,9.849775,10.607714,10.88551,10.604284,11.118723,9.863494,8.213862,6.9346256,6.1629686,5.346727,5.0140567,5.209543,5.7651367,6.3001523,7.377043,8.083538,8.241299,8.001227,7.8434668,8.100685,7.486789,7.5210853,8.196714,7.963502,8.049242,7.8434668,7.7577267,7.970361,8.423067,8.508806,8.676856,8.700864,8.625413,8.759167,8.831187,9.187865,9.407358,9.750318,11.153018,11.948683,11.633161,11.561139,12.055,12.421966,0.6036074,0.78537554,0.8848336,0.9534253,1.0254467,1.1283343,0.939707,0.8779744,0.8745448,0.8745448,0.84024894,0.9431366,0.980862,0.9911508,1.0117283,1.0666018,1.1077567,1.2483698,1.4232788,1.5844694,1.6942163,1.8039631,1.7799559,1.6942163,1.6667795,1.8759843,2.7711067,3.426158,3.7142432,3.8274195,4.280125,5.096367,5.219832,4.99005,4.605936,4.105216,3.7108135,3.4021509,3.1620796,3.100347,3.4638834,3.1895163,2.952875,2.9048605,2.9906003,2.959734,3.1277838,3.2581081,3.4638834,3.649081,3.4707425,3.5016088,3.0111778,2.551613,2.2909644,2.0097382,1.7971039,1.7319417,1.7696671,1.8485477,1.8862731,1.8313997,1.9754424,2.0063086,1.8382589,1.6221949,1.2895249,1.0597426,0.89855194,0.764798,0.607037,0.52815646,0.47671264,0.4046913,0.29837412,0.18176813,0.13032432,0.106317215,0.08573969,0.058302987,0.034295876,0.024007112,0.0274367,0.030866288,0.0274367,0.030866288,0.037725464,0.037725464,0.044584636,0.044584636,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.037725464,0.09602845,0.35324752,0.9877212,2.194936,3.0729103,3.998899,4.9180284,5.576509,5.528495,2.7230926,1.0357354,0.25721905,0.07545093,0.06516216,0.14061308,0.29837412,0.5727411,1.0185875,1.7216529,2.7951138,2.6545007,1.4472859,0.048014224,0.058302987,0.030866288,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.08573969,0.017147938,0.010288762,0.010288762,0.0034295875,0.01371835,0.020577524,0.041155048,0.09602845,0.18519773,0.28808534,0.29151493,0.36696586,0.490431,0.64476246,0.83338976,0.88826317,1.1763484,1.471293,1.704505,1.9823016,2.4452958,2.9494452,3.4673128,4.149801,5.3227196,6.0806584,6.6293926,7.1369715,7.654839,8.114404,8.519095,8.796892,8.855195,8.81747,9.012956,9.56512,9.935514,10.566559,11.588576,12.840376,12.792361,13.337666,13.567448,13.241637,12.816368,12.212761,11.814929,11.996697,12.377381,11.8115,12.408247,12.864383,12.857523,12.312219,11.393089,12.401388,12.994707,13.162757,13.077017,13.070158,11.4754,11.986408,12.600305,12.5145645,12.120162,13.241637,13.762935,14.3974085,15.37827,16.475739,15.6526375,14.534592,13.567448,13.063298,13.210771,13.900118,14.208781,14.599753,15.086755,15.234227,15.96816,16.616352,17.110212,17.274832,16.832415,16.822126,16.47231,16.20137,16.256245,16.743246,16.239098,15.199932,14.579176,14.273943,13.114742,13.039291,13.059869,13.38225,14.181344,15.635489,15.913286,15.885849,16.081335,16.287111,15.580616,15.268523,15.014734,15.196502,15.96816,17.254255,18.269413,18.30028,18.053349,17.717249,16.983316,15.649208,14.479718,14.092175,14.153908,13.392539,11.852654,11.005547,10.926665,11.197603,10.906088,8.920357,7.641121,6.893471,6.8214493,7.8674736,8.762596,8.354475,7.7268605,7.4936485,7.7920227,9.832627,11.122152,12.003556,12.768354,13.656617,14.438563,15.4742985,15.165636,13.71492,13.138749,14.027013,14.013294,14.147048,14.733508,15.350834,15.645778,16.191082,17.346853,18.728977,19.198832,20.7833,20.845032,20.063087,20.069946,23.43094,23.732746,20.52951,19.325726,21.637268,24.987974,22.168854,13.978998,7.7714453,5.8543057,5.504488,4.5270553,2.4247184,1.0151579,0.7133542,0.5555932,2.085189,2.6956558,2.8877127,2.976882,3.083199,7.0203657,7.6342616,8.1212635,9.273604,9.47595,9.537683,8.512236,8.30646,8.594546,6.807731,8.64599,9.671436,9.345626,8.285883,8.2481575,7.864044,8.628842,8.628842,7.56224,6.715132,6.7665763,7.1198235,7.130112,6.416758,4.835718,3.3952916,2.8980014,2.976882,3.2992632,3.549623,3.3644254,3.4467354,3.9508848,4.6093655,4.73969,5.1238036,5.4496145,5.593657,5.576509,5.5833683,5.0106273,4.5922174,4.3349986,4.1120753,3.6696587,3.5839188,3.316411,3.3438478,3.683377,3.8685746,3.974892,4.623084,4.7979927,4.3349986,3.9063,4.232111,4.2526884,4.1292233,3.9063,3.5461934,3.3884325,3.415869,3.4913201,3.6593697,4.1463714,4.6127954,5.2026844,5.8062916,6.3035817,6.584808,6.7631464,7.010077,7.157549,7.2295704,7.442205,7.56224,7.4524937,7.3050213,7.191845,7.034084,7.1369715,7.1232533,6.975781,6.807731,6.8557453,7.2295704,7.0786686,7.0032177,7.15069,7.208993,7.099246,6.9963584,6.948344,6.989499,7.1198235,6.893471,6.39961,6.0154963,5.909179,6.0497923,6.3447366,6.852316,7.016936,6.725421,6.3138704,5.9880595,5.686256,5.610805,5.686256,5.597087,5.768566,5.7994323,6.0532217,6.4990683,6.7185616,7.2947326,8.385342,9.338767,10.076128,11.087856,10.731179,10.834066,11.159878,11.653738,12.459691,13.440554,14.263655,14.5585985,14.277372,13.666906,13.293081,13.173045,12.847235,12.154458,11.252477,11.399949,12.6929035,12.902108,11.849225,11.399949,11.375941,10.521975,10.161868,10.031544,8.279024,7.9292064,6.948344,5.2815647,3.8034124,4.3109913,4.15666,2.4487255,1.313532,1.5330256,2.5241764,6.2864337,6.6636887,6.8385973,7.7440085,8.073249,5.439326,4.400161,4.636802,5.3090014,5.07236,5.103226,4.4550343,5.329579,7.4284863,7.963502,7.449064,8.868914,10.209882,11.005547,12.346515,12.487128,12.55229,11.729189,10.405369,10.182446,11.183885,11.780633,12.109874,11.8115,10.028113,10.401938,9.517105,8.786603,8.827758,9.465661,8.255017,8.018375,7.6514096,6.927767,6.495639,6.715132,6.5196457,6.3721733,6.334448,6.0532217,6.444195,7.610255,7.966932,8.453933,12.521424,9.054111,9.472521,9.132992,7.7440085,9.362774,10.333347,10.714031,10.943813,11.214751,11.499407,12.30536,13.337666,13.564018,12.960411,12.535142,10.717461,11.012405,11.351934,11.019264,10.652299,6.5710897,3.8377085,2.318401,2.452155,5.2472687,8.577398,6.101236,7.431916,11.146159,4.7602673,5.1683884,4.787704,3.6182148,1.9342873,0.28808534,0.41498008,0.2194936,0.37382504,0.7922347,0.65162164,3.3369887,3.8137012,2.8088322,1.8245405,3.1415021,2.5241764,2.8534167,2.9906003,2.7093742,2.702515,2.8294096,2.7779658,3.5359046,4.4104495,3.0626216,3.8274195,3.9165888,4.1120753,4.756838,5.7377,4.9488945,5.288424,5.7068334,5.9743414,6.6705475,6.9689217,7.160979,7.750868,8.532814,8.601405,9.448513,9.884071,10.247607,10.583707,10.6488695,10.89237,11.499407,12.044711,12.428825,12.857523,12.71691,12.939834,12.857523,12.397959,12.092726,12.507706,12.487128,12.4974165,12.487128,11.893809,11.605724,10.381361,9.781183,10.244178,11.101575,11.015835,11.814929,12.710052,13.498857,14.55174,14.592895,14.822677,15.001016,14.846684,14.054449,12.528283,12.085866,11.670886,11.091286,11.036412,11.163307,10.854645,10.487679,10.521975,11.482259,11.835506,10.827208,10.295622,10.744898,11.345076,11.612583,10.813489,10.048691,9.822338,10.038403,10.604284,11.818358,12.600305,12.445972,11.434244,10.830637,10.655728,10.501397,10.117283,9.3936405,9.880642,10.659158,11.201033,11.365653,11.399949,10.88551,10.010965,9.129561,8.200144,6.7871537,6.0086374,5.4084597,5.535354,6.324159,7.0958166,7.5725293,7.4970784,7.010077,6.6293926,7.233,7.5279446,7.407909,7.781734,8.515666,8.440215,7.8434668,7.6274023,7.829748,8.275595,8.570539,8.625413,8.200144,8.244728,8.659708,8.296172,9.15014,9.619993,10.079557,10.751757,11.71547,12.840376,12.830087,12.281353,11.684605,11.406808,0.6001778,0.6927767,0.8128122,0.94656616,1.0837497,1.2037852,1.1729189,1.0700313,1.0048691,0.9774324,0.89169276,0.9842916,0.980862,0.9945804,1.0597426,1.1420527,1.2963841,1.4061309,1.6016173,1.8348293,1.8965619,1.920569,1.879414,1.9102802,2.136633,2.6647894,3.4638834,3.899441,4.1360826,4.338428,4.6573796,4.8905916,4.8254294,4.5682106,4.184097,3.6868064,3.223812,2.9665933,2.9322972,3.059192,3.192946,3.3369887,3.4021509,3.3815732,3.3301294,3.357566,3.6456516,3.6147852,3.666229,3.782835,3.542764,2.9631636,2.5310357,2.1640697,1.8759843,1.7662375,1.6016173,1.646202,1.6530612,1.5536032,1.4369972,1.546744,1.6633499,1.6153357,1.4198492,1.2758065,1.0734608,0.96714365,0.83338976,0.64476246,0.48357183,0.42183927,0.38754338,0.32924038,0.24007112,0.16804978,0.12689474,0.09602845,0.06516216,0.037725464,0.020577524,0.017147938,0.01371835,0.020577524,0.0274367,0.020577524,0.020577524,0.017147938,0.041155048,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.14061308,0.44584638,0.9328478,1.529596,2.7333813,4.187526,5.8508763,7.040943,6.420188,2.9288676,1.1420527,2.3081124,5.0586414,5.40503,2.2806756,1.2415106,0.97400284,0.9259886,1.3169615,1.8554068,2.0749004,1.2929544,0.044584636,0.06859175,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.044584636,0.11317638,0.18519773,0.24350071,0.30866286,0.4081209,0.53844523,0.6790583,0.72021335,0.89169276,1.097468,1.2895249,1.4541451,1.8725548,2.352697,2.7128036,3.1449318,4.2218223,4.7602673,5.188966,5.6176643,6.0806584,6.5539417,7.4113383,8.176137,8.546532,8.615124,8.858624,9.102125,9.534253,10.233889,11.245617,12.562579,12.689473,12.665466,12.517994,12.312219,12.168177,11.22161,11.105004,11.506266,11.938394,11.749766,12.627741,12.648318,12.264205,11.691463,10.9198065,11.729189,12.528283,12.452832,11.670886,11.351934,10.405369,10.998687,11.862943,12.281353,12.082437,13.101024,14.102464,15.193072,16.146498,16.420864,15.776102,14.678635,13.742357,13.371962,13.766364,14.088745,14.174485,14.579176,15.172495,15.151917,16.019604,16.63007,16.760393,16.691803,17.21653,16.7844,16.170506,15.769243,15.707511,15.854982,15.138199,14.222499,13.570878,13.004995,11.701753,12.30193,12.339656,12.7272,13.7938,15.278812,15.666355,15.899568,16.067617,15.964729,15.097044,14.71636,14.490007,14.949572,16.101913,17.429163,18.61923,18.79414,18.238546,17.271402,16.252815,15.278812,14.452282,14.160767,14.2533655,14.030442,13.193623,12.528283,12.13731,11.986408,11.910957,10.882081,9.81205,8.875772,8.357904,8.666568,9.510246,9.606275,9.126132,8.495089,8.40249,8.656279,9.72288,11.194174,12.542002,13.118172,13.684054,14.099034,13.958421,13.430264,13.262215,13.786942,13.687484,13.574307,13.80066,14.441993,14.832966,16.153357,17.682953,18.982767,19.895037,22.048819,22.648996,22.830763,23.719027,26.448978,26.658184,25.505842,24.665592,24.284908,22.981665,17.20281,10.576848,5.5079174,3.40901,4.695105,3.474172,2.0097382,1.0871792,0.8196714,0.65848076,1.546744,3.3987212,5.4804807,6.999788,7.130112,7.390761,7.208993,8.584257,10.947243,11.166737,10.525404,10.271614,9.89093,9.078118,7.740579,8.543102,8.923786,8.611694,7.9943686,8.1041155,7.764586,8.7145815,8.875772,7.915488,7.2707253,7.442205,6.8591747,6.4304767,6.135532,5.0277753,3.4192986,2.8739944,2.7882545,2.8739944,3.1689389,2.9220085,3.1552205,3.4776018,3.7691166,4.166949,4.5099077,4.698535,4.7019644,4.5990767,4.588788,4.5682106,4.5990767,4.4756117,4.187526,3.923448,4.057202,3.6627994,3.5153272,3.7759757,4.0057583,4.0606318,4.4584637,4.633373,4.4550343,4.249259,4.3658648,4.2698364,4.0777793,3.765687,3.1689389,3.2443898,3.4878905,3.7279615,3.9508848,4.307562,4.804852,5.504488,6.111525,6.461343,6.5299344,6.5470824,6.7219915,6.869464,7.0203657,7.4353456,7.671987,7.6445503,7.414768,7.143831,7.0889573,7.0958166,6.941485,6.7665763,6.725421,6.9723516,7.2192817,7.284444,7.2535777,7.157549,6.9792104,6.910619,6.883182,6.869464,6.90033,7.06495,7.1369715,6.776865,6.341307,6.060081,6.046363,6.262427,6.543653,6.5642304,6.324159,6.135532,5.919468,5.6656785,5.586798,5.675967,5.672538,5.641671,5.597087,5.7102633,5.9914894,6.307011,7.016936,8.1212635,9.235879,10.199594,11.084427,11.094715,11.434244,11.64345,11.873232,12.905538,13.169616,13.63261,13.906977,13.872682,13.680624,13.512574,12.956982,12.274493,11.646879,11.153018,10.926665,11.982979,12.490558,11.958971,11.231899,11.293632,10.31277,9.692014,9.506817,8.501947,7.5759587,6.6053853,5.4941993,4.616225,4.8117113,4.57164,3.093488,1.704505,1.1523414,1.6256244,3.3301294,3.6216443,3.4810312,3.5633414,4.173808,3.9200184,3.9646032,4.431027,4.9660425,4.7671266,5.686256,5.844017,6.3035817,7.2878733,8.179566,8.577398,9.3764925,10.30934,11.197603,11.914387,11.406808,11.681175,10.998687,9.609704,9.757176,9.877212,10.326488,11.0981455,11.650309,10.8958,10.388221,9.832627,9.345626,9.006097,8.827758,8.632272,8.06296,7.459353,7.1129646,7.2535777,7.473071,7.2467184,6.9346256,6.7494283,6.7700057,7.1781263,8.375052,8.903209,8.450503,7.8366075,8.381912,9.105555,8.776315,7.9292064,8.875772,11.153018,11.852654,11.838936,11.770344,12.079007,11.897239,13.395968,14.263655,13.738928,12.614022,11.543991,12.133881,12.548861,12.21962,11.852654,8.916927,5.1238036,2.4555845,2.3595562,5.7754254,6.615674,5.6039457,7.257007,9.770895,5.0174866,4.7808447,2.9460156,1.5193073,0.97057325,0.22635277,0.17490897,0.08916927,0.22292319,0.48014224,0.41840968,1.6016173,1.3684053,0.8162418,0.7339317,1.6153357,1.5261664,1.9823016,2.3801336,2.417859,2.0886188,2.5824795,2.5138876,3.1243541,3.9886103,2.9906003,3.981751,4.3041325,4.3624353,4.6745276,5.892031,5.3090014,5.377593,5.5113473,5.751418,6.7459984,7.675417,8.213862,8.772884,9.15014,8.522525,8.673427,9.455373,10.323058,10.827208,10.621432,10.967821,11.252477,11.489118,11.739478,12.096155,11.938394,12.445972,12.88496,12.987847,12.939834,13.522863,13.320518,12.915827,12.610593,12.445972,12.284782,11.766914,11.30049,11.019264,10.799771,10.981539,12.003556,13.152468,14.13676,15.066177,15.731518,16.002455,15.772673,15.12448,14.30481,13.238208,12.943263,12.524854,11.921246,11.897239,11.664027,11.050131,10.381361,10.082987,10.696883,11.619442,11.177026,10.847785,11.087856,11.338216,10.9541025,10.110424,9.592556,9.6817255,10.120712,10.4705305,10.491108,10.978109,11.63659,11.074138,10.326488,10.155008,10.347065,10.549411,10.261326,10.271614,11.002116,11.543991,11.808069,12.511135,12.123591,11.324498,10.371073,9.318189,8.014946,7.099246,6.667118,6.8591747,7.4970784,8.107545,8.093826,7.4799304,6.728851,6.2418494,6.375603,6.6431108,6.944915,7.514226,8.110974,8.038953,7.8846216,7.8091707,7.9463544,8.282454,8.64256,8.903209,8.752307,8.800322,9.0369625,8.827758,9.554831,10.034973,10.621432,11.321068,11.8115,13.149038,13.265644,12.562579,11.550851,10.823778,0.5453044,0.71678376,0.9328478,1.138623,1.2998136,1.4129901,1.4267083,1.2895249,1.1763484,1.138623,1.0940384,1.1351935,1.0871792,1.1283343,1.2620882,1.3238207,1.5604624,1.6599203,1.8073926,2.0028791,2.0714707,1.9857311,1.9514352,2.1126258,2.4967396,3.0317552,3.6627994,4.0366244,4.341858,4.616225,4.7431192,4.465323,4.4413157,4.214963,3.6696587,3.0077481,2.6922262,2.503599,2.5550427,2.750529,2.784825,3.3850029,3.758828,3.8274195,3.707384,3.7108135,3.7485392,3.508468,3.3061223,3.199805,3.0077481,2.3595562,2.1469216,1.9720128,1.7593783,1.7353712,1.6290541,1.6976458,1.6290541,1.3786942,1.1797781,1.2723769,1.4061309,1.4129901,1.2826657,1.1592005,0.9945804,0.8711152,0.7133542,0.5418748,0.44927597,0.4046913,0.35324752,0.2777966,0.1920569,0.15090185,0.12346515,0.082310095,0.044584636,0.024007112,0.01371835,0.010288762,0.024007112,0.030866288,0.020577524,0.010288762,0.01371835,0.006859175,0.024007112,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.05144381,0.1371835,0.45956472,0.9534253,1.2895249,2.6613598,4.180667,6.5230756,8.961512,9.338767,5.24041,2.411,3.2581081,7.0923867,10.134431,4.4550343,2.7162333,1.9857311,1.2449403,1.3958421,0.939707,1.0700313,0.7579388,0.044584636,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.05144381,0.082310095,0.15090185,0.20920484,0.28465575,0.37725464,0.48700142,0.53844523,0.65848076,0.8093826,0.97057325,1.1249046,1.4164196,1.8999915,2.2429502,2.5310357,3.275256,3.4192986,3.7519686,4.180667,4.6402316,5.096367,6.2898636,7.222711,7.8091707,8.182996,8.694004,8.711152,9.242738,9.880642,10.528833,11.372512,11.756626,11.509696,11.255906,11.204462,11.14273,10.861504,11.492548,12.106443,12.260776,11.993267,12.843805,12.761495,12.30536,11.80121,11.345076,11.996697,12.5145645,12.161317,11.091286,10.371073,9.853205,10.065839,10.628291,11.252477,11.732618,12.277924,13.581166,15.169065,16.314548,16.050468,15.902997,15.090185,14.345964,14.092175,14.46257,14.579176,14.345964,14.404267,14.7026415,14.510585,15.179354,15.741806,15.885849,15.927004,16.798119,16.348843,15.590904,15.004445,14.812388,14.96329,14.174485,13.354814,12.593445,11.821788,10.820349,11.660598,11.739478,12.30193,13.529722,14.538021,15.481158,17.065628,16.763824,14.767803,13.954991,14.459141,14.562028,15.234227,16.619781,18.063637,18.728977,18.993055,18.612371,17.645227,16.492886,15.4742985,14.953001,14.812388,14.826107,14.678635,14.404267,14.0750265,13.708061,13.37882,13.227919,12.9809885,12.336226,11.561139,10.840926,10.285333,10.484249,10.734609,10.539123,9.897789,9.294182,8.783174,9.431366,10.796341,12.113303,12.30536,12.7272,12.421966,12.116733,12.271064,13.066729,13.577737,13.821238,13.910407,14.023583,14.3974085,15.0250225,16.606062,18.115082,19.404606,21.187992,22.53925,23.876787,25.231476,26.531288,27.577312,29.449867,30.50961,28.359259,23.839062,21.067955,13.817808,8.618553,4.437886,1.9445761,3.4981792,2.318401,1.4781522,1.0220171,0.88826317,0.89855194,1.08032,3.7931237,6.3207297,7.534804,7.8674736,7.6857057,7.7714453,9.3079,11.447963,11.324498,10.295622,10.268185,9.9698105,9.023245,7.9600725,7.891481,7.6925645,7.349606,7.0375133,7.133542,7.675417,8.81061,9.06097,8.340756,7.98065,8.1487,6.944915,5.953764,5.5902276,5.0757895,3.3987212,3.1586502,3.083199,2.8465576,3.0386145,2.7470996,3.1586502,3.4810312,3.5599117,3.8788633,4.046913,4.0846386,4.016047,3.858286,3.642222,4.046913,4.3795834,4.4584637,4.3109913,4.149801,4.2938433,4.091498,3.940596,4.012617,4.2526884,4.197815,4.3349986,4.413879,4.40359,4.4687524,4.57507,4.506478,4.3178506,4.0057583,3.4913201,3.7485392,4.0880685,4.372724,4.5819287,4.804852,5.144381,5.6313825,6.077229,6.3653145,6.475061,6.2967224,6.468202,6.800872,7.1884155,7.5931067,7.740579,7.795452,7.610255,7.3393173,7.442205,7.2535777,7.0032177,6.866034,6.931196,7.181556,7.301592,7.191845,6.9689217,6.7802944,6.807731,6.9071894,6.931196,6.8557453,6.728851,6.711703,6.7974424,6.4887795,6.108095,5.8645945,5.8508763,6.0223556,6.018926,5.909179,5.7651367,5.6348124,5.9160385,5.7925735,5.6999745,5.754848,5.751418,5.7411294,5.720552,5.7925735,5.9400454,6.046363,6.910619,7.9943686,9.012956,9.832627,10.436234,10.587136,11.118723,11.447963,11.660598,12.504276,12.655178,13.193623,13.540011,13.564018,13.564018,13.96871,13.5503,12.524854,11.454823,11.2593355,11.22161,11.835506,12.346515,12.298501,11.537132,11.303921,10.569988,9.935514,9.455373,8.659708,7.7783046,6.835168,5.874883,5.219832,5.4770513,5.096367,3.806842,2.3218307,1.3992717,1.8416885,2.6887965,2.8945718,2.702515,2.4727325,2.6853669,4.139512,4.15323,4.262977,4.715683,4.4550343,5.662249,6.433906,6.8626046,7.250148,8.1041155,9.194724,9.97324,10.542552,10.967821,11.266195,10.573419,10.762046,10.124143,8.968371,9.602845,9.369633,9.493098,10.257896,11.341646,11.828648,10.645439,10.024684,9.568549,8.992378,8.1384115,8.64256,8.014946,7.377043,7.2604365,7.630832,7.798882,7.98408,7.7028537,7.160979,7.233,7.7542973,8.721441,9.31133,8.711152,6.1458206,7.2295704,6.6876955,6.601956,7.466212,8.186425,10.686595,11.825217,11.893809,11.650309,12.291641,11.55771,12.987847,13.954991,13.615462,12.905538,13.13532,13.577737,13.728639,12.929544,10.377932,9.218731,5.4907694,2.435007,2.085189,5.254128,4.5990767,5.6142344,7.1781263,7.8777623,6.0223556,4.355576,2.2052248,1.0563129,0.939707,0.42183927,0.2777966,0.3566771,0.6927767,0.99801,0.66191036,0.6241849,0.7099246,0.6927767,0.6207553,0.8265306,1.1008976,1.371835,1.8313997,2.2326615,1.8931323,2.8911421,2.976882,3.3266997,3.9440255,3.649081,4.0057583,4.3452873,4.48933,4.7328305,5.8371577,5.4599032,5.4736214,5.5147767,5.6999745,6.6396813,7.9943686,8.906639,9.541112,9.729739,8.992378,8.831187,9.9698105,11.170166,11.705182,11.369082,11.749766,11.790922,11.633161,11.38623,11.132441,10.933525,11.273054,11.821788,12.373952,12.840376,13.443983,13.653188,13.313659,12.761495,12.836946,12.542002,12.456262,11.852654,10.89237,10.604284,11.0981455,11.993267,13.169616,14.38026,15.237658,16.13278,16.424294,16.084764,15.343974,14.675205,13.810948,13.701202,13.526293,13.066729,12.71691,12.312219,11.355364,10.429376,10.000677,10.398509,11.540562,11.808069,11.818358,11.873232,11.958971,11.482259,10.755186,10.189304,9.925226,9.832627,10.652299,9.705732,9.3079,9.825768,9.671436,9.033533,9.434795,10.278474,10.981539,10.9541025,10.669447,11.321068,11.893809,12.343085,13.591455,13.965281,13.419975,12.343085,11.019264,9.619993,8.594546,8.501947,8.937505,9.530824,9.928656,9.352485,8.519095,7.5862474,6.7700057,6.355026,6.210983,6.392751,6.7974424,7.1712675,7.130112,7.56224,7.764586,7.970361,8.2653055,8.618553,9.026674,9.451943,9.592556,9.431366,9.256456,9.836057,10.179015,10.744898,11.482259,11.797781,12.878101,12.9981365,12.336226,11.283342,10.446524,0.59674823,0.90541106,1.1763484,1.3821237,1.4987297,1.4987297,1.4438564,1.3615463,1.3066728,1.2998136,1.3169615,1.3238207,1.3203912,1.4507155,1.6633499,1.7010754,1.8759843,1.9548649,2.0063086,2.054323,2.085189,1.9514352,2.0097382,2.2669573,2.609916,2.8088322,3.4433057,3.899441,4.2766957,4.537344,4.496189,4.0057583,3.9783216,3.765687,3.1723683,2.4555845,2.3286898,2.1674993,2.1503513,2.3252604,2.5961976,3.2992632,3.7211025,3.8720043,3.7862647,3.5564823,3.1415021,2.8499873,2.6167753,2.4144297,2.2120838,2.0303159,1.9651536,1.9137098,1.8416885,1.7936742,1.6633499,1.6324836,1.5090185,1.2963841,1.1763484,1.1111864,1.3375391,1.4678634,1.3546871,1.1008976,0.89169276,0.6824879,0.5212973,0.4389872,0.48014224,0.42183927,0.33266997,0.24007112,0.16119061,0.12003556,0.10288762,0.0548734,0.024007112,0.01371835,0.01371835,0.0034295875,0.044584636,0.048014224,0.010288762,0.010288762,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08916927,0.061732575,0.37382504,1.0151579,1.5158776,2.760818,3.9646032,6.252138,9.294182,11.290202,7.840037,4.0537724,2.5824795,4.7534084,10.556271,5.312431,4.2183924,3.3712845,1.8862731,1.8862731,1.1249046,0.7990939,0.4424168,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.07888051,0.15433143,0.22978236,0.2777966,0.30866286,0.42526886,0.5658819,0.72707254,0.9431366,1.08032,1.4575747,1.8279701,2.1297739,2.4795918,2.452155,2.6887965,3.1243541,3.6559403,4.1635194,5.5559316,6.2555676,6.5813785,6.927767,7.750868,8.038953,8.752307,9.177576,9.235879,9.445084,9.97667,10.155008,10.237319,10.192734,9.6817255,10.587136,12.037852,12.919256,12.850664,12.171606,13.011855,13.015285,12.651748,12.346515,12.476839,13.05301,12.943263,12.308789,11.396519,10.545981,10.244178,10.14472,10.275044,10.796341,12.006986,11.862943,12.912396,14.417986,15.618341,15.731518,15.830976,15.477728,15.175924,15.110763,15.110763,15.011304,14.493437,14.171056,14.081886,13.687484,13.653188,14.0750265,14.654627,15.169065,15.481158,15.323397,14.623761,13.965281,13.711491,14.006435,13.282792,12.428825,11.63659,11.087856,10.9369545,11.622872,11.797781,12.562579,13.7697935,14.003006,16.29397,19.46291,17.809847,12.542002,11.760056,14.270514,15.155347,15.906426,17.168514,18.763273,18.595222,18.506054,18.420315,18.159666,17.463459,16.163645,15.512024,15.402277,15.532601,15.374841,15.251375,15.117621,15.110763,15.182784,15.117621,15.086755,14.685493,14.105893,13.437123,12.686044,12.377381,12.027563,11.63659,11.111863,10.264755,10.213311,10.240748,10.635151,11.207891,11.317638,12.055,11.447963,10.731179,10.81006,12.247057,13.13532,13.906977,14.610043,15.179354,15.440002,16.362562,17.528622,18.739265,20.2037,22.52896,22.62156,24.586712,26.565584,27.580742,27.52587,31.891733,33.465916,28.880556,21.28059,20.316875,12.315649,7.7542973,4.173808,1.5570327,2.3389788,1.7971039,1.2003556,0.8745448,0.9602845,1.3958421,1.7525192,4.6127954,6.166398,5.8474464,6.3173003,7.857185,8.992378,10.573419,12.127021,11.825217,10.446524,9.760606,9.349055,8.824328,7.81603,7.281014,7.0135064,6.5882373,6.0395036,5.8543057,7.099246,8.285883,8.676856,8.412778,8.519095,8.790032,8.049242,7.023795,6.166398,5.689686,3.7862647,3.57363,3.5221863,3.2683969,3.590778,3.0043187,3.2032347,3.4913201,3.6216443,3.799983,3.8857226,3.8171308,3.7794054,3.74168,3.4192986,3.666229,3.899441,4.2183924,4.4756117,4.2595477,4.266407,4.338428,4.307562,4.245829,4.4584637,4.5030484,4.6608095,4.6745276,4.5990767,4.8014226,4.9248877,4.8734436,4.722542,4.5339146,4.341858,4.705394,4.8940215,5.0586414,5.302142,5.6519604,5.703404,5.826869,6.0566516,6.327589,6.461343,6.2247014,6.3310184,6.824879,7.438775,7.596536,7.5725293,7.7097125,7.7714453,7.7920227,8.080108,7.8091707,7.5931067,7.500508,7.517656,7.5519514,7.740579,7.239859,6.694555,6.5196457,6.883182,6.9826403,7.06838,6.9517736,6.6293926,6.2967224,6.101236,5.6965446,5.4153185,5.3981705,5.5730796,5.672538,5.535354,5.470192,5.4736214,5.24041,6.0223556,6.0154963,5.885172,5.892031,5.90232,6.142391,6.2487082,6.3481665,6.368744,6.036074,6.9723516,7.8091707,8.488229,8.985519,9.31133,9.314759,9.956093,10.840926,11.619442,11.979549,12.157887,13.101024,13.824667,13.900118,13.440554,14.003006,14.520873,13.9138365,12.442543,11.705182,11.8869505,12.21962,12.517994,12.566009,12.099585,11.602294,11.317638,10.947243,10.288762,9.235879,8.827758,8.038953,6.869464,5.761707,5.610805,5.751418,4.856296,3.3369887,2.1297739,2.6956558,4.201245,3.549623,2.7573884,2.5310357,2.2841053,4.5853586,4.4721823,4.297273,4.616225,4.190956,5.007198,5.878313,6.64997,7.3084507,7.9737906,9.15014,10.326488,10.748327,10.419086,10.096705,10.172156,10.278474,9.534253,8.543102,9.373062,9.678296,10.000677,10.611144,11.543991,12.600305,11.526843,10.515115,9.716022,8.992378,7.939495,8.371623,7.9875093,7.6959944,7.7851634,7.932636,8.255017,8.97866,8.916927,8.131552,7.939495,8.217292,8.553391,8.820899,8.762596,7.956643,6.0326443,4.0949273,4.48933,6.725421,7.466212,9.263316,11.050131,11.619442,11.393089,12.411677,11.986408,12.80265,13.186764,12.953552,13.38225,14.160767,14.325387,14.452282,13.241637,7.5107965,7.281014,4.4927597,2.3904223,2.510458,4.650521,4.8185706,7.390761,8.855195,8.707723,9.441654,5.1169443,2.609916,1.8176813,2.3458378,3.508468,1.2380811,1.3272504,1.961724,2.9288676,5.593657,2.3767042,1.6496316,1.2689474,0.6036074,0.53158605,0.82996017,0.7442205,1.0837497,1.8142518,2.085189,3.2443898,3.6044965,3.7965534,4.0674906,4.2698364,3.8891523,4.1463714,4.461893,4.7774153,5.5559316,5.360445,5.528495,5.7308407,5.9640527,6.5642304,7.9875093,9.191295,10.017825,10.343636,10.096705,9.853205,11.077567,12.188754,12.4974165,12.178465,12.4974165,12.343085,11.821788,11.063849,10.220171,10.055551,9.880642,10.017825,10.587136,11.519984,11.941824,12.874671,13.080446,12.593445,12.7272,12.682614,12.542002,11.698323,10.717461,11.314209,11.616013,12.072148,12.953552,14.061309,14.7095,15.412566,15.738377,15.79325,15.63206,15.247946,14.38026,14.466,14.544881,14.147048,13.293081,12.97413,11.739478,10.645439,10.240748,10.569988,11.55771,12.500846,12.857523,12.7272,12.836946,12.946692,12.435684,11.794352,11.146159,10.240748,11.492548,10.30591,9.030104,8.584257,8.467651,8.196714,9.431366,10.9369545,11.838936,11.64345,11.444533,12.055,12.590015,13.073587,14.445422,15.505165,15.3302555,14.441993,13.1593275,11.578287,10.4533825,10.422516,11.026124,11.742908,11.979549,10.984968,10.127572,9.074688,7.9429245,7.3118806,6.5162163,6.094377,5.9812007,6.0395036,6.0566516,6.8283086,7.3701835,7.805741,8.186425,8.491658,8.796892,9.750318,10.189304,9.860064,9.407358,9.836057,9.962952,10.436234,11.187314,11.458252,11.88352,11.965831,11.612583,10.926665,10.206452,0.91569984,1.039165,1.0871792,1.1660597,1.2415106,1.1454822,1.1694894,1.1934965,1.2415106,1.2655178,1.1454822,1.1797781,1.3821237,1.6770682,1.978872,2.2120838,2.2600982,2.2738166,2.1640697,1.9754424,1.8759843,1.9514352,2.2052248,2.4624438,2.6236343,2.6853669,3.2821152,3.4878905,3.642222,3.8102717,3.799983,3.8960114,3.6936657,3.3815732,3.0557625,2.6990852,2.311542,2.037175,2.0268862,2.2909644,2.7299516,2.9151495,3.069481,2.9117198,2.4315774,1.9068506,1.7971039,1.8416885,2.1057668,2.335549,1.9685832,2.0303159,1.9171394,1.8485477,1.8554068,1.7696671,1.8931323,1.6770682,1.430138,1.2758065,1.1283343,1.1283343,1.2929544,1.3066728,1.0666018,0.6859175,0.61389613,0.548734,0.48700142,0.4664239,0.5658819,0.42869842,0.31552204,0.22978236,0.16804978,0.106317215,0.06859175,0.034295876,0.01371835,0.01371835,0.0,0.01371835,0.006859175,0.0,0.010288762,0.044584636,0.034295876,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.26407823,0.8711152,1.9068506,2.6167753,4.4584637,6.258997,7.2364297,7.0032177,6.5642304,4.057202,2.534465,3.1586502,5.171818,4.098357,4.8837323,4.266407,2.2635276,2.1674993,1.5330256,0.9877212,0.45613512,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.017147938,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.106317215,0.22978236,0.16804978,0.16804978,0.20577525,0.28465575,0.42869842,0.6859175,0.881404,1.1043272,1.371835,1.7010754,2.0920484,2.335549,2.3424082,2.4555845,2.8945718,3.724532,5.127233,5.504488,5.456474,5.470192,5.919468,6.677407,7.4970784,7.881192,7.870903,8.042382,8.309891,8.669997,9.352485,9.877212,9.047252,10.1481495,11.125582,11.952112,12.377381,11.962401,12.939834,12.634601,12.092726,12.175035,13.564018,13.749216,13.529722,12.723769,11.609154,10.926665,11.657167,11.979549,12.332796,13.059869,14.390549,13.718349,13.732068,13.807519,13.975569,14.939283,14.4145565,14.79524,15.302819,15.37827,14.695783,14.205351,13.63604,13.725209,14.188204,13.687484,12.929544,13.063298,13.660047,14.112752,13.625751,12.9809885,12.295071,11.862943,11.760056,11.869802,11.077567,10.367643,9.829198,9.887501,11.290202,12.281353,12.792361,13.622321,14.586036,14.527733,19.641247,22.9508,19.03421,10.600855,8.515666,13.834956,16.019604,16.684942,17.175373,18.554068,18.396307,17.62465,17.141079,17.134218,17.058767,16.715809,16.0539,15.518884,15.422854,15.9613,15.837835,15.395418,15.402277,15.913286,16.266533,16.839275,16.561478,15.87213,15.199932,14.970149,14.503725,13.059869,12.061859,12.010415,12.511135,11.427385,10.401938,9.897789,10.257896,11.732618,12.723769,11.869802,11.05356,10.964391,11.122152,11.269625,12.295071,13.858963,15.254805,15.426285,16.6335,17.652086,18.969048,20.7833,22.978235,23.540688,26.658184,28.67135,28.870268,29.480734,35.094967,35.876915,29.796255,20.19341,15.762384,8.964942,4.5339146,2.153781,1.4472859,1.9823016,1.6290541,1.4953002,1.3855534,1.4541451,2.2120838,3.566771,6.6876955,9.606275,11.297061,11.688034,11.039842,12.024134,13.519434,14.839825,15.731518,14.363112,12.823228,11.204462,9.657719,8.378482,7.606825,7.3701835,7.2775846,7.2192817,7.3530354,6.40304,6.1458206,6.3893213,7.0443726,8.117833,9.019815,9.5033865,9.1981535,8.31332,7.630832,5.051782,3.6319332,3.234101,3.690236,4.7774153,3.590778,3.3061223,3.1586502,3.0557625,3.5564823,3.8479972,3.9303071,4.0229063,4.139512,4.0880685,3.5770597,3.642222,4.2389703,4.822,4.3349986,4.4550343,4.4756117,4.3795834,4.3109913,4.5922174,5.2026844,5.576509,5.861165,6.108095,6.2418494,5.4976287,5.0346346,4.804852,4.880303,5.4770513,6.025785,5.761707,5.5490727,5.785714,6.4098988,6.420188,6.6053853,6.8385973,6.910619,6.5470824,6.48535,6.3138704,6.468202,6.8283086,6.728851,6.800872,7.1061053,7.5862474,8.165848,8.7283,8.875772,8.690575,8.453933,8.285883,8.162418,8.567109,8.628842,8.354475,7.98408,7.9943686,7.798882,7.9909387,7.8846216,7.2364297,6.210983,5.4907694,5.0620713,4.928317,5.0483527,5.3398676,5.206114,5.137522,5.295283,5.56965,5.56965,6.3618846,6.385892,6.0703697,5.802862,5.950334,6.6225333,6.90033,6.9071894,6.7700057,6.6225333,7.099246,7.4181976,7.6376915,7.8331776,8.1041155,8.076678,9.033533,10.820349,12.665466,13.152468,12.809509,13.375391,14.46257,15.086755,13.670336,12.977559,14.4317045,15.542891,15.110763,13.245067,12.977559,13.200482,13.114742,12.710052,12.771784,12.332796,12.185325,11.97269,11.592006,11.214751,10.532263,9.455373,7.9772205,6.5230756,5.950334,6.3790326,6.914048,5.2987127,2.5241764,2.8534167,5.552502,4.5682106,3.1826572,2.7128036,2.5173173,4.5442033,4.9420357,5.038064,5.0449233,4.0434837,4.715683,4.9831905,5.6176643,6.680836,7.5210853,8.512236,10.103564,10.604284,9.849775,9.2153015,10.096705,10.261326,9.575408,8.711152,9.139851,9.349055,10.679735,11.80464,12.367092,13.015285,12.723769,11.650309,10.357354,9.246168,8.573969,8.049242,7.874333,8.2653055,8.958082,9.201583,9.736599,10.456812,10.563129,10.113853,10.041832,9.235879,8.923786,9.22216,9.091836,6.3310184,7.0786686,3.8479972,3.673088,6.7322803,6.3790326,7.5519514,10.360784,11.996697,12.168177,13.107883,13.862392,14.116182,13.725209,13.173045,13.564018,12.528283,13.138749,15.018164,14.908417,6.667118,4.9351764,2.6716487,2.5721905,4.173808,3.8445675,7.0786686,10.864933,12.38424,12.641459,16.448301,6.742569,4.3281393,5.3158607,8.3922,14.79867,4.2286816,3.3644254,3.806842,6.8866115,23.633287,8.669997,3.8479972,1.9754424,0.26407823,0.33609957,0.116605975,0.14404267,0.6379033,1.5364552,2.486451,2.620205,3.0043187,3.1620796,3.1449318,3.525616,4.647091,5.3330083,5.178677,4.602506,4.822,5.0655007,5.346727,5.6210938,5.9160385,6.3310184,7.8331776,9.592556,10.690024,10.960961,10.984968,10.216741,11.132441,11.814929,11.825217,12.1921835,12.120162,11.4033785,10.847785,10.587136,10.086417,9.9869585,9.489669,9.194724,9.407358,10.117283,9.932085,11.122152,11.784062,11.592006,11.8115,12.775213,12.394529,11.965831,12.133881,12.878101,12.377381,12.21619,12.284782,12.500846,12.816368,13.450842,14.023583,14.784951,15.470869,15.275383,15.028452,14.977009,14.836395,14.476289,13.917266,13.588025,11.948683,10.995257,11.108434,11.046701,12.024134,13.073587,13.526293,13.238208,12.603734,13.018714,12.617453,12.442543,12.620882,12.3911,12.339656,11.540562,10.55284,9.554831,8.347616,9.043822,10.744898,12.452832,13.375391,12.922686,12.812939,13.639469,14.057879,14.081886,15.0456,15.789821,15.498305,15.049029,14.692352,14.068168,12.590015,11.756626,11.876661,12.531713,12.542002,11.859513,10.844356,9.97324,9.290752,8.423067,7.373613,6.433906,5.675967,5.2026844,5.1409516,6.2041235,6.9826403,7.4284863,7.720001,8.268735,8.1487,9.417647,10.515115,10.703742,10.055551,9.458802,9.489669,9.942374,10.347065,9.993818,9.860064,9.97324,10.48082,10.912948,10.192734,1.2929544,1.6393428,1.6359133,1.4987297,1.3512574,1.2037852,1.2380811,1.3238207,1.3341095,1.3101025,1.4610043,1.4610043,1.6290541,1.8725548,2.0886188,2.1640697,1.978872,1.8519772,1.7353712,1.6804979,1.8142518,1.937717,2.0028791,2.136633,2.352697,2.551613,2.6887965,2.568761,2.5241764,2.5481834,2.2600982,2.417859,2.6956558,2.668219,2.3664153,2.2841053,2.1194851,2.2258022,2.16064,2.020027,2.4384367,2.8465576,2.9254382,2.9563043,2.9151495,2.469303,2.486451,2.2566686,2.020027,1.8485477,1.6393428,1.9342873,2.1126258,2.253239,2.311542,2.1469216,2.0474637,1.8828435,1.7456601,1.5947582,1.2620882,1.155771,1.0666018,0.922559,0.7339317,0.58988905,0.65162164,0.59331864,0.5453044,0.5521636,0.5521636,0.41840968,0.28808534,0.18862732,0.12003556,0.058302987,0.030866288,0.020577524,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06859175,0.216064,0.52815646,1.1763484,2.0303159,2.8328393,3.7691166,4.5853586,4.5990767,3.806842,2.253239,1.214074,1.0906088,1.3752645,1.1900668,1.670209,1.9651536,1.7422304,1.1660597,1.6942163,1.0528834,0.36353627,0.08916927,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.006859175,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0274367,0.06516216,0.082310095,0.09259886,0.12346515,0.17490897,0.25378948,0.3806842,0.607037,0.7922347,1.0117283,1.2998136,1.6496316,1.7593783,1.9411465,2.218943,2.5584722,2.8808534,3.8925817,4.0949273,4.0263357,4.170378,4.945465,5.8371577,5.9880595,5.8817425,5.9983487,6.831738,7.500508,7.7783046,7.997798,8.210432,8.169277,9.033533,9.956093,10.748327,11.365653,11.876661,12.627741,12.686044,13.032433,13.817808,14.369971,13.858963,13.402828,13.046151,12.689473,12.072148,12.298501,12.953552,13.622321,14.174485,14.743796,13.485138,13.443983,13.934414,14.366542,14.2190695,13.584596,13.917266,14.644339,15.059319,14.315098,13.114742,12.723769,12.874671,13.241637,13.443983,13.673765,13.3033695,13.505715,14.2533655,14.321958,13.725209,13.169616,12.614022,12.394529,13.227919,12.6586075,11.592006,10.521975,10.22703,11.766914,12.415107,13.3033695,14.417986,15.453721,15.830976,20.584383,21.757303,16.475739,8.330468,7.366754,13.039291,14.270514,14.764374,15.9750185,17.103354,16.232237,15.96816,15.673215,15.230798,15.069608,15.29596,14.949572,14.740367,14.946142,15.422854,15.477728,15.54632,15.745236,16.04018,16.266533,16.410576,16.558048,16.53747,16.259674,15.724659,15.193072,13.951562,12.380811,11.4376745,12.672326,10.823778,9.757176,9.160428,9.184435,10.429376,10.947243,11.166737,10.964391,10.580277,10.611144,11.1393,12.147599,13.560589,14.953001,15.573756,17.103354,17.943602,19.257133,21.109112,22.467228,24.209457,26.531288,27.611609,28.637054,33.778008,36.216442,30.890295,24.408375,18.893597,11.941824,5.329579,2.726522,1.937717,1.6942163,1.6667795,1.4472859,1.8245405,2.6819375,4.1155047,6.4236174,6.6568294,9.407358,12.113303,13.924125,15.741806,15.22051,15.590904,16.242527,16.743246,16.842705,15.484588,13.704632,12.205902,11.129011,10.062409,8.491658,7.870903,7.798882,7.7680154,7.160979,6.8900414,6.557371,6.4064693,6.7631464,8.032094,8.505377,8.471081,8.375052,8.172707,7.3255987,5.9880595,5.0586414,4.32128,3.923448,4.386442,4.0023284,3.8925817,3.7862647,3.5633414,3.275256,3.6147852,3.673088,3.5839188,3.5359046,3.758828,3.82399,4.184097,4.383013,4.338428,4.3590055,4.996909,5.051782,5.051782,5.1992545,5.3741636,5.6828265,5.919468,6.1149545,6.2864337,6.447624,6.2898636,6.142391,6.142391,6.351596,6.783724,6.776865,6.6122446,6.492209,6.526505,6.7391396,6.8763227,6.9346256,6.9963584,7.023795,6.8626046,6.989499,6.9380555,6.824879,6.759717,6.8385973,6.5230756,6.6396813,7.0135064,7.490219,7.936065,7.8091707,7.7028537,7.4044795,7.058091,7.15069,7.671987,8.107545,8.608265,9.098696,9.277034,9.335337,9.3764925,9.054111,8.2653055,7.160979,6.3447366,5.950334,5.689686,5.5079174,5.5833683,5.6348124,5.874883,6.077229,6.2041235,6.39961,6.6053853,6.615674,6.5127864,6.39961,6.3893213,6.584808,6.7357097,6.90033,7.133542,7.466212,7.658269,7.5553813,7.466212,7.6033955,8.076678,8.522525,9.424506,10.6488695,12.082437,13.666906,14.369971,14.057879,13.978998,14.496866,15.110763,15.217079,16.602633,17.494326,17.161655,15.916716,14.486577,13.073587,12.442543,12.445972,12.037852,12.185325,12.017275,11.64345,11.369082,11.701753,10.686595,10.340206,9.537683,8.056101,6.584808,7.3255987,7.6033955,6.9346256,5.6793966,5.051782,5.2472687,4.7602673,4.664239,4.9351764,4.4447455,5.3981705,6.2967224,6.81802,6.6431108,5.446185,5.7377,5.8165803,6.125243,6.852316,7.949784,8.097256,8.625413,9.345626,9.80862,9.290752,9.006097,8.632272,8.632272,8.803751,8.272165,8.999237,10.813489,12.010415,12.421966,13.430264,13.63604,12.243628,10.772334,9.719451,8.539673,8.872343,8.450503,8.2653055,8.721441,9.626852,10.254466,10.847785,11.074138,11.094715,11.578287,10.587136,10.456812,9.47595,7.4044795,5.4667625,3.2032347,3.0729103,3.5016088,4.636802,8.344186,8.371623,10.347065,11.914387,12.483699,13.227919,13.38911,13.320518,12.956982,12.641459,13.101024,11.790922,12.257345,14.363112,15.21022,9.156999,6.701414,4.712253,4.184097,4.770556,4.773986,5.7136927,7.936065,9.160428,9.575408,11.821788,5.1238036,3.1380725,2.8980014,5.003768,13.629181,4.5990767,4.938606,4.479041,4.2698364,16.606062,7.3701835,3.8788633,2.0028791,0.30866286,0.07888051,0.034295876,0.048014224,0.53844523,1.471293,2.3664153,2.3149714,3.8788633,4.40359,3.666229,3.8788633,5.0414934,5.425607,5.6210938,5.7308407,5.394741,6.2727156,6.5882373,7.1026754,7.881192,8.285883,7.9120584,8.694004,9.290752,9.3593445,9.55826,9.510246,10.045261,10.367643,10.374502,10.64201,10.978109,10.542552,10.254466,10.209882,9.657719,9.208443,8.834618,8.64256,8.604835,8.543102,8.906639,9.513676,9.740028,9.853205,11.029553,11.55428,11.657167,11.574858,11.664027,12.3911,12.895248,12.686044,12.542002,12.528283,11.986408,11.900668,12.905538,14.30138,15.54632,16.239098,16.365992,15.937293,15.450292,15.110763,14.843254,14.112752,12.63117,11.677745,11.526843,11.427385,12.130451,12.950122,13.646329,14.033872,13.996146,13.581166,12.775213,12.788932,13.738928,14.661487,14.318527,14.88098,14.942713,13.828096,11.592006,10.549411,10.779194,11.399949,11.660598,10.933525,11.478829,12.445972,13.231348,13.88297,15.083325,15.4742985,15.21365,14.894698,14.740367,14.606613,13.958421,12.809509,12.161317,12.048141,11.55428,11.993267,11.47197,10.9369545,10.525404,9.568549,8.2653055,7.349606,6.5162163,5.7719955,5.446185,5.9640527,6.5470824,7.1952744,7.7371492,7.8194594,7.932636,9.177576,10.539123,11.269625,10.88551,10.209882,9.623423,9.421077,9.510246,9.421077,9.530824,9.56512,9.846346,10.209882,9.997248,1.3341095,1.471293,1.3649758,1.1832076,1.0528834,1.0460242,1.155771,1.1866373,1.2175035,1.2620882,1.2758065,1.4987297,1.6976458,1.7971039,1.8039631,1.8039631,1.6324836,1.5398848,1.4610043,1.4198492,1.5364552,1.5741806,1.6256244,1.7971039,2.0131679,2.0337453,1.9171394,1.7010754,1.5501735,1.5124481,1.5090185,1.8416885,2.1503513,2.2841053,2.277246,2.3389788,2.5721905,2.6716487,2.4658735,2.153781,2.318401,2.527606,2.4967396,2.527606,2.585909,2.287535,2.3972816,2.2600982,2.1503513,2.1434922,2.1434922,2.218943,2.2635276,2.2155135,2.1229146,2.1503513,2.0817597,1.9480057,1.786815,1.5570327,1.1420527,1.0014396,0.90198153,0.7990939,0.6893471,0.61046654,0.58988905,0.5590228,0.5178677,0.4698535,0.39440256,0.3018037,0.22292319,0.15433143,0.08916927,0.037725464,0.01371835,0.006859175,0.006859175,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.11317638,0.34638834,1.0288762,1.6942163,2.1743584,2.6373527,3.059192,3.2203827,2.4590142,1.4438564,0.65848076,0.28122616,0.18176813,0.216064,0.65848076,1.1729189,1.3889829,0.90541106,1.2346514,0.89512235,0.41498008,0.09602845,0.030866288,0.034295876,0.020577524,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0274367,0.116605975,0.06859175,0.07888051,0.10288762,0.14747226,0.26064864,0.39783216,0.5453044,0.69963586,0.8711152,1.0666018,1.1832076,1.4369972,1.7353712,2.037175,2.386993,2.7951138,3.0900583,3.3026927,3.5290456,3.9303071,4.681387,4.870014,4.9248877,5.161529,5.778855,6.279575,6.708273,7.1369715,7.548522,7.829748,8.255017,9.084977,9.640571,10.05898,11.290202,11.982979,11.982979,11.945253,12.253916,12.9981365,13.039291,12.367092,12.05157,12.092726,11.406808,11.880091,12.9638405,13.759505,14.044161,14.291091,13.481709,13.488567,13.845244,13.951562,13.077017,12.96727,14.040731,15.162207,15.587475,14.953001,13.690913,13.035862,12.881531,13.169616,13.876111,14.688923,14.483148,14.428274,14.802099,14.973578,14.490007,14.147048,13.814379,13.9138365,15.422854,15.46744,14.270514,13.029003,12.476839,12.895248,12.847235,13.29994,14.335675,15.584045,16.194511,19.161106,18.056778,13.262215,8.042382,8.543102,12.620882,13.094165,13.642899,15.199932,15.923574,14.802099,14.863832,14.956431,14.784951,14.911846,15.261664,14.778092,14.531162,14.819247,15.189643,15.433144,15.680074,15.940722,16.256245,16.678083,16.671225,16.729528,16.750105,16.510035,15.649208,15.151917,14.270514,13.227919,12.445972,12.528283,11.2593355,10.768905,10.189304,9.575408,9.918367,10.278474,10.597425,11.029553,11.406808,11.2593355,11.72233,12.535142,13.807519,15.268523,16.276823,17.734396,18.766703,20.169403,21.897917,23.087982,25.35494,27.141756,28.3524,30.334702,35.876915,30.389574,26.719915,21.808746,15.278812,9.458802,3.4981792,1.7559488,1.6633499,1.7902447,1.8519772,2.153781,2.6613598,3.9680326,6.135532,8.694004,10.124143,11.540562,13.13189,15.12448,17.778982,18.564358,18.69811,18.523201,18.423744,18.821575,17.96761,16.221949,14.589465,13.402828,12.332796,10.861504,9.791472,9.040393,8.340756,7.2467184,6.9963584,6.948344,7.016936,7.2364297,7.764586,8.004657,7.781734,7.4010496,6.9346256,6.2144127,6.0737996,6.094377,5.6793966,4.9077396,4.5167665,4.3178506,4.1360826,4.07435,4.046913,3.7622573,4.064061,4.098357,4.0674906,4.064061,4.081209,4.1772375,4.417309,4.540774,4.5647807,4.7842746,5.113515,5.377593,5.6210938,5.8543057,6.046363,6.2555676,6.416758,6.5230756,6.5882373,6.6293926,6.8591747,7.0889573,7.3050213,7.5725293,8.045813,7.963502,7.8434668,7.7268605,7.6514096,7.6445503,7.81603,7.6857057,7.6033955,7.613684,7.473071,7.623973,7.7542973,7.5931067,7.2604365,7.2775846,6.7665763,6.64997,6.9963584,7.4936485,7.4353456,7.3118806,7.1849856,6.9346256,6.6636887,6.6876955,7.1129646,7.781734,8.532814,9.259886,9.918367,10.134431,10.206452,9.908078,9.163857,8.042382,7.1781263,6.324159,5.8474464,5.7719955,5.8200097,6.262427,6.7700057,6.9654922,6.917478,7.1369715,6.9792104,6.8214493,6.8385973,6.992929,7.0306544,6.9860697,6.8626046,6.883182,7.1129646,7.4456344,7.349606,7.3427467,7.3084507,7.3564653,7.8537555,8.347616,9.513676,11.228469,13.090735,14.424845,14.627191,14.651197,14.730078,14.853543,14.778092,15.244516,16.88729,18.084215,18.04649,16.815268,15.182784,13.107883,12.109874,12.212761,11.928105,11.650309,11.30049,10.978109,10.844356,11.1393,10.244178,9.993818,9.400499,8.162418,6.6705475,7.2707253,7.5382333,8.083538,8.618553,7.970361,7.373613,5.6142344,4.787704,5.3878818,6.2830043,6.924337,7.720001,8.327039,8.416207,7.675417,7.438775,7.5759587,8.200144,9.1810055,10.14472,9.81205,9.788043,9.880642,9.801761,9.1981535,8.477941,8.152129,8.093826,8.069819,7.7268605,8.484799,9.932085,11.166737,12.017275,13.011855,12.764925,11.413667,10.189304,9.263316,7.750868,7.764586,8.014946,8.189855,8.381912,9.067829,9.911508,10.573419,10.923236,11.235329,12.202472,11.235329,11.691463,10.199594,6.56766,3.7553983,2.5653315,5.645101,6.0703697,4.5819287,9.585697,10.508256,10.823778,11.928105,13.742357,14.723219,13.690913,13.416546,12.96727,12.312219,12.325937,11.845795,11.47197,13.05301,15.306249,13.828096,11.183885,8.186425,6.8385973,6.910619,5.9469047,5.579939,5.895461,6.948344,8.491658,9.952662,5.785714,3.0454736,1.5227368,2.9665933,11.084427,3.9268777,3.292404,2.7745364,2.3321195,8.282454,4.9934793,3.549623,3.4295874,3.234101,0.7099246,0.9602845,1.1900668,2.5070283,4.705394,6.279575,4.3658648,5.2747054,5.6965446,5.15467,5.9983487,6.5059276,6.715132,6.7940125,6.5539417,5.446185,6.9380555,7.449064,7.9463544,8.611694,8.800322,8.368194,8.879202,9.078118,8.827758,9.098696,8.64256,8.820899,9.047252,9.2153015,9.685155,10.117283,10.240748,10.484249,10.549411,9.386781,8.80718,8.351046,8.038953,7.9086285,8.011517,8.224151,8.755736,9.266746,9.791472,10.72432,11.108434,11.012405,10.693454,10.63858,11.5645685,12.9707,13.371962,13.570878,13.536582,12.428825,12.46998,13.197053,14.517444,16.249386,18.156237,18.571217,17.62808,16.259674,15.241087,15.175924,14.726648,13.978998,13.214201,12.511135,11.712041,11.46854,11.797781,12.507706,13.344524,13.996146,14.325387,14.270514,14.342535,14.71636,15.227368,15.237658,16.907866,18.04306,17.566347,15.498305,14.167625,13.2862215,12.778643,12.21962,10.813489,10.957532,12.188754,13.145609,13.536582,14.147048,14.232788,14.5414505,14.688923,14.514014,14.061309,13.762935,13.049581,12.490558,12.061859,11.132441,11.201033,10.871792,10.302481,9.578837,8.7145815,8.056101,7.8194594,7.2775846,6.324159,5.442755,5.627953,6.3138704,7.0923867,7.582818,7.421627,7.548522,8.378482,9.534253,10.4533825,10.415657,9.801761,9.115844,8.536243,8.330468,8.882631,9.801761,10.1481495,9.993818,9.695444,9.866923,1.0597426,1.0425946,0.94656616,0.8848336,0.89512235,0.9431366,1.0494537,1.0425946,1.08032,1.1694894,1.1592005,1.3924125,1.5501735,1.5913286,1.5501735,1.5090185,1.4472859,1.4061309,1.3272504,1.2346514,1.2483698,1.1934965,1.2860953,1.4541451,1.5707511,1.4541451,1.2929544,1.1008976,1.0048691,1.0940384,1.4267083,1.7902447,1.937717,2.1572106,2.4384367,2.435007,2.6407824,2.5996273,2.3595562,2.1091962,2.177788,2.136633,2.07833,2.0817597,2.0749004,1.8485477,1.9582944,1.9480057,2.0063086,2.177788,2.3732746,2.2052248,2.1469216,2.0303159,1.9068506,2.0474637,1.9342873,1.8108221,1.6496316,1.4027013,1.0117283,0.8779744,0.805953,0.7407909,0.64819205,0.53844523,0.4938606,0.4938606,0.44584638,0.33952916,0.26407823,0.20920484,0.16119061,0.1097468,0.058302987,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.05144381,0.20577525,0.7339317,1.2106444,1.6667795,1.9514352,2.0886188,2.3046827,2.6407824,2.0508933,1.0254467,0.13375391,0.01371835,0.048014224,0.5041494,0.97400284,1.1866373,1.0357354,1.1900668,1.0666018,0.6241849,0.09945804,0.024007112,0.034295876,0.020577524,0.030866288,0.05144381,0.0,0.0,0.0,0.0034295875,0.017147938,0.0548734,0.010288762,0.0,0.0,0.010288762,0.0548734,0.010288762,0.0,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.034295876,0.14061308,0.07888051,0.08916927,0.09602845,0.09602845,0.17490897,0.23664154,0.35324752,0.4629943,0.548734,0.6241849,0.7339317,0.9431366,1.1832076,1.4507155,1.8176813,1.9548649,2.3218307,2.7745364,3.1586502,3.3198407,3.8685746,4.1463714,4.3761535,4.6676683,5.0277753,5.2335505,5.813151,6.4064693,6.924337,7.5690994,7.596536,8.107545,8.371623,8.56025,9.72631,10.30591,10.261326,9.935514,9.80519,10.501397,11.4205265,10.978109,10.611144,10.666017,10.419086,11.228469,11.821788,12.229909,12.603734,13.210771,12.596875,12.634601,12.984418,13.162757,12.535142,13.13189,14.291091,15.021593,15.069608,14.911846,13.937843,13.063298,12.55229,12.634601,13.533153,14.973578,15.265094,15.162207,15.254805,15.995596,15.769243,15.429714,15.172495,15.46401,17.058767,16.859852,15.4742985,14.30138,13.862392,13.821238,13.358243,13.612033,14.678635,16.023033,16.46888,17.089634,15.0078745,11.88352,9.767465,11.063849,12.795791,12.809509,13.279363,14.3974085,14.3974085,13.7526455,14.037301,14.503725,14.942713,15.673215,15.841265,15.374841,15.097044,15.217079,15.340545,15.419425,15.638919,16.002455,16.46545,16.938732,16.835844,16.80155,16.86671,16.832415,16.266533,15.54632,14.586036,13.80066,13.193623,12.363663,11.780633,11.605724,11.231899,10.799771,11.194174,10.88894,11.029553,11.701753,12.439114,12.195613,12.984418,13.371962,14.153908,15.498305,16.96617,18.53692,19.853882,21.325174,22.86163,23.883648,26.35981,27.84825,30.218096,32.454185,30.663942,22.810186,22.957659,20.20027,12.425395,6.307011,2.534465,1.4815818,1.5398848,1.8382589,2.2120838,3.4295874,4.57507,6.279575,8.47451,10.408798,11.948683,12.4974165,13.433694,15.385129,18.231688,19.963629,20.484926,20.087093,19.490345,19.843594,19.795578,18.53692,16.681513,14.79867,13.423406,12.795791,11.8869505,10.823778,9.668007,8.405919,7.798882,7.5416627,7.466212,7.4627824,7.507367,7.56224,7.143831,6.6431108,6.327589,6.3173003,6.711703,6.759717,6.186976,5.2335505,4.650521,4.232111,4.046913,4.1360826,4.3109913,4.1360826,4.180667,4.3178506,4.4996185,4.7259717,5.038064,4.722542,4.5339146,4.629943,4.9523244,5.2301207,5.4907694,5.936616,6.3035817,6.5127864,6.6739774,6.7219915,6.842027,6.9826403,7.130112,7.3290286,7.6685576,7.9429245,8.193284,8.519095,9.071259,9.0369625,8.831187,8.632272,8.512236,8.4264965,8.591117,8.333898,8.220721,8.351046,8.327039,8.378482,8.419638,8.117833,7.6514096,7.682276,7.250148,7.016936,7.1952744,7.459353,6.9654922,6.989499,6.7871537,6.6053853,6.5470824,6.5950966,6.9792104,7.7714453,8.64599,9.482809,10.371073,10.714031,10.566559,10.065839,9.304471,8.357904,7.641121,6.660259,6.121814,6.1492505,6.2898636,7.0546613,7.723431,8.028665,8.001227,7.949784,7.5862474,7.274155,7.274155,7.5210853,7.6171136,7.500508,7.3427467,7.281014,7.332458,7.3839016,7.1541195,7.2021337,7.1884155,7.164408,7.5725293,8.124693,9.314759,11.118723,13.145609,14.627191,14.21564,14.514014,15.073037,15.343974,14.654627,14.500296,15.776102,17.192522,17.686382,16.431154,15.241087,13.4474125,12.171606,11.80464,11.982979,11.519984,11.05699,10.542552,10.172156,10.412228,9.791472,9.517105,9.084977,8.258447,7.06838,7.1884155,7.3084507,8.042382,9.040393,8.985519,8.553391,6.125243,4.835718,5.6656785,7.407909,8.217292,8.786603,9.263316,9.599416,9.547972,8.8929205,9.006097,9.750318,10.765475,11.46854,11.149589,10.912948,10.569988,9.997248,9.112414,8.285883,8.131552,7.888051,7.548522,7.891481,8.676856,9.290752,10.045261,10.8958,11.46854,11.4376745,10.161868,8.961512,8.114404,6.8728933,6.4579134,7.281014,7.9943686,8.241299,8.64599,9.3593445,10.079557,10.618003,11.231899,12.651748,12.082437,12.435684,11.2593355,7.7714453,2.8534167,4.389872,6.8454566,6.783724,5.5250654,9.177576,11.657167,11.605724,12.367092,14.21564,14.352823,13.162757,13.557159,13.066729,11.540562,11.159878,11.701753,11.180455,12.264205,15.014734,16.87357,14.459141,10.693454,9.119273,9.098696,5.802862,4.3761535,3.6936657,4.636802,6.6396813,7.716572,7.486789,4.338428,1.5741806,1.7319417,6.56766,3.9954693,2.2086544,1.2758065,1.3958421,2.8877127,2.6990852,2.603057,3.7005248,4.746549,2.1572106,1.4850113,3.4981792,4.8768735,5.3158607,7.5245147,6.2658563,7.2467184,7.2775846,6.3310184,7.5245147,7.723431,7.6033955,7.5931067,7.4524937,6.2830043,8.069819,8.279024,8.543102,9.2153015,9.379922,9.640571,10.041832,9.846346,9.218731,9.205012,8.594546,8.748878,8.940934,9.078118,9.709162,9.966381,10.463672,10.991828,11.029553,9.760606,9.119273,8.484799,8.049242,7.905199,8.042382,7.7783046,8.440215,9.47938,10.542552,11.4754,11.578287,10.861504,10.117283,10.021255,11.159878,13.262215,14.359683,14.96329,14.826107,12.953552,13.512574,14.335675,15.402277,16.87014,19.082224,19.901896,19.010202,17.192522,15.488017,15.21365,15.29253,15.22051,14.644339,13.536582,12.202472,11.170166,10.923236,11.345076,12.195613,13.118172,14.164196,14.836395,15.241087,15.29596,14.7095,15.306249,17.055338,18.660385,19.13024,17.782412,16.753534,15.618341,14.760944,13.910407,12.130451,11.413667,12.487128,13.618892,13.920695,13.317088,12.926115,13.673765,14.527733,14.71636,13.725209,12.905538,12.490558,12.343085,12.103014,11.204462,10.576848,10.254466,9.654288,8.694004,7.8263187,7.795452,8.080108,7.675417,6.478491,5.295283,5.336438,5.9880595,6.725421,7.2192817,7.3290286,7.5450926,8.272165,9.15014,9.801761,9.836057,9.366203,8.930646,8.357904,8.035523,8.882631,10.017825,10.4705305,10.405369,10.024684,9.592556,0.6790583,0.6790583,0.6824879,0.7956643,0.9568549,0.94999576,0.97057325,0.9911508,0.9911508,1.0151579,1.1660597,1.1866373,1.255229,1.3478279,1.4095604,1.3684053,1.3821237,1.3272504,1.214074,1.0871792,1.0254467,0.9534253,1.0528834,1.138623,1.1317638,1.039165,0.97400284,0.84024894,0.90884066,1.2346514,1.6873571,1.9651536,1.9480057,2.1743584,2.534465,2.2635276,2.1263442,2.0165975,1.8725548,1.7765263,1.9274281,1.8108221,1.8691251,1.8965619,1.7799559,1.4953002,1.5330256,1.5227368,1.5741806,1.7456601,2.054323,1.8313997,1.8313997,1.8313997,1.7936742,1.845118,1.5947582,1.5193073,1.4404267,1.2655178,0.9842916,0.85739684,0.7682276,0.66533995,0.52815646,0.37382504,0.39440256,0.41498008,0.35324752,0.24350071,0.2194936,0.16804978,0.1097468,0.058302987,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.041155048,0.07888051,0.22635277,0.607037,1.0940384,1.3581166,1.4404267,1.7559488,3.350707,2.9974594,1.6084765,0.22635277,0.01371835,0.041155048,0.4698535,0.8711152,1.0666018,1.1283343,1.5638919,1.3478279,0.72707254,0.09602845,0.01371835,0.0034295875,0.0,0.044584636,0.08916927,0.0,0.0,0.0,0.0034295875,0.030866288,0.11317638,0.07545093,0.058302987,0.041155048,0.05144381,0.15090185,0.05144381,0.010288762,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0034295875,0.006859175,0.0,0.0034295875,0.0,0.006859175,0.034295876,0.10288762,0.08573969,0.1097468,0.11317638,0.09259886,0.08916927,0.12689474,0.20920484,0.29151493,0.36010668,0.42526886,0.4698535,0.5761707,0.72707254,0.91912943,1.1454822,1.3409687,1.6427724,2.1332035,2.6990852,3.0351849,3.5187566,3.7519686,3.9268777,4.1463714,4.4447455,4.6093655,5.1855364,5.610805,5.9743414,7.023795,6.910619,7.040943,7.140401,7.2604365,7.7577267,8.035523,8.008087,7.8949103,7.905199,8.22758,9.554831,9.692014,9.3079,9.050681,9.544542,10.316199,9.884071,9.644,10.216741,11.417097,10.89237,11.129011,11.705182,12.277924,12.590015,13.629181,14.126471,13.88983,13.402828,13.824667,13.320518,12.38767,11.780633,11.893809,12.754636,14.664916,15.340545,15.333686,15.553179,17.264544,17.511473,16.79469,16.235666,16.441442,17.501184,16.386568,14.932424,13.9481325,13.759505,14.212211,13.88297,14.30138,15.3817,16.571766,16.856422,15.642348,13.951562,12.764925,12.624311,13.642899,13.296511,13.317088,13.642899,13.80409,12.950122,12.96727,13.317088,14.105893,15.22051,16.338554,16.362562,16.204802,16.064188,15.947581,15.697222,15.398848,15.5085945,15.933864,16.448301,16.684942,16.575195,16.722668,17.051908,17.408587,17.556059,16.492886,15.097044,13.937843,13.1421795,12.415107,12.243628,12.020704,11.931535,12.281353,13.491997,12.247057,12.425395,12.946692,13.275933,13.430264,14.733508,14.712931,14.96329,16.067617,17.610931,19.442331,20.855322,22.347193,23.839062,24.672453,27.038868,28.544456,31.895163,32.924038,20.580954,17.29884,20.100813,18.598652,10.80663,3.1415021,2.0920484,1.8862731,2.1126258,2.5550427,3.1826572,5.1409516,7.226141,9.523964,11.561139,12.308789,12.38767,12.857523,13.790371,15.357693,17.830425,19.322296,20.433481,20.70099,20.220848,19.641247,20.145397,19.500635,17.679523,15.306249,13.653188,13.533153,13.145609,12.466551,11.492548,10.251037,9.355915,8.512236,7.764586,7.2432885,7.174697,6.9826403,6.5230756,6.3653145,6.7528577,7.599966,7.9737906,7.1781263,5.9571934,4.9660425,4.7534084,4.033195,4.033195,4.331569,4.530485,4.262977,4.091498,4.3933015,4.756838,5.1580997,5.9571934,5.360445,4.9077396,4.996909,5.5113473,5.8200097,6.3653145,6.8214493,7.0718093,7.1232533,7.130112,6.9723516,7.0203657,7.2124224,7.56224,8.131552,8.361334,8.519095,8.786603,9.22216,9.753747,9.753747,9.451943,9.15014,8.988949,8.951223,8.995808,8.7283,8.656279,8.868914,9.043822,9.019815,8.793462,8.309891,7.8023114,7.798882,7.579388,7.449064,7.3839016,7.2158523,6.6225333,6.7459984,6.4887795,6.3653145,6.5230756,6.756287,7.208993,8.032094,8.968371,9.860064,10.645439,11.019264,10.518545,9.654288,8.766026,8.032094,7.6205435,7.0375133,6.6293926,6.56766,6.8283086,7.682276,8.399059,8.964942,9.249598,9.012956,8.40249,7.8949103,7.7542973,7.963502,8.217292,8.1487,8.217292,8.220721,8.073249,7.7885933,7.425057,7.2878733,7.1884155,7.1541195,7.4456344,8.405919,9.386781,10.504827,11.921246,13.841815,13.622321,13.951562,14.812388,15.683503,15.525743,14.273943,14.428274,15.398848,16.173935,15.306249,14.901558,13.9481325,12.665466,11.7086115,12.144169,11.907528,11.47197,10.6488695,9.80862,9.880642,9.506817,9.287323,9.112414,8.776315,8.014946,7.5759587,7.39762,7.407909,7.613684,8.083538,8.258447,6.574519,5.6965446,6.4064693,7.610255,8.838047,9.4862385,9.884071,10.240748,10.628291,9.757176,9.602845,9.997248,10.645439,11.14273,11.266195,11.118723,10.902658,10.487679,9.427936,8.639131,8.553391,8.162418,7.6342616,8.323608,9.1981535,9.129561,9.208443,9.606275,9.592556,10.508256,9.47595,8.052671,6.975781,6.1629686,5.8405876,6.7940125,7.7714453,8.333898,8.858624,9.146709,9.798331,10.5597,11.499407,13.008426,13.186764,12.737488,12.325937,10.521975,3.8137012,6.9552035,6.23499,5.809721,6.7974424,7.274155,11.255906,12.483699,12.984418,13.272504,12.343085,11.921246,13.022143,12.418536,10.261326,10.103564,11.094715,11.279913,12.037852,13.87954,16.47231,14.589465,11.509696,10.72432,10.782623,5.288424,2.6167753,1.6667795,2.527606,4.2835546,5.0277753,8.865483,6.1972647,2.585909,0.9774324,1.6976458,5.0312047,2.719663,0.805953,1.1008976,1.1900668,1.2929544,1.4987297,2.6133456,3.998899,3.5599117,1.3203912,5.0449233,5.593657,2.8156912,5.5662203,6.8626046,8.772884,8.690575,7.164408,7.9257765,8.31675,7.932636,8.155559,8.824328,8.203573,9.901219,9.547972,9.506817,10.371073,10.971251,11.581717,11.7257595,11.2593355,10.408798,9.774324,9.592556,9.918367,9.9869585,9.818909,10.216741,10.192734,10.676306,11.159878,11.2250395,10.539123,9.904649,9.321619,9.050681,9.006097,8.748878,8.128122,8.7283,9.914937,11.334786,12.898679,12.936404,11.862943,10.765475,10.487679,11.650309,13.790371,15.275383,16.173935,16.005884,13.745787,14.387119,15.470869,16.324837,17.089634,18.739265,19.723558,19.53836,18.169954,16.338554,15.498305,15.830976,16.04018,15.553179,14.335675,12.905538,11.602294,10.854645,10.741467,11.122152,11.640019,13.015285,14.027013,14.987297,15.604623,14.990726,15.282242,16.091625,17.436022,18.608942,18.169954,17.549198,16.842705,16.300829,15.6526375,14.112752,12.346515,12.614022,13.797231,14.520873,13.162757,12.061859,12.521424,13.88983,14.922135,13.7697935,12.027563,11.543991,11.681175,11.88352,11.646879,10.679735,10.271614,9.72631,8.858624,7.9943686,7.98408,8.025234,7.4010496,6.166398,5.113515,5.206114,5.6142344,6.2247014,6.910619,7.548522,7.9943686,8.964942,9.630281,9.709162,9.47595,9.434795,9.445084,9.235879,8.97523,9.266746,10.086417,10.511685,10.909517,10.899229,9.373062,0.59674823,0.53501564,0.51100856,0.6310441,0.84024894,0.90198153,0.91227025,0.9877212,0.89169276,0.70306545,0.823101,0.8711152,0.9945804,1.0940384,1.1351935,1.1592005,1.1351935,0.9911508,0.88826317,0.85396725,0.7922347,0.82996017,0.8676856,0.90884066,0.9431366,0.9294182,0.9294182,0.84024894,1.0048691,1.430138,1.786815,2.1400626,2.0989075,2.1846473,2.277246,1.6187652,1.6667795,1.7319417,1.6530612,1.5021594,1.587899,1.6359133,1.9685832,2.085189,1.8382589,1.4335675,1.4335675,1.2963841,1.3032433,1.5055889,1.7250825,1.6393428,1.6736387,1.605047,1.4198492,1.2963841,1.1146159,1.2312219,1.2758065,1.1454822,1.0220171,0.864256,0.72364295,0.5761707,0.4355576,0.34981793,0.3018037,0.29151493,0.26064864,0.20920484,0.18176813,0.12346515,0.061732575,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.041155048,0.09259886,0.33609957,0.8265306,1.0700313,1.1934965,1.937717,2.452155,1.7079345,0.84367853,0.33266997,0.01371835,0.041155048,0.4115505,0.78537554,0.922559,0.70306545,1.313532,0.7613684,0.18519773,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.26064864,0.29151493,0.21263443,0.14061308,0.21263443,0.15090185,0.0548734,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.017147938,0.037725464,0.0,0.01371835,0.006859175,0.006859175,0.017147938,0.030866288,0.030866288,0.030866288,0.07888051,0.1371835,0.07545093,0.07545093,0.10288762,0.15090185,0.22978236,0.34981793,0.38754338,0.45956472,0.5144381,0.5693115,0.71678376,0.764798,0.91569984,1.2689474,1.8279701,2.486451,3.2306714,3.5461934,3.5873485,3.5393343,3.6010668,4.2835546,4.6402316,4.729401,4.938606,5.950334,6.108095,6.3138704,6.5813785,6.8557453,6.989499,6.7700057,6.4407654,6.5127864,7.0786686,7.8126,8.399059,8.848335,8.464222,7.7028537,8.179566,8.275595,8.052671,7.716572,7.682276,8.56025,9.599416,10.707172,11.238758,11.396519,12.236768,12.9809885,13.334236,12.929544,12.260776,12.665466,12.775213,11.667457,11.567999,12.778643,13.656617,15.059319,15.412566,15.470869,16.067617,18.080786,19.13024,17.580065,16.365992,16.46545,16.890718,15.803539,15.038741,14.239647,13.673765,14.2362175,14.493437,14.647768,15.021593,15.769243,16.890718,15.608052,14.438563,14.260224,14.815818,14.695783,13.38911,14.085316,14.726648,14.342535,13.059869,12.562579,12.617453,13.821238,15.5085945,15.776102,16.276823,16.365992,16.45859,16.46888,15.806969,15.587475,15.608052,15.758954,15.87899,15.731518,16.026463,16.674654,17.29884,17.71382,17.960749,17.031332,15.62863,14.143619,13.049581,12.878101,13.293081,13.334236,13.3033695,13.516005,14.29795,13.101024,13.862392,14.2190695,14.126471,15.885849,16.63007,16.743246,17.408587,18.526632,18.722118,20.310017,21.345753,22.847912,24.7822,26.078583,27.652763,29.683079,31.449318,29.089762,15.6252,16.307688,19.572655,16.822126,8.327039,3.2512488,2.3972816,3.0866287,4.2526884,5.271276,5.967482,7.3084507,9.355915,12.493987,15.285671,14.479718,14.003006,14.38026,14.990726,15.854982,17.62465,17.562918,18.3723,20.172834,21.544668,19.5315,19.37374,18.663815,17.686382,16.595774,15.412566,13.495427,12.80608,12.775213,12.593445,11.214751,10.703742,9.997248,8.7145815,7.174697,6.392751,5.8200097,6.142391,6.7219915,7.2947326,7.963502,8.625413,7.5519514,6.3378778,5.658819,5.2781353,4.5956473,4.8905916,5.2644167,5.24041,4.7774153,5.0826488,5.3501563,5.562791,5.6519604,5.4941993,5.8337283,6.0840883,6.4098988,6.8214493,7.1884155,7.517656,7.7097125,7.630832,7.3358874,7.0786686,6.9826403,6.800872,6.7974424,7.0786686,7.630832,7.764586,8.375052,9.126132,9.753747,10.069269,10.168727,10.082987,9.791472,9.499957,9.657719,9.242738,9.112414,8.947794,8.762596,8.89635,9.078118,8.97866,8.628842,8.100685,7.4936485,7.284444,7.4696417,7.466212,7.14726,6.866034,6.8043017,6.5985265,6.5539417,6.7700057,7.1095347,7.56224,8.344186,9.019815,9.55826,10.316199,10.436234,10.093276,9.328478,8.323608,7.3839016,7.239859,7.130112,6.8557453,6.5813785,6.852316,7.5210853,8.220721,9.0644,9.938945,10.511685,9.266746,8.251588,7.915488,8.340756,9.23245,9.328478,9.517105,9.517105,9.253027,8.848335,7.874333,7.500508,7.4353456,7.5210853,7.750868,9.716022,10.840926,11.204462,11.303921,12.024134,13.22106,14.222499,15.189643,16.13621,16.96617,15.6869335,14.651197,13.992717,13.783512,14.037301,14.441993,14.167625,13.629181,13.107883,12.740917,12.240198,11.8869505,11.362224,10.515115,9.369633,9.15014,8.958082,8.992378,9.174147,9.126132,8.453933,8.193284,8.076678,7.9737906,7.888051,8.81747,8.536243,7.8503256,7.2947326,7.1095347,8.80718,10.230459,11.005547,11.177026,11.214751,10.275044,9.626852,9.489669,9.798331,10.237319,10.957532,11.348505,11.478829,11.317638,10.7586155,10.196163,10.055551,9.31133,8.1041155,7.750868,8.447074,8.656279,9.023245,9.482809,9.263316,10.323058,10.323058,9.047252,7.016936,5.4770513,5.977771,6.944915,7.750868,8.405919,9.568549,9.736599,10.1481495,11.050131,12.168177,12.679185,13.7526455,12.88839,12.874671,12.614022,7.1095347,7.5759587,7.6342616,8.1041155,8.114404,5.113515,10.4705305,13.193623,12.919256,11.379372,12.404818,11.794352,11.249047,10.052121,8.968371,10.237319,10.494537,11.173596,11.245617,11.149589,12.771784,11.622872,11.612583,12.47341,12.367092,7.888051,3.6525106,1.5227368,2.3595562,4.7088237,4.804852,8.433355,6.6739774,3.2203827,0.6241849,0.30523327,5.6999745,3.1140654,0.45270553,0.42183927,0.5178677,1.2277923,1.4232788,2.3389788,3.6079261,3.2649672,1.2998136,2.0646117,2.2086544,2.1469216,6.042933,6.3721733,7.764586,8.783174,8.903209,8.498518,8.851766,8.968371,9.873782,11.06042,10.497967,11.900668,11.821788,11.688034,12.325937,13.96185,13.4474125,13.138749,12.857523,12.30193,11.032983,11.105004,11.214751,10.995257,10.425946,9.825768,9.705732,9.81205,10.30591,10.878652,10.7586155,10.329918,10.580277,11.129011,11.447963,10.847785,10.518545,10.336777,10.542552,11.495977,13.656617,15.011304,14.918706,13.673765,12.432255,13.214201,13.9481325,15.302819,16.523752,17.017612,16.355703,15.46744,15.470869,16.023033,16.993607,18.509483,18.547209,19.140528,19.109661,18.149376,16.828985,16.523752,16.585485,16.105343,14.908417,13.564018,12.367092,11.345076,10.6317215,10.151579,9.613133,11.797781,13.241637,14.455711,16.149927,19.226267,16.492886,16.11906,16.856422,17.802988,18.403166,18.169954,17.754974,17.168514,16.441442,15.6252,12.55915,11.530273,12.147599,13.419975,13.749216,11.808069,10.707172,11.650309,13.588025,13.245067,11.523414,10.984968,10.971251,11.303921,12.267634,11.537132,11.005547,10.425946,9.801761,9.400499,8.570539,7.1712675,6.138962,5.6142344,4.945465,5.346727,5.593657,6.245279,7.233,7.8434668,8.501947,9.417647,9.784613,9.427936,8.803751,9.914937,10.477389,10.7757635,10.593996,9.2153015,10.497967,11.478829,11.698323,11.05699,9.81205,0.4355576,0.47328308,0.5521636,0.6173257,0.6344737,0.607037,0.61046654,0.64133286,0.65848076,0.6276145,0.50757897,0.5555932,0.6859175,0.823101,0.9259886,0.9877212,0.9534253,0.99801,0.9534253,0.8128122,0.7339317,0.7305021,0.8676856,1.0117283,1.0734608,1.0048691,0.9842916,1.0700313,1.1523414,1.2346514,1.4438564,1.6016173,1.8142518,1.9685832,1.9342873,1.5673214,1.4918705,1.3512574,1.255229,1.2655178,1.3924125,1.4404267,1.6324836,1.5947582,1.3306799,1.2517995,1.1729189,1.1763484,1.2860953,1.4781522,1.6873571,1.5810398,1.5158776,1.371835,1.1660597,1.0666018,1.0288762,1.1111864,1.1043272,0.980862,0.88826317,0.66191036,0.51100856,0.41840968,0.36010668,0.31552204,0.28465575,0.2709374,0.24007112,0.18176813,0.09602845,0.0548734,0.030866288,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.020577524,0.07888051,0.17833854,0.45613512,0.7442205,1.0288762,1.4507155,1.1111864,0.59674823,0.2194936,0.06516216,0.0034295875,0.006859175,0.28122616,0.7339317,1.0871792,0.8471081,1.313532,0.6927767,0.12346515,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.274367,0.548734,0.0034295875,0.30523327,0.24350071,0.2777966,0.490431,0.6036074,0.5521636,0.6173257,0.4938606,0.31895164,0.6756287,0.490431,0.2194936,0.082310095,0.07888051,0.024007112,0.048014224,0.034295876,0.024007112,0.024007112,0.017147938,0.0274367,0.037725464,0.048014224,0.06859175,0.12346515,0.09602845,0.08573969,0.10288762,0.14404267,0.216064,0.31209245,0.45956472,0.5555932,0.58645946,0.607037,0.65505123,0.75450927,0.9431366,1.2655178,1.7662375,2.435007,3.2203827,3.5153272,3.333559,3.309552,3.7965534,3.8685746,3.957744,4.32471,5.0346346,5.360445,5.504488,5.751418,6.186976,6.684266,6.619104,6.6293926,6.4064693,6.307011,7.3598948,7.1369715,7.366754,7.4284863,7.5039372,8.604835,8.05953,7.9017696,8.090397,8.378482,8.340756,9.4862385,10.600855,10.940384,10.878652,11.897239,12.377381,12.809509,12.936404,12.788932,12.665466,13.371962,12.449403,12.178465,13.029003,13.642899,14.678635,15.244516,15.724659,16.45173,17.703531,17.425734,16.45173,15.621771,15.309678,15.415996,14.534592,14.706071,14.284232,13.231348,13.101024,13.495427,13.742357,14.13333,14.743796,15.426285,15.618341,15.29253,14.891269,14.534592,14.023583,13.478279,14.088745,14.472859,14.099034,13.306799,13.029003,12.836946,13.05301,13.567448,13.838386,14.942713,15.820687,16.427725,16.55119,15.7966795,15.498305,15.364552,15.29253,15.450292,16.280252,16.338554,16.595774,16.986746,17.436022,17.837284,16.314548,15.038741,14.126471,13.54687,13.121602,13.478279,13.584596,13.9309845,14.424845,14.393978,14.87755,15.542891,15.71094,15.62863,16.45859,15.46401,16.300829,17.95046,19.243416,18.845583,21.095392,22.2786,23.866499,26.10602,28.006012,29.00402,31.34643,30.214666,23.585274,12.21962,16.359133,17.237106,14.0750265,8.251588,3.2992632,2.8739944,4.3487167,5.8474464,7.0546613,9.225591,10.168727,12.065289,14.2362175,15.909856,16.225378,15.71094,15.570327,15.6526375,15.6869335,15.278812,15.824117,16.45516,17.54234,18.996485,20.262003,19.829874,18.410025,17.357141,16.993607,16.619781,15.193072,14.733508,14.63062,14.068168,12.034423,11.430815,11.255906,10.882081,9.897789,8.100685,7.157549,6.824879,6.6705475,6.543653,6.560801,7.0443726,6.8728933,6.601956,6.3035817,5.5833683,5.576509,5.627953,5.7102633,5.7891436,5.861165,5.7274113,5.689686,5.7822843,5.895461,5.785714,6.2830043,6.677407,7.0923867,7.5245147,7.8331776,8.06639,7.932636,7.613684,7.2295704,6.835168,6.807731,7.157549,7.531374,7.7920227,8.018375,8.213862,8.289313,8.803751,9.589127,9.729739,9.561689,9.623423,9.571979,9.369633,9.294182,8.779744,8.961512,8.971801,8.491658,7.747438,8.028665,8.320179,8.464222,8.354475,7.9189177,7.5862474,7.257007,6.9963584,6.931196,7.2432885,7.301592,7.1232533,7.006647,7.133542,7.56224,7.7611566,8.1487,8.519095,8.831187,9.2153015,9.0369625,8.97523,8.7145815,8.207003,7.6788464,7.208993,7.0546613,7.1266828,7.191845,6.8626046,7.349606,8.05953,8.608265,9.06097,9.928656,9.657719,9.1810055,8.790032,8.687145,8.961512,9.578837,9.788043,9.959522,9.897789,8.851766,7.970361,7.56567,7.3564653,7.380472,7.98408,9.119273,11.074138,12.181894,12.168177,12.147599,12.912396,14.225929,15.426285,16.263103,16.907866,15.6252,14.164196,13.461131,13.615462,13.893259,13.893259,13.900118,13.598314,13.186764,13.375391,13.2862215,12.521424,11.619442,10.796341,9.942374,9.517105,9.026674,8.769455,8.827758,9.050681,9.006097,8.80718,8.440215,8.176137,8.56025,9.644,9.760606,9.156999,8.340756,8.100685,9.39707,10.233889,11.115293,12.212761,13.351384,12.490558,11.187314,10.511685,10.456812,9.959522,9.585697,10.076128,10.419086,10.31277,10.172156,10.518545,10.772334,10.696883,10.203023,9.349055,9.225591,9.23245,9.22216,9.325048,9.945804,10.930096,11.094715,10.528833,9.342196,7.6376915,6.8900414,7.3255987,7.949784,8.385342,8.872343,9.637141,9.97667,10.600855,11.46854,11.777204,12.528283,12.181894,12.154458,12.600305,12.394529,8.573969,8.89635,8.182996,6.1629686,7.466212,9.321619,10.851214,10.803201,10.343636,13.087306,11.893809,11.245617,11.235329,11.4033785,10.738038,11.170166,11.825217,12.065289,12.024134,12.614022,9.15014,8.172707,7.2467184,5.562791,3.9337368,3.1346428,5.3227196,6.310441,6.7219915,11.996697,9.283894,5.2609873,2.0303159,0.48357183,0.29151493,3.1483612,1.8245405,0.36696586,0.26064864,0.39783216,0.4424168,0.6756287,1.6530612,2.7368107,2.0920484,0.65505123,2.311542,2.6476414,1.978872,5.346727,4.0263357,4.3590055,6.433906,8.937505,9.170717,9.671436,9.815479,10.55284,11.543991,11.156448,11.986408,11.931535,11.996697,12.600305,13.570878,13.13532,13.063298,12.596875,11.478829,9.945804,9.990388,10.377932,10.161868,9.242738,8.361334,9.06097,9.678296,10.028113,10.172156,10.439664,10.031544,9.949233,10.319629,10.858074,10.88551,11.482259,12.264205,12.614022,12.624311,13.094165,15.0078745,15.765814,15.594335,15.097044,15.251375,15.985307,17.243965,18.403166,18.506054,16.283682,14.874121,15.343974,16.558048,17.679523,18.166525,18.838724,19.87789,19.86074,18.931322,18.78385,18.108221,17.724108,16.942162,15.666355,14.369971,13.046151,11.766914,10.666017,9.935514,9.80862,11.465111,12.960411,14.105893,14.634049,14.184773,8.48137,13.05301,17.137648,17.4566,18.183672,19.630959,20.169403,19.733847,18.526632,17.017612,15.525743,13.941273,12.960411,12.614022,12.257345,11.47197,11.046701,11.650309,12.751206,12.634601,11.351934,10.569988,10.39165,10.748327,11.399949,11.293632,10.566559,9.938945,9.568549,9.057541,8.570539,7.1095347,5.885172,5.3330083,5.137522,5.336438,5.562791,6.23156,7.3839016,8.697433,9.403929,9.609704,9.362774,8.820899,8.217292,8.539673,8.865483,8.920357,8.752307,8.738589,10.518545,11.996697,12.569438,12.055,10.703742,0.5418748,0.7579388,0.7339317,0.7442205,0.8162418,0.71678376,0.58645946,0.6859175,0.70649505,0.5761707,0.48357183,0.53844523,0.61046654,0.6756287,0.7476501,0.8711152,0.8128122,0.8848336,0.9568549,0.9877212,1.0185875,0.939707,0.86082643,0.89169276,1.0082988,1.039165,1.0666018,1.1934965,1.3032433,1.3615463,1.430138,1.3889829,1.5261664,1.5741806,1.4541451,1.2620882,1.196926,1.0494537,0.97400284,1.0666018,1.3615463,1.4095604,1.4198492,1.2963841,1.1043272,1.0666018,0.9911508,1.0323058,1.138623,1.2963841,1.5398848,1.5055889,1.4198492,1.2963841,1.1694894,1.1077567,1.1214751,1.1317638,1.0185875,0.8128122,0.69963586,0.6001778,0.48357183,0.40126175,0.34981793,0.26750782,0.24350071,0.23321195,0.19548649,0.12346515,0.041155048,0.024007112,0.017147938,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.11317638,0.31895164,0.58645946,0.8505377,1.0254467,0.6001778,0.24007112,0.041155048,0.0,0.0,0.0,0.12003556,0.5521636,1.0631721,0.9945804,0.97400284,0.4938606,0.11317638,0.017147938,0.006859175,0.006859175,0.010288762,0.037725464,0.058302987,0.0,0.0,0.0,0.1371835,0.274367,0.0,0.14061308,0.17147937,0.2503599,0.39097297,0.44584638,0.823101,0.9568549,0.72707254,0.36696586,0.490431,0.4629943,0.4081209,0.48700142,0.5727411,0.24007112,0.17147937,0.09602845,0.0548734,0.05144381,0.061732575,0.05144381,0.10288762,0.116605975,0.082310095,0.072021335,0.058302987,0.08916927,0.13375391,0.17833854,0.23664154,0.29494452,0.4046913,0.50757897,0.5761707,0.607037,0.6036074,0.6344737,0.71678376,0.90198153,1.2483698,1.6153357,2.153781,2.5241764,2.6956558,2.9322972,3.1586502,3.2889743,3.457024,3.7108135,4.0091877,4.187526,4.2046742,4.307562,4.57164,4.931747,5.411889,5.7994323,5.7925735,5.645101,6.159539,6.368744,6.468202,6.680836,7.1884155,8.14527,7.64798,7.5245147,7.98065,8.752307,9.098696,9.897789,10.971251,11.492548,11.530273,12.065289,12.048141,12.3533745,13.039291,13.824667,14.102464,14.2533655,13.214201,12.895248,13.557159,13.807519,14.1299,14.246507,14.243076,14.29452,14.661487,14.740367,14.640909,14.46257,14.435134,14.946142,14.640909,14.733508,14.3974085,13.711491,13.670336,13.992717,14.366542,15.014734,15.601193,15.217079,15.484588,15.0250225,14.369971,13.745787,13.077017,13.426835,13.433694,13.279363,13.097594,12.991278,13.029003,13.251926,13.327377,13.310229,13.653188,14.448852,15.090185,15.481158,15.549749,15.244516,15.035312,14.754086,14.743796,15.083325,15.584045,15.4742985,15.405707,15.5085945,15.848124,16.441442,15.4742985,14.764374,14.246507,13.872682,13.605173,13.896688,14.044161,14.3974085,14.88098,14.987297,15.824117,15.902997,16.091625,16.513464,16.54776,15.515453,17.737827,19.397747,19.435472,19.552078,21.44178,22.419212,24.425522,28.712505,35.839188,30.886866,28.390125,24.391226,18.132229,12.044711,16.383139,14.610043,10.374502,6.217842,3.5393343,2.877424,3.7931237,4.8288593,6.025785,8.89635,10.97468,13.004995,14.637479,16.023033,17.816708,17.226818,17.658945,17.70696,16.87014,15.573756,14.928994,15.278812,16.510035,18.30028,20.11796,19.967058,18.653526,17.847572,17.71039,16.894148,16.050468,15.601193,15.391989,15.031882,13.9138365,13.38568,12.830087,12.264205,11.478829,10.048691,8.858624,7.953213,7.1781263,6.660259,6.8043017,7.507367,7.73372,7.699424,7.4627824,6.9071894,6.509357,6.4304767,6.5333643,6.6876955,6.756287,6.4990683,6.3138704,6.324159,6.468202,6.4819202,6.7185616,6.7528577,6.8557453,7.0375133,7.0443726,7.442205,7.500508,7.517656,7.507367,7.205563,7.0032177,7.39762,7.8537555,8.1487,8.381912,8.416207,8.279024,8.632272,9.325048,9.414218,9.5205345,9.729739,9.829198,9.764035,9.630281,9.3593445,9.349055,9.239308,8.865483,8.275595,8.244728,8.31675,8.309891,8.1487,7.8606143,7.699424,7.394191,7.1712675,7.14726,7.301592,7.548522,7.6376915,7.455923,7.233,7.548522,7.5416627,7.6376915,7.7611566,7.888051,8.035523,7.888051,7.723431,7.6274023,7.6685576,7.870903,7.891481,7.874333,7.8949103,7.805741,7.2432885,7.6514096,8.107545,8.543102,8.992378,9.578837,10.089847,9.767465,9.283894,8.964942,8.786603,9.39021,9.445084,9.496528,9.613133,9.362774,8.625413,7.9086285,7.390761,7.250148,7.675417,8.200144,10.179015,11.845795,12.579727,12.926115,13.323947,14.308239,15.422854,16.228807,16.314548,15.134769,14.102464,13.423406,13.179905,13.306799,13.214201,13.13532,13.258785,13.6086035,14.009865,14.0750265,13.087306,11.996697,11.204462,10.563129,9.73317,9.448513,9.613133,10.021255,10.343636,10.655728,10.487679,10.179015,10.028113,10.257896,10.844356,11.465111,11.345076,10.405369,9.263316,9.938945,11.043272,12.130451,13.032433,13.876111,13.540011,12.322508,11.080997,10.347065,10.319629,9.414218,9.568549,9.750318,9.654288,9.705732,10.110424,10.357354,10.669447,10.9369545,10.683165,10.597425,10.539123,10.569988,10.734609,11.06042,11.71547,11.619442,11.197603,10.542552,9.39707,7.939495,7.723431,8.2310095,8.89635,9.119273,9.952662,10.247607,10.539123,10.906088,10.957532,11.283342,11.574858,11.952112,12.939834,15.440002,12.271064,12.79922,10.580277,6.7357097,9.942374,8.838047,10.261326,11.732618,12.408247,13.077017,12.370522,11.351934,10.967821,11.105004,10.569988,11.948683,12.127021,11.218181,10.628291,13.059869,8.745448,6.118384,4.314421,3.1209247,2.9906003,3.4776018,14.366542,15.597764,7.8194594,12.394529,10.089847,5.7651367,2.2600982,0.69963586,0.52815646,4.0091877,2.3595562,0.6927767,0.7339317,0.8162418,0.69963586,0.8093826,1.3169615,1.7250825,0.85739684,0.28465575,2.2978237,2.5996273,1.5261664,4.029765,2.6545007,4.0229063,6.574519,8.652849,8.488229,9.537683,9.839486,10.532263,11.595435,11.852654,12.089295,12.000127,11.88352,12.065289,12.915827,13.087306,12.380811,11.701753,11.077567,9.654288,9.602845,9.880642,9.781183,9.283894,9.047252,9.1981535,9.554831,9.777754,9.9698105,10.672876,11.447963,11.067279,10.676306,10.652299,10.593996,11.399949,12.157887,12.6586075,12.881531,13.018714,13.80409,14.544881,15.227368,15.755525,15.954441,16.702091,17.991615,19.44919,20.186552,18.773561,16.365992,16.029892,16.688372,17.432592,17.54234,18.28313,19.044498,19.078794,18.663815,19.078794,17.761833,17.525192,17.144508,16.143068,14.808959,13.38911,12.140739,11.129011,10.48082,10.405369,11.413667,13.272504,14.925565,15.367981,13.656617,10.820349,13.430264,16.077906,16.811838,17.130789,18.067066,19.600092,20.498644,20.207129,18.866161,18.814716,17.562918,15.999025,14.472859,12.809509,11.965831,12.109874,12.332796,12.109874,11.30049,10.618003,10.367643,10.295622,10.353925,10.672876,10.991828,10.4705305,9.945804,9.575408,8.824328,8.241299,6.9723516,5.8543057,5.302142,5.3158607,5.456474,5.761707,6.2692857,7.1369715,8.663138,9.273604,9.256456,9.012956,8.711152,8.282454,8.779744,9.321619,9.191295,8.659708,8.995808,10.995257,11.8869505,12.401388,12.579727,11.760056,0.7133542,0.939707,0.78537554,0.7373613,0.86082643,0.7956643,0.65848076,0.7579388,0.7510797,0.6036074,0.59331864,0.6036074,0.66533995,0.6859175,0.6824879,0.7922347,0.7682276,0.8471081,0.9534253,1.039165,1.08032,1.0151579,0.8676856,0.86082643,0.9877212,1.0048691,1.1146159,1.2758065,1.4129901,1.4678634,1.4198492,1.214074,1.2380811,1.2003556,1.039165,0.9294182,0.91912943,0.83338976,0.823101,0.9568549,1.2037852,1.2723769,1.2312219,1.1351935,1.0288762,0.9568549,0.9259886,0.9911508,1.1043272,1.2586586,1.5055889,1.5364552,1.4953002,1.4164196,1.3375391,1.2860953,1.3443983,1.2380811,0.980862,0.6824879,0.5590228,0.548734,0.47671264,0.39783216,0.32238123,0.22635277,0.19548649,0.17490897,0.13032432,0.06516216,0.01371835,0.01371835,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.07888051,0.22292319,0.41840968,0.5761707,0.5555932,0.31552204,0.12689474,0.024007112,0.0,0.0,0.0034295875,0.17147937,0.5624523,0.9774324,0.96371406,0.6893471,0.3566771,0.12003556,0.024007112,0.0,0.0,0.006859175,0.07545093,0.1371835,0.0,0.020577524,0.020577524,0.010288762,0.0,0.0,0.01371835,0.12003556,0.20577525,0.23664154,0.2503599,0.8265306,0.9294182,0.7373613,0.4424168,0.23664154,0.37382504,0.52472687,0.70306545,0.78194594,0.48014224,0.4115505,0.22635277,0.1097468,0.09945804,0.07888051,0.0548734,0.106317215,0.12346515,0.08573969,0.061732575,0.06516216,0.11317638,0.16119061,0.19891608,0.2503599,0.2503599,0.29837412,0.38754338,0.48014224,0.5144381,0.5178677,0.5418748,0.58302987,0.67219913,0.864256,1.0082988,1.255229,1.5776103,1.9720128,2.4315774,2.5138876,2.7573884,3.018037,3.1826572,3.1620796,3.1655092,3.1380725,3.1415021,3.234101,3.4673128,4.15323,4.770556,5.0620713,5.1066556,5.3158607,5.830299,5.9297566,6.111525,6.492209,6.831738,6.9860697,7.2604365,7.870903,8.759167,9.619993,9.918367,10.830637,11.530273,11.760056,11.845795,11.873232,12.05157,12.740917,13.780083,14.476289,14.044161,13.094165,12.936404,13.540011,13.519434,13.80409,13.96871,13.814379,13.4474125,13.251926,13.680624,13.944703,14.150477,14.455711,15.066177,15.090185,14.997586,14.654627,14.21564,14.126471,14.870691,15.518884,16.499744,17.027903,15.117621,14.88441,14.225929,13.622321,13.183334,12.648318,13.114742,12.857523,12.634601,12.734058,12.97413,13.190193,13.543441,13.485138,13.173045,13.502286,14.081886,14.623761,14.894698,14.839825,14.603184,14.623761,14.2362175,14.195063,14.486577,14.339106,14.13333,14.030442,14.05102,14.2533655,14.750656,14.4145565,14.239647,14.078457,13.934414,13.958421,14.479718,14.747226,15.100473,15.522313,15.62863,16.46888,16.400288,16.811838,17.576635,17.034761,17.19938,20.460918,20.53637,17.487467,17.744686,19.997925,21.798458,25.001692,30.633076,38.89152,30.725674,24.617579,18.969048,14.201921,12.754636,15.241087,12.243628,7.7268605,4.2938433,3.192946,2.4658735,2.452155,3.1106358,4.5990767,7.274155,10.22703,12.644889,14.225929,15.419425,17.425734,16.599203,17.367432,17.573206,16.839275,16.575195,15.542891,15.889278,16.7844,17.809847,18.934752,19.356592,18.900457,18.386019,17.947031,16.997036,16.20137,15.741806,15.549749,15.481158,15.3302555,15.083325,14.335675,13.516005,12.710052,11.677745,10.329918,9.294182,8.368194,7.7851634,8.213862,8.659708,8.779744,8.597976,8.128122,7.377043,7.099246,7.140401,7.2432885,7.3050213,7.3530354,7.3050213,7.2775846,7.2878733,7.3221693,7.349606,7.407909,7.3050213,7.233,7.2192817,7.099246,7.438775,7.7268605,7.970361,8.05953,7.7714453,7.5588107,7.870903,8.381912,8.89635,9.335337,9.108984,8.875772,8.97866,9.321619,9.3764925,9.630281,9.962952,10.230459,10.38479,10.48082,10.521975,10.281903,9.97324,9.619993,9.057541,8.368194,7.9120584,7.582818,7.3118806,7.06838,7.1061053,6.9792104,6.9517736,7.0786686,7.181556,7.500508,7.5931067,7.394191,7.1026754,7.181556,7.040943,7.06838,7.1987042,7.3221693,7.301592,7.160979,7.058091,7.160979,7.500508,7.966932,8.327039,8.484799,8.48137,8.368194,8.224151,8.457363,8.621983,8.844906,9.177576,9.616563,10.302481,10.1481495,9.818909,9.469091,8.748878,9.102125,8.968371,8.844906,8.940934,9.1981535,8.934075,8.440215,7.7680154,7.2295704,7.3839016,7.7714453,9.235879,10.834066,12.096155,13.056439,13.694343,14.424845,15.429714,16.362562,16.352274,15.241087,14.229359,13.409687,12.88496,12.761495,12.370522,12.13731,12.555719,13.454271,14.003006,14.140189,13.29994,12.271064,11.482259,10.984968,10.007536,9.8429165,10.353925,11.187314,11.756626,12.312219,12.425395,12.538571,12.627741,12.202472,11.72233,11.996697,12.295071,12.089295,11.036412,10.89237,11.893809,13.05301,13.828096,14.119612,13.999576,13.13532,11.835506,10.7586155,10.916377,10.216741,9.877212,9.757176,9.853205,10.295622,10.398509,10.556271,11.077567,11.770344,11.928105,11.876661,11.681175,11.674315,11.825217,11.749766,11.794352,11.598865,11.22161,10.710602,10.093276,8.803751,8.182996,8.491658,9.297611,9.472521,10.288762,10.463672,10.449953,10.463672,10.48082,10.494537,11.327928,12.212761,13.54687,16.921585,16.146498,12.977559,8.604835,6.138962,10.569988,9.736599,9.407358,10.134431,11.358793,11.434244,11.780633,10.827208,10.22703,10.89237,13.001566,13.330807,12.47341,10.518545,9.0369625,11.063849,7.208993,4.262977,2.726522,2.386993,2.3081124,3.0660512,12.521424,14.023583,8.4264965,14.095605,9.482809,6.036074,3.457024,1.920569,2.061182,7.675417,4.8597255,2.1880767,2.3492675,2.1332035,2.16064,1.8416885,1.9171394,1.920569,0.19891608,0.3018037,2.8019729,3.357566,2.0303159,3.2718265,2.3458378,4.139512,6.245279,7.366754,7.301592,9.095266,9.547972,10.31277,11.561139,11.962401,12.068718,12.243628,12.30536,12.3911,12.932974,12.991278,11.924676,11.207891,11.05699,10.425946,10.323058,10.206452,9.901219,9.530824,9.530824,9.383351,9.530824,9.942374,10.597425,11.495977,12.651748,12.319078,11.571428,11.036412,10.88551,11.660598,12.30536,12.912396,13.330807,13.190193,12.956982,13.536582,14.472859,15.340545,15.758954,16.341984,17.37772,19.054789,20.598103,20.29287,17.689812,16.660936,16.592344,16.835844,16.698662,17.240536,17.422304,17.20967,17.014183,17.682953,16.86671,16.973028,17.017612,16.475739,15.275383,13.780083,12.583157,11.739478,11.231899,10.981539,11.399949,13.097594,14.843254,15.566897,14.328816,13.87954,13.903547,14.740367,15.954441,16.328266,16.431154,17.580065,18.530062,18.591793,17.604073,18.410025,18.389448,17.847572,16.558048,13.762935,11.849225,11.821788,11.80121,11.022695,9.818909,10.072699,10.360784,10.398509,10.22703,10.182446,10.607714,10.326488,9.870353,9.39707,8.697433,7.9292064,6.927767,6.012067,5.4736214,5.5490727,5.768566,6.0806584,6.509357,7.2638664,8.755736,8.97866,9.0369625,9.22902,9.386781,8.875772,9.4862385,10.299051,10.319629,9.73317,9.873782,10.912948,11.180455,11.547421,11.945253,11.38623,0.8128122,0.83338976,0.6824879,0.6379033,0.7373613,0.7888051,0.764798,0.7339317,0.6962063,0.67219913,0.6824879,0.6241849,0.71678376,0.764798,0.72707254,0.7373613,0.77165717,0.8745448,0.9328478,0.91912943,0.8848336,0.9431366,0.94656616,1.0117283,1.0940384,0.9911508,1.1420527,1.3238207,1.4061309,1.3546871,1.2346514,0.97400284,0.97057325,0.9259886,0.77851635,0.72707254,0.75450927,0.7476501,0.823101,0.94999576,0.9568549,1.0563129,1.0563129,1.0323058,1.0014396,0.939707,1.0048691,1.1317638,1.2792361,1.4404267,1.6427724,1.704505,1.728512,1.670209,1.5536032,1.4815818,1.5604624,1.3169615,0.9328478,0.6001778,0.48357183,0.48014224,0.4389872,0.36696586,0.274367,0.19548649,0.15090185,0.106317215,0.061732575,0.0274367,0.01371835,0.01371835,0.006859175,0.0034295875,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.07888051,0.048014224,0.106317215,0.20234565,0.2469303,0.12689474,0.058302987,0.030866288,0.017147938,0.0,0.0034295875,0.116605975,0.50757897,0.82996017,0.91912943,0.8128122,0.5761707,0.31552204,0.12003556,0.024007112,0.0,0.0,0.0034295875,0.09945804,0.19548649,0.017147938,0.07545093,0.06859175,0.034295876,0.0,0.0,0.0,0.07888051,0.14747226,0.16462019,0.17147937,0.58988905,0.5796003,0.548734,0.5418748,0.20920484,0.34295875,0.5007198,0.5624523,0.53501564,0.5555932,0.59674823,0.4046913,0.26064864,0.21263443,0.09259886,0.061732575,0.061732575,0.058302987,0.058302987,0.116605975,0.1097468,0.12346515,0.14061308,0.16119061,0.20577525,0.16462019,0.17833854,0.24007112,0.31552204,0.33609957,0.37382504,0.44927597,0.50757897,0.548734,0.6207553,0.70649505,0.864256,1.0666018,1.3478279,1.8142518,1.9102802,2.1846473,2.4795918,2.6545007,2.585909,2.5961976,2.5996273,2.585909,2.620205,2.860276,3.2992632,3.981751,4.465323,4.698535,5.0140567,5.2644167,5.3501563,5.3981705,5.3913116,5.1512403,6.0497923,6.914048,7.6514096,8.323608,9.15014,9.191295,10.007536,10.875222,11.369082,11.372512,11.677745,11.766914,12.000127,12.55229,13.419975,12.929544,12.555719,12.823228,13.454271,13.361672,13.972139,14.596324,14.88098,14.778092,14.5585985,14.616901,14.640909,14.874121,15.265094,15.477728,15.254805,15.247946,15.004445,14.493437,14.092175,15.676644,16.750105,17.580065,17.484037,14.836395,13.876111,13.38911,13.152468,13.008426,12.843805,13.104454,13.056439,13.111313,13.351384,13.502286,13.649758,13.574307,13.101024,12.593445,12.950122,13.728639,14.479718,14.853543,14.726648,14.21564,14.376831,13.965281,13.725209,13.701202,13.234778,13.080446,13.152468,13.241637,13.310229,13.495427,13.423406,13.560589,13.72178,13.858963,14.037301,14.932424,15.433144,15.868701,16.245956,16.242527,17.21653,17.28512,17.79613,18.547209,17.778982,19.936192,23.458378,20.992504,14.339106,14.448852,17.960749,21.836184,26.421541,31.044626,34.01465,27.17605,21.098822,15.927004,12.607163,12.908967,13.042721,10.621432,6.848886,3.3781435,2.3046827,1.8965619,1.3478279,1.9171394,3.7519686,5.8988905,8.920357,11.592006,13.416546,14.490007,15.525743,14.592895,14.904987,14.904987,14.791811,16.520323,16.62321,17.28169,17.394867,17.014183,17.364002,18.094503,18.46147,18.187103,17.511473,17.2131,16.11906,15.6697855,15.590904,15.734947,16.091625,16.023033,15.477728,14.627191,13.673765,12.840376,11.578287,10.748327,10.05898,9.626852,9.9869585,9.757176,9.47595,9.009526,8.261876,7.1781263,7.5519514,7.747438,7.7440085,7.682276,7.8537555,8.128122,8.40249,8.443645,8.258447,8.097256,8.23444,8.375052,8.429926,8.399059,8.364764,8.23444,8.443645,8.64256,8.625413,8.351046,8.3922,8.673427,9.287323,10.124143,10.868362,10.446524,10.017825,9.743458,9.647429,9.623423,9.692014,10.089847,10.467101,10.72432,11.012405,11.30049,11.022695,10.580277,10.062409,9.249598,7.9463544,7.0546613,6.560801,6.3001523,5.9743414,6.0395036,5.994919,6.1149545,6.433906,6.7665763,7.0135064,6.8866115,6.756287,6.7185616,6.5813785,6.451054,6.5813785,6.8900414,7.1884155,7.181556,7.0478024,7.250148,7.613684,7.970361,8.117833,8.31675,8.515666,8.56368,8.628842,9.191295,9.030104,9.006097,8.937505,8.947794,9.458802,9.89436,10.100135,10.22703,10.048691,8.961512,8.838047,8.488229,8.285883,8.344186,8.519095,8.745448,8.913498,8.40249,7.466212,7.239859,7.8537555,8.7283,9.80519,10.984968,12.109874,13.365103,14.191633,15.182784,16.280252,16.756964,15.645778,14.232788,13.306799,12.9638405,12.590015,11.667457,11.290202,11.664027,12.535142,13.200482,13.502286,13.1593275,12.439114,11.667457,11.22161,10.563129,10.275044,10.662587,11.629731,12.682614,13.306799,13.876111,14.603184,14.953001,13.642899,11.331357,10.786053,11.640019,12.898679,12.926115,12.109874,12.415107,13.443983,14.5243025,14.7095,14.417986,13.756075,12.88839,12.106443,11.845795,11.581717,10.984968,10.693454,10.971251,11.712041,11.664027,11.941824,12.63803,13.409687,13.46799,13.169616,12.644889,12.319078,12.22648,12.027563,11.410237,11.252477,10.9369545,10.367643,9.97324,9.403929,8.690575,8.625413,9.170717,9.431366,10.429376,10.573419,10.412228,10.288762,10.336777,10.271614,11.30735,12.415107,13.762935,16.729528,17.700102,9.661148,3.6353626,4.139512,9.1810055,10.957532,8.361334,6.461343,7.023795,8.519095,9.510246,9.043822,8.755736,10.744898,17.573206,15.268523,13.272504,10.353925,7.301592,6.917478,4.6848164,3.2958336,3.1723683,3.3644254,1.5638919,2.1915064,2.2806756,3.7691166,9.414218,22.793037,11.928105,7.8606143,5.761707,3.9440255,3.8445675,10.878652,8.364764,5.809721,6.1149545,5.552502,4.245829,2.9563043,3.223812,3.7039545,0.1920569,1.3958421,3.8308492,4.8014226,4.2595477,4.8151407,3.3747141,4.2595477,5.312431,5.7651367,6.23156,8.296172,9.012956,9.9801,11.252477,11.321068,11.869802,12.346515,12.826657,13.190193,13.121602,12.55229,11.876661,11.365653,11.245617,11.660598,11.55428,11.146159,10.501397,9.822338,9.469091,9.523964,9.685155,10.47396,11.746337,12.6929035,13.334236,13.426835,12.912396,12.151029,11.928105,12.843805,13.471419,13.989287,14.21564,13.615462,13.166186,13.773223,14.325387,14.627191,15.388559,15.772673,16.273392,17.62122,19.325726,19.672113,17.806417,16.643787,16.012743,15.6697855,15.29939,15.741806,15.645778,15.182784,14.894698,15.676644,16.050468,16.311117,16.338554,16.084764,15.577187,14.435134,13.296511,12.456262,11.914387,11.345076,11.447963,12.404818,13.63604,14.596324,14.784951,14.774663,14.208781,14.284232,15.182784,16.064188,15.951012,15.738377,15.4742985,15.042171,14.157337,14.822677,15.9750185,17.185663,17.343424,14.668345,11.712041,10.847785,10.535692,9.9698105,9.081548,10.093276,10.635151,10.672876,10.319629,9.832627,9.97324,9.829198,9.462232,8.995808,8.628842,7.891481,7.1541195,6.433906,5.909179,5.919468,6.217842,6.4133286,6.866034,7.7714453,9.156999,9.191295,9.383351,9.932085,10.405369,9.716022,9.863494,10.765475,11.231899,11.05699,11.022695,10.436234,10.39508,10.521975,10.477389,9.959522,0.7613684,0.53158605,0.6379033,0.8025235,0.90884066,1.0082988,0.94656616,0.72021335,0.61046654,0.64819205,0.61046654,0.5624523,0.61389613,0.72364295,0.7990939,0.70306545,0.6790583,0.7339317,0.8093826,0.8711152,0.94656616,1.1420527,1.2003556,1.2312219,1.2586586,1.2346514,1.2483698,1.2895249,1.1832076,0.96714365,0.8711152,0.7339317,0.7579388,0.72021335,0.64133286,0.7613684,0.7613684,0.8711152,0.97057325,1.0082988,1.0082988,1.1043272,0.97400284,0.89512235,0.939707,0.9774324,1.2586586,1.4644338,1.5913286,1.6907866,1.862266,1.9239986,1.9925903,1.8965619,1.6770682,1.6187652,1.5673214,1.2175035,0.8265306,0.5418748,0.39783216,0.48357183,0.45613512,0.37725464,0.28122616,0.18176813,0.1097468,0.06516216,0.041155048,0.0274367,0.01371835,0.01371835,0.01371835,0.01371835,0.024007112,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.09259886,0.030866288,0.024007112,0.030866288,0.030866288,0.030866288,0.017147938,0.01371835,0.010288762,0.0034295875,0.01371835,0.52815646,1.0494537,1.1660597,0.922559,0.823101,0.48357183,0.22292319,0.07545093,0.024007112,0.0,0.0,0.010288762,0.09945804,0.20234565,0.09259886,0.17833854,0.13375391,0.0548734,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.0,0.29151493,0.14747226,0.14747226,0.34638834,0.26064864,0.18519773,0.2503599,0.26750782,0.22635277,0.274367,0.33609957,0.5521636,0.6241849,0.4698535,0.21263443,0.16462019,0.106317215,0.06516216,0.06859175,0.15090185,0.07888051,0.061732575,0.06859175,0.09602845,0.16804978,0.12003556,0.106317215,0.12346515,0.17833854,0.274367,0.21263443,0.31895164,0.44584638,0.53501564,0.59674823,0.6790583,0.764798,0.8025235,0.864256,1.1454822,1.3272504,1.529596,1.7113642,1.8999915,2.1812177,2.486451,2.4898806,2.411,2.3972816,2.5173173,2.760818,3.4810312,4.122364,4.4413157,4.5030484,4.4275975,4.125794,4.0091877,4.1017866,4.029765,4.8597255,5.744559,6.6465406,7.3427467,7.414768,7.915488,9.15014,10.528833,11.55428,11.8115,11.249047,11.173596,11.207891,11.502836,12.710052,12.648318,13.392539,14.376831,15.093615,15.107333,14.788382,14.956431,15.518884,16.184223,16.46545,15.683503,15.498305,15.721229,16.04018,15.9921665,14.928994,15.110763,15.241087,14.911846,14.616901,16.6335,18.142517,17.405157,15.217079,14.922135,12.895248,12.912396,13.059869,12.8197975,13.077017,14.627191,14.658057,14.352823,14.249936,14.2362175,14.040731,13.395968,12.517994,12.010415,12.864383,13.876111,14.321958,14.448852,14.421415,14.311668,14.092175,13.790371,13.423406,13.090735,12.953552,13.149038,13.21763,13.149038,13.056439,13.152468,13.190193,13.491997,13.814379,13.989287,13.917266,14.733508,15.553179,15.971589,16.21852,17.1205,18.327715,17.61436,17.439453,18.073925,17.607502,22.148275,25.300066,21.246294,13.485138,14.815818,19.089085,25.327503,29.85113,30.290117,25.6053,20.124819,16.143068,14.198492,13.505715,11.993267,11.149589,10.124143,7.1849856,3.2203827,1.7559488,1.6221949,1.4850113,1.8108221,3.0317552,5.56965,8.56025,10.624862,12.535142,14.243076,14.87755,14.658057,13.96185,12.576297,11.674315,13.810948,15.395418,16.396858,16.664366,16.54776,16.877,16.815268,16.479168,16.441442,16.832415,17.333136,16.61292,16.05733,15.971589,16.444872,17.350283,16.664366,16.047039,14.922135,13.708061,13.7938,13.183334,12.380811,11.787492,11.4376745,10.984968,10.669447,10.103564,9.407358,8.790032,8.546532,8.570539,8.375052,8.337327,8.536243,8.742019,8.999237,9.256456,9.263316,8.937505,8.378482,8.683716,9.06097,9.31133,9.366203,9.294182,8.40249,7.9943686,8.220721,8.793462,8.988949,9.328478,9.6817255,10.30934,11.2593355,12.343085,12.003556,11.067279,10.347065,10.072699,9.901219,9.709162,10.062409,10.264755,10.086417,9.781183,10.182446,10.072699,9.647429,9.091836,8.591117,7.442205,6.7185616,6.385892,6.2075534,5.7068334,5.48734,5.3227196,5.254128,5.3501563,5.693115,5.861165,5.8680243,5.9228973,6.0086374,5.874883,6.046363,6.217842,6.540223,7.010077,7.4627824,7.7783046,8.1041155,8.495089,8.790032,8.604835,8.433355,8.327039,8.176137,8.141841,8.666568,7.8606143,7.7714453,7.671987,7.4936485,7.798882,8.323608,9.047252,9.750318,10.086417,9.599416,8.536243,7.7680154,7.682276,8.213862,8.834618,8.652849,8.954653,8.886061,8.141841,6.958633,7.689135,8.543102,9.445084,10.216741,10.5597,11.756626,12.860953,13.896688,14.891269,15.854982,14.743796,13.687484,13.334236,13.457702,12.9707,11.773774,11.108434,11.015835,11.382801,11.931535,12.651748,12.9707,12.72034,12.075578,11.550851,11.63659,11.255906,11.039842,11.523414,13.121602,13.416546,14.157337,15.29939,15.841265,13.838386,8.467651,8.354475,10.782623,13.255356,13.488567,12.816368,12.63117,13.406258,14.781522,15.563468,15.319967,14.342535,13.831526,13.920695,13.701202,12.908967,12.809509,12.775213,12.603734,12.542002,13.032433,13.9138365,14.956431,15.786391,15.885849,15.371411,14.308239,13.478279,13.087306,12.771784,11.928105,11.30735,10.830637,10.460241,10.192734,9.887501,9.1810055,8.525954,8.309891,8.834618,10.347065,10.97468,10.998687,10.679735,10.237319,10.360784,10.957532,11.581717,12.346515,13.9481325,14.448852,9.719451,5.137522,3.9680326,7.3839016,9.6817255,9.266746,7.208993,5.284994,5.9812007,5.7994323,5.48734,5.07236,7.795452,20.111101,17.130789,14.932424,9.671436,3.4398763,4.256118,4.6608095,5.7754254,7.9600725,8.755736,2.884283,3.0420442,4.7945633,5.422178,12.075578,41.762085,27.724785,16.973028,9.880642,5.7377,2.7470996,7.6925645,10.813489,12.696333,13.536582,13.121602,5.6519604,2.49331,4.190956,6.492209,0.34981793,4.804852,4.619654,5.4153185,8.515666,10.9541025,6.193835,6.094377,6.478491,5.90232,5.645101,6.40304,7.881192,9.184435,9.918367,10.2236,11.55428,11.482259,11.588576,12.024134,11.537132,11.4754,11.742908,11.646879,11.355364,11.917816,11.72233,11.784062,11.482259,10.847785,10.542552,10.179015,10.05898,10.875222,12.459691,13.780083,14.791811,15.440002,15.134769,14.054449,13.138749,14.7369375,14.898128,14.874121,14.970149,14.5414505,14.260224,15.031882,14.891269,14.239647,15.837835,16.496315,16.55119,16.578627,16.997036,18.097933,16.877,15.656067,14.232788,12.929544,12.590015,13.491997,14.212211,14.417986,14.445422,15.275383,15.189643,15.055889,14.335675,13.684054,14.953001,15.405707,14.575747,13.481709,12.542002,11.5645685,11.821788,12.22648,12.915827,13.992717,15.518884,17.37429,17.178804,15.96816,15.014734,15.806969,16.12592,15.830976,15.529172,15.158776,13.96185,13.083877,13.440554,14.778092,16.21852,16.280252,14.181344,12.603734,11.382801,10.545981,10.316199,10.679735,11.375941,11.345076,10.419086,9.3079,8.796892,8.759167,8.796892,8.711152,8.529384,8.272165,7.8606143,7.3050213,6.7631464,6.5299344,6.6053853,6.632822,7.016936,7.9120584,9.23245,10.377932,10.47396,10.467101,10.593996,10.374502,9.448513,10.206452,11.022695,11.375941,11.842365,10.912948,10.508256,10.017825,9.534253,9.825768,0.7373613,1.0734608,0.7339317,0.4664239,0.48700142,0.50757897,0.5144381,0.52472687,0.5521636,0.5796003,0.5624523,0.90198153,0.7956643,0.71678376,0.7888051,0.7888051,0.65505123,0.7682276,0.91227025,1.0048691,1.0666018,1.0768905,1.0220171,1.0597426,1.1626302,1.138623,1.1214751,1.0082988,0.96714365,0.9431366,0.65162164,0.58302987,0.70306545,0.7888051,0.7956643,0.8471081,0.8471081,0.922559,0.97057325,0.9568549,0.90884066,1.1146159,0.97400284,0.84367853,0.91227025,1.1832076,1.5227368,1.7147937,1.8485477,1.978872,2.1297739,2.0063086,1.9274281,1.7525192,1.5364552,1.5433143,1.2998136,0.9362774,0.6790583,0.5658819,0.45613512,0.5624523,0.490431,0.36696586,0.25721905,0.17147937,0.106317215,0.072021335,0.048014224,0.030866288,0.0274367,0.017147938,0.024007112,0.030866288,0.034295876,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.006859175,0.0034295875,0.006859175,0.006859175,0.006859175,0.0034295875,0.0034295875,0.0034295875,0.024007112,0.12346515,1.3512574,1.8588364,1.5433143,0.7956643,0.5418748,0.30866286,0.13375391,0.048014224,0.0274367,0.01371835,0.01371835,0.01371835,0.037725464,0.06859175,0.0548734,0.10288762,0.106317215,0.12689474,0.12689474,0.0,0.15776102,0.20234565,0.15090185,0.09259886,0.19548649,0.14747226,0.37725464,0.3841138,0.22978236,0.5144381,0.35324752,0.28808534,0.22292319,0.20234565,0.39783216,0.41840968,0.48014224,0.5041494,0.4424168,0.274367,0.432128,0.30866286,0.20577525,0.22978236,0.28808534,0.22292319,0.23664154,0.2709374,0.29837412,0.31552204,0.274367,0.20577525,0.16119061,0.15776102,0.17833854,0.17490897,0.25721905,0.33609957,0.39440256,0.48357183,0.61046654,0.6824879,0.7922347,0.94656616,1.0700313,1.1180456,1.1454822,1.1626302,1.2037852,1.3272504,1.5638919,1.7182233,1.8725548,2.061182,2.2600982,2.3801336,2.7230926,3.2032347,3.673088,3.940596,3.426158,3.350707,3.508468,3.7691166,4.0777793,4.839148,5.346727,5.7479887,6.0223556,5.9880595,7.0443726,9.242738,10.47396,10.329918,10.124143,9.517105,9.331907,10.014396,11.31078,12.295071,13.55373,14.1299,14.201921,14.184773,14.7026415,14.239647,14.634049,14.96329,15.035312,15.415996,14.983868,14.455711,14.229359,14.21564,13.807519,14.774663,15.436573,15.453721,15.388559,16.70552,18.475187,19.850452,19.312008,16.345413,11.430815,11.622872,12.46312,12.682614,12.572867,13.992717,15.247946,15.193072,14.46257,13.749216,13.783512,13.169616,12.4802685,12.181894,12.363663,12.740917,13.656617,14.538021,15.066177,14.973578,14.030442,13.498857,13.337666,13.152468,12.891819,12.843805,12.826657,13.001566,13.104454,13.101024,13.190193,13.402828,14.181344,14.421415,13.965281,13.598314,14.486577,15.553179,16.263103,16.588915,17.021042,18.36887,18.193962,18.650097,19.857311,19.891607,23.437801,26.740494,24.878227,19.411465,18.36887,23.520111,32.3513,34.08667,27.090311,18.879879,14.092175,15.865272,14.479718,9.506817,9.80862,13.049581,11.050131,6.7219915,2.7745364,1.7319417,1.214074,0.97057325,1.313532,2.2429502,3.4467354,5.6073756,6.8145905,8.539673,10.875222,12.535142,12.891819,13.245067,12.943263,12.439114,13.296511,13.361672,14.507155,15.868701,16.894148,17.353712,16.45173,15.854982,15.944152,16.619781,17.28512,16.976458,16.894148,16.609491,16.444872,17.484037,17.024471,16.242527,15.738377,15.5085945,14.942713,14.291091,13.224489,12.397959,11.924676,11.365653,10.998687,10.738038,10.484249,10.131001,9.534253,9.431366,9.47595,9.575408,9.688584,9.818909,9.80862,9.582268,9.551401,9.750318,9.853205,9.798331,9.822338,9.818909,9.73317,9.571979,8.632272,7.8503256,7.675417,8.107545,8.694004,9.97324,11.05699,11.910957,12.504276,12.809509,12.319078,11.441104,10.676306,10.288762,10.2921915,10.275044,10.460241,10.323058,9.911508,9.829198,9.6645775,9.767465,9.657719,9.256456,8.872343,8.738589,7.606825,6.5470824,5.9228973,5.4016004,5.103226,4.98662,5.0895076,5.3913116,5.802862,6.118384,5.919468,5.6828265,5.501058,5.0929375,5.254128,5.658819,6.0052075,6.327589,6.9860697,7.4799304,7.7748747,8.083538,8.351046,8.2653055,8.152129,7.8331776,7.6376915,7.7748747,8.337327,7.7371492,7.3393173,7.1952744,7.2878733,7.517656,7.798882,8.412778,8.995808,9.331907,9.342196,8.700864,7.7131424,7.3118806,7.7131424,8.443645,8.347616,8.467651,8.738589,8.992378,8.971801,8.433355,8.923786,9.458802,9.849775,10.731179,11.749766,12.504276,13.049581,13.5503,14.280802,13.704632,13.341095,13.176475,13.056439,12.6757555,12.164746,11.427385,11.032983,11.14273,11.506266,12.000127,12.600305,13.066729,13.176475,12.710052,12.768354,12.415107,12.020704,12.027563,12.950122,13.203912,14.092175,15.0456,14.79524,11.348505,10.432805,11.664027,12.6757555,12.792361,13.025573,13.183334,13.762935,14.843254,15.916716,15.868701,14.579176,13.766364,13.732068,14.328816,14.946142,14.514014,14.332246,13.869251,13.193623,12.946692,13.951562,14.918706,15.875561,16.616352,16.715809,16.084764,15.021593,13.900118,13.306799,14.054449,13.992717,13.190193,12.493987,12.157887,11.842365,10.285333,9.89436,9.352485,8.47451,8.200144,10.388221,11.965831,12.586586,12.229909,11.204462,11.207891,11.358793,11.543991,11.814929,12.408247,14.198492,12.620882,9.047252,6.1492505,7.8983397,5.6999745,7.5382333,8.3922,7.1369715,6.543653,6.0669403,5.844017,8.069819,10.960961,8.745448,12.349944,13.927555,9.578837,2.301253,1.9857311,2.5961976,4.5819287,7.140401,8.927217,8.083538,10.086417,10.257896,9.318189,10.508256,19.572655,24.586712,20.443771,12.723769,5.977771,3.7108135,5.638242,12.092726,18.866161,22.26831,19.140528,12.55915,7.953213,6.927767,7.2432885,2.7916842,3.9474552,3.8377085,5.586798,9.0644,10.871792,9.342196,8.525954,7.3084507,5.8817425,5.744559,7.2432885,7.98408,8.553391,9.091836,9.321619,10.55284,10.398509,10.72775,11.492548,10.741467,10.847785,11.852654,11.849225,10.960961,11.355364,12.0309925,11.327928,10.597425,10.247607,9.72631,9.253027,9.589127,10.504827,11.698323,12.80265,14.195063,16.314548,16.997036,16.074476,15.385129,15.772673,14.994157,14.243076,14.057879,14.335675,15.138199,16.187653,16.931873,16.94902,15.9613,14.891269,16.095055,18.084215,19.69955,20.135109,17.418875,14.88098,12.943263,11.928105,12.065289,12.4974165,12.939834,13.282792,13.817808,15.223939,15.364552,15.46401,15.100473,14.592895,15.001016,15.738377,15.827546,15.477728,14.730078,13.471419,13.656617,13.927555,13.625751,13.3033695,14.712931,18.746124,19.21255,18.115082,16.88386,16.355703,16.527182,16.37971,16.462019,16.324837,14.5243025,14.181344,13.814379,13.46799,13.341095,13.790371,14.280802,13.574307,12.627741,11.856084,11.146159,11.091286,11.002116,10.545981,9.688584,8.683716,8.320179,8.018375,8.128122,8.436785,8.176137,8.340756,8.477941,7.9772205,7.1369715,7.1781263,7.1061053,7.3084507,7.7611566,8.303031,8.632272,9.887501,10.038403,10.024684,10.264755,10.679735,10.525404,10.696883,10.97468,11.516555,12.878101,12.116733,11.465111,10.525404,9.410788,8.766026,0.65162164,0.9362774,0.78537554,0.7133542,0.7990939,0.6824879,0.6859175,0.6859175,0.8162418,0.9568549,0.7339317,1.4507155,0.9945804,0.5796003,0.61389613,0.6893471,0.764798,0.8848336,1.1351935,1.3375391,1.0254467,0.9877212,0.97400284,0.9877212,0.980862,0.84024894,0.82996017,0.8025235,0.84367853,0.90541106,0.7956643,0.70306545,0.6927767,0.72364295,0.78537554,0.8779744,0.8779744,0.9877212,1.0700313,1.0631721,0.9568549,1.0597426,0.9877212,0.90541106,0.91569984,1.0631721,1.4678634,1.7010754,1.8245405,1.8519772,1.7593783,1.6221949,1.5124481,1.3752645,1.255229,1.2895249,1.0837497,0.8471081,0.65505123,0.5418748,0.51100856,0.53158605,0.48357183,0.38754338,0.28122616,0.19548649,0.12689474,0.07888051,0.05144381,0.041155048,0.041155048,0.041155048,0.07545093,0.072021335,0.030866288,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12346515,0.2503599,0.0,0.030866288,0.020577524,0.010288762,0.006859175,0.0,0.006859175,0.010288762,0.017147938,0.072021335,0.24350071,1.4267083,1.8073926,1.5261664,0.91569984,0.490431,0.20920484,0.16119061,0.1097468,0.010288762,0.006859175,0.006859175,0.010288762,0.017147938,0.024007112,0.037725464,0.12346515,0.09602845,0.07888051,0.10288762,0.082310095,0.12346515,0.116605975,0.09259886,0.1097468,0.23664154,0.15090185,0.32238123,0.36353627,0.29494452,0.5418748,0.490431,0.4972902,0.36010668,0.16462019,0.28122616,0.30866286,0.29837412,0.33266997,0.41498008,0.47328308,0.65162164,0.50757897,0.41840968,0.4629943,0.42869842,0.26750782,0.30523327,0.37039545,0.3841138,0.37725464,0.3566771,0.31209245,0.22292319,0.14747226,0.20920484,0.17490897,0.21263443,0.28122616,0.35324752,0.42183927,0.51100856,0.61389613,0.6790583,0.7305021,0.86082643,0.90198153,0.9602845,0.9568549,0.9568549,1.1489118,1.1592005,1.2380811,1.3272504,1.4267083,1.611906,1.937717,2.0680413,2.2498093,2.5173173,2.6750782,2.5721905,2.7916842,3.0797696,3.3781435,3.82399,4.4447455,4.5647807,4.619654,4.73969,4.7602673,5.9126086,8.080108,9.328478,9.15014,8.450503,8.663138,8.838047,9.788043,11.406808,12.648318,13.203912,13.330807,13.104454,12.840376,13.090735,12.812939,13.152468,13.193623,13.1421795,14.335675,13.673765,12.950122,12.737488,12.782072,11.986408,13.310229,14.695783,15.278812,15.662926,17.940172,18.245405,18.608942,18.362011,16.79126,13.1421795,12.46312,12.679185,12.662037,12.46312,13.279363,13.701202,13.985858,13.735497,13.111313,12.840376,12.024134,12.010415,12.133881,12.103014,12.0138445,12.994707,13.749216,14.359683,14.5414505,13.649758,13.056439,12.939834,12.956982,12.929544,12.843805,13.371962,13.526293,13.570878,13.687484,13.975569,14.284232,14.997586,15.217079,14.898128,14.846684,15.103903,15.649208,16.252815,16.739817,16.96274,18.317427,18.87645,19.857311,21.208569,21.623549,25.814505,31.26412,30.814844,24.548986,19.78872,25.049707,32.848587,31.658522,22.069395,16.811838,12.775213,13.831526,13.660047,11.019264,9.746887,17.412016,12.607163,5.8165803,2.2223728,1.704505,1.5570327,1.0048691,1.0460242,1.7422304,2.2360911,4.0949273,5.099797,6.210983,7.7542973,9.421077,10.63858,12.185325,12.915827,12.843805,13.1421795,13.203912,14.037301,14.647768,14.870691,15.364552,15.206791,15.042171,15.505165,16.328266,16.338554,16.650646,17.645227,18.187103,18.019053,17.744686,17.117071,16.750105,16.578627,16.331696,15.539461,15.415996,14.771234,14.267084,13.858963,12.795791,12.264205,12.116733,12.096155,11.828648,10.823778,10.652299,10.6488695,10.611144,10.528833,10.569988,10.755186,10.48082,10.398509,10.672876,11.002116,10.686595,10.573419,10.621432,10.618003,10.192734,9.451943,8.858624,8.64942,8.903209,9.527394,10.607714,11.712041,12.394529,12.600305,12.6586075,12.274493,11.255906,10.316199,9.798331,9.678296,9.863494,9.959522,9.97667,9.952662,9.952662,9.273604,9.091836,9.054111,8.988949,8.913498,8.597976,7.56224,6.550512,5.8988905,5.5250654,5.2472687,5.055212,5.2026844,5.6793966,6.2212715,6.3653145,6.39961,6.0875177,5.5079174,5.099797,5.360445,5.7136927,6.0875177,6.433906,6.7391396,7.3187394,7.5862474,7.675417,7.73029,7.8949103,7.781734,7.5725293,7.6171136,7.9189177,8.128122,7.723431,7.421627,7.2467184,7.2535777,7.5210853,7.5107965,7.932636,8.361334,8.615124,8.7283,8.453933,7.706283,7.164408,7.1232533,7.4765005,7.5862474,7.8091707,8.309891,8.930646,9.191295,8.608265,8.659708,9.016385,9.602845,10.580277,11.293632,12.034423,12.648318,12.991278,12.960411,13.145609,13.354814,13.365103,13.104454,12.641459,12.144169,11.444533,11.06042,11.050131,11.022695,11.485688,11.97269,12.583157,13.248496,13.742357,13.9309845,13.855534,13.7526455,13.732068,13.780083,14.088745,14.767803,15.343974,15.316538,14.160767,14.7369375,14.1299,13.265644,12.71691,12.699762,12.850664,13.536582,14.88441,16.400288,16.942162,15.7795315,14.706071,14.030442,13.858963,14.085316,14.126471,14.191633,14.174485,14.157337,14.428274,15.189643,16.12935,17.154797,17.96761,18.067066,17.099922,16.146498,14.994157,13.893259,13.560589,13.780083,13.87954,13.906977,13.924125,14.009865,12.274493,11.331357,10.569988,9.938945,9.945804,11.63659,13.097594,13.745787,13.471419,12.651748,12.356804,12.277924,12.212761,12.127021,12.161317,13.416546,13.780083,12.0309925,9.132992,8.237869,6.7391396,7.6788464,7.7885933,7.486789,10.88551,9.860064,7.891481,8.697433,10.405369,5.5490727,8.2481575,8.429926,5.5490727,1.5913286,1.0528834,1.2072148,2.6819375,4.5510626,7.6616983,14.63062,18.890167,18.44775,15.21022,12.843805,16.78783,15.515453,12.953552,10.299051,8.1041155,6.2487082,8.001227,11.015835,14.0750265,16.417435,17.744686,15.573756,12.38767,9.709162,7.6376915,4.8322887,5.453044,5.2438393,6.7357097,9.338767,9.349055,8.275595,8.570539,7.822889,6.3378778,7.15069,6.9654922,7.630832,8.279024,8.735159,9.513676,10.203023,9.818909,9.962952,10.72432,10.652299,10.72089,11.962401,12.46998,11.945253,11.701753,11.506266,10.347065,9.489669,9.325048,9.366203,9.2153015,10.288762,11.595435,12.545431,12.943263,14.315098,16.12592,16.901007,16.561478,16.393429,16.492886,15.484588,14.819247,14.805529,14.613472,15.906426,17.096493,18.019053,18.38259,17.785841,16.077906,16.513464,18.62609,20.958208,21.057667,17.837284,14.308239,11.955542,11.266195,11.749766,12.644889,13.101024,12.9809885,13.066729,15.055889,16.005884,15.738377,15.121051,14.781522,15.114192,15.848124,16.074476,15.923574,15.539461,15.073037,14.754086,15.271953,14.651197,13.21763,13.588025,15.350834,16.616352,17.758404,18.639809,18.581505,17.230247,16.019604,15.683503,15.690363,14.243076,14.472859,14.061309,13.395968,12.994707,13.471419,13.251926,12.439114,11.80121,11.495977,11.067279,10.618003,10.477389,10.079557,9.280463,8.347616,7.9429245,7.7131424,7.8126,7.997798,7.6205435,7.8434668,8.001227,7.8503256,7.5245147,7.531374,7.56224,7.881192,8.337327,8.776315,9.050681,10.268185,10.542552,10.449953,10.360784,10.436234,10.38479,10.436234,10.48082,10.772334,11.910957,11.578287,11.0981455,10.247607,9.177576,8.405919,0.65162164,0.65162164,0.66876954,0.78194594,0.90884066,0.8128122,0.72707254,0.70649505,0.84367853,1.0014396,0.805953,1.3169615,1.0871792,0.9259886,0.97057325,0.65848076,0.89512235,0.9568549,1.1146159,1.2723769,0.94656616,0.9534253,0.91227025,0.8676856,0.83338976,0.78537554,0.7956643,0.7682276,0.764798,0.7888051,0.77851635,0.7442205,0.70649505,0.7305021,0.8265306,0.96371406,0.91569984,1.0220171,1.1008976,1.0871792,1.039165,1.0288762,1.0014396,0.9568549,0.90541106,0.86082643,1.1934965,1.3889829,1.4747226,1.4575747,1.313532,1.2106444,1.0940384,1.0117283,0.99801,1.0494537,0.91912943,0.78537554,0.6379033,0.5212973,0.5521636,0.50757897,0.47328308,0.39440256,0.28122616,0.18862732,0.13032432,0.082310095,0.058302987,0.06859175,0.12003556,0.16119061,0.14404267,0.08916927,0.030866288,0.010288762,0.0034295875,0.0,0.034295876,0.07545093,0.041155048,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12346515,0.2503599,0.0,0.0548734,0.037725464,0.01371835,0.017147938,0.017147938,0.024007112,0.034295876,0.07545093,0.30866286,1.0185875,1.4267083,1.3821237,1.1111864,0.7510797,0.34638834,0.1371835,0.17147937,0.14061308,0.0034295875,0.0,0.0,0.006859175,0.01371835,0.024007112,0.037725464,0.14404267,0.07888051,0.0548734,0.1371835,0.22978236,0.22292319,0.08916927,0.041155048,0.116605975,0.18519773,0.216064,0.33952916,0.4115505,0.4389872,0.5693115,0.53158605,0.5727411,0.48014224,0.28808534,0.26407823,0.20234565,0.15090185,0.2194936,0.40126175,0.5521636,0.5555932,0.53844523,0.5041494,0.45956472,0.40126175,0.3841138,0.41840968,0.432128,0.4046913,0.37382504,0.32581082,0.32238123,0.2777966,0.21263443,0.2503599,0.21263443,0.1920569,0.2503599,0.34981793,0.36010668,0.41498008,0.53501564,0.5624523,0.5555932,0.7922347,0.7407909,0.8162418,0.83338976,0.823101,1.0597426,1.0528834,1.1008976,1.1043272,1.0734608,1.1351935,1.4815818,1.5364552,1.5776103,1.6976458,1.8073926,1.9720128,2.2052248,2.4418662,2.719663,3.1723683,3.625074,3.8342788,3.99204,4.1326528,4.15666,5.144381,6.5882373,7.4524937,7.3839016,6.711703,7.3530354,7.9257765,8.97866,10.4705305,11.80121,11.5645685,11.55771,11.38623,11.022695,10.786053,10.792912,11.30049,11.427385,11.4754,12.956982,12.274493,11.561139,11.465111,11.760056,11.327928,12.4802685,14.092175,15.079896,15.724659,17.655516,16.986746,16.149927,15.772673,15.621771,14.592895,13.457702,13.011855,12.80265,12.63803,12.576297,12.4974165,12.542002,12.442543,12.144169,11.808069,11.153018,11.461681,11.688034,11.585147,11.677745,12.555719,13.282792,13.841815,14.033872,13.478279,13.13189,12.72034,12.6586075,12.953552,13.224489,13.978998,14.188204,14.198492,14.263655,14.544881,14.894698,15.395418,15.601193,15.501736,15.525743,15.251375,15.367981,15.930434,16.681513,17.034761,18.45461,19.342873,20.52951,22.055677,23.163433,28.064314,35.73973,35.774025,28.132906,23.142857,25.042849,29.415571,26.579304,17.562918,14.109323,11.982979,12.339656,12.325937,11.8115,13.419975,21.887627,14.013294,5.127233,1.7147937,1.4267083,1.6290541,1.0185875,0.8196714,1.2449403,1.4987297,2.9494452,3.7725463,4.4756117,5.4667625,7.0478024,7.963502,9.712592,11.118723,11.897239,12.641459,13.245067,13.584596,13.371962,12.994707,13.516005,13.718349,13.807519,14.459141,15.385129,15.337115,16.266533,17.497755,18.45461,18.674105,17.78927,17.274832,17.326277,17.240536,16.852993,16.510035,16.506605,16.184223,15.885849,15.494876,14.407697,13.865822,13.581166,13.495427,13.3033695,12.435684,12.439114,12.240198,12.003556,11.852654,11.852654,11.880091,11.72233,11.7086115,11.948683,12.325937,12.041282,11.650309,11.523414,11.5645685,11.2250395,10.463672,10.096705,10.000677,10.22703,11.005547,11.567999,12.05157,12.072148,11.667457,11.286773,11.118723,10.319629,9.637141,9.373062,9.366203,9.551401,9.386781,9.438225,9.764035,9.904649,9.554831,9.108984,8.738589,8.525954,8.443645,8.200144,7.606825,6.927767,6.351596,5.9914894,5.826869,5.6485305,5.7136927,6.0223556,6.276145,6.3035817,6.461343,6.2864337,5.826869,5.6313825,5.8680243,6.046363,6.3893213,6.8043017,6.8900414,7.140401,7.298162,7.2535777,7.226141,7.7783046,7.7542973,7.6342616,7.747438,8.008087,7.9086285,7.6376915,7.394191,7.2124224,7.181556,7.4456344,7.298162,7.517656,7.740579,7.915488,8.296172,8.196714,7.6342616,7.0786686,6.773435,6.7391396,7.058091,7.438775,7.9772205,8.56368,8.886061,8.604835,8.368194,8.553391,9.22216,10.110424,10.4705305,11.156448,12.000127,12.614022,12.356804,12.764925,13.087306,13.152468,12.926115,12.507706,12.0309925,11.454823,11.012405,10.80663,10.803201,11.235329,11.47197,11.893809,12.706621,13.954991,14.544881,14.915276,15.2033615,15.326826,14.970149,15.402277,15.9613,16.37285,16.62321,16.94902,18.087645,17.412016,15.858413,14.263655,13.38911,13.6086035,13.869251,14.692352,16.009314,17.158226,16.516893,15.484588,14.407697,13.649758,13.591455,13.934414,14.153908,14.373401,14.7369375,15.391989,16.060759,16.945591,17.730967,18.262554,18.54378,17.823566,16.955881,15.920145,14.812388,13.838386,13.845244,14.284232,14.832966,15.313108,15.683503,14.260224,12.713481,11.626302,11.341646,11.979549,12.939834,14.057879,14.647768,14.654627,14.654627,14.315098,14.171056,14.057879,13.9138365,13.790371,14.143619,14.712931,14.400838,12.908967,10.731179,9.949233,9.606275,8.656279,8.31332,12.068718,10.906088,7.8949103,7.596536,8.947794,5.23698,5.3741636,12.397959,11.423956,2.6819375,1.5227368,1.728512,2.3904223,3.549623,6.3721733,13.149038,18.78042,19.507494,17.161655,14.407697,14.760944,8.457363,5.950334,7.130112,9.9801,10.576848,14.232788,13.6086035,12.6757555,13.2862215,15.148488,16.324837,13.845244,10.425946,7.6514096,5.98463,5.8405876,5.9331865,7.390761,9.194724,8.176137,6.385892,6.742569,6.543653,5.970912,8.076678,6.694555,6.8728933,7.5862474,8.453933,9.764035,9.757176,9.194724,9.2153015,9.897789,10.251037,10.744898,11.746337,12.404818,12.373952,11.814929,11.197603,10.209882,9.448513,9.239308,9.647429,9.932085,11.249047,12.607163,13.423406,13.529722,13.958421,14.802099,15.738377,16.578627,17.261114,17.302269,16.88386,16.45859,16.149927,15.752095,16.499744,17.806417,19.075365,19.977346,20.464348,18.890167,17.988186,18.962189,20.903336,20.793589,17.916164,14.764374,12.411677,11.454823,12.017275,13.001566,13.443983,13.296511,13.258785,14.764374,16.033321,15.422854,14.46257,13.96871,14.054449,14.342535,14.54831,14.846684,15.29253,15.810398,15.549749,16.177364,15.858413,14.466,13.612033,12.929544,13.924125,15.827546,17.916164,19.480057,17.487467,15.446862,14.287662,13.992717,13.615462,14.040731,13.718349,13.426835,13.540011,14.057879,12.71691,11.667457,11.194174,11.1393,10.899229,10.041832,9.788043,9.534253,8.954653,8.021805,7.675417,7.5862474,7.599966,7.5588107,7.31531,7.455923,7.6925645,7.9600725,8.186425,8.268735,8.40249,8.666568,8.98209,9.349055,9.846346,10.683165,10.926665,10.772334,10.446524,10.209882,10.285333,10.30591,10.209882,10.131001,10.398509,10.388221,10.127572,9.523964,8.704293,8.018375,0.6859175,0.4972902,0.48014224,0.5624523,0.65848076,0.6790583,0.52472687,0.53844523,0.59674823,0.64133286,0.6859175,0.6173257,0.9534253,1.371835,1.4610043,0.7099246,0.94656616,0.922559,0.85739684,0.8471081,0.864256,0.91569984,0.8196714,0.7579388,0.805953,0.9362774,0.9431366,0.805953,0.6927767,0.6344737,0.5555932,0.7099246,0.7682276,0.8128122,0.8848336,0.9877212,0.90541106,1.0048691,1.0494537,1.0185875,1.1146159,1.0837497,1.0220171,0.94999576,0.85739684,0.7305021,0.881404,0.9568549,0.9842916,0.9877212,0.99801,0.9431366,0.83681935,0.7956643,0.8505377,0.91227025,0.805953,0.69963586,0.59674823,0.53844523,0.6001778,0.53158605,0.48357183,0.38754338,0.2503599,0.16119061,0.13032432,0.09259886,0.082310095,0.14404267,0.31209245,0.36353627,0.2503599,0.12346515,0.05144381,0.0034295875,0.0,0.0,0.06859175,0.16119061,0.116605975,0.082310095,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.0548734,0.037725464,0.037725464,0.07545093,0.12346515,0.20920484,0.24350071,0.2777966,0.6893471,2.1469216,1.5227368,0.97057325,0.5693115,0.31209245,0.09945804,0.09259886,0.12689474,0.12003556,0.058302987,0.0034295875,0.0,0.0034295875,0.020577524,0.05144381,0.0548734,0.1371835,0.09602845,0.13032432,0.26407823,0.33609957,0.44927597,0.216064,0.116605975,0.20920484,0.09602845,0.2777966,0.47328308,0.607037,0.65848076,0.64819205,0.5624523,0.490431,0.4698535,0.4629943,0.3566771,0.23664154,0.13032432,0.19548649,0.38754338,0.44584638,0.26407823,0.39783216,0.4355576,0.31209245,0.29837412,0.5590228,0.5418748,0.4664239,0.41840968,0.36353627,0.29151493,0.28122616,0.30523327,0.32238123,0.26750782,0.26407823,0.18862732,0.22978236,0.3566771,0.31895164,0.34638834,0.4664239,0.52472687,0.58302987,0.89512235,0.6756287,0.71678376,0.7510797,0.7407909,0.8848336,1.0768905,1.1934965,1.1832076,1.0906088,1.0425946,1.1351935,1.2003556,1.2689474,1.3752645,1.5501735,1.5981878,1.6256244,1.7113642,1.9171394,2.2806756,2.585909,3.216953,3.7313912,3.9474552,3.9440255,4.602506,5.195825,5.4496145,5.3570156,5.1821065,5.528495,6.2727156,7.301592,8.440215,9.455373,9.14328,9.280463,9.277034,8.947794,8.512236,8.841476,9.705732,10.192734,10.357354,11.218181,10.902658,10.456812,10.528833,11.105004,11.526843,12.421966,13.629181,14.534592,15.069608,15.724659,15.110763,13.670336,12.97413,13.317088,13.708061,13.375391,12.88496,12.6586075,12.651748,12.370522,12.240198,11.499407,10.984968,10.912948,10.88551,10.604284,10.738038,10.861504,11.002116,11.622872,12.30536,13.296511,13.88983,13.9138365,13.725209,13.749216,12.943263,12.572867,13.046151,13.900118,14.38369,14.685493,14.757515,14.699212,14.778092,14.983868,15.326826,15.494876,15.3817,15.097044,14.613472,14.726648,15.46744,16.54433,17.346853,18.79414,19.480057,20.742146,22.762173,24.583282,29.43615,37.98268,37.82492,29.782537,27.909983,23.76361,23.835632,20.817596,14.160767,10.065839,10.508256,11.605724,10.89237,10.978109,19.524641,23.52354,13.972139,4.773986,1.4404267,1.1008976,1.2072148,0.88826317,0.7922347,1.0425946,1.255229,2.0268862,2.4795918,3.1209247,4.249259,5.9160385,5.830299,7.0615206,8.611694,10.065839,11.592006,12.569438,12.699762,12.46998,12.3533745,12.79922,12.55229,12.476839,12.88839,13.684054,14.345964,15.536031,16.355703,17.2131,17.895588,17.573206,17.53891,17.799559,17.761833,17.511473,17.799559,17.28169,17.137648,16.918156,16.441442,15.7966795,15.361122,14.850114,14.514014,14.335675,14.040731,14.496866,14.177915,13.855534,13.7697935,13.63261,13.22106,13.22106,13.371962,13.529722,13.677195,13.581166,12.915827,12.466551,12.415107,12.312219,11.413667,11.177026,11.231899,11.547421,12.445972,12.572867,12.205902,11.441104,10.456812,9.537683,9.647429,9.421077,9.3079,9.448513,9.650859,9.72631,9.290752,9.081548,9.273604,9.458802,9.983529,9.589127,8.858624,8.196714,7.8537555,8.131552,7.9943686,7.599966,7.0923867,6.5985265,6.478491,6.324159,6.2075534,6.0875177,5.796003,5.892031,5.9400454,5.967482,6.0086374,6.111525,6.279575,6.3207297,6.5813785,7.016936,7.1987042,6.944915,6.9620624,6.948344,7.0306544,7.7680154,7.98065,7.81603,7.7440085,7.7851634,7.531374,7.3839016,7.0786686,6.914048,6.9723516,7.1266828,6.927767,7.006647,7.0718093,7.239859,8.008087,8.011517,7.490219,6.9860697,6.7048435,6.5127864,6.989499,7.4181976,7.8194594,8.2310095,8.721441,8.683716,8.405919,8.423067,8.858624,9.39021,9.582268,10.2236,11.238758,12.21619,12.394529,12.569438,12.624311,12.586586,12.439114,12.113303,11.917816,11.55771,11.067279,10.700313,10.9541025,11.231899,11.262765,11.461681,12.140739,13.505715,14.575747,15.470869,16.143068,16.462019,16.21509,16.61292,17.007324,17.442883,17.816708,17.885298,19.301718,20.827885,20.03222,17.117071,14.942713,15.162207,15.059319,15.093615,15.522313,16.393429,15.9613,15.402277,14.589465,13.810948,13.80066,14.150477,14.424845,14.668345,14.990726,15.590904,16.516893,17.439453,17.7927,17.700102,17.974468,17.936743,17.106783,16.232237,15.638919,15.22051,14.970149,14.887839,15.343974,16.13621,16.496315,15.522313,13.845244,12.511135,12.185325,13.118172,13.848674,14.874121,15.481158,15.786391,16.743246,16.780972,16.70552,16.63007,16.55119,16.355703,16.321407,15.954441,16.143068,16.489456,15.319967,13.992717,12.987847,11.80121,10.686595,10.669447,8.093826,5.3261495,5.5662203,7.3873315,4.7534084,4.091498,19.826445,20.004784,3.9611735,2.287535,3.5976372,3.8925817,4.4756117,5.4016004,5.470192,10.463672,13.080446,14.38026,13.680624,8.532814,5.857735,3.724532,5.586798,10.439664,12.816368,19.185112,18.338005,16.918156,16.479168,13.516005,15.659496,13.365103,9.952662,7.490219,6.7802944,5.219832,5.645101,7.0306544,8.110974,7.377043,4.9214582,4.3349986,4.355576,4.9934793,7.548522,6.584808,6.183546,6.7940125,8.2310095,9.674867,8.954653,8.467651,8.755736,9.534253,9.668007,10.858074,11.4205265,11.876661,12.21619,11.88352,11.646879,11.321068,10.72775,10.192734,10.573419,11.2250395,12.127021,13.111313,13.893259,14.071597,13.344524,13.4645605,14.668345,16.513464,17.87158,17.748116,18.231688,17.940172,17.058767,17.333136,17.37772,18.770132,20.522652,21.921923,22.52553,21.318316,19.661825,19.329155,20.11453,19.833303,17.923023,15.9578705,13.958421,12.528283,12.881531,13.344524,13.762935,14.064738,14.2533655,14.387119,15.316538,14.760944,13.876111,13.183334,12.576297,12.199042,12.195613,13.049581,14.527733,15.693792,16.023033,16.424294,16.359133,15.707511,14.79524,13.63604,13.7526455,14.417986,15.645778,18.190533,17.223389,15.3302555,13.440554,12.394529,12.950122,13.265644,12.9809885,13.097594,13.80066,14.455711,13.063298,12.017275,11.492548,11.327928,11.046701,9.870353,9.235879,8.9100685,8.519095,7.5588107,7.3358874,7.3290286,7.3393173,7.332458,7.455923,7.517656,7.9875093,8.536243,8.995808,9.362774,9.633711,9.760606,9.949233,10.288762,10.751757,11.077567,11.135871,10.923236,10.587136,10.429376,10.755186,10.696883,10.419086,9.9801,9.321619,9.211872,8.999237,8.604835,8.028665,7.3358874,0.5041494,0.48014224,0.5178677,0.61046654,0.6790583,0.59674823,0.59674823,0.5693115,0.53844523,0.5144381,0.5041494,0.45613512,0.48014224,0.5453044,0.61389613,0.6241849,0.8196714,0.7888051,0.7339317,0.7305021,0.71678376,0.6927767,0.7888051,0.91569984,0.9602845,0.77851635,0.70649505,0.6310441,0.58988905,0.5796003,0.5796003,0.9568549,0.9328478,0.7888051,0.67219913,0.61046654,0.6824879,0.9294182,1.0528834,1.0528834,1.2346514,1.2243627,1.0734608,0.90198153,0.77851635,0.71678376,0.7888051,0.8162418,0.78194594,0.70649505,0.65505123,0.7305021,0.7099246,0.7339317,0.8162418,0.84024894,0.75450927,0.65162164,0.59674823,0.61389613,0.6859175,0.58988905,0.5178677,0.39783216,0.2469303,0.19891608,0.18519773,0.1371835,0.15090185,0.29837412,0.64133286,0.5693115,0.45613512,0.29151493,0.11317638,0.01371835,0.0034295875,0.0,0.0,0.030866288,0.15090185,0.07888051,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.106317215,0.034295876,0.024007112,0.12346515,0.29151493,0.42869842,0.8676856,0.9568549,0.7990939,0.9362774,2.3664153,1.3992717,0.8676856,0.4698535,0.15090185,0.07545093,0.1371835,0.07888051,0.13375391,0.23664154,0.01371835,0.0034295875,0.010288762,0.058302987,0.116605975,0.09259886,0.16462019,0.22978236,0.3018037,0.33609957,0.21263443,0.4938606,0.34638834,0.37039545,0.5007198,0.0,0.31895164,0.48014224,0.7888051,1.0734608,0.67219913,0.84367853,0.5178677,0.28808534,0.29494452,0.26064864,0.48014224,0.30523327,0.22635277,0.32238123,0.274367,0.28808534,0.2709374,0.34981793,0.4938606,0.5178677,0.59331864,0.4629943,0.42869842,0.51100856,0.47328308,0.51100856,0.37382504,0.32238123,0.37725464,0.30523327,0.28122616,0.1920569,0.22978236,0.36696586,0.36696586,0.31895164,0.45956472,0.6379033,0.78537554,0.9294182,0.7099246,0.8196714,0.91912943,0.89855194,0.8848336,1.1180456,1.2209331,1.1729189,1.08032,1.1900668,1.1180456,1.1900668,1.1900668,1.1214751,1.2209331,1.2586586,1.3478279,1.3992717,1.4267083,1.5707511,1.7799559,2.369845,2.8465576,3.0626216,3.234101,3.4055803,3.841138,4.184097,4.338428,4.4859004,4.413879,4.972902,5.7651367,6.4990683,6.989499,6.989499,6.8969,6.9346256,7.1061053,7.2158523,7.9875093,8.827758,9.366203,9.472521,9.277034,9.266746,9.407358,9.932085,10.696883,11.183885,11.465111,12.130451,12.620882,12.723769,12.590015,12.394529,11.849225,11.619442,11.766914,11.780633,11.732618,11.691463,11.526843,11.444533,11.993267,11.626302,10.63858,9.89436,9.750318,10.055551,9.921797,10.206452,10.367643,10.353925,10.635151,11.502836,12.788932,13.7526455,14.201921,14.496866,14.555169,13.996146,13.519434,13.594885,14.448852,14.863832,15.031882,15.138199,15.268523,15.426285,14.973578,15.237658,15.340545,15.0250225,14.634049,13.924125,14.225929,15.22051,16.588915,18.005335,19.092514,19.408035,21.174273,24.154585,25.680752,29.648783,36.75489,36.370773,29.535606,28.959436,20.378609,17.072487,14.263655,10.686595,8.573969,10.151579,9.767465,9.630281,12.932974,23.832203,18.770132,10.683165,4.338428,1.6016173,1.4198492,0.8711152,0.9534253,1.4644338,2.0097382,1.9994495,2.1091962,2.2463799,2.8328393,3.9886103,5.5387836,6.125243,7.7714453,8.882631,9.297611,10.299051,11.019264,11.8869505,12.428825,12.566009,12.603734,12.202472,11.924676,11.616013,11.588576,12.648318,13.272504,14.829536,16.311117,17.182234,17.364002,17.63151,18.094503,18.430603,18.509483,18.386019,17.21653,17.837284,18.20425,17.676094,17.027903,16.46888,16.033321,15.54632,15.079896,14.970149,16.029892,15.995596,15.824117,15.693792,14.997586,14.791811,15.042171,15.261664,15.083325,14.2533655,14.068168,13.766364,13.529722,13.279363,12.679185,12.178465,12.264205,12.5145645,12.737488,12.9707,12.7272,12.034423,11.177026,10.367643,9.719451,10.182446,10.336777,10.288762,10.100135,9.794902,10.089847,9.925226,9.424506,8.81061,8.4093485,8.934075,9.009526,8.790032,8.450503,8.193284,8.378482,8.186425,7.8674736,7.514226,7.051232,6.550512,6.094377,5.717122,5.40503,5.1100855,5.3570156,5.381023,5.3432975,5.3913116,5.662249,6.101236,6.210983,6.385892,6.7219915,7.0032177,6.9071894,6.910619,7.0375133,7.2158523,7.2775846,7.864044,7.6171136,7.390761,7.3255987,6.835168,6.9689217,6.7665763,6.625963,6.636252,6.5779486,6.125243,6.166398,6.3618846,6.6533995,7.2638664,7.6651278,7.3564653,6.914048,6.6465406,6.560801,7.133542,7.407909,7.6274023,8.014946,8.759167,8.964942,8.834618,8.906639,9.071259,8.56025,9.122703,10.261326,11.317638,12.0138445,12.466551,12.857523,12.788932,12.535142,12.147599,11.489118,11.684605,11.688034,11.664027,11.612583,11.369082,11.30735,11.262765,11.574858,12.332796,13.38225,14.5414505,15.9578705,17.141079,17.741257,17.532051,17.326277,16.815268,16.993607,17.899017,18.629519,19.301718,21.356041,21.644127,19.384027,16.173935,15.138199,15.765814,16.571766,16.722668,16.0539,14.867262,14.7369375,14.321958,13.409687,12.908967,13.004995,13.670336,14.750656,15.810398,16.12935,17.141079,18.355152,18.77699,18.241976,17.425734,17.37772,16.6335,15.88242,15.553179,15.806969,16.163645,15.755525,15.810398,16.45859,16.739817,16.225378,15.110763,13.773223,12.826657,13.107883,14.596324,15.902997,16.444872,16.643787,17.912735,18.646667,18.773561,18.591793,18.173384,17.38115,17.806417,17.072487,16.907866,17.909306,19.5315,19.054789,17.250826,15.584045,14.771234,14.771234,5.456474,2.8808534,3.5599117,4.5099077,3.2649672,4.5956473,4.729401,3.069481,0.83681935,1.0666018,4.437886,5.223262,4.650521,4.0023284,4.6402316,6.018926,8.303031,11.228469,12.30536,6.835168,4.6402316,3.4021509,5.90575,9.277034,5.003768,13.111313,16.13621,16.935303,15.896138,10.940384,13.649758,14.970149,12.147599,7.5759587,8.759167,7.2947326,6.7631464,6.0806584,5.2164025,5.2026844,2.9940298,3.457024,4.5030484,5.120374,5.4016004,5.8543057,6.4407654,7.3221693,8.429926,9.489669,8.038953,8.042382,9.201583,10.497967,10.192734,11.266195,11.7086115,12.428825,13.347955,13.395968,12.895248,13.128461,12.542002,11.441104,11.979549,12.895248,13.149038,13.797231,14.644339,14.267084,14.095605,14.390549,15.117621,16.077906,16.907866,16.527182,17.110212,16.976458,16.503176,18.1288,19.517782,20.845032,22.28546,23.146286,21.86705,20.522652,19.637817,19.435472,19.589804,19.21255,18.588364,16.499744,14.743796,14.030442,13.992717,14.150477,14.904987,15.179354,14.7026415,14.006435,14.7026415,14.712931,14.805529,14.774663,13.443983,12.771784,11.677745,12.113303,14.009865,15.306249,15.6697855,15.642348,14.527733,13.512574,15.6869335,16.050468,16.80155,16.7844,16.081335,16.005884,17.021042,16.311117,14.407697,12.483699,12.373952,12.840376,12.672326,12.644889,13.063298,13.749216,13.419975,12.531713,11.780633,11.4754,11.537132,10.340206,9.434795,8.628842,7.8023114,6.910619,6.5710897,6.584808,6.975781,7.56567,7.98065,8.052671,8.512236,9.006097,9.458802,10.069269,10.840926,11.039842,11.492548,12.106443,11.8869505,12.144169,12.106443,11.753197,11.334786,11.382801,11.592006,11.485688,10.960961,10.100135,9.184435,8.296172,7.8434668,7.6342616,7.3598948,6.591667,0.5144381,0.5007198,0.4698535,0.44927597,0.4424168,0.4355576,0.61046654,0.7099246,0.6241849,0.45270553,0.48014224,0.58645946,0.5761707,0.5418748,0.5418748,0.61389613,0.90541106,0.90541106,0.78537554,0.66533995,0.59674823,0.5212973,0.5590228,0.6001778,0.61389613,0.64476246,0.65848076,0.59331864,0.59331864,0.65848076,0.6276145,0.75450927,0.67219913,0.6241849,0.66191036,0.65848076,0.7922347,0.89855194,1.0048691,1.1214751,1.2346514,1.155771,1.0460242,0.939707,0.8505377,0.7888051,0.78537554,0.7339317,0.6927767,0.7133542,0.84024894,0.9328478,0.9568549,0.96371406,0.9568549,0.864256,0.7579388,0.7099246,0.65505123,0.607037,0.65162164,0.53158605,0.4355576,0.33266997,0.2503599,0.26064864,0.20920484,0.20920484,0.4115505,0.7133542,0.7510797,1.155771,1.1660597,0.70306545,0.082310095,0.0034295875,0.0,0.0,0.0,0.006859175,0.030866288,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.06516216,0.034295876,0.048014224,0.18176813,0.4629943,0.5212973,0.67219913,1.0837497,1.5913286,1.6804979,1.1763484,0.6241849,0.25378948,0.116605975,0.11317638,0.07545093,0.1097468,0.11317638,0.058302987,0.01371835,0.01371835,0.01371835,0.061732575,0.17147937,0.32238123,0.5727411,0.432128,0.4355576,0.6001778,0.42183927,0.53501564,0.5212973,0.5590228,0.6207553,0.45270553,0.48700142,0.5555932,0.7922347,1.0151579,0.72021335,0.66533995,0.65162164,0.5418748,0.42183927,0.58988905,0.31895164,0.15776102,0.16119061,0.25721905,0.23664154,0.24007112,0.31209245,0.34981793,0.34295875,0.34638834,0.45956472,0.45270553,0.37725464,0.3566771,0.58302987,0.45270553,0.274367,0.274367,0.39097297,0.26750782,0.29151493,0.20234565,0.18862732,0.26064864,0.23321195,0.2709374,0.4664239,0.5418748,0.48700142,0.5658819,0.65848076,0.70649505,0.7305021,0.77851635,0.922559,1.0151579,1.0563129,1.0220171,1.0254467,1.313532,1.4232788,1.5090185,1.4575747,1.313532,1.2449403,1.3101025,1.3821237,1.4335675,1.4781522,1.546744,1.6873571,1.9754424,2.352697,2.7368107,3.0146074,3.1072063,3.2032347,3.5118976,4.0229063,4.5099077,4.897451,5.1238036,5.446185,5.9160385,6.355026,6.540223,6.451054,6.433906,6.5642304,6.6568294,7.1712675,7.606825,7.864044,7.9189177,7.798882,7.689135,8.23444,8.680285,9.023245,10.000677,11.080997,11.14273,10.912948,10.792912,10.844356,10.813489,10.628291,10.364213,9.9801,9.290752,9.661148,9.644,9.801761,10.316199,10.991828,10.840926,10.374502,10.010965,9.925226,10.041832,9.897789,9.9801,10.072699,10.230459,10.744898,11.825217,12.905538,13.834956,14.448852,14.555169,14.4317045,14.126471,13.872682,13.841815,14.119612,14.712931,15.158776,15.309678,15.127911,14.668345,15.165636,15.782962,16.269962,16.554619,16.719238,15.680074,16.03675,16.664366,17.357141,18.811287,19.95677,19.94305,21.657845,24.651875,25.142305,31.980904,40.414257,40.249638,32.220974,27.995722,17.463459,11.996697,10.374502,9.990388,6.8557453,7.6959944,8.097256,13.430264,22.316326,26.606739,14.928994,7.2021337,2.9494452,1.3443983,1.2106444,1.3958421,1.2209331,1.1763484,1.4232788,1.7902447,2.0268862,2.6064866,3.5153272,4.5922174,5.5250654,7.596536,8.934075,9.534253,10.000677,11.55771,11.612583,12.298501,12.823228,12.80265,12.260776,12.006986,11.8115,11.910957,12.418536,13.334236,14.064738,14.846684,15.892709,16.911295,17.134218,17.741257,18.427174,18.759844,18.680964,18.509483,17.679523,18.02934,18.608942,18.917604,18.897026,18.608942,18.420315,18.135658,17.748116,17.436022,17.597214,17.586924,18.187103,17.923023,13.046151,14.802099,15.724659,16.191082,16.21166,15.46058,14.856973,14.390549,13.982429,13.454271,12.535142,12.072148,12.151029,12.504276,13.032433,13.80066,13.049581,12.075578,11.478829,11.255906,10.792912,10.7586155,10.940384,11.118723,11.194174,11.201033,10.906088,9.9869585,9.009526,8.241299,7.6616983,7.8263187,8.1212635,8.2310095,8.158989,8.193284,8.299602,8.292743,7.8983397,7.2878733,7.085528,6.6431108,6.1458206,5.552502,4.972902,4.6608095,4.7979927,5.1100855,5.394741,5.5902276,5.7719955,5.9469047,6.036074,6.2555676,6.4887795,6.2727156,6.526505,6.5642304,6.667118,6.883182,7.023795,7.4113383,7.291303,7.15069,7.1129646,6.944915,6.9037595,7.1026754,7.31531,7.3290286,6.9552035,6.893471,6.776865,6.7974424,7.023795,7.4113383,7.939495,7.73372,7.3393173,7.0272245,6.8043017,7.085528,7.298162,7.5382333,7.8091707,8.025234,8.117833,8.388771,8.632272,8.718011,8.584257,8.951223,9.97324,11.105004,11.989838,12.490558,12.617453,12.696333,12.72034,12.507706,11.72233,11.72233,12.175035,12.439114,12.415107,12.55229,12.754636,12.617453,12.600305,13.004995,13.96871,15.069608,16.170506,17.384579,18.386019,18.410025,18.674105,18.338005,18.163095,18.259123,18.094503,18.11165,20.975357,21.057667,17.322845,13.330807,12.936404,12.202472,12.109874,12.936404,14.246507,13.05301,12.603734,12.699762,12.871242,12.360233,12.926115,14.140189,15.896138,17.669235,18.533491,18.38259,18.656956,19.253704,19.709839,19.1954,18.091074,17.134218,16.393429,15.940722,15.844694,16.393429,16.46888,16.78783,17.28169,17.093063,16.47231,15.481158,14.352823,13.409687,13.094165,14.174485,15.758954,16.736387,17.168514,18.293419,18.564358,19.092514,19.027351,18.28313,17.53891,18.091074,18.019053,17.754974,17.669235,18.053349,18.485476,18.132229,16.822126,15.405707,15.748666,11.1393,7.449064,7.500508,9.259886,5.8165803,5.1340923,3.9371665,2.901431,2.5996273,3.4981792,3.9165888,4.496189,3.875434,2.819121,4.187526,3.9440255,7.4970784,9.932085,9.407358,7.140401,3.9954693,4.383013,8.244728,12.607163,11.595435,16.832415,12.984418,8.940934,8.31332,9.451943,10.676306,10.48082,9.818909,10.055551,12.956982,12.370522,9.993818,7.4010496,5.597087,5.007198,3.9714622,3.4878905,4.40702,5.7377,4.681387,5.593657,6.3035817,6.824879,7.291303,7.953213,7.9463544,8.858624,9.719451,10.100135,10.106995,11.074138,12.55915,13.9138365,14.79867,15.179354,14.472859,14.970149,14.544881,13.073587,12.428825,14.037301,14.953001,15.206791,14.956431,14.46257,15.326826,15.361122,15.488017,15.985307,16.503176,16.654078,16.94902,17.075916,17.250826,18.248835,19.805868,21.102251,21.973368,21.85676,19.802439,18.187103,17.562918,17.658945,18.338005,19.589804,18.663815,16.098484,14.565458,14.596324,14.579176,15.086755,15.659496,16.420864,16.846134,15.741806,15.556609,15.1862135,15.100473,15.391989,15.748666,15.978448,14.5243025,13.443983,13.694343,15.145059,16.79126,17.141079,15.889278,14.466,16.0539,17.1205,18.084215,18.646667,18.687822,18.252264,18.015623,16.739817,15.172495,13.7526455,12.617453,12.878101,13.509145,13.786942,13.395968,12.428825,12.178465,11.279913,10.882081,11.194174,11.499407,10.401938,9.455373,8.663138,7.9772205,7.291303,6.615674,6.667118,7.06495,7.599966,8.200144,8.525954,8.800322,9.194724,9.866923,10.9369545,11.921246,12.277924,12.363663,12.356804,12.264205,12.178465,12.284782,12.46312,12.507706,12.116733,12.089295,11.742908,10.789482,9.342196,7.9292064,7.514226,7.2707253,7.3221693,7.377043,6.725421,0.34638834,0.32581082,0.28122616,0.26407823,0.29494452,0.36010668,0.41840968,0.4629943,0.432128,0.36353627,0.4081209,0.4389872,0.44584638,0.4629943,0.50757897,0.59331864,0.6962063,0.64476246,0.6241849,0.6310441,0.4629943,0.5761707,0.5555932,0.50757897,0.5212973,0.66533995,0.70306545,0.6173257,0.5693115,0.58645946,0.5590228,0.7133542,0.66533995,0.6001778,0.58988905,0.58988905,0.70649505,0.83338976,0.939707,1.0288762,1.1351935,1.0082988,1.0082988,0.9294182,0.7990939,0.85396725,0.823101,0.8128122,0.8505377,0.91569984,0.939707,0.9945804,1.0048691,1.0151579,1.0117283,0.9259886,0.77165717,0.65162164,0.5590228,0.52472687,0.6036074,0.45956472,0.39440256,0.33952916,0.30866286,0.3841138,0.29494452,0.607037,0.90541106,1.0906088,1.3924125,3.4776018,3.1209247,1.5501735,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.0274367,0.017147938,0.07545093,0.25378948,0.30523327,0.5007198,0.91569984,1.2723769,0.97057325,0.72707254,0.34981793,0.106317215,0.05144381,0.048014224,0.037725464,0.0548734,0.041155048,0.006859175,0.006859175,0.006859175,0.034295876,0.08916927,0.2469303,0.64819205,0.823101,0.52815646,0.34295875,0.4424168,0.6276145,0.48357183,0.50757897,0.6756287,0.77851635,0.4081209,0.42526886,0.4938606,0.7373613,1.0117283,0.89855194,1.08032,0.9602845,0.6790583,0.42526886,0.432128,0.2469303,0.24007112,0.22978236,0.16804978,0.15433143,0.16462019,0.2503599,0.29151493,0.274367,0.30523327,0.31895164,0.3566771,0.34295875,0.32924038,0.48357183,0.4355576,0.36010668,0.33266997,0.33952916,0.2777966,0.37382504,0.23664154,0.16462019,0.21263443,0.18862732,0.20577525,0.33609957,0.42183927,0.45270553,0.5658819,0.64819205,0.6276145,0.5796003,0.6036074,0.8025235,0.805953,0.90884066,1.0117283,1.1180456,1.3238207,1.4541451,1.5261664,1.4575747,1.3786942,1.6256244,1.5913286,1.5947582,1.6530612,1.7353712,1.7593783,2.037175,2.2292318,2.4624438,2.7882545,3.1792276,3.3129816,3.2855449,3.3609958,3.6696587,4.214963,4.8322887,5.055212,5.254128,5.562791,5.8645945,6.433906,6.5059276,6.3618846,6.23156,6.2864337,6.540223,6.680836,6.8591747,7.0615206,7.1095347,7.058091,7.4456344,7.9086285,8.405919,9.211872,10.39508,10.47396,10.189304,9.908078,9.609704,9.9801,10.062409,9.836057,9.314759,8.519095,9.523964,9.822338,10.014396,10.353925,10.762046,10.984968,11.043272,11.029553,10.967821,10.799771,10.703742,10.779194,10.679735,10.569988,11.129011,11.897239,12.826657,13.687484,14.212211,14.105893,13.920695,13.886399,13.591455,13.282792,13.855534,14.805529,15.498305,15.899568,16.064188,16.12935,16.393429,16.750105,17.151367,17.607502,18.176813,17.580065,17.79613,18.152807,18.687822,20.138538,21.489796,22.501524,24.4461,26.483274,25.660173,34.971504,41.07274,40.290794,34.052376,28.890844,16.726099,10.028113,9.328478,11.0981455,7.740579,8.460793,8.724871,14.044161,21.575535,20.104242,9.592556,4.2115335,2.568761,2.4967396,1.0494537,1.0048691,0.9328478,1.1454822,1.8828435,3.3129816,3.9851806,4.5442033,5.1821065,5.9640527,6.831738,8.899779,10.456812,11.660598,12.576297,13.179905,12.682614,12.895248,13.193623,13.337666,13.502286,13.402828,13.810948,14.267084,14.562028,14.757515,15.536031,15.885849,15.995596,16.307688,17.504614,17.799559,18.005335,18.104792,18.303709,19.044498,18.818146,18.355152,18.499195,19.339443,20.21399,20.923914,20.272291,19.70641,19.661825,19.54179,18.821575,18.70154,17.580065,14.891269,11.101575,11.444533,12.939834,14.29795,15.021593,15.388559,14.891269,14.733508,14.448852,13.862392,13.118172,12.932974,13.214201,13.536582,13.862392,14.538021,14.04759,13.22106,12.843805,12.860953,12.370522,11.691463,11.664027,11.585147,11.204462,10.72775,9.818909,9.246168,8.663138,8.100685,7.9909387,7.8503256,7.7783046,7.7885933,7.8606143,7.9086285,8.1041155,8.025234,7.8366075,7.623973,7.3873315,6.8591747,6.39961,5.8543057,5.271276,4.90431,5.0586414,5.3501563,5.65539,5.8474464,5.778855,5.6999745,5.6039457,5.658819,5.874883,6.0978065,6.5127864,6.385892,6.228131,6.2212715,6.2247014,6.5024977,6.7974424,6.999788,7.1849856,7.6033955,7.4970784,7.4456344,7.4044795,7.377043,7.425057,7.1987042,6.7494283,6.6122446,6.883182,7.2364297,7.73029,7.8434668,7.682276,7.3255987,6.8111606,6.8591747,6.927767,7.174697,7.4284863,7.1849856,7.3118806,7.6651278,8.097256,8.457363,8.628842,8.687145,9.445084,10.340206,11.129011,11.845795,12.487128,12.63117,12.699762,12.662037,12.034423,12.127021,12.373952,12.404818,12.336226,12.764925,12.991278,13.05301,12.977559,13.066729,13.903547,15.004445,15.738377,16.54776,17.439453,18.008764,18.320856,18.005335,17.826996,18.084215,18.602083,18.056778,20.587814,20.11453,16.955881,17.799559,11.80464,8.707723,7.298162,6.9517736,7.613684,7.6274023,7.840037,8.224151,8.855195,9.914937,11.622872,13.330807,15.412566,17.70696,19.52807,19.922474,19.949911,20.107672,20.310017,19.884748,19.397747,18.550638,17.511473,16.695232,16.760393,16.88386,17.12736,17.326277,17.29884,16.859852,16.763824,15.580616,14.284232,13.402828,13.018714,14.009865,15.419425,16.619781,17.422304,18.073925,18.190533,18.821575,18.989626,18.54378,18.156237,18.197392,18.708399,18.907316,18.653526,18.46147,19.517782,19.582945,18.12537,15.896138,14.901558,12.569438,10.093276,9.095266,8.827758,6.1629686,3.2409601,2.6887965,3.2855449,4.3590055,5.778855,5.0449233,4.1292233,4.3349986,5.456474,5.813151,4.1772375,8.522525,9.863494,6.852316,5.751418,2.4967396,6.0840883,8.851766,8.783174,9.510246,11.338216,8.309891,5.178677,4.5922174,7.0923867,7.720001,6.9071894,6.245279,6.9792104,10.024684,11.204462,11.454823,9.692014,6.8111606,5.693115,4.976331,4.616225,4.65395,4.866585,4.7945633,5.3570156,5.6656785,6.0635104,6.728851,7.6788464,8.032094,8.625413,8.927217,8.98209,9.39021,9.962952,11.4205265,13.107883,14.472859,15.083325,15.148488,15.673215,15.46058,14.342535,13.183334,15.676644,16.283682,15.88242,15.258235,15.114192,16.420864,16.811838,16.70895,16.582056,16.925014,16.311117,16.160215,15.927004,15.920145,17.326277,18.972477,20.11453,20.978786,21.236006,20.028791,17.346853,17.117071,17.79613,18.499195,18.989626,20.131678,17.412016,14.994157,14.445422,14.723219,14.435134,14.994157,16.273392,17.758404,18.526632,17.809847,16.496315,15.415996,15.172495,16.153357,17.638369,17.147938,15.8138275,14.870691,15.656067,16.479168,17.062197,16.86671,16.383139,17.113642,16.997036,17.473747,17.86815,17.607502,16.232237,15.193072,14.249936,13.780083,13.684054,13.38568,13.056439,13.430264,13.920695,13.80066,12.202472,11.763485,11.080997,10.837497,11.087856,11.269625,10.487679,9.688584,8.951223,8.23444,7.4044795,6.931196,6.824879,6.90033,7.1952744,7.98065,8.289313,8.519095,8.872343,9.650859,11.235329,12.229909,12.782072,12.555719,11.581717,10.254466,10.024684,10.041832,10.666017,11.629731,12.0138445,11.952112,11.211322,10.021255,8.666568,7.4936485,7.363324,7.205563,7.421627,7.7714453,7.390761,0.216064,0.20577525,0.18176813,0.18176813,0.2194936,0.29151493,0.26407823,0.28122616,0.30866286,0.32924038,0.34638834,0.3566771,0.37382504,0.4081209,0.45613512,0.5178677,0.4972902,0.44584638,0.5178677,0.6379033,0.50757897,0.5761707,0.5796003,0.5521636,0.5453044,0.64819205,0.66533995,0.5658819,0.5212973,0.5453044,0.48357183,0.59674823,0.5727411,0.53844523,0.53158605,0.5144381,0.61389613,0.7442205,0.805953,0.8025235,0.8745448,0.805953,0.8711152,0.8196714,0.69963586,0.8471081,0.8162418,0.82996017,0.90198153,0.9842916,0.9568549,0.9568549,0.91912943,0.91912943,0.939707,0.864256,0.6962063,0.5453044,0.4698535,0.47328308,0.53158605,0.42526886,0.39097297,0.39783216,0.44584638,0.5727411,0.72364295,1.1934965,1.4369972,1.5090185,2.0577524,5.4976287,4.2218223,1.7216529,0.082310095,0.0,0.020577524,0.010288762,0.0,0.006859175,0.037725464,0.07545093,0.0548734,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.01371835,0.017147938,0.010288762,0.01371835,0.07545093,0.42869842,0.47671264,0.7305021,1.0082988,0.42183927,0.30866286,0.14061308,0.034295876,0.01371835,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.030866288,0.07545093,0.22292319,0.4938606,0.83681935,0.8162418,0.5144381,0.30523327,0.36353627,0.66533995,0.4081209,0.39097297,0.5658819,0.6962063,0.35324752,0.29151493,0.432128,0.72707254,0.97057325,0.8162418,1.1146159,1.0048691,0.7682276,0.5418748,0.36010668,0.22978236,0.26064864,0.28808534,0.2469303,0.18519773,0.16804978,0.26407823,0.28808534,0.22978236,0.26407823,0.18519773,0.24007112,0.2709374,0.26407823,0.33609957,0.38754338,0.33266997,0.28808534,0.2709374,0.20920484,0.32581082,0.21263443,0.14061308,0.17833854,0.17833854,0.22292319,0.26750782,0.31895164,0.40126175,0.5521636,0.5178677,0.5624523,0.59331864,0.6207553,0.7613684,0.7339317,0.83338976,0.94999576,1.0528834,1.1832076,1.3924125,1.4267083,1.3821237,1.4129901,1.7353712,1.704505,1.7079345,1.8313997,1.978872,1.8965619,2.2086544,2.335549,2.503599,2.8019729,3.1552205,3.2443898,3.2066643,3.1312134,3.2032347,3.707384,4.3692946,4.756838,5.0449233,5.295283,5.4633327,6.0497923,6.307011,6.2555676,6.0566516,5.9983487,5.809721,5.8680243,6.0497923,6.2487082,6.385892,6.5539417,6.948344,7.5690994,8.309891,8.961512,9.860064,10.065839,9.918367,9.599416,9.122703,9.561689,9.647429,9.445084,9.122703,8.961512,10.124143,10.576848,10.786053,10.984968,11.156448,11.502836,11.629731,11.619442,11.595435,11.7086115,11.842365,11.808069,11.698323,11.674315,11.979549,12.332796,13.025573,13.594885,13.858963,13.917266,13.725209,13.7697935,13.564018,13.358243,14.13676,15.402277,16.105343,16.691803,17.29198,17.720678,17.864721,18.190533,18.533491,18.989626,19.915615,19.929333,20.262003,20.52951,20.855322,21.87048,23.211449,24.895376,26.76107,27.872257,26.531288,36.56969,41.07274,42.90757,41.371113,32.196968,17.909306,10.542552,9.650859,11.495977,9.043822,9.14328,8.937505,12.3533745,16.606062,12.178465,5.4941993,2.7470996,2.843128,3.4947495,1.2277923,1.0014396,0.9568549,1.1934965,1.8554068,3.1072063,4.0949273,4.99005,5.693115,6.392751,7.582818,9.115844,11.2593355,13.111313,14.109323,14.016724,13.529722,13.337666,13.272504,13.433694,14.198492,14.417986,15.37827,16.252815,16.595774,16.331696,16.856422,17.161655,17.189093,17.271402,18.139088,18.217968,18.187103,18.351723,18.965618,20.234566,20.505503,19.973917,20.001354,20.759293,21.222288,21.808746,20.958208,20.395756,20.591244,20.728426,20.505503,20.930773,18.37573,13.509145,11.303921,10.55284,11.180455,11.849225,12.325937,13.481709,13.855534,14.054449,13.958421,13.687484,13.63261,13.728639,13.934414,14.188204,14.435134,14.637479,14.308239,13.944703,13.865822,13.896688,13.402828,12.644889,12.343085,11.718901,10.714031,9.959522,9.030104,8.779744,8.495089,8.086967,8.100685,7.9737906,7.658269,7.5039372,7.5759587,7.658269,7.963502,8.069819,8.207003,8.289313,7.9017696,7.133542,6.7494283,6.4373355,6.1046658,5.885172,5.844017,5.9400454,6.025785,5.9434752,5.5422134,5.470192,5.353586,5.31929,5.48734,5.9640527,6.276145,6.2041235,6.1321025,6.159539,6.108095,6.3035817,6.526505,6.636252,6.7322803,7.14726,7.226141,7.291303,7.191845,7.0718093,7.3839016,7.222711,6.869464,6.7322803,6.869464,6.9860697,7.5553813,7.8537555,7.8194594,7.507367,7.0615206,6.7631464,6.6533995,6.7802944,6.931196,6.636252,6.776865,7.1266828,7.781734,8.515666,8.793462,8.776315,9.352485,10.017825,10.593996,11.2421875,12.055,12.370522,12.6586075,12.926115,12.713481,12.627741,12.79922,12.836946,12.778643,13.083877,13.210771,13.13189,12.984418,13.046151,13.725209,14.592895,14.977009,15.347404,15.927004,16.702091,17.343424,17.343424,17.086205,16.983316,17.501184,17.007324,19.133669,19.497204,18.3723,20.656404,11.238758,6.667118,4.695105,3.9303071,3.8377085,3.4433057,4.7019644,6.334448,7.7714453,9.139851,11.303921,13.207341,15.162207,17.079346,18.495766,19.775002,20.70099,21.0268,20.851892,20.594673,20.52951,19.823015,18.70497,17.63151,17.29884,17.003895,17.178804,17.271402,17.055338,16.616352,17.1205,15.913286,14.363112,13.238208,12.730629,14.020154,15.536031,16.96274,17.87158,17.71039,17.566347,17.809847,18.022482,18.084215,18.187103,18.118511,18.831865,19.507494,19.819586,19.922474,20.958208,20.642687,19.137098,17.089634,15.6526375,14.325387,12.63117,10.696883,8.759167,7.160979,4.139512,3.093488,3.3198407,4.355576,5.9812007,6.40304,4.972902,5.212973,6.9826403,6.492209,6.193835,9.414218,8.824328,4.7088237,4.9831905,2.0886188,4.7842746,6.5779486,6.3378778,8.299602,5.874883,4.2183924,3.1483612,2.9940298,4.5956473,5.994919,7.016936,6.2487082,5.1066556,7.8263187,10.690024,12.034423,10.875222,8.594546,8.937505,9.5033865,8.251588,6.125243,4.434457,4.8425775,5.0312047,5.020916,5.579939,6.574519,6.9826403,7.7268605,8.2481575,8.385342,8.405919,8.992378,9.373062,10.882081,12.476839,13.567448,14.016724,15.21365,15.601193,15.227368,14.29452,13.152468,15.367981,15.512024,14.935853,14.613472,15.165636,16.739817,17.78927,18.03963,17.737827,17.62808,16.564907,15.937293,15.282242,14.928994,16.026463,17.525192,18.763273,20.145397,21.260014,20.913624,18.28313,17.87158,17.995045,17.837284,17.480608,19.294859,17.655516,15.803539,15.165636,15.37827,14.411126,14.483148,15.621771,17.665806,20.262003,20.03908,18.293419,16.300829,15.199932,15.988737,17.662374,17.672665,16.859852,16.108772,16.331696,15.920145,16.506605,17.405157,18.12537,18.341434,16.13278,15.402277,15.29253,14.935853,13.450842,12.236768,11.664027,11.873232,12.758065,13.941273,13.474849,13.152468,13.293081,13.426835,12.281353,11.670886,11.180455,10.9541025,10.9541025,10.971251,10.624862,10.22703,9.72288,9.054111,8.155559,7.630832,7.010077,6.6876955,6.8728933,7.589677,7.805741,8.117833,8.501947,9.266746,11.05356,11.934964,12.493987,12.000127,10.576848,9.205012,9.400499,9.386781,9.884071,10.864933,11.567999,11.286773,10.065839,8.964942,8.31332,7.7028537,7.3564653,7.2158523,7.3598948,7.6171136,7.56224,0.20920484,0.2194936,0.21263443,0.20234565,0.19891608,0.23321195,0.22635277,0.274367,0.31552204,0.32581082,0.31552204,0.4081209,0.42183927,0.41840968,0.42526886,0.432128,0.4389872,0.4664239,0.53501564,0.61389613,0.6276145,0.48357183,0.548734,0.58988905,0.5418748,0.50757897,0.5178677,0.4355576,0.4424168,0.5178677,0.432128,0.39783216,0.37382504,0.42526886,0.50757897,0.48357183,0.5693115,0.64133286,0.6310441,0.5761707,0.6276145,0.64476246,0.6859175,0.67219913,0.64819205,0.7888051,0.7579388,0.7510797,0.7956643,0.8676856,0.89169276,0.8505377,0.75450927,0.7407909,0.78194594,0.6790583,0.5624523,0.48700142,0.4938606,0.53844523,0.5041494,0.4629943,0.4389872,0.490431,0.6276145,0.8471081,1.3992717,1.7799559,1.9342873,2.0440342,2.5413244,5.6073756,3.5359046,1.0494537,0.12346515,0.0034295875,0.041155048,0.020577524,0.0,0.030866288,0.15090185,0.20577525,0.16462019,0.07888051,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.01371835,0.01371835,0.010288762,0.006859175,0.030866288,0.72707254,0.5555932,0.6893471,1.0185875,0.13375391,0.072021335,0.041155048,0.024007112,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.1097468,0.37382504,0.764798,0.84367853,0.6756287,0.45270553,0.39783216,0.51100856,0.5693115,0.38754338,0.3018037,0.33266997,0.4115505,0.4115505,0.17147937,0.39440256,0.72364295,0.8779744,0.6344737,0.7133542,0.8128122,0.85396725,0.7613684,0.47328308,0.25721905,0.18519773,0.28122616,0.4115505,0.31552204,0.24350071,0.32581082,0.30866286,0.1920569,0.2194936,0.14061308,0.18176813,0.20577525,0.1920569,0.22978236,0.274367,0.17833854,0.16119061,0.21263443,0.09602845,0.16462019,0.13375391,0.116605975,0.15090185,0.17490897,0.28465575,0.2777966,0.24350071,0.26407823,0.4115505,0.33266997,0.5418748,0.7373613,0.8025235,0.805953,0.805953,0.8265306,0.83338976,0.86082643,1.0014396,1.2895249,1.3101025,1.3306799,1.4164196,1.4610043,1.6016173,1.7079345,1.8759843,2.0028791,1.7902447,1.9994495,2.0680413,2.2566686,2.5584722,2.6887965,2.6990852,2.7402403,2.6990852,2.7299516,3.2443898,3.8137012,4.314421,4.681387,4.931747,5.1340923,5.4667625,5.7754254,5.9400454,5.9126086,5.7239814,5.195825,5.336438,5.4976287,5.504488,5.638242,6.1629686,6.8043017,7.56567,8.337327,8.89635,9.510246,9.760606,9.740028,9.537683,9.235879,9.277034,9.119273,8.934075,8.97523,9.592556,10.405369,10.81006,11.166737,11.540562,11.712041,11.89038,11.794352,11.605724,11.622872,12.271064,12.699762,12.627741,12.80265,13.224489,13.169616,13.173045,13.560589,13.72178,13.642899,13.920695,13.738928,13.831526,14.009865,14.2533655,14.726648,16.064188,16.702091,17.38115,18.169954,18.4649,18.811287,19.507494,20.069946,20.587814,21.702429,22.330044,23.160004,23.571554,23.571554,23.811626,24.6896,26.016851,27.361248,28.10204,27.460707,36.055252,40.73664,47.602673,51.515835,36.08955,20.539799,13.145609,10.80663,10.419086,8.89635,8.872343,8.080108,9.582268,11.516555,7.1095347,3.590778,2.767677,3.2135234,3.3815732,1.6084765,1.6084765,1.4369972,1.313532,1.3443983,1.5193073,2.534465,3.8960114,4.979761,5.8817425,7.4113383,8.676856,11.125582,12.932974,13.540011,13.653188,13.797231,13.560589,13.255356,13.258785,14.003006,14.805529,15.985307,17.058767,17.62808,17.38115,17.45317,18.015623,18.828436,19.428614,19.154245,19.517782,19.819586,20.189981,20.834743,22.007662,22.426073,22.340332,22.53239,22.751883,21.719578,21.246294,20.652975,20.416334,20.62897,20.989075,22.258022,23.722456,20.752434,14.675205,12.775213,12.21962,11.231899,10.024684,9.362774,10.5597,12.113303,12.8197975,13.121602,13.419975,14.092175,14.38026,14.349394,14.496866,14.781522,14.647768,14.160767,14.1299,14.212211,14.126471,13.63261,13.13189,12.569438,11.516555,10.199594,9.527394,9.006097,8.683716,8.385342,8.05953,7.7714453,7.8777623,7.6514096,7.431916,7.377043,7.486789,7.8777623,8.495089,8.944365,8.954653,8.3922,7.4627824,7.160979,7.082098,7.0272245,6.9860697,6.5642304,6.4407654,6.307011,5.9812007,5.4084597,5.435896,5.4633327,5.4804807,5.545643,5.754848,5.857735,6.012067,6.279575,6.5539417,6.5642304,6.660259,6.385892,6.046363,5.8234396,5.7719955,6.1286726,6.6533995,6.7802944,6.5710897,6.7048435,6.8763227,7.0546613,7.157549,7.130112,6.958633,7.5862474,7.795452,7.723431,7.534804,7.425057,6.773435,6.5539417,6.5024977,6.4819202,6.4887795,6.5985265,7.0032177,7.8331776,8.759167,8.97866,9.026674,9.489669,10.079557,10.590566,10.88551,11.417097,12.010415,12.614022,13.121602,13.37882,12.878101,13.210771,13.63604,13.797231,13.728639,13.762935,13.203912,12.891819,13.104454,13.560589,13.985858,14.13676,14.267084,14.5585985,15.127911,16.2974,16.88386,16.499744,15.498305,14.973578,14.939283,16.78783,18.897026,19.997925,19.147387,10.875222,6.111525,4.2835546,4.4721823,5.394741,3.1826572,4.99005,7.970361,10.240748,10.861504,12.524854,14.147048,15.806969,17.089634,17.069057,18.440891,20.406046,21.45207,21.4555,21.69214,21.349182,20.814167,19.991066,18.890167,17.604073,17.000465,16.808409,16.753534,16.691803,16.63007,17.418875,16.46888,14.781522,13.227919,12.548861,14.239647,15.995596,17.549198,18.36887,17.652086,17.130789,16.815268,16.811838,17.158226,17.802988,18.101362,18.632948,19.486916,20.502073,21.239435,21.911634,21.143406,20.011642,18.975908,17.854433,16.55119,14.393978,12.037852,9.956093,8.440215,6.8900414,4.547633,3.1483612,3.3541365,4.7774153,6.8626046,6.4236174,6.090947,6.3378778,5.4496145,8.628842,9.626852,6.958633,3.0729103,4.3349986,2.3424082,1.2106444,3.3061223,7.589677,9.599416,3.799983,1.7730967,1.6016173,2.1469216,3.0420442,5.2506986,9.160428,8.80718,5.6073756,8.371623,12.147599,12.068718,10.401938,9.777754,13.214201,14.96672,12.483699,8.354475,4.9660425,4.4996185,4.6127954,4.588788,5.435896,6.6293926,6.0875177,7.291303,8.217292,8.625413,8.7145815,9.132992,9.6645775,11.592006,12.792361,12.751206,12.583157,14.726648,14.79524,14.037301,13.1593275,12.319078,13.4645605,13.505715,13.262215,13.368532,14.260224,16.21509,17.881868,18.770132,18.842154,18.495766,17.556059,16.606062,15.830976,15.354263,15.258235,16.383139,17.730967,19.579515,21.37662,21.747015,20.220848,19.263992,17.947031,16.37285,15.676644,16.448301,16.338554,16.204802,16.328266,16.414005,15.584045,14.946142,15.350834,17.1205,20.052797,21.27716,20.244854,18.001905,15.96816,15.9578705,17.03819,16.80498,16.530611,16.640358,16.715809,15.817257,16.173935,17.398296,18.677534,18.770132,14.987297,12.991278,12.367092,12.240198,11.266195,10.467101,10.103564,10.408798,11.5645685,13.735497,13.817808,13.032433,12.500846,12.442543,12.175035,11.519984,11.084427,10.782623,10.611144,10.63858,10.796341,10.943813,10.844356,10.374502,9.547972,8.573969,7.3358874,6.7459984,6.9552035,7.377043,7.442205,7.8263187,8.31675,9.081548,10.64201,11.427385,11.835506,11.115293,9.832627,9.866923,10.820349,11.015835,10.88894,10.799771,11.012405,10.401938,8.632272,7.6925645,7.8777623,7.81603,7.1061053,6.9826403,6.9723516,6.958633,7.174697,0.26064864,0.2469303,0.216064,0.20920484,0.23321195,0.24350071,0.2194936,0.20577525,0.216064,0.25378948,0.29151493,0.36353627,0.41840968,0.47328308,0.50757897,0.45613512,0.48357183,0.58988905,0.53844523,0.3841138,0.45613512,0.5178677,0.48700142,0.42869842,0.36010668,0.274367,0.3841138,0.34638834,0.31209245,0.32238123,0.33609957,0.34638834,0.36010668,0.41498008,0.48357183,0.45613512,0.50757897,0.51100856,0.52815646,0.6173257,0.823101,0.70306545,0.65162164,0.6824879,0.75450927,0.77851635,0.70649505,0.6962063,0.7579388,0.8162418,0.7339317,0.67219913,0.5658819,0.5693115,0.64476246,0.53501564,0.5212973,0.59331864,0.70306545,0.77165717,0.6859175,0.5761707,0.5693115,0.6173257,0.7888051,1.2517995,1.862266,2.1332035,2.4315774,2.7985435,2.9460156,2.5927682,1.2860953,0.31895164,0.07545093,0.01371835,0.01371835,0.006859175,0.0,0.07888051,0.39783216,0.7133542,0.48357183,0.18176813,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.061732575,0.041155048,0.010288762,0.006859175,0.030866288,0.64133286,0.6276145,0.66533995,0.7339317,0.12346515,0.061732575,0.0274367,0.0274367,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.06859175,0.274367,0.59674823,0.7922347,0.7442205,0.48357183,0.47328308,0.6790583,0.59674823,0.51100856,0.4046913,0.32581082,0.3018037,0.34981793,0.06859175,0.28465575,0.5693115,0.78194594,1.039165,0.7442205,0.85396725,0.9568549,0.8265306,0.4115505,0.34981793,0.26407823,0.24350071,0.3018037,0.34981793,0.24007112,0.19548649,0.18176813,0.20920484,0.30523327,0.30523327,0.26750782,0.29151493,0.32581082,0.16804978,0.09602845,0.17833854,0.21263443,0.15433143,0.106317215,0.106317215,0.08916927,0.08916927,0.12346515,0.19891608,0.20920484,0.23321195,0.20920484,0.18176813,0.29151493,0.38754338,0.64133286,0.83681935,0.8676856,0.7339317,0.78194594,0.8196714,0.864256,0.9294182,1.039165,1.0631721,1.2243627,1.3169615,1.2792361,1.2037852,1.5604624,1.821111,1.8039631,1.5707511,1.4507155,1.6084765,1.7765263,1.9411465,2.0165975,1.845118,2.0406046,2.318401,2.4418662,2.5619018,3.2203827,3.6353626,3.9028704,4.0366244,4.2423997,4.914599,5.4496145,5.5113473,5.528495,5.5902276,5.4324665,5.4187484,5.610805,5.638242,5.5422134,5.7377,6.6533995,7.2295704,7.7611566,8.200144,8.162418,8.992378,9.31133,9.451943,9.527394,9.431366,8.906639,8.453933,8.375052,8.639131,8.89635,9.445084,9.97667,10.611144,11.2593355,11.626302,11.688034,11.876661,11.979549,11.989838,12.099585,12.528283,13.145609,13.817808,14.308239,14.280802,13.893259,14.095605,14.119612,13.725209,13.214201,13.032433,13.680624,14.46257,14.887839,14.678635,15.656067,16.678083,17.576635,18.21111,18.478617,18.502625,19.459478,20.522652,21.3629,22.155134,23.671013,25.19375,25.996273,25.985985,25.680752,25.52299,25.831654,26.531288,27.495003,28.534168,34.062664,38.356506,46.933903,52.77792,36.346767,23.931662,17.686382,13.207341,8.858624,5.7822843,9.177576,7.5725293,7.31531,8.625413,5.5833683,3.069481,3.1380725,2.8980014,1.8039631,1.6324836,1.9754424,1.821111,1.670209,1.8862731,2.7162333,3.5461934,4.2389703,5.06893,6.1561093,7.4627824,9.39021,10.714031,11.355364,11.664027,12.421966,13.481709,13.766364,13.783512,13.903547,14.342535,16.026463,17.12736,17.480608,17.29884,17.151367,17.017612,17.916164,19.065077,20.104242,21.1194,22.302607,23.211449,23.101702,22.655855,23.986534,24.072275,23.214878,22.806757,22.673002,21.071384,20.803877,20.334024,20.03565,20.172834,20.903336,22.515242,24.391226,20.70099,13.275933,11.626302,10.81006,10.1652975,8.937505,7.7885933,8.790032,10.693454,12.689473,14.123041,14.874121,15.350834,15.765814,16.050468,15.971589,15.782962,16.235666,15.71094,15.066177,14.658057,14.363112,13.594885,12.507706,11.705182,10.9198065,10.041832,9.126132,8.464222,8.073249,7.98065,8.025234,7.8434668,7.939495,7.8366075,7.6342616,7.4010496,7.157549,7.6925645,8.752307,9.379922,9.211872,8.453933,7.905199,7.675417,7.5588107,7.363324,6.910619,6.3138704,6.108095,6.2247014,6.4098988,6.2247014,5.8337283,5.830299,5.90232,5.888602,5.768566,5.9400454,5.9640527,6.0532217,6.1972647,6.1492505,6.0875177,5.7891436,5.5079174,5.40503,5.5387836,5.8062916,6.0395036,6.0703697,5.9126086,5.751418,5.7754254,6.351596,6.9620624,7.349606,7.507367,7.6788464,7.5759587,7.4524937,7.363324,7.157549,6.5333643,6.433906,6.3961806,6.341307,6.560801,6.7185616,7.291303,8.052671,8.711152,8.879202,8.635701,8.738589,9.448513,10.374502,10.484249,11.177026,11.976119,12.425395,12.586586,13.001566,12.452832,12.624311,13.334236,14.085316,14.085316,14.143619,13.419975,12.953552,13.025573,13.121602,13.231348,13.416546,13.557159,13.725209,14.174485,15.237658,16.12592,16.064188,15.083325,14.006435,13.9481325,14.96672,17.024471,18.598652,16.691803,10.491108,5.7102633,3.4878905,4.6265135,9.582268,7.3598948,8.049242,9.55826,11.094715,13.169616,14.2190695,14.928994,16.815268,19.181683,19.11995,18.900457,19.596663,20.546658,21.544668,22.827333,22.326614,22.302607,21.959648,20.923914,19.226267,17.981327,16.945591,16.170506,15.9578705,16.859852,17.384579,16.691803,15.141628,13.560589,13.245067,14.819247,15.944152,17.099922,18.152807,18.3723,17.724108,17.508043,17.20967,17.134218,18.403166,18.670673,18.931322,19.54522,20.399187,20.872469,21.78817,21.688711,21.43835,20.676983,17.806417,14.939283,12.205902,10.216741,8.673427,6.3790326,4.3761535,3.7108135,3.9371665,4.6402316,5.446185,5.5833683,6.4407654,6.9380555,6.3310184,4.180667,9.283894,10.028113,6.773435,2.037175,0.48700142,0.4389872,0.5178677,3.9474552,8.625413,7.1095347,2.568761,1.0048691,0.5658819,1.039165,3.8617156,3.7622573,7.2707253,7.016936,4.0366244,7.798882,11.30049,11.351934,9.259886,8.30646,13.762935,12.713481,12.085866,9.5033865,5.597087,3.998899,4.2286816,4.314421,5.212973,6.64997,7.1266828,7.822889,8.601405,9.14328,9.342196,9.294182,10.1481495,12.264205,13.101024,12.178465,11.094715,13.509145,12.987847,12.3533745,12.370522,11.732618,13.114742,13.622321,13.533153,13.138749,12.771784,15.371411,17.2131,18.214539,18.79071,19.850452,18.519772,17.62122,17.19938,16.942162,16.173935,16.856422,17.494326,18.656956,20.488356,22.734735,21.356041,20.591244,18.910746,16.396858,14.723219,15.896138,15.265094,14.867262,15.484588,16.6335,16.88729,16.438013,16.335125,17.000465,18.235117,20.992504,22.021381,20.433481,17.398296,16.12935,17.813278,17.857862,17.096493,16.335125,16.37285,16.383139,16.352274,16.688372,17.185663,17.014183,14.009865,12.068718,11.149589,10.545981,8.9100685,8.81404,9.009526,9.668007,10.830637,12.404818,13.358243,13.073587,12.487128,12.041282,11.688034,11.039842,10.549411,10.124143,9.89436,10.2236,10.957532,11.513125,11.787492,11.598865,10.696883,9.39021,8.083538,7.466212,7.5725293,7.7680154,7.4627824,7.641121,8.323608,9.3593445,10.422516,11.324498,11.698323,10.80663,9.537683,10.39165,11.598865,12.30536,11.7257595,10.425946,10.316199,9.815479,7.390761,6.025785,6.327589,6.5470824,6.327589,6.307011,6.495639,6.8214493,7.1266828,0.30866286,0.28465575,0.274367,0.30866286,0.36353627,0.36696586,0.3018037,0.29151493,0.30866286,0.33952916,0.37382504,0.40126175,0.34638834,0.31552204,0.32924038,0.34638834,0.31209245,0.34638834,0.37039545,0.36353627,0.34638834,0.34981793,0.34295875,0.32924038,0.31895164,0.31209245,0.30523327,0.274367,0.2709374,0.30523327,0.33609957,0.39783216,0.3566771,0.34638834,0.4115505,0.4938606,0.58302987,0.53501564,0.5590228,0.6790583,0.7373613,0.7922347,0.82996017,0.8093826,0.7407909,0.71678376,0.6241849,0.6036074,0.59674823,0.58988905,0.61046654,0.607037,0.5521636,0.5521636,0.59674823,0.5453044,0.7476501,0.78537554,0.8505377,0.9362774,0.8196714,0.83681935,0.91227025,0.94999576,1.1214751,1.8485477,2.3218307,2.6133456,2.7882545,2.9974594,3.4467354,2.0749004,0.9328478,0.2503599,0.048014224,0.12346515,0.16462019,0.16462019,0.17490897,0.20577525,0.2503599,0.35324752,0.31552204,0.20234565,0.07888051,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.072021335,0.06516216,0.024007112,0.01371835,0.010288762,0.0,0.0,0.1097468,0.09259886,0.106317215,0.15090185,0.07888051,0.45613512,0.53844523,0.42526886,0.216064,0.037725464,0.01371835,0.006859175,0.010288762,0.017147938,0.0,0.0,0.006859175,0.017147938,0.020577524,0.0,0.0548734,0.2194936,0.37039545,0.4698535,0.59674823,0.45270553,0.4389872,0.44584638,0.4424168,0.48357183,0.41840968,0.5624523,0.6241849,0.4938606,0.24007112,0.22292319,0.31895164,0.53844523,0.72364295,0.548734,0.70649505,0.83338976,0.7990939,0.65162164,0.607037,0.5178677,0.3566771,0.36696586,0.4938606,0.37382504,0.29494452,0.3806842,0.38754338,0.28465575,0.24350071,0.36010668,0.25721905,0.24350071,0.33266997,0.24007112,0.14747226,0.19548649,0.16804978,0.06859175,0.12003556,0.08916927,0.09945804,0.106317215,0.12346515,0.2469303,0.2503599,0.28465575,0.3018037,0.34981793,0.5453044,0.4972902,0.64819205,0.7407909,0.6859175,0.5624523,0.6001778,0.59331864,0.6756287,0.8093826,0.7922347,0.8676856,0.922559,1.0185875,1.1214751,1.0940384,1.4404267,1.4953002,1.4129901,1.3409687,1.4267083,1.605047,1.7182233,1.7422304,1.728512,1.821111,2.0474637,2.177788,2.270387,2.5310357,3.316411,3.5187566,3.6216443,3.940596,4.431027,4.681387,5.1409516,5.284994,5.2506986,5.147811,5.0655007,5.562791,5.754848,5.895461,6.142391,6.543653,6.9689217,7.5862474,8.128122,8.344186,8.004657,9.2153015,9.400499,9.126132,8.9100685,9.22216,9.781183,9.547972,9.177576,8.971801,8.89635,9.582268,10.065839,10.556271,11.039842,11.31078,11.547421,11.705182,11.821788,11.763485,11.2593355,12.133881,13.203912,14.088745,14.7369375,15.405707,14.925565,14.640909,14.366542,14.092175,13.958421,13.581166,13.865822,14.531162,15.326826,16.047039,17.031332,17.501184,18.056778,18.86959,19.675543,20.19684,20.913624,21.544668,22.103691,22.875349,23.588703,24.675882,25.34122,25.43725,25.471546,25.540138,25.375517,25.505842,26.284359,27.885975,31.699677,31.548775,40.932125,51.824497,34.710854,25.27606,20.052797,13.845244,6.5813785,3.3301294,7.349606,6.8145905,6.927767,8.570539,8.296172,4.9214582,5.885172,4.770556,1.2826657,1.2655178,1.3649758,1.8382589,2.8328393,3.8960114,3.974892,4.5990767,5.2987127,6.0806584,7.0272245,8.303031,9.9801,11.585147,12.782072,13.505715,13.972139,13.392539,13.560589,14.177915,14.970149,15.673215,17.271402,17.586924,17.288551,16.88043,16.674654,17.322845,18.550638,20.025362,21.558388,23.118849,24.665592,26.26721,27.241213,27.35096,26.805656,26.579304,26.126596,25.787067,25.43382,24.490685,23.557837,21.956219,21.009653,21.256582,22.419212,24.079134,24.984545,20.971928,13.783512,11.091286,10.693454,9.750318,8.718011,7.9189177,7.531374,8.879202,11.005547,13.056439,14.507155,15.165636,16.324837,17.154797,17.165085,16.383139,15.3817,15.364552,14.743796,14.160767,13.824667,13.533153,13.375391,12.542002,11.701753,10.816919,9.15014,8.275595,7.8434668,7.6857057,7.641121,7.5245147,7.438775,7.3084507,7.298162,7.4696417,7.7920227,7.956643,8.820899,9.541112,9.616563,8.879202,8.292743,8.375052,8.131552,7.4456344,7.0718093,6.6396813,6.1972647,6.060081,6.1149545,5.8337283,6.108095,5.953764,5.8165803,5.8645945,5.9880595,6.101236,6.0497923,5.977771,5.9640527,6.0532217,6.1286726,5.9126086,5.6176643,5.3981705,5.3570156,5.439326,5.6245236,5.6793966,5.638242,5.802862,5.7377,5.967482,6.3618846,6.8866115,7.5931067,7.5279446,7.2638664,6.8626046,6.4304767,6.108095,5.8645945,5.6176643,5.381023,5.394741,6.121814,6.8557453,7.1541195,7.407909,7.6857057,7.7097125,7.805741,8.1212635,8.81404,9.654288,10.007536,10.779194,11.492548,11.897239,12.116733,12.6586075,12.919256,12.908967,13.094165,13.481709,13.618892,13.876111,13.718349,13.543441,13.498857,13.488567,13.179905,12.662037,12.569438,12.994707,13.516005,14.441993,15.347404,15.745236,15.498305,14.812388,13.512574,14.147048,15.861842,18.084215,20.526081,15.261664,8.577398,4.389872,3.5564823,3.8342788,5.2644167,6.48535,7.099246,7.377043,8.261876,10.882081,11.7086115,13.296511,16.071047,18.313997,18.866161,19.089085,19.150816,19.44919,20.604961,21.356041,21.246294,20.587814,19.682402,18.835295,17.933313,17.254255,16.431154,15.824117,16.54433,16.952452,16.640358,15.741806,14.620332,13.855534,14.668345,15.0456,15.570327,16.317978,16.87014,16.53404,16.654078,16.396858,16.098484,17.230247,18.094503,18.598652,19.384027,20.20027,19.884748,21.239435,21.35947,21.393766,21.225718,19.480057,12.343085,9.108984,7.0443726,5.5662203,6.217842,3.0454736,1.7662375,1.5947582,1.9994495,2.6887965,4.0537724,5.195825,5.8543057,6.2041235,6.866034,11.794352,10.868362,6.852316,2.5310357,0.70649505,0.4046913,0.30523327,1.0768905,3.2032347,6.9654922,4.3658648,2.2909644,0.90884066,1.1934965,4.9214582,3.8479972,5.4599032,5.0929375,3.4467354,6.550512,6.228131,6.8385973,6.7322803,6.914048,11.039842,8.155559,7.0375133,6.077229,4.664239,3.192946,4.763697,4.962613,5.7994323,7.449064,8.2481575,8.848335,9.72631,10.213311,10.233889,10.281903,10.803201,12.281353,13.056439,12.627741,11.667457,12.521424,11.958971,11.646879,12.037852,12.367092,14.003006,14.575747,14.205351,13.690913,14.503725,15.172495,16.654078,17.79613,18.54035,19.925903,19.45262,18.643238,17.96761,17.662374,17.71382,17.545769,16.976458,16.592344,17.003895,18.828436,19.157675,19.054789,18.38259,17.089634,15.199932,14.723219,13.618892,13.173045,13.7938,15.021593,15.62863,16.204802,16.715809,17.278261,18.149376,20.008213,22.213438,22.432932,20.800447,19.901896,19.46634,19.236557,18.636377,17.86815,17.936743,17.576635,17.099922,17.04848,16.938732,15.244516,13.255356,11.592006,10.185875,9.139851,8.704293,8.529384,8.375052,8.81404,10.014396,11.732618,13.097594,13.450842,13.169616,12.576297,11.921246,10.998687,10.367643,9.993818,9.962952,10.467101,11.084427,11.89038,12.277924,11.976119,11.063849,9.825768,8.601405,8.152129,8.354475,8.217292,7.8949103,7.9429245,8.460793,9.338767,10.275044,10.583707,10.923236,10.316199,9.122703,9.047252,9.6988735,10.14129,10.268185,10.271614,10.621432,9.427936,7.438775,6.2212715,6.0532217,5.9126086,5.3501563,5.7068334,6.619104,7.5245147,7.675417,0.31209245,0.34638834,0.432128,0.41498008,0.30866286,0.2777966,0.25721905,0.26407823,0.31895164,0.36353627,0.26750782,0.28122616,0.2469303,0.22635277,0.24007112,0.2469303,0.21263443,0.20920484,0.23321195,0.26064864,0.2469303,0.23664154,0.26064864,0.26064864,0.22978236,0.22978236,0.22292319,0.20577525,0.2194936,0.26407823,0.29837412,0.29151493,0.26064864,0.31895164,0.4355576,0.42183927,0.4972902,0.53844523,0.6001778,0.66876954,0.66191036,0.7373613,0.7922347,0.75450927,0.64133286,0.5727411,0.52815646,0.48700142,0.44927597,0.42869842,0.4698535,0.44584638,0.4938606,0.58302987,0.67219913,0.6859175,1.0014396,1.1797781,1.2312219,1.1934965,1.138623,1.1660597,1.1283343,1.1900668,1.4541451,1.9514352,2.5310357,3.4021509,3.7142432,3.625074,4.3041325,3.6525106,1.9480057,0.5590228,0.061732575,0.24350071,0.36010668,0.29151493,0.22635277,0.20577525,0.13032432,0.12003556,0.28465575,0.3841138,0.31209245,0.07888051,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.12689474,0.34638834,0.52815646,0.4424168,0.09259886,0.006859175,0.0034295875,0.0034295875,0.010288762,0.058302987,0.061732575,0.09259886,0.13375391,0.1097468,0.26750782,0.28808534,0.18519773,0.034295876,0.006859175,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.0034295875,0.0034295875,0.030866288,0.06516216,0.06516216,0.16119061,0.274367,0.32238123,0.33952916,0.48357183,0.64476246,0.48357183,0.33952916,0.33266997,0.3841138,0.881404,0.7510797,0.5590228,0.4664239,0.23321195,0.33266997,0.30866286,0.4081209,0.5693115,0.42869842,0.7099246,0.7133542,0.7682276,0.8676856,0.6824879,0.8265306,0.6962063,0.4972902,0.34295875,0.28122616,0.3018037,0.34638834,0.29151493,0.18519773,0.22978236,0.4115505,0.28465575,0.2194936,0.28808534,0.2503599,0.30523327,0.30866286,0.22978236,0.116605975,0.09602845,0.072021335,0.09602845,0.09945804,0.106317215,0.20577525,0.29151493,0.31895164,0.33266997,0.3806842,0.490431,0.42869842,0.48014224,0.5007198,0.47671264,0.5453044,0.4938606,0.548734,0.66533995,0.7888051,0.8505377,0.77508676,0.8196714,0.90198153,0.9362774,0.85739684,0.9877212,1.0288762,1.0768905,1.1626302,1.2826657,1.3855534,1.5158776,1.670209,1.8142518,1.8691251,2.0131679,2.1023371,2.2326615,2.4658735,2.8396983,3.1312134,3.3129816,3.5942078,3.974892,4.2766957,4.7088237,5.113515,5.3330083,5.3570156,5.305572,6.169828,6.327589,6.351596,6.4304767,6.3790326,6.608815,6.992929,7.5279446,8.021805,8.073249,9.050681,9.098696,8.525954,7.9292064,8.189855,8.838047,8.769455,8.556821,8.40249,8.128122,8.971801,9.448513,10.065839,10.799771,11.101575,11.039842,11.094715,11.30049,11.447963,11.067279,11.958971,13.066729,13.87954,14.3974085,15.138199,15.155347,15.227368,15.412566,15.704081,16.050468,15.4742985,15.501736,15.7966795,16.194511,16.70895,17.425734,17.802988,18.20768,18.890167,19.984205,21.229147,21.921923,22.288889,22.43979,22.350622,22.745024,23.225166,23.773901,24.288338,24.579853,24.466677,24.473536,24.494114,24.905664,26.572443,30.098059,32.220974,42.88356,55.346684,46.182823,32.15581,21.60983,12.2093315,4.619654,2.486451,4.290414,4.530485,4.722542,5.6176643,7.205563,4.605936,3.981751,3.199805,1.8862731,1.4404267,1.1900668,1.8519772,2.7573884,3.549623,4.149801,5.662249,7.0443726,8.347616,9.554831,10.583707,11.893809,12.867812,13.430264,13.886399,14.935853,15.367981,15.645778,15.913286,16.321407,17.031332,18.019053,18.602083,18.646667,18.327715,18.12194,17.741257,18.54035,19.888178,21.482935,23.35549,24.919382,26.754211,28.654203,30.019178,29.864847,30.152933,30.379286,30.324413,29.782537,28.541027,26.93598,25.334362,24.343212,23.983105,23.69502,24.919382,25.999702,22.710728,15.837835,11.183885,10.131001,9.208443,8.903209,9.078118,8.97523,7.750868,7.953213,9.599416,12.144169,14.46257,15.916716,16.657507,16.6335,15.999025,15.13134,14.623761,13.989287,13.313659,12.723769,12.394529,12.123591,11.540562,11.026124,10.412228,8.98209,8.549961,8.172707,8.162418,8.320179,7.922347,7.7885933,7.7131424,7.9189177,8.340756,8.635701,8.988949,9.235879,9.513676,9.616563,8.988949,8.375052,8.193284,7.7542973,7.06838,6.8454566,6.4407654,6.029215,5.8817425,5.895461,5.5833683,5.9983487,6.0497923,6.186976,6.420188,6.327589,6.293293,6.2247014,6.1801167,6.0703697,5.689686,5.535354,5.5113473,5.5422134,5.5319247,5.3741636,5.329579,5.3398676,5.329579,5.3570156,5.6313825,5.802862,5.9434752,6.276145,6.8385973,7.4765005,7.421627,7.2535777,6.800872,6.166398,5.717122,5.518206,5.2266912,5.06893,5.271276,6.0669403,6.5299344,6.8454566,6.9037595,6.842027,7.051232,7.1952744,7.8434668,8.546532,9.078118,9.448513,10.264755,10.80663,11.166737,11.540562,12.260776,12.542002,12.843805,13.1593275,13.488567,13.841815,13.927555,13.7938,13.622321,13.443983,13.121602,12.620882,11.934964,11.876661,12.593445,13.560589,14.198492,15.076467,15.6697855,15.580616,14.5585985,13.245067,13.29994,14.417986,16.359133,18.95876,18.79071,13.876111,8.697433,5.3913116,3.7691166,6.0326443,7.1129646,6.5710897,5.096367,4.5270553,6.8969,8.632272,10.120712,11.567999,12.994707,15.042171,15.830976,16.21509,16.846134,18.145947,19.068506,19.823015,19.888178,19.37031,19.013634,17.53548,16.818697,16.39,16.21166,16.691803,16.808409,16.438013,15.892709,15.268523,14.455711,14.706071,15.011304,15.46058,15.9750185,16.338554,16.221949,16.513464,16.482597,16.263103,16.863281,17.267973,18.139088,18.862732,19.161106,19.089085,20.423193,20.402617,22.264881,24.682741,21.78474,11.931535,6.4407654,3.7759757,2.8877127,3.1963756,1.8588364,0.94656616,0.64133286,0.9294182,1.587899,2.9220085,4.32128,5.079219,5.830299,8.553391,10.295622,7.6274023,4.1600895,1.8108221,0.8162418,0.42183927,0.26750782,0.45613512,1.7902447,5.7925735,6.5950966,3.998899,3.9268777,5.9331865,3.210094,5.672538,5.164959,4.0091877,4.245829,7.641121,3.7451096,6.258997,7.0443726,4.9180284,5.645101,4.6436615,4.012617,3.957744,4.0194764,3.100347,5.6142344,5.813151,6.193835,7.274155,7.6033955,8.282454,9.599416,9.9698105,9.3936405,9.47595,9.489669,10.714031,11.691463,11.934964,11.928105,11.893809,11.495977,11.430815,11.766914,11.958971,13.399398,14.102464,14.143619,14.143619,15.241087,14.610043,15.79325,17.072487,17.96418,19.21255,19.167965,18.62609,17.820137,17.223389,17.53891,17.730967,16.969599,16.386568,16.21852,15.79325,15.436573,15.340545,15.326826,15.3302555,15.412566,14.733508,13.690913,13.083877,13.289652,14.280802,15.319967,16.45173,17.353712,17.95389,18.44775,19.716698,22.011093,23.084553,22.673002,22.52896,21.973368,21.428062,20.6907,19.95677,19.809298,18.440891,17.134218,16.88386,17.117071,15.707511,13.642899,11.746337,9.983529,8.594546,8.093826,8.014946,7.7851634,8.172707,9.362774,10.988399,12.425395,12.88496,12.586586,11.856084,11.146159,10.573419,10.213311,10.131001,10.364213,10.923236,11.499407,12.243628,12.421966,11.797781,10.597425,9.654288,8.680285,8.289313,8.361334,8.045813,8.237869,8.573969,9.246168,10.185875,11.05356,11.108434,11.297061,10.583707,9.095266,8.117833,8.1487,8.680285,9.517105,10.319629,10.6145735,8.7283,6.5230756,5.4941993,5.645101,5.5250654,5.1992545,5.686256,6.5162163,7.3393173,7.932636,0.2503599,0.29837412,0.37725464,0.33952916,0.21263443,0.20577525,0.216064,0.23664154,0.28465575,0.30866286,0.20920484,0.216064,0.19891608,0.18862732,0.18862732,0.1920569,0.18176813,0.17147937,0.17490897,0.18519773,0.18176813,0.16804978,0.1920569,0.19548649,0.16804978,0.15433143,0.16462019,0.16804978,0.18176813,0.21263443,0.2503599,0.22978236,0.21263443,0.28465575,0.39440256,0.35324752,0.40126175,0.5041494,0.5658819,0.58302987,0.6379033,0.58645946,0.6173257,0.6173257,0.5624523,0.53158605,0.4389872,0.3841138,0.3566771,0.35324752,0.36696586,0.33609957,0.48014224,0.6790583,0.84024894,0.89512235,1.2723769,1.4575747,1.5124481,1.5124481,1.5364552,1.4404267,1.3478279,1.4815818,1.8588364,2.2841053,2.8019729,3.8377085,4.3933015,4.3692946,4.557922,4.8768735,2.7230926,0.75450927,0.06859175,0.20234565,0.4046913,0.33266997,0.2194936,0.15776102,0.082310095,0.024007112,0.4664239,0.75450927,0.6173257,0.18176813,0.09602845,0.041155048,0.010288762,0.030866288,0.15776102,0.07888051,0.19891608,0.4046913,0.58302987,0.6001778,0.13032432,0.017147938,0.020577524,0.024007112,0.0274367,0.037725464,0.09259886,0.10288762,0.07545093,0.08573969,0.14404267,0.116605975,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.037725464,0.12003556,0.20920484,0.36353627,0.36010668,0.35324752,0.38754338,0.41840968,0.7579388,0.4629943,0.3018037,0.42869842,0.37382504,1.0528834,0.9259886,0.6344737,0.45956472,0.31895164,0.432128,0.30523327,0.30523327,0.4698535,0.52472687,0.77508676,0.6824879,0.75450927,0.9568549,0.7373613,0.89855194,0.864256,0.6379033,0.39440256,0.51100856,0.45613512,0.33952916,0.1920569,0.09602845,0.18176813,0.35324752,0.32238123,0.26750782,0.26407823,0.274367,0.39097297,0.4115505,0.31895164,0.16462019,0.08916927,0.08573969,0.09602845,0.09259886,0.09259886,0.1371835,0.24007112,0.274367,0.30523327,0.34638834,0.33952916,0.32924038,0.3841138,0.41840968,0.4389872,0.5521636,0.4424168,0.5521636,0.72021335,0.84367853,0.85739684,0.7956643,0.84024894,0.89169276,0.8711152,0.72364295,0.7442205,0.8128122,0.88826317,0.96371406,1.0425946,1.1317638,1.2860953,1.5810398,1.9137098,2.0234566,1.8828435,1.9171394,2.0749004,2.253239,2.2841053,2.6785078,2.9734523,3.192946,3.4398763,3.9200184,4.40702,4.866585,5.2506986,5.48734,5.4804807,6.1732574,6.385892,6.4579134,6.4716315,6.2384195,6.358455,6.5642304,6.9963584,7.5553813,7.9086285,8.875772,8.865483,8.141841,7.390761,7.689135,7.829748,7.5588107,7.486789,7.6651278,7.606825,8.385342,8.89635,9.469091,10.086417,10.388221,10.460241,10.4705305,10.645439,10.9369545,11.012405,11.880091,12.922686,13.72178,14.177915,14.527733,15.347404,16.074476,16.743246,17.37429,17.95389,17.480608,17.261114,17.29884,17.508043,17.69667,17.926455,18.001905,18.115082,18.557497,19.744135,21.232576,21.908205,22.086544,21.942501,21.52066,21.78131,21.661274,21.959648,22.758743,23.424082,23.44809,23.917942,24.065414,24.11343,25.282919,29.076042,32.721695,42.657207,54.36925,52.404095,34.940636,20.495214,10.017825,4.461893,4.756838,3.8445675,3.175798,3.0420442,3.6559403,5.137522,3.8548563,3.0111778,2.9151495,3.0077481,1.879414,1.8759843,2.8225505,3.6147852,4.180667,5.470192,7.2192817,8.371623,9.712592,11.2421875,12.188754,13.059869,13.7526455,14.030442,14.311668,15.656067,16.80155,17.662374,18.005335,18.063637,18.564358,18.948471,19.03764,18.969048,18.852442,18.766703,17.95389,18.392878,19.325726,20.502073,22.196291,23.732746,25.392666,27.206917,28.774239,29.240664,29.532177,30.10149,30.242102,29.614489,28.252941,26.527859,25.416672,24.919382,24.665592,23.900795,24.627867,26.18147,23.26975,16.846134,14.109323,11.266195,10.350495,10.13786,10.13786,10.587136,8.56368,7.2638664,7.1129646,8.330468,10.923236,11.866373,13.502286,14.441993,14.393978,14.13676,13.094165,12.295071,11.417097,10.64201,10.6488695,10.587136,10.401938,10.161868,9.73317,8.762596,8.584257,8.05953,8.06296,8.591117,8.735159,8.512236,8.303031,8.429926,8.834618,9.074688,9.462232,9.571979,9.6645775,9.702303,9.342196,8.700864,8.165848,7.5416627,6.90033,6.5882373,6.2041235,5.90575,5.720552,5.675967,5.802862,6.1149545,6.262427,6.591667,7.0032177,6.941485,6.526505,6.23499,5.9126086,5.552502,5.267846,5.0449233,5.051782,5.206114,5.3707337,5.336438,5.1855364,5.137522,5.2164025,5.40503,5.65539,5.967482,6.1904054,6.5470824,6.9826403,7.1712675,7.0718093,7.040943,6.7322803,6.1492505,5.638242,5.2644167,5.0586414,5.0483527,5.346727,6.1458206,6.4990683,6.7459984,6.715132,6.56766,6.8043017,6.9620624,7.6171136,8.196714,8.591117,9.14328,9.822338,10.034973,10.131001,10.425946,11.231899,11.516555,12.185325,12.79922,13.200482,13.519434,13.63261,13.519434,13.375391,13.179905,12.706621,12.38424,11.849225,11.773774,12.3533745,13.29994,14.061309,15.055889,15.79325,15.683503,14.037301,12.823228,12.703192,13.560589,15.028452,16.479168,18.989626,17.559488,14.356253,10.738038,7.2604365,8.831187,8.718011,6.6122446,4.383013,6.0497923,4.245829,5.1512403,7.222711,9.325048,10.72432,13.37882,14.634049,15.450292,16.393429,17.645227,18.512913,19.750994,20.306587,20.045938,19.733847,17.95732,16.983316,16.62321,16.70552,17.089634,17.257685,17.103354,16.897577,16.554619,15.614912,15.29939,15.179354,15.37827,15.79325,16.11906,16.071047,16.21852,16.37285,16.61292,17.267973,17.28512,18.077356,18.516342,18.406595,18.4649,19.891607,18.54378,21.177702,25.300066,19.154245,9.692014,5.2815647,3.666229,2.860276,1.1317638,0.9842916,0.6824879,1.3889829,2.7368107,2.8259802,3.40901,5.0655007,6.101236,6.701414,8.89635,8.110974,4.9660425,2.393852,1.4644338,1.371835,0.7888051,0.6036074,0.77508676,2.2086544,6.773435,7.514226,4.5167665,5.4633327,8.320179,1.3169615,4.506478,3.8102717,3.2203827,4.5819287,7.6171136,2.9631636,5.844017,6.5642304,3.316411,2.2086544,2.609916,2.3458378,2.6750782,3.391862,2.8396983,4.9694724,5.2438393,5.5730796,6.355026,6.475061,7.1952744,8.309891,8.467651,7.8949103,8.39563,7.98065,8.971801,10.034973,10.618003,10.947243,11.293632,11.321068,11.410237,11.657167,11.869802,13.430264,14.092175,14.435134,14.802099,15.302819,14.531162,15.282242,16.29054,17.03819,17.741257,17.984756,17.826996,17.058767,16.204802,16.496315,16.828985,16.698662,16.835844,16.671225,14.321958,13.351384,13.059869,13.029003,13.481709,15.302819,14.668345,14.273943,14.081886,14.147048,14.613472,15.536031,16.856422,17.96418,18.608942,18.924463,19.919044,21.976797,23.386356,23.482386,22.645567,22.642136,22.645567,22.645567,22.570116,22.28546,20.255144,18.03963,16.990177,16.973028,16.365992,14.126471,12.127021,10.408798,8.985519,7.829748,7.630832,7.5450926,7.9189177,8.879202,10.329918,11.622872,11.89038,11.540562,10.930096,10.347065,10.158438,10.041832,10.264755,10.820349,11.434244,12.085866,12.648318,12.442543,11.423956,10.175586,9.31133,8.48137,8.117833,8.1487,7.9875093,8.532814,9.105555,9.925226,10.909517,11.664027,11.742908,11.691463,10.707172,9.030104,7.9292064,7.98065,8.303031,8.930646,9.582268,9.661148,7.6616983,5.744559,5.0620713,5.425607,5.2987127,5.411889,5.8337283,6.355026,6.924337,7.6616983,0.17833854,0.18519773,0.15776102,0.14404267,0.15776102,0.19891608,0.20577525,0.22292319,0.2194936,0.20234565,0.22292319,0.22292319,0.19548649,0.16119061,0.14404267,0.16462019,0.17833854,0.17147937,0.16462019,0.15433143,0.14747226,0.1371835,0.1371835,0.14061308,0.14747226,0.13375391,0.1371835,0.15433143,0.16804978,0.17833854,0.20577525,0.22978236,0.2194936,0.22635277,0.2709374,0.31895164,0.33952916,0.41840968,0.4629943,0.48014224,0.5796003,0.39783216,0.4046913,0.45956472,0.5007198,0.5418748,0.39097297,0.33266997,0.32924038,0.33952916,0.33266997,0.36353627,0.5418748,0.7922347,1.0254467,1.138623,1.5227368,1.546744,1.6016173,1.7662375,1.8313997,1.6564908,1.6187652,1.8313997,2.311542,3.018037,3.210094,3.865145,4.605936,4.9077396,4.0949273,4.746549,2.7951138,0.8745448,0.09945804,0.061732575,0.33952916,0.32581082,0.20920484,0.106317215,0.08573969,0.044584636,0.7099246,1.0666018,0.83681935,0.48357183,0.32581082,0.16462019,0.0548734,0.07545093,0.32238123,0.16119061,0.14747226,0.15433143,0.18862732,0.3841138,0.10288762,0.05144381,0.072021335,0.07888051,0.0548734,0.06859175,0.15090185,0.1371835,0.034295876,0.024007112,0.082310095,0.06859175,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0274367,0.020577524,0.061732575,0.17490897,0.30866286,0.51100856,0.42869842,0.4355576,0.5521636,0.42869842,0.6173257,0.34295875,0.29494452,0.52472687,0.42183927,0.84024894,1.0871792,0.9842916,0.65162164,0.51100856,0.52472687,0.33266997,0.28122616,0.4424168,0.61389613,0.8025235,0.72364295,0.7305021,0.8471081,0.77508676,0.7407909,0.7682276,0.7099246,0.64819205,0.89169276,0.6927767,0.42869842,0.22292319,0.12689474,0.12003556,0.22292319,0.33609957,0.34981793,0.3018037,0.36353627,0.38754338,0.4389872,0.35324752,0.17147937,0.116605975,0.1371835,0.12346515,0.12346515,0.1371835,0.116605975,0.14061308,0.17833854,0.24007112,0.29151493,0.25721905,0.29837412,0.39440256,0.48700142,0.53158605,0.51100856,0.41840968,0.548734,0.7579388,0.8779744,0.7339317,0.84024894,0.83681935,0.84024894,0.8505377,0.72021335,0.78194594,0.8471081,0.8505377,0.8196714,0.8745448,1.0357354,1.1866373,1.4953002,1.920569,2.2120838,1.8073926,1.8142518,1.9925903,2.1332035,2.0646117,2.5001693,2.8568463,3.018037,3.1483612,3.7176728,4.3041325,4.6093655,4.9351764,5.2644167,5.2815647,5.470192,5.8062916,6.121814,6.3138704,6.351596,6.447624,6.601956,6.8283086,7.140401,7.5382333,8.666568,8.738589,8.182996,7.6445503,7.9909387,7.5450926,6.9654922,6.824879,7.1712675,7.531374,8.080108,8.628842,8.98209,9.160428,9.39707,9.9869585,10.172156,10.281903,10.539123,11.05699,11.928105,12.878101,13.697772,14.208781,14.239647,15.728088,16.983316,17.916164,18.560926,19.078794,18.845583,18.410025,18.313997,18.560926,18.629519,18.416885,18.001905,17.758404,18.04306,19.188541,20.361462,21.019941,21.229147,21.160555,21.112541,21.191422,20.728426,20.70442,21.410915,22.474087,22.998814,23.887077,24.27119,24.209457,24.658733,28.568464,30.958885,37.440807,46.320007,48.62126,31.648233,18.053349,9.091836,5.545643,7.7028537,5.844017,3.6353626,2.976882,3.8342788,4.2183924,4.389872,5.0655007,5.6313825,5.2575574,2.8637056,3.0386145,4.40359,5.809721,7.0032177,8.625413,9.877212,9.932085,10.532263,11.8869505,12.6586075,13.049581,13.9481325,14.658057,15.199932,16.300829,17.267973,18.564358,19.250275,19.36688,19.912186,20.248285,19.408035,18.71526,18.584934,18.509483,18.331144,18.684393,19.11309,19.555508,20.344313,21.541239,22.741594,23.756752,24.579853,25.382378,25.553856,26.1849,26.298077,25.51613,24.075705,22.679861,21.993944,22.052248,22.508383,22.60441,22.957659,24.7822,21.880768,16.0539,17.117071,12.922686,12.065289,11.351934,10.216741,10.717461,10.2236,8.872343,6.7185616,5.086078,6.5779486,6.3961806,8.961512,11.101575,11.705182,11.7086115,10.686595,9.901219,8.944365,8.203573,8.868914,9.482809,9.56512,9.386781,9.023245,8.351046,8.251588,7.689135,7.6274023,8.296172,9.225591,8.796892,8.529384,8.491658,8.669997,8.97866,9.153569,9.575408,9.846346,9.880642,9.925226,9.445084,8.676856,7.840037,7.0923867,6.5162163,6.258997,6.036074,5.7136927,5.5319247,6.108095,6.2555676,6.358455,6.6739774,7.140401,7.3873315,6.632822,6.1046658,5.4016004,4.7328305,4.9214582,4.852866,4.7362604,4.7328305,4.8768735,5.0620713,4.99005,5.0655007,5.3707337,5.802862,6.0703697,6.3447366,6.615674,6.9071894,7.0923867,6.883182,6.6396813,6.6396813,6.5333643,6.1972647,5.7479887,5.2335505,5.1238036,5.1340923,5.302142,6.0086374,6.6465406,6.800872,6.790583,6.800872,6.8969,7.1026754,7.425057,7.73029,8.114404,8.903209,9.328478,9.218731,9.009526,9.112414,9.925226,10.439664,11.238758,11.955542,12.367092,12.394529,12.655178,12.737488,12.809509,12.850664,12.63803,12.734058,12.507706,12.336226,12.397959,12.662037,13.666906,14.778092,15.721229,15.765814,13.725209,12.38424,12.319078,13.162757,14.373401,15.247946,16.918156,18.293419,18.663815,17.195951,12.926115,12.898679,10.422516,6.5985265,4.7945633,10.624862,4.616225,3.216953,5.593657,9.770895,12.644889,15.110763,16.602633,17.737827,18.746124,19.469769,20.255144,21.242865,21.558388,21.102251,20.553518,18.969048,17.737827,17.072487,17.007324,17.388008,17.929884,18.468328,18.811287,18.612371,17.37772,16.39,15.422854,15.103903,15.5085945,16.13621,15.954441,15.865272,16.088194,16.756964,17.909306,18.094503,18.495766,18.636377,18.516342,18.602083,20.183123,17.237106,18.550638,21.558388,12.339656,5.528495,4.605936,4.979761,4.0091877,0.99801,0.8265306,1.1763484,3.3198407,6.0395036,5.658819,5.8165803,7.5107965,8.776315,8.97866,8.81747,7.606825,5.2301207,3.2718265,2.4075704,2.3972816,1.4644338,1.4850113,2.037175,3.8617156,8.831187,6.7700057,3.649081,4.2355404,6.3653145,0.94999576,1.2689474,1.7765263,2.6476414,4.0023284,5.9126086,3.3438478,4.616225,4.5853586,2.4658735,1.8348293,1.9068506,1.6804979,2.0749004,2.7916842,2.3081124,3.2306714,3.5564823,4.122364,4.98662,5.453044,6.018926,6.5059276,6.5230756,6.4579134,7.490219,6.883182,7.5931067,8.543102,9.105555,9.095266,10.569988,11.077567,11.293632,11.660598,12.38767,14.315098,14.891269,15.179354,15.405707,14.96329,14.79524,15.151917,15.642348,16.029892,16.242527,16.561478,16.585485,15.9750185,15.179354,15.46744,15.560039,16.149927,17.021042,17.065628,14.280802,13.375391,12.778643,12.295071,12.456262,14.5243025,14.054449,14.417986,14.997586,15.409137,15.501736,16.029892,17.28512,18.468328,19.198832,19.54179,20.36832,22.223726,23.873358,23.989964,21.146837,21.417774,22.501524,23.571554,24.291767,24.802776,23.218307,20.673553,18.344864,16.818697,16.081335,14.105893,12.517994,11.293632,10.093276,8.296172,7.781734,7.8503256,8.152129,8.721441,9.959522,10.912948,10.8958,10.593996,10.285333,9.8429165,9.877212,9.884071,10.271614,11.022695,11.677745,12.38767,12.847235,12.339656,11.046701,10.031544,9.047252,8.217292,7.81603,7.8537555,8.076678,8.700864,9.345626,10.206452,11.149589,11.718901,11.852654,11.626302,10.535692,8.954653,8.134981,8.735159,8.639131,8.433355,8.330468,8.179566,6.5710897,5.4804807,5.209543,5.439326,5.24041,5.5559316,5.8508763,6.276145,6.81802,7.3255987,0.21263443,0.20234565,0.17147937,0.14747226,0.1371835,0.1371835,0.12346515,0.12346515,0.12689474,0.1371835,0.1371835,0.1371835,0.1097468,0.09259886,0.09259886,0.09259886,0.10288762,0.106317215,0.106317215,0.1097468,0.12346515,0.12346515,0.13032432,0.1371835,0.13375391,0.12346515,0.13375391,0.14747226,0.16462019,0.18176813,0.16804978,0.15433143,0.16119061,0.18176813,0.20920484,0.26064864,0.26064864,0.26750782,0.36696586,0.45613512,0.274367,0.2503599,0.28122616,0.30523327,0.31209245,0.33609957,0.4081209,0.40126175,0.34981793,0.31895164,0.3806842,0.53844523,0.6173257,0.7922347,1.1008976,1.4198492,1.6770682,1.6496316,1.6427724,1.7319417,1.7696671,1.9171394,1.9239986,2.095478,2.6647894,3.799983,3.5804894,4.0366244,4.722542,4.914599,3.6319332,3.7176728,2.867135,1.4953002,0.26750782,0.12346515,0.4389872,0.40126175,0.22292319,0.072021335,0.061732575,0.14747226,0.6241849,0.8196714,0.7888051,1.3272504,0.97400284,0.490431,0.16119061,0.0548734,0.030866288,0.006859175,0.010288762,0.020577524,0.030866288,0.030866288,0.041155048,0.09259886,0.14747226,0.16462019,0.09259886,0.06859175,0.041155048,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.1371835,0.09602845,0.1371835,0.23664154,0.07545093,0.30866286,0.2469303,0.29151493,0.5007198,0.61046654,0.4389872,0.21263443,0.07888051,0.12689474,0.39783216,0.8848336,1.2826657,1.371835,1.155771,0.84024894,0.5693115,0.37382504,0.31552204,0.3566771,0.3806842,0.58988905,0.6036074,0.7373613,0.922559,0.70306545,0.77508676,0.6379033,0.5418748,0.5624523,0.61046654,0.6962063,0.5144381,0.36353627,0.3018037,0.16804978,0.1920569,0.2709374,0.34981793,0.42526886,0.53501564,0.45956472,0.33266997,0.23664154,0.18862732,0.15090185,0.20234565,0.20577525,0.26064864,0.32238123,0.21263443,0.18862732,0.16462019,0.18176813,0.25721905,0.36696586,0.37725464,0.33609957,0.37725464,0.47328308,0.4115505,0.38754338,0.5727411,0.7133542,0.72021335,0.67219913,0.72021335,0.5761707,0.51100856,0.58645946,0.67219913,0.6824879,0.7510797,0.84367853,0.94999576,1.0837497,1.3032433,1.3958421,1.6153357,1.9823016,2.2738166,2.1503513,2.3767042,2.633923,2.7128036,2.5173173,3.0797696,3.4776018,3.415869,3.1792276,3.6319332,4.266407,4.5990767,4.804852,4.90431,4.746549,4.90431,5.2918534,5.693115,5.9983487,6.1801167,6.5710897,6.5779486,6.5882373,6.8557453,7.4765005,8.001227,8.361334,8.580828,8.601405,8.285883,7.8091707,7.6274023,7.332458,7.0203657,7.2638664,7.798882,8.309891,8.718011,9.006097,9.201583,9.6645775,10.449953,10.851214,10.957532,11.64345,12.288212,12.953552,13.4474125,13.862392,14.555169,15.995596,17.364002,18.53692,19.384027,19.775002,19.288,18.825006,18.362011,17.943602,17.700102,17.576635,17.189093,17.021042,17.384579,18.434032,19.312008,20.11796,20.958208,21.637268,21.637268,21.342323,21.10568,20.954779,21.153696,22.216867,22.998814,23.924803,24.658733,25.073713,25.269201,28.650774,30.42044,31.76484,35.022945,43.70323,27.930561,18.825006,11.351934,5.23698,4.945465,6.1046658,5.212973,4.3452873,4.557922,5.888602,7.9292064,8.7317295,10.062409,10.4533825,5.219832,3.508468,4.931747,7.98408,11.125582,12.785502,14.373401,14.1299,13.690913,13.574307,13.183334,13.087306,13.694343,14.712931,15.858413,16.859852,18.533491,18.612371,18.241976,18.46147,20.217419,21.647556,21.894485,21.393766,20.570665,19.850452,19.936192,20.087093,20.152256,19.8676,18.828436,18.512913,19.21255,20.162544,21.266872,23.087982,25.162884,26.284359,26.212337,24.77191,21.86705,20.512363,19.713268,19.476627,19.613811,19.761284,19.809298,21.551527,19.641247,14.5414505,12.528283,10.597425,10.336777,9.774324,8.690575,8.604835,9.301042,8.906639,7.298162,5.9160385,7.795452,6.601956,6.64997,7.56567,8.436785,7.829748,7.6445503,7.8091707,7.534804,7.0752387,7.720001,8.405919,8.217292,7.9875093,7.864044,7.3393173,7.997798,8.457363,8.676856,8.615124,8.224151,7.5039372,8.056101,8.495089,8.477941,8.697433,8.940934,9.177576,9.39707,9.668007,10.131001,10.425946,9.455373,8.22758,7.284444,6.697984,6.783724,6.5230756,6.101236,5.6793966,5.3878818,5.3981705,5.7308407,6.1286726,6.4373355,6.608815,6.252138,6.1458206,5.830299,5.24041,4.715683,4.616225,4.530485,4.4687524,4.4413157,4.4413157,5.0003386,5.2781353,5.6656785,6.252138,6.852316,7.143831,7.099246,6.975781,6.9346256,7.0203657,6.715132,6.5813785,6.492209,6.358455,6.1492505,5.9297566,5.638242,5.336438,5.1409516,5.2026844,5.9469047,6.5196457,6.848886,7.0203657,7.2638664,7.459353,7.5450926,7.514226,7.548522,8.011517,8.340756,8.323608,8.347616,8.7145815,9.644,10.316199,10.875222,11.2593355,11.393089,11.183885,10.978109,11.228469,11.763485,12.418536,13.015285,13.358243,13.505715,13.433694,13.114742,12.528283,12.723769,13.485138,14.706071,15.409137,13.749216,12.528283,11.8115,12.085866,13.341095,15.076467,16.7844,17.466888,18.248835,19.360022,20.141968,17.566347,11.712041,6.632822,5.329579,9.736599,9.369633,7.3084507,7.298162,10.096705,13.488567,16.774113,19.123379,21.143406,22.546108,22.155134,22.36434,23.009102,22.6147,21.260014,20.61525,18.941612,17.717249,17.051908,16.911295,17.1205,17.778982,19.188541,20.409475,20.649546,19.257133,17.497755,16.163645,15.601193,15.902997,16.890718,16.328266,16.520323,16.739817,16.942162,17.761833,18.492336,19.023922,19.250275,19.5315,20.6907,21.801888,19.689262,18.108221,16.184223,8.4093485,3.2683969,1.2963841,0.9911508,1.155771,0.90198153,2.0474637,3.4227283,5.07236,6.7459984,7.905199,9.527394,10.593996,11.331357,11.526843,10.511685,10.182446,8.48137,6.5196457,4.839148,3.3884325,2.0920484,3.059192,5.562791,7.7440085,6.6225333,5.4016004,2.651071,1.845118,3.0489032,2.9151495,2.510458,2.393852,2.668219,3.4467354,4.835718,4.7019644,4.386442,3.3472774,2.07833,2.0920484,1.821111,1.9548649,2.2978237,2.527606,2.1983654,3.0043187,2.9940298,3.0317552,3.525616,4.4413157,4.5270553,5.4084597,5.7068334,5.4633327,6.135532,5.645101,6.2487082,7.0889573,7.716572,8.056101,9.777754,10.336777,10.782623,11.605724,12.740917,14.363112,15.29253,15.512024,15.145059,14.448852,14.291091,14.829536,15.278812,15.532601,16.143068,15.885849,15.3302555,14.829536,14.733508,15.3817,15.940722,16.064188,16.2974,16.269962,14.695783,13.3033695,12.010415,11.444533,11.71547,12.435684,13.21763,13.430264,13.985858,14.977009,15.6869335,16.71238,17.7927,18.982767,20.04251,20.4472,20.762722,22.419212,24.590141,25.258911,21.19485,20.899906,22.017952,22.244305,22.299177,25.924252,26.448978,25.18003,22.089973,18.008764,14.603184,13.419975,12.902108,12.408247,11.410237,9.506817,8.934075,8.81747,8.89635,9.2153015,10.131001,10.449953,10.281903,10.069269,9.853205,9.294182,9.571979,9.846346,10.199594,10.652299,11.153018,11.619442,12.229909,11.897239,10.679735,9.750318,8.934075,8.152129,7.4936485,7.1952744,7.658269,8.549961,9.342196,10.268185,11.180455,11.537132,11.327928,11.2593355,10.666017,9.379922,7.720001,8.429926,8.577398,8.419638,8.093826,7.630832,6.1766872,5.411889,5.2781353,5.470192,5.446185,5.2164025,5.552502,6.39961,7.4353456,8.073249,0.20234565,0.2194936,0.22292319,0.19548649,0.14061308,0.11317638,0.1097468,0.1097468,0.116605975,0.12346515,0.11317638,0.10288762,0.09602845,0.09602845,0.1097468,0.12689474,0.12003556,0.11317638,0.116605975,0.14061308,0.17147937,0.16119061,0.15433143,0.14061308,0.13032432,0.15776102,0.16119061,0.16462019,0.15776102,0.14404267,0.13032432,0.17833854,0.1920569,0.22292319,0.26064864,0.20920484,0.20234565,0.1920569,0.19891608,0.20920484,0.20234565,0.18519773,0.20577525,0.23321195,0.2709374,0.33609957,0.4081209,0.4081209,0.39783216,0.42183927,0.5041494,0.6036074,0.7305021,0.96714365,1.2415106,1.3341095,1.6770682,1.7662375,1.9068506,2.1023371,2.0508933,1.8073926,2.1194851,2.9082901,3.7519686,3.9097297,3.690236,4.0606318,4.73969,5.3981705,5.658819,3.0283258,1.728512,0.85739684,0.17490897,0.08573969,0.14747226,0.17833854,0.16804978,0.11317638,0.01371835,0.037725464,0.26750782,0.5624523,0.8711152,1.2415106,1.2895249,0.8265306,0.39440256,0.18519773,0.0548734,0.030866288,0.061732575,0.1097468,0.12003556,0.030866288,0.09259886,0.09259886,0.08573969,0.12003556,0.2503599,0.1097468,0.0548734,0.034295876,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.08916927,0.07545093,0.11317638,0.20920484,0.26064864,0.05144381,0.20577525,0.2503599,0.24350071,0.24007112,0.28122616,0.16804978,0.19891608,0.22635277,0.2469303,0.39783216,0.72021335,1.0871792,1.2106444,1.0700313,0.94999576,0.67219913,0.48700142,0.30866286,0.22292319,0.490431,0.5144381,0.5555932,0.59674823,0.6001778,0.50757897,0.72707254,0.5727411,0.66191036,0.91912943,0.59674823,0.8676856,0.6927767,0.4355576,0.29151493,0.26407823,0.24007112,0.3018037,0.34981793,0.36696586,0.38754338,0.3841138,0.25721905,0.17833854,0.19548649,0.22635277,0.20577525,0.22292319,0.2777966,0.32238123,0.26407823,0.2194936,0.2709374,0.2777966,0.29494452,0.5624523,0.45613512,0.31895164,0.30866286,0.3841138,0.3018037,0.47328308,0.51100856,0.48357183,0.53158605,0.85396725,0.7682276,0.70649505,0.65505123,0.6207553,0.64819205,0.805953,0.864256,1.0014396,1.2655178,1.5844694,1.5398848,1.7559488,1.9514352,2.0063086,1.9685832,2.0406046,2.1023371,2.194936,2.335549,2.5310357,2.9734523,3.093488,3.0077481,2.901431,3.0214665,3.8137012,4.5647807,4.9351764,4.8837323,4.695105,5.079219,5.31929,5.5147767,5.754848,6.094377,6.2418494,6.2967224,6.4236174,6.759717,7.390761,7.9737906,8.31332,8.464222,8.529384,8.652849,8.838047,8.89635,8.508806,7.932636,7.970361,8.381912,8.7283,9.218731,9.80862,10.189304,10.593996,11.101575,11.417097,11.612583,12.130451,13.011855,13.495427,13.660047,13.7938,14.363112,15.481158,16.582056,17.429163,18.053349,18.773561,18.999914,18.9519,18.605513,18.070496,17.590355,17.720678,17.55263,17.250826,17.086205,17.432592,18.30028,19.089085,19.764713,20.145397,19.891607,19.901896,20.025362,20.241425,20.731855,21.86362,23.297188,23.907654,24.669024,25.725336,26.380386,27.827673,30.218096,31.58307,35.972942,53.491276,42.454865,27.302946,13.88983,5.967482,5.1752477,5.9743414,4.290414,3.340418,4.1600895,5.597087,8.241299,10.175586,12.874671,15.028452,12.566009,7.548522,8.052671,10.851214,13.749216,15.594335,17.689812,17.929884,17.799559,17.837284,17.652086,17.20281,16.88043,17.137648,18.04649,19.29143,20.601532,21.44521,20.941061,19.425184,18.44775,18.588364,19.346302,20.141968,20.61182,20.632399,20.35803,19.630959,19.339443,19.346302,18.523201,18.674105,18.70154,18.897026,19.761284,22.000803,23.499533,23.94195,23.78419,23.11542,21.69557,21.297739,20.937632,20.666695,20.714708,21.506943,20.968498,21.085104,19.493774,15.858413,11.880091,10.401938,10.264755,9.904649,9.1810055,9.386781,9.97667,10.278474,9.585697,8.615124,9.517105,10.089847,9.966381,9.616563,8.505377,5.0826488,5.267846,5.967482,6.2830043,6.279575,6.975781,7.2021337,7.390761,7.4970784,7.4627824,7.2295704,7.2638664,7.5279446,7.8606143,8.073249,7.956643,8.06639,8.289313,8.344186,8.279024,8.477941,8.584257,8.501947,8.505377,8.639131,8.690575,8.711152,8.31675,7.6514096,6.914048,6.358455,6.001778,5.857735,5.861165,5.826869,5.446185,5.312431,5.192395,5.113515,5.2266912,5.7891436,5.3878818,5.456474,5.5250654,5.2987127,4.6676683,4.605936,4.506478,4.417309,4.32128,4.1360826,4.619654,5.470192,6.2658563,6.7322803,6.7665763,6.776865,6.835168,6.632822,6.2487082,6.1286726,5.9400454,6.0635104,6.3138704,6.4579134,6.210983,5.970912,5.6793966,5.422178,5.254128,5.2266912,5.8165803,6.444195,6.831738,7.0032177,7.274155,7.363324,7.4524937,7.3118806,7.034084,7.010077,7.0958166,7.082098,7.2535777,7.846896,9.057541,9.866923,10.329918,10.587136,10.618003,10.244178,10.155008,10.501397,11.091286,11.996697,13.55373,13.766364,14.023583,13.989287,13.653188,13.320518,12.950122,13.203912,13.63604,13.773223,13.138749,12.826657,12.05843,11.543991,11.787492,13.063298,15.755525,17.4566,18.36887,19.03764,20.337454,20.272291,16.05733,10.251037,5.802862,6.060081,5.4324665,5.65539,5.8200097,6.660259,10.569988,14.527733,16.753534,18.910746,21.006224,21.386908,21.993944,22.288889,22.021381,21.19485,20.04251,17.820137,16.365992,16.03675,16.585485,17.144508,18.45804,20.347742,21.61669,21.630407,20.306587,18.763273,16.87357,15.515453,15.29253,16.523752,16.208231,16.671225,17.134218,17.508043,18.38259,18.814716,19.078794,19.891607,21.187992,22.144846,17.754974,12.46998,11.941824,13.786942,7.5519514,3.2443898,2.6064866,4.029765,4.8117113,1.155771,1.0837497,2.5584722,4.0880685,5.830299,9.589127,14.201921,14.692352,14.1299,12.88839,8.683716,7.64798,6.6122446,5.689686,5.2026844,5.693115,2.8465576,4.5922174,7.870903,9.472521,6.025785,2.5378947,1.039165,1.0425946,1.587899,1.2175035,1.4781522,1.8348293,2.3561265,2.9974594,3.5804894,3.7176728,3.6147852,2.9734523,2.1846473,2.335549,1.920569,2.2669573,2.510458,2.4967396,2.7711067,3.216953,2.9563043,2.9117198,3.3301294,3.7553983,4.4859004,5.055212,5.4839106,5.8337283,6.183546,5.7822843,6.464772,7.2124224,7.699424,8.275595,9.674867,10.336777,11.012405,11.869802,12.4974165,13.426835,13.917266,14.212211,14.2533655,13.694343,13.622321,14.400838,15.018164,15.158776,15.193072,14.692352,14.071597,13.872682,14.2190695,14.805529,14.774663,15.193072,15.611482,15.645778,15.001016,13.9481325,13.125031,12.864383,13.251926,14.109323,14.13676,14.119612,14.057879,14.13676,14.695783,16.386568,18.344864,19.696121,20.364891,21.081675,20.169403,20.467777,22.77589,25.629307,25.282919,23.585274,23.835632,22.926792,21.215427,22.556396,24.888515,24.94682,23.20802,20.28258,16.935303,15.182784,14.143619,12.723769,10.734609,8.906639,8.676856,8.615124,8.666568,8.875772,9.410788,10.062409,10.1652975,9.788043,9.14328,8.621983,8.666568,9.071259,9.489669,9.777754,9.993818,10.086417,10.5597,10.628291,10.120712,9.506817,8.971801,8.416207,7.846896,7.5039372,7.829748,8.594546,9.170717,9.482809,9.695444,10.206452,10.700313,10.412228,9.280463,7.7714453,6.842027,7.2364297,7.7542973,7.9772205,7.5416627,6.138962,5.360445,5.0929375,5.0620713,5.0483527,4.897451,4.7259717,4.863155,5.90575,7.4799304,8.2310095,0.23664154,0.18519773,0.15433143,0.13032432,0.106317215,0.106317215,0.12003556,0.12346515,0.1371835,0.15090185,0.12346515,0.106317215,0.12346515,0.12346515,0.11317638,0.1371835,0.14747226,0.14061308,0.15776102,0.18862732,0.17490897,0.14747226,0.14747226,0.14747226,0.14747226,0.17833854,0.17833854,0.16462019,0.15433143,0.14747226,0.15776102,0.21263443,0.20234565,0.19891608,0.20920484,0.18176813,0.16804978,0.18862732,0.18176813,0.15433143,0.1920569,0.19548649,0.21263443,0.26750782,0.33609957,0.37382504,0.3806842,0.39097297,0.42869842,0.48357183,0.53501564,0.70649505,0.96714365,1.1866373,1.3409687,1.5227368,1.7490896,1.9068506,2.1057668,2.2909644,2.2395205,1.9925903,2.4075704,3.0317552,3.4364467,3.2135234,3.858286,4.5030484,5.888602,7.7542973,8.848335,3.9063,1.5124481,0.490431,0.09945804,0.041155048,0.030866288,0.048014224,0.061732575,0.048014224,0.0,0.01371835,0.15776102,0.51100856,0.881404,0.8093826,0.69963586,0.42869842,0.23321195,0.14747226,0.034295876,0.017147938,0.030866288,0.05144381,0.0548734,0.01371835,0.041155048,0.044584636,0.048014224,0.09602845,0.24350071,0.19891608,0.15776102,0.13032432,0.1097468,0.06516216,0.01371835,0.0,0.017147938,0.044584636,0.044584636,0.010288762,0.0,0.017147938,0.0548734,0.08916927,0.106317215,0.22635277,0.24007112,0.1371835,0.09945804,0.16804978,0.14747226,0.11317638,0.12346515,0.19891608,0.19548649,0.25378948,0.26750782,0.28122616,0.4972902,0.8505377,1.1180456,1.2792361,1.2758065,1.0048691,0.8025235,0.5624523,0.30866286,0.18176813,0.40126175,0.34638834,0.39440256,0.5796003,0.69963586,0.29151493,0.8505377,0.6859175,0.64476246,0.8196714,0.5590228,0.5624523,0.50757897,0.4046913,0.30866286,0.35324752,0.22978236,0.25721905,0.33266997,0.37382504,0.32238123,0.2469303,0.17833854,0.16462019,0.19548649,0.20920484,0.23664154,0.25378948,0.28122616,0.3018037,0.28465575,0.2709374,0.29151493,0.30523327,0.32924038,0.44584638,0.34638834,0.31552204,0.42526886,0.53501564,0.31209245,0.47328308,0.4629943,0.45956472,0.5590228,0.7990939,0.65505123,0.7305021,0.8025235,0.8128122,0.8711152,1.138623,1.039165,1.0220171,1.2483698,1.6084765,1.4610043,1.5501735,1.6256244,1.6153357,1.6187652,1.9823016,2.020027,2.0097382,2.1126258,2.3767042,2.551613,2.7539587,2.901431,2.9563043,2.9322972,3.4467354,3.9097297,4.149801,4.201245,4.3007026,4.835718,5.120374,5.3673043,5.675967,6.0532217,6.368744,6.468202,6.550512,6.7528577,7.160979,7.6925645,8.124693,8.543102,8.992378,9.458802,9.606275,9.626852,9.39707,9.088407,9.153569,9.342196,9.561689,9.949233,10.504827,11.087856,11.38966,11.561139,11.739478,12.116733,12.956982,13.574307,14.006435,14.291091,14.579176,15.138199,15.6697855,16.12592,16.53404,16.911295,17.233677,17.892159,17.995045,17.878439,17.703531,17.45317,17.473747,17.484037,17.449741,17.412016,17.466888,17.78927,18.416885,18.800999,18.814716,18.732407,18.972477,19.37031,19.833303,20.37175,21.12283,22.77589,23.832203,24.970827,26.171183,26.719915,27.584171,29.583622,30.948597,35.218433,51.2689,50.809338,35.31103,18.091074,7.181556,5.3330083,4.4756117,3.0523329,2.6785078,3.6387923,4.8905916,7.3427467,9.331907,11.924676,14.452282,14.503725,10.041832,10.518545,13.073587,15.954441,18.512913,19.401176,19.37031,19.78529,20.831314,21.53438,20.460918,20.045938,20.183123,20.79016,21.812176,22.971376,24.171732,24.202599,22.885637,21.064526,18.410025,17.62122,18.252264,19.401176,19.709839,19.161106,18.509483,18.053349,18.008764,18.485476,19.339443,19.281141,18.86959,18.653526,19.174824,20.399187,21.139977,21.53438,21.506943,20.762722,20.53294,20.351171,20.104242,19.87789,19.963629,19.5315,19.905325,19.167965,16.283682,11.105004,10.323058,10.206452,10.168727,10.0041065,9.901219,10.463672,11.245617,10.755186,9.283894,8.886061,8.844906,9.129561,8.580828,6.9380555,4.8254294,4.482471,4.73969,4.979761,5.178677,5.90232,6.4373355,6.56766,6.5642304,6.632822,6.927767,7.39762,7.531374,7.805741,8.165848,8.045813,8.237869,8.47451,8.519095,8.378482,8.340756,8.134981,8.032094,7.953213,7.8606143,7.7542973,7.7714453,7.5759587,7.1026754,6.4716315,5.9983487,5.48734,5.3570156,5.518206,5.7136927,5.5079174,5.2266912,4.931747,4.6608095,4.5270553,4.722542,4.4275975,4.5990767,4.712253,4.605936,4.48933,4.4550343,4.523626,4.5339146,4.4721823,4.4996185,5.2781353,6.1972647,6.9071894,7.239859,7.2021337,7.0306544,6.8969,6.7459984,6.5059276,6.0703697,5.809721,5.9297566,6.108095,6.2487082,6.492209,6.0635104,5.669108,5.442755,5.40503,5.442755,5.802862,6.4133286,6.7528577,6.8557453,7.3050213,7.5210853,7.4284863,7.157549,6.8763227,6.7871537,6.475061,6.427047,6.5333643,6.9517736,8.124693,8.971801,9.438225,9.8429165,10.103564,9.72631,10.089847,10.751757,11.379372,12.116733,13.605173,13.71492,13.687484,13.574307,13.471419,13.54687,13.011855,13.344524,13.481709,13.094165,12.590015,12.895248,12.466551,12.068718,12.05843,12.421966,14.315098,16.331696,17.638369,18.37916,19.654966,19.86417,18.969048,15.522313,10.443094,7.010077,6.217842,5.079219,4.7774153,5.950334,8.680285,11.859513,13.533153,14.973578,16.540901,17.669235,18.37916,18.317427,18.001905,17.730967,17.590355,16.2974,15.388559,15.165636,15.776102,17.21653,19.819586,21.253153,21.69214,21.273731,20.093952,19.305147,17.638369,16.317978,15.865272,16.105343,16.317978,16.828985,17.19938,17.556059,18.584934,19.013634,19.36688,20.711279,22.079683,20.464348,14.366542,9.146709,9.73317,13.152468,8.529384,4.1635194,3.3747141,4.180667,4.461893,1.9342873,1.2037852,2.2155135,5.4941993,10.494537,15.577187,13.7938,16.149927,14.476289,8.237869,4.5442033,3.8788633,4.1600895,4.9488945,5.9126086,6.8385973,3.9851806,6.989499,9.239308,7.8503256,3.6593697,1.2758065,0.9294182,1.5090185,1.8691251,0.8128122,1.0768905,1.8965619,2.8225505,3.40901,3.199805,3.357566,3.2032347,2.760818,2.4075704,2.8637056,2.153781,2.3972816,2.760818,2.952875,3.2272418,3.8960114,3.7211025,3.5359046,3.6044965,3.6216443,4.695105,5.284994,5.662249,6.001778,6.3961806,6.5882373,6.9792104,7.486789,7.9943686,8.323608,9.441654,10.14129,10.768905,11.355364,11.585147,12.459691,12.854094,13.183334,13.522863,13.615462,13.097594,14.109323,14.826107,14.874121,15.3302555,15.361122,14.836395,14.493437,14.38369,13.858963,13.756075,14.081886,14.445422,14.675205,14.836395,14.428274,14.157337,14.356253,15.031882,15.87213,15.80011,15.29253,14.634049,14.287662,14.870691,16.300829,18.097933,19.764713,20.721567,20.306587,19.750994,19.740705,21.664703,24.85422,26.59988,26.10945,25.649885,24.422092,22.892496,22.820475,23.68473,23.125708,21.829325,20.028791,17.518333,15.728088,14.068168,12.250486,10.38479,8.988949,8.803751,8.591117,8.601405,8.841476,9.074688,9.403929,9.369633,9.019815,8.529384,8.179566,8.47451,8.9100685,9.153569,9.170717,9.239308,9.39021,9.736599,10.089847,10.185875,9.692014,9.22902,8.9100685,8.577398,8.309891,8.412778,9.057541,9.026674,8.831187,8.81061,9.112414,9.73317,9.325048,8.110974,6.708273,6.1561093,6.392751,7.267296,7.798882,7.366754,5.7308407,5.223262,5.120374,4.870014,4.413879,4.201245,4.4550343,5.0620713,6.15268,7.2432885,7.2535777,0.20920484,0.14061308,0.09945804,0.08573969,0.09259886,0.106317215,0.13032432,0.1371835,0.14747226,0.14747226,0.106317215,0.106317215,0.12346515,0.12346515,0.11317638,0.1371835,0.16804978,0.17147937,0.17833854,0.18176813,0.14404267,0.12689474,0.13375391,0.14061308,0.14747226,0.17147937,0.19891608,0.17833854,0.16462019,0.18176813,0.20234565,0.19548649,0.17490897,0.16119061,0.17147937,0.1920569,0.19548649,0.22978236,0.23321195,0.20577525,0.216064,0.25378948,0.29837412,0.36010668,0.4046913,0.37382504,0.39783216,0.4664239,0.5453044,0.61046654,0.64476246,0.91569984,1.1283343,1.3272504,1.5536032,1.8416885,1.9411465,2.07833,2.3081124,2.534465,2.503599,2.2909644,2.5584722,2.9974594,3.2992632,3.175798,4.2252517,5.456474,7.2535777,9.136421,9.764035,4.650521,1.6770682,0.35324752,0.05144381,0.010288762,0.017147938,0.010288762,0.0034295875,0.034295876,0.16462019,0.1371835,0.14747226,0.33952916,0.59674823,0.52815646,0.36010668,0.216064,0.20577525,0.26064864,0.1371835,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.06516216,0.14747226,0.19891608,0.19548649,0.17490897,0.15433143,0.1371835,0.0274367,0.0,0.030866288,0.07545093,0.07545093,0.01371835,0.0034295875,0.034295876,0.072021335,0.058302987,0.1371835,0.274367,0.2503599,0.09602845,0.09602845,0.16804978,0.1371835,0.09945804,0.116605975,0.20920484,0.28465575,0.42526886,0.5521636,0.61046654,0.5658819,0.864256,1.1832076,1.4164196,1.4335675,1.0906088,1.0494537,0.70649505,0.32924038,0.1371835,0.28465575,0.26064864,0.3566771,0.5796003,0.71678376,0.35324752,0.8265306,0.72364295,0.58988905,0.59331864,0.5212973,0.52472687,0.53844523,0.47328308,0.39440256,0.52472687,0.33266997,0.4046913,0.45270553,0.3841138,0.30523327,0.216064,0.16804978,0.15433143,0.15776102,0.14747226,0.1920569,0.2194936,0.2469303,0.2709374,0.2709374,0.26064864,0.32238123,0.34638834,0.31209245,0.31209245,0.26750782,0.32238123,0.45270553,0.5453044,0.41498008,0.48700142,0.44584638,0.5453044,0.7373613,0.6893471,0.7305021,0.8745448,0.9294182,0.91227025,1.039165,1.2415106,1.1454822,1.097468,1.2312219,1.4747226,1.5193073,1.6153357,1.6530612,1.6221949,1.605047,1.9239986,1.9239986,1.937717,2.1023371,2.3458378,2.335549,2.510458,2.719663,2.8534167,2.836269,3.07634,3.2889743,3.5153272,3.7965534,4.184097,4.6745276,5.0346346,5.3913116,5.809721,6.2864337,6.550512,6.8557453,7.0615206,7.1541195,7.239859,7.671987,8.093826,8.64599,9.225591,9.506817,9.798331,9.846346,9.767465,9.736599,9.990388,10.031544,10.220171,10.487679,10.813489,11.204462,11.423956,11.417097,11.499407,11.934964,12.956982,13.505715,14.092175,14.664916,15.227368,15.827546,16.04018,16.149927,16.403717,16.671225,16.427725,16.774113,16.894148,16.986746,17.075916,16.990177,16.839275,17.034761,17.429163,17.737827,17.549198,17.439453,17.86815,18.053349,17.981327,18.389448,18.629519,19.301718,20.141968,20.930773,21.496655,22.703869,24.260902,25.680752,26.805656,27.820814,29.405283,30.444448,31.0069,34.32674,46.80358,51.35121,38.84694,21.657845,8.790032,5.885172,4.2046742,2.884283,2.750529,3.7451096,4.9351764,7.205563,9.057541,11.029553,12.96727,14.033872,11.211322,11.523414,13.7938,16.835844,19.45262,19.905325,19.572655,19.826445,20.70785,20.934202,20.714708,21.513802,22.055677,22.079683,22.347193,23.643576,25.042849,25.9414,25.93111,24.792488,21.44178,18.993055,18.149376,18.54035,18.69811,17.782412,17.463459,17.175373,17.110212,18.214539,19.45262,19.977346,19.857311,19.322296,18.752985,19.222837,19.987637,20.61868,20.851892,20.574095,20.488356,20.183123,19.70641,19.089085,18.341434,17.432592,17.929884,18.235117,16.808409,12.168177,10.281903,9.685155,9.822338,10.22703,10.539123,11.290202,12.168177,11.598865,9.801761,8.831187,6.9209075,7.1129646,6.8626046,5.6485305,4.9831905,3.474172,3.3747141,3.5564823,3.7725463,4.6436615,5.360445,5.5319247,5.8645945,6.375603,6.40304,7.205563,7.596536,8.196714,8.865483,8.680285,8.666568,8.985519,9.084977,8.844906,8.56025,8.237869,8.001227,7.7611566,7.531374,7.4181976,7.5107965,7.2124224,6.6705475,6.0703697,5.638242,5.3878818,5.3844523,5.4084597,5.329579,5.1066556,5.195825,4.8254294,4.413879,4.07435,3.6079261,3.6456516,3.8685746,3.9680326,3.9165888,3.974892,4.064061,4.4447455,4.623084,4.681387,5.2747054,6.1732574,6.835168,7.2535777,7.4524937,7.4696417,7.3050213,7.016936,6.927767,6.9209075,6.4373355,6.0532217,6.0635104,6.186976,6.368744,6.800872,6.492209,5.9743414,5.535354,5.353586,5.4976287,5.888602,6.375603,6.574519,6.591667,7.023795,7.191845,6.9826403,6.7185616,6.56766,6.560801,6.108095,6.111525,6.2830043,6.632822,7.48336,8.2310095,8.800322,9.352485,9.760606,9.609704,10.120712,10.981539,11.784062,12.487128,13.395968,13.166186,13.059869,12.987847,12.946692,13.022143,12.7272,13.197053,13.361672,12.977559,12.644889,12.908967,12.586586,12.397959,12.542002,12.706621,13.419975,15.196502,16.849564,18.101362,19.569225,18.825006,19.342873,18.499195,15.484588,11.276484,9.225591,5.586798,4.07435,5.435896,7.4353456,9.866923,10.899229,11.547421,12.291641,13.087306,13.711491,13.738928,13.776653,14.092175,14.606613,14.712931,14.544881,14.637479,15.433144,17.271402,20.169403,21.236006,21.109112,20.306587,19.21255,19.164536,18.056778,17.055338,16.54433,16.105343,16.369421,16.523752,16.640358,17.051908,18.334574,18.739265,19.510923,20.735287,21.36633,19.233126,12.010415,8.4264965,11.1393,15.361122,8.851766,4.770556,3.3198407,3.391862,3.8548563,3.5393343,1.9102802,2.0234566,4.8185706,9.644,14.2533655,10.902658,12.521424,11.115293,6.101236,4.3349986,4.016047,4.623084,5.545643,6.5059276,7.5519514,7.1987042,9.784613,9.962952,6.7802944,3.6970954,2.085189,2.1400626,2.2326615,1.6633499,0.65848076,0.7922347,1.4267083,2.4007113,3.340418,3.666229,3.5633414,3.1826572,2.8739944,2.7916842,2.9048605,2.201795,2.5173173,2.8637056,3.0386145,3.642222,4.3692946,4.180667,3.8685746,3.7862647,3.8617156,4.911169,5.5730796,6.046363,6.351596,6.3481665,7.082098,7.3187394,7.579388,8.076678,8.707723,9.81205,10.535692,11.091286,11.427385,11.211322,11.753197,11.852654,12.085866,12.644889,13.351384,13.008426,13.701202,14.160767,14.363112,15.505165,16.11906,15.9921665,15.851553,15.553179,14.078457,13.680624,13.725209,13.886399,14.140189,14.757515,15.244516,15.337115,15.4914465,15.8138275,16.067617,16.173935,15.721229,15.206791,14.977009,15.22051,16.345413,17.412016,19.288,20.86904,19.068506,19.19197,19.757853,21.12283,23.44809,26.716486,28.040308,27.364677,25.982555,24.682741,23.729315,22.919933,21.397196,19.812727,18.252264,16.221949,14.723219,13.138749,11.622872,10.429376,9.897789,9.788043,9.462232,9.266746,9.273604,9.277034,9.112414,8.855195,8.309891,7.7268605,7.798882,8.40249,8.992378,9.174147,8.97866,8.889491,9.297611,9.633711,9.997248,10.213311,9.839486,9.469091,9.266746,9.0369625,8.848335,9.054111,9.414218,8.7145815,8.289313,8.491658,8.697433,9.078118,8.491658,7.390761,6.293293,5.7582774,6.1458206,7.06495,7.5588107,7.0375133,5.254128,4.99005,5.051782,4.8494368,4.417309,4.3795834,4.976331,5.8405876,6.697984,7.2192817,7.0203657,0.12689474,0.106317215,0.09259886,0.09259886,0.10288762,0.106317215,0.13032432,0.13375391,0.12689474,0.1097468,0.06859175,0.10288762,0.10288762,0.1097468,0.12689474,0.15090185,0.17147937,0.18176813,0.16462019,0.12346515,0.106317215,0.116605975,0.12346515,0.12346515,0.13032432,0.15090185,0.21263443,0.1920569,0.17833854,0.20234565,0.20920484,0.14404267,0.13375391,0.15433143,0.18862732,0.23321195,0.26064864,0.29494452,0.30866286,0.3018037,0.29151493,0.36696586,0.42526886,0.4629943,0.45270553,0.37382504,0.5007198,0.6241849,0.72707254,0.8025235,0.84367853,1.1317638,1.2277923,1.5055889,1.9548649,2.201795,2.253239,2.3595562,2.585909,2.8225505,2.7539587,2.6922262,2.7299516,3.1517909,3.765687,3.9303071,4.5956473,6.3207297,7.98408,8.707723,7.840037,4.2423997,1.6256244,0.30866286,0.041155048,0.0,0.030866288,0.024007112,0.01371835,0.09602845,0.432128,0.35324752,0.18862732,0.12003556,0.22292319,0.4629943,0.48014224,0.3566771,0.37725464,0.48700142,0.3018037,0.14747226,0.048014224,0.006859175,0.01371835,0.06516216,0.01371835,0.0,0.0034295875,0.017147938,0.037725464,0.09602845,0.13032432,0.12689474,0.11317638,0.17147937,0.0548734,0.010288762,0.0274367,0.061732575,0.061732575,0.01371835,0.006859175,0.034295876,0.058302987,0.0274367,0.116605975,0.20234565,0.20920484,0.14061308,0.058302987,0.16804978,0.23321195,0.22978236,0.20234565,0.26407823,0.48700142,0.77165717,1.0940384,1.2483698,0.8196714,0.922559,1.3478279,1.5844694,1.4781522,1.2312219,1.2655178,0.8265306,0.34638834,0.11317638,0.26750782,0.26407823,0.39440256,0.4972902,0.53158605,0.59674823,0.607037,0.6173257,0.548734,0.4629943,0.53844523,0.78537554,0.83338976,0.6962063,0.5453044,0.7099246,0.5727411,0.66876954,0.61389613,0.3841138,0.29151493,0.28465575,0.2194936,0.14747226,0.106317215,0.09945804,0.106317215,0.14747226,0.20577525,0.2503599,0.25721905,0.216064,0.3566771,0.39097297,0.28122616,0.26407823,0.28465575,0.32238123,0.36010668,0.4081209,0.5212973,0.53158605,0.4972902,0.66876954,0.89512235,0.6173257,0.94656616,1.0563129,0.9877212,0.90198153,1.0768905,1.0494537,1.1214751,1.1934965,1.2655178,1.4232788,1.7833855,2.0406046,2.1263442,2.0406046,1.8862731,1.8725548,1.8382589,1.9582944,2.2155135,2.428148,2.4007113,2.4247184,2.4898806,2.568761,2.6064866,2.74367,2.9631636,3.2615378,3.6387923,4.0880685,4.4447455,4.856296,5.3261495,5.8645945,6.478491,6.5642304,7.1232533,7.5553813,7.6445503,7.5245147,7.795452,8.069819,8.508806,8.951223,8.930646,9.499957,9.592556,9.551401,9.637141,10.017825,10.189304,10.532263,10.803201,10.882081,10.789482,10.779194,10.734609,10.840926,11.293632,12.30536,13.200482,14.068168,14.781522,15.340545,15.87899,16.11906,16.355703,16.770683,17.086205,16.55119,16.21166,16.239098,16.39,16.475739,16.369421,16.160215,16.520323,17.178804,17.689812,17.422304,17.29884,17.638369,17.88873,18.084215,18.821575,19.102802,20.015072,21.187992,22.264881,22.913074,23.1943,24.816494,26.226055,27.289227,29.271528,32.210686,31.730543,30.228384,32.255272,44.512615,49.48895,38.89838,23.043398,10.155008,6.3824625,5.3330083,3.8479972,3.3884325,4.262977,5.6245236,8.032094,9.942374,11.297061,12.229909,13.073587,11.873232,11.866373,13.615462,16.431154,18.406595,19.812727,19.586374,19.154245,18.756414,17.446312,19.03421,21.19828,22.086544,21.558388,21.20514,22.659285,24.041409,25.564144,26.77479,26.569014,24.795918,22.079683,19.932762,18.962189,18.852442,17.607502,17.425734,17.401728,17.415445,18.142517,19.267422,20.484926,20.999365,20.742146,20.382038,20.248285,20.676983,21.112541,21.36633,21.630407,21.78817,21.304598,20.430052,19.29143,17.926455,16.2974,16.434584,17.686382,18.423744,16.050468,11.859513,9.901219,9.373062,9.925226,11.646879,12.531713,12.871242,12.075578,10.532263,9.589127,6.4304767,6.0326443,6.0737996,5.5490727,4.7671266,2.5584722,2.2978237,2.4041407,2.5241764,3.542764,4.2526884,4.671098,5.6005163,6.6636887,6.307011,6.776865,7.3530354,8.333898,9.342196,9.335337,9.270175,9.616563,9.702303,9.349055,8.851766,8.755736,8.423067,8.052671,7.7542973,7.548522,7.507367,6.9963584,6.3207297,5.7136927,5.31929,5.377593,5.442755,5.1580997,4.6127954,4.3590055,4.8185706,4.420738,3.9646032,3.5702004,2.6853669,3.0729103,3.2203827,3.309552,3.350707,3.1826572,3.4192986,4.057202,4.482471,4.7979927,5.8200097,6.7048435,7.0786686,7.2192817,7.274155,7.250148,7.222711,6.9517736,6.8969,7.006647,6.7048435,6.3447366,6.245279,6.420188,6.759717,7.058091,7.082098,6.5059276,5.7377,5.209543,5.3878818,5.888602,6.210983,6.2830043,6.23499,6.3893213,6.334448,6.1286726,5.9812007,5.9640527,6.0154963,5.7925735,5.909179,6.2658563,6.7974424,7.4627824,8.165848,8.851766,9.349055,9.613133,9.740028,10.038403,10.89237,11.921246,12.795791,13.251926,12.768354,12.785502,12.768354,12.555719,12.356804,12.343085,12.723769,12.977559,12.991278,13.046151,12.902108,12.449403,12.30536,12.620882,13.073587,13.125031,14.582606,16.441442,18.20425,19.898466,18.509483,18.224829,18.643238,18.722118,16.780972,13.430264,7.73029,4.506478,4.955754,6.660259,8.447074,9.112414,9.225591,9.208443,9.318189,9.8429165,10.326488,10.988399,11.746337,12.22305,13.282792,13.63261,14.373401,15.817257,17.494326,19.62067,20.666695,20.416334,19.243416,18.12194,18.423744,17.95389,17.394867,17.024471,16.702091,16.599203,16.208231,16.064188,16.53747,17.833855,18.149376,19.37031,19.997925,19.442331,18.005335,10.690024,8.951223,13.817808,18.526632,8.515666,5.0312047,3.1072063,2.9082901,4.091498,5.8234396,3.3747141,2.6750782,2.784825,3.7451096,6.560801,7.4284863,6.711703,6.914048,8.038953,7.5931067,6.910619,7.085528,7.3873315,7.7680154,8.844906,12.298501,12.394529,9.798331,6.7357097,7.0032177,4.6265135,3.6010668,2.3732746,0.94999576,0.8779744,0.607037,0.7407909,1.5638919,2.9288676,4.273266,3.841138,3.3678548,3.2478194,3.2992632,2.7642474,2.4144297,2.8019729,2.860276,2.7470996,3.8377085,4.262977,4.07435,3.882293,3.9611735,4.249259,4.98662,5.593657,6.2658563,6.7391396,6.276145,7.099246,7.5450926,7.7885933,8.2310095,9.510246,10.912948,11.64345,12.075578,12.185325,11.561139,11.348505,11.180455,11.372512,12.0138445,12.953552,13.368532,13.440554,13.437123,13.783512,15.059319,15.765814,16.184223,16.811838,17.189093,15.916716,14.928994,14.572317,14.363112,14.376831,15.234227,16.341984,16.492886,16.156786,15.618341,14.973578,15.100473,15.223939,15.422854,15.563468,15.285671,16.317978,16.674654,18.293419,20.124819,18.11165,18.807858,20.165974,21.150267,22.288889,25.680752,27.913412,27.724785,26.383816,24.85079,23.773901,22.590693,20.738716,18.728977,16.780972,14.808959,13.337666,12.298501,11.434244,10.851214,11.026124,11.05699,10.909517,10.6317215,10.323058,10.127572,9.668007,9.177576,8.237869,7.284444,7.610255,8.275595,9.0644,9.366203,9.15014,8.97523,9.493098,9.887501,10.045261,9.97324,9.801761,9.582268,9.39021,9.174147,9.102125,9.544542,9.482809,8.453933,8.018375,8.460793,8.793462,8.882631,8.042382,7.157549,6.5196457,5.830299,6.451054,7.0752387,7.31531,6.6739774,4.5647807,4.465323,4.650521,4.791134,4.870014,5.192395,5.919468,6.6533995,7.157549,7.4353456,7.7268605,0.09259886,0.07888051,0.07545093,0.07545093,0.082310095,0.106317215,0.13032432,0.12003556,0.106317215,0.10288762,0.09259886,0.116605975,0.13032432,0.15433143,0.18519773,0.19891608,0.16119061,0.14404267,0.12003556,0.09602845,0.106317215,0.106317215,0.12346515,0.1371835,0.14061308,0.15090185,0.16462019,0.15776102,0.14747226,0.1371835,0.1371835,0.15090185,0.17833854,0.20577525,0.2194936,0.24350071,0.29151493,0.36010668,0.40126175,0.42869842,0.48700142,0.5624523,0.53501564,0.5144381,0.53158605,0.5178677,0.66533995,0.7305021,0.83338976,0.96714365,0.9911508,1.1146159,1.5193073,2.0680413,2.5310357,2.5790498,2.651071,2.8705647,2.9871707,2.8980014,2.6545007,3.3747141,3.4638834,3.683377,4.139512,4.273266,4.431027,5.8062916,7.291303,7.6205435,5.3878818,2.3458378,0.71678376,0.11317638,0.061732575,0.0,0.0,0.010288762,0.034295876,0.15090185,0.5178677,0.45613512,0.34295875,0.34638834,0.41498008,0.24350071,0.31895164,0.29837412,0.35324752,0.42526886,0.22978236,0.22978236,0.12003556,0.034295876,0.07545093,0.31895164,0.06516216,0.0,0.0,0.0,0.0,0.0,0.037725464,0.037725464,0.024007112,0.12346515,0.12346515,0.058302987,0.010288762,0.0,0.0,0.0,0.0,0.01371835,0.0274367,0.01371835,0.0274367,0.041155048,0.034295876,0.044584636,0.16804978,0.13032432,0.23321195,0.34295875,0.39783216,0.39783216,1.1283343,1.3478279,1.5570327,1.8348293,1.845118,1.7730967,1.9102802,1.8725548,1.611906,1.4027013,1.0734608,0.6241849,0.30866286,0.24350071,0.42869842,0.20920484,0.15090185,0.24350071,0.4115505,0.53501564,0.40126175,0.4664239,0.5212973,0.53844523,0.67219913,0.64819205,0.9328478,0.9774324,0.7339317,0.6859175,0.8196714,0.6241849,0.45956472,0.40126175,0.24350071,0.30523327,0.2469303,0.16804978,0.12346515,0.1371835,0.16119061,0.19548649,0.23321195,0.26750782,0.30523327,0.30523327,0.28808534,0.32238123,0.36353627,0.22978236,0.32581082,0.29494452,0.3566771,0.4972902,0.47328308,0.5212973,0.67219913,0.77508676,0.7510797,0.5796003,0.86082643,0.89512235,0.91912943,1.0151579,1.1146159,0.881404,0.9534253,1.0254467,1.1283343,1.6187652,1.9582944,2.1915064,2.2155135,2.0817597,1.9823016,1.862266,2.0131679,2.1674993,2.2326615,2.318401,2.369845,2.5721905,2.6407824,2.5447538,2.534465,2.644212,2.7813954,2.7813954,2.7059445,2.8534167,3.3301294,3.841138,4.48933,5.209543,5.7822843,6.358455,6.8385973,7.133542,7.257007,7.3530354,7.281014,7.4284863,7.7885933,8.368194,9.184435,9.211872,8.934075,8.848335,9.030104,9.139851,9.945804,10.768905,11.262765,11.314209,11.046701,10.254466,10.065839,10.374502,11.170166,12.511135,13.917266,14.990726,15.306249,15.097044,15.244516,15.4742985,15.964729,16.554619,16.955881,16.722668,16.527182,16.276823,16.204802,16.283682,16.235666,16.112202,16.496315,16.88386,17.154797,17.532051,17.799559,18.351723,19.071936,19.678972,19.713268,20.776442,21.764162,22.594122,23.242313,23.743034,23.204588,24.19574,25.3618,26.538147,28.746801,32.361588,29.381275,24.408375,25.3618,43.487167,57.671944,41.453423,21.462358,10.093276,5.4770513,5.610805,4.6848164,3.8788633,4.0263357,5.6005163,8.261876,10.30934,11.149589,11.317638,12.452832,13.426835,13.937843,14.589465,15.731518,17.439453,19.94305,20.385468,20.056227,19.425184,18.142517,19.730417,20.62211,20.731855,20.53637,21.071384,22.134558,22.875349,23.94538,24.761621,23.5304,22.381487,21.85676,21.380049,20.941061,21.088533,19.977346,19.514353,19.270851,19.19197,19.60695,20.351171,21.187992,20.797018,19.490345,19.21255,20.639257,21.482935,22.011093,22.546108,23.437801,23.389786,23.228596,22.264881,20.392326,18.097933,17.425734,18.073925,19.95677,22.127699,22.751883,18.307138,13.735497,10.587136,10.168727,13.5503,13.831526,12.617453,11.338216,10.295622,8.697433,7.548522,7.133542,7.023795,6.5230756,4.6676683,4.180667,3.1346428,2.3835633,2.369845,3.1277838,4.420738,4.9660425,5.4839106,6.4304767,7.98065,7.4936485,6.958633,7.1232533,7.98065,8.772884,9.239308,9.582268,9.599416,9.194724,8.378482,8.766026,9.112414,9.071259,8.56368,7.781734,7.0375133,6.5024977,5.9126086,5.31929,5.1100855,4.671098,4.1600895,3.6593697,3.4433057,3.9680326,3.234101,2.952875,2.8465576,2.6853669,2.2566686,2.4795918,2.2498093,2.1812177,2.3767042,2.4247184,2.585909,3.0900583,3.9028704,4.746549,5.1100855,6.468202,6.941485,6.9620624,6.800872,6.591667,6.6533995,6.475061,6.475061,6.5813785,6.2418494,6.2898636,6.118384,6.2041235,6.667118,7.2775846,7.205563,6.691125,5.9983487,5.4496145,5.4633327,5.4633327,5.720552,5.895461,5.8543057,5.645101,5.610805,5.3707337,5.2438393,5.2815647,5.295283,5.501058,5.610805,5.909179,6.6568294,8.073249,9.242738,9.866923,9.97667,9.815479,9.825768,10.096705,10.902658,11.842365,12.7272,13.581166,13.862392,13.584596,13.155897,12.881531,12.953552,12.538571,12.528283,12.614022,12.668896,12.740917,12.754636,12.572867,12.590015,12.696333,12.267634,12.572867,14.46257,16.499744,17.95732,18.79757,19.12681,18.825006,18.821575,19.490345,20.676983,19.308577,12.63117,7.7542973,6.694555,6.3790326,6.293293,7.2432885,6.9792104,6.0223556,7.6445503,8.268735,9.016385,9.712592,10.401938,11.369082,12.075578,12.490558,14.023583,16.530611,18.324286,20.107672,20.975357,20.231136,18.37916,17.1205,17.21653,17.408587,17.62122,17.775553,17.775553,17.751545,17.233677,16.952452,17.137648,17.518333,17.919594,19.044498,19.576086,17.943602,12.329367,10.034973,9.277034,13.395968,17.806417,9.993818,6.135532,4.3487167,3.275256,3.625074,8.179566,6.444195,5.9297566,5.329579,4.8151407,6.012067,4.5853586,6.9552035,8.872343,8.64256,7.140401,5.0895076,6.1972647,9.0369625,11.736049,11.993267,17.20624,14.123041,7.970361,4.7328305,11.153018,7.7714453,3.3678548,1.2860953,1.9274281,2.7470996,0.9877212,1.611906,2.9117198,3.7725463,3.6627994,3.2718265,3.3472774,3.5976372,3.8034124,3.8137012,3.8274195,3.4192986,3.0043187,2.9082901,3.3712845,3.5050385,4.0057583,4.5613513,4.846007,4.5167665,4.8940215,5.219832,5.7754254,6.5230756,7.0958166,7.291303,8.2653055,9.0644,9.544542,10.374502,12.267634,12.922686,12.881531,12.46312,11.780633,11.012405,11.595435,12.298501,12.734058,13.38225,13.893259,14.112752,14.023583,13.780083,13.718349,13.680624,14.332246,15.923574,17.87158,18.739265,17.4566,16.55119,15.659496,15.258235,16.660936,17.12736,17.04848,16.54433,15.741806,14.802099,14.311668,14.658057,15.073037,15.21365,15.151917,15.920145,16.304258,16.739817,17.357141,17.991615,19.565796,20.755863,21.891056,22.642136,22.017952,23.228596,24.336353,23.924803,22.590693,22.919933,22.6147,21.428062,19.86074,18.276272,16.921585,14.249936,12.977559,12.21962,11.550851,11.002116,11.002116,11.550851,12.044711,12.130451,11.701753,11.410237,10.477389,9.431366,8.587687,8.025234,8.320179,8.988949,9.39021,9.427936,9.537683,9.585697,9.901219,9.904649,9.644,9.764035,9.595985,9.451943,9.547972,9.801761,9.825768,9.410788,8.858624,8.388771,8.23444,8.635701,8.783174,7.7680154,7.222711,7.298162,6.636252,6.941485,7.2192817,7.48336,7.0443726,4.5167665,4.016047,3.9200184,4.125794,4.557922,5.1409516,5.960623,6.715132,7.1849856,7.4456344,7.874333,0.20234565,0.18862732,0.1920569,0.20920484,0.22635277,0.24007112,0.216064,0.17833854,0.15433143,0.14747226,0.116605975,0.13032432,0.12003556,0.13032432,0.15433143,0.1371835,0.1097468,0.10288762,0.09602845,0.09602845,0.12003556,0.1371835,0.14747226,0.15090185,0.15090185,0.16462019,0.16804978,0.14404267,0.14061308,0.16462019,0.17490897,0.19548649,0.26407823,0.35324752,0.4355576,0.5007198,0.48014224,0.52472687,0.52815646,0.5041494,0.5727411,0.58988905,0.5624523,0.5624523,0.6001778,0.6276145,0.83338976,0.86082643,0.9877212,1.2689474,1.5158776,1.6496316,2.1091962,2.4418662,2.5413244,2.627064,3.2683969,3.4364467,3.4947495,3.5187566,3.3129816,3.450165,3.426158,3.6182148,3.9851806,4.0880685,4.3452873,5.3501563,7.2947326,9.1810055,8.851766,3.4227283,1.1351935,0.94656616,1.5124481,1.196926,0.25721905,0.06859175,0.12003556,0.25378948,0.6893471,0.4046913,0.2469303,0.26407823,0.33952916,0.20920484,0.4355576,0.48014224,0.4115505,0.32581082,0.31552204,0.26407823,0.1371835,0.13032432,0.20577525,0.08916927,0.017147938,0.2503599,0.26750782,0.037725464,0.0,0.34981793,0.18176813,0.006859175,0.017147938,0.08573969,0.14404267,0.07888051,0.020577524,0.010288762,0.0,0.020577524,0.017147938,0.010288762,0.006859175,0.01371835,0.017147938,0.12346515,0.18862732,0.18519773,0.17833854,0.14404267,0.22978236,0.31895164,0.4389872,0.7510797,1.0837497,1.2106444,1.5776103,2.0165975,1.7353712,1.8279701,1.7525192,1.5981878,1.4232788,1.2449403,1.0425946,0.764798,0.4629943,0.22978236,0.20920484,0.17490897,0.20920484,0.29494452,0.36696586,0.31552204,0.18176813,0.47328308,0.5590228,0.45270553,0.82996017,0.7476501,0.83681935,1.0151579,1.1043272,0.8196714,1.0837497,0.82996017,0.59674823,0.52815646,0.37725464,0.33266997,0.2469303,0.21263443,0.22635277,0.20920484,0.18519773,0.19891608,0.20920484,0.21263443,0.26750782,0.31895164,0.29494452,0.32924038,0.39097297,0.31552204,0.34295875,0.3841138,0.41498008,0.432128,0.4355576,0.4355576,0.6756287,0.7407909,0.5693115,0.44584638,0.6001778,0.64476246,0.77165717,1.0117283,1.2346514,1.471293,1.3169615,1.2243627,1.3341095,1.471293,1.6667795,1.8965619,2.020027,1.99602,1.8965619,1.8142518,1.9102802,2.0749004,2.3321195,2.8568463,2.8156912,2.6407824,2.4384367,2.301253,2.287535,2.3286898,2.6853669,2.8945718,2.884283,2.9631636,3.0969174,3.6216443,4.1017866,4.5030484,5.1855364,5.98463,6.3173003,6.5127864,6.636252,6.4990683,6.8763227,6.8728933,7.006647,7.442205,7.9772205,7.9429245,7.966932,7.905199,7.939495,8.567109,9.547972,10.2921915,10.868362,11.187314,10.998687,10.693454,10.772334,11.1393,11.718901,12.476839,13.773223,14.973578,15.426285,15.37827,15.964729,16.263103,16.63007,16.911295,16.969599,16.698662,16.931873,17.19938,17.429163,17.562918,17.55263,16.993607,17.079346,17.45317,17.885298,18.313997,18.650097,18.903887,19.46291,20.186552,20.399187,20.78673,21.644127,22.745024,23.832203,24.583282,24.144297,24.03455,24.312346,24.915953,25.670462,27.625326,25.821363,24.072275,26.85024,39.265347,39.014988,32.958336,22.237446,10.703742,4.866585,5.188966,4.4447455,4.0194764,4.482471,5.586798,7.7131424,9.616563,10.878652,11.266195,10.741467,11.358793,12.30536,13.440554,14.870691,16.938732,18.886738,19.46634,19.61038,19.713268,19.644676,19.912186,19.816156,19.637817,19.562366,19.668684,20.467777,20.975357,21.668133,22.43979,22.6147,22.374628,22.419212,22.607841,22.823904,22.978235,22.727877,22.930222,22.94394,22.44322,21.414345,21.0268,21.301168,21.578964,21.726437,22.127699,21.993944,22.158566,22.662714,22.957659,21.935642,19.222837,18.893597,18.78042,18.04992,17.230247,17.995045,18.818146,18.756414,18.331144,19.54179,15.673215,13.166186,11.729189,11.423956,12.644889,12.46998,11.0981455,9.966381,9.640571,9.80862,8.584257,8.06639,7.4353456,6.2418494,4.4241676,4.307562,3.7794054,3.4364467,3.2786856,2.6887965,3.865145,4.8322887,5.669108,6.574519,7.870903,8.093826,8.076678,8.045813,7.891481,7.160979,7.822889,8.412778,8.934075,9.23245,8.999237,8.882631,8.4264965,7.596536,6.591667,5.8405876,5.2438393,5.2644167,4.911169,4.1463714,3.8788633,3.5187566,3.0317552,2.6545007,2.452155,2.3321195,1.8348293,1.8725548,1.920569,1.7833855,1.611906,1.6736387,1.6942163,1.7216529,1.7936742,1.8999915,2.4590142,2.8534167,3.7005248,4.791134,5.086078,6.6465406,7.233,7.222711,6.927767,6.591667,6.416758,6.0737996,5.844017,5.8200097,5.885172,6.0223556,6.1732574,6.392751,6.715132,7.1678376,6.831738,6.142391,5.453044,5.020916,5.0243454,5.1512403,5.2918534,5.254128,5.07236,5.0106273,5.0414934,5.120374,5.130663,5.127233,5.3570156,5.6210938,6.169828,6.711703,7.1987042,7.8023114,9.081548,10.1481495,10.494537,10.281903,10.364213,10.535692,11.129011,11.869802,12.548861,13.032433,13.351384,13.536582,13.399398,12.860953,11.965831,12.264205,12.9638405,13.529722,13.577737,12.898679,12.679185,12.439114,12.432255,12.555719,12.3533745,12.562579,14.167625,15.906426,17.195951,18.176813,18.78042,19.263992,19.219408,18.818146,18.821575,20.11796,18.825006,17.267973,15.29253,10.247607,6.0806584,4.976331,4.5819287,4.6608095,7.0958166,9.613133,12.133881,13.951562,14.71636,14.4317045,14.143619,14.222499,16.060759,19.356592,22.096832,21.644127,21.723007,21.112541,19.692692,18.46147,18.080786,18.307138,18.87645,19.62753,20.484926,20.27572,19.761284,19.486916,19.37374,18.739265,18.62266,18.9519,19.078794,18.550638,17.113642,14.613472,13.5503,14.891269,16.245956,11.862943,8.47451,5.593657,3.8891523,3.8788633,5.9331865,5.312431,6.6568294,5.7479887,3.391862,5.439326,8.083538,8.577398,7.9120584,6.931196,6.3481665,5.672538,6.7391396,8.591117,9.921797,9.0644,11.279913,8.488229,4.6745276,3.974892,10.679735,9.650859,4.2938433,1.3684053,2.2258022,2.819121,2.3492675,4.3933015,5.127233,4.0709205,4.0777793,4.9660425,4.996909,5.055212,5.288424,5.096367,5.0106273,4.5784993,4.5201964,4.8597255,4.9351764,5.2164025,5.8200097,6.2041235,6.2898636,6.468202,6.416758,6.5333643,6.927767,7.3530354,7.205563,8.131552,9.040393,9.880642,10.439664,10.350495,11.979549,12.562579,12.418536,11.924676,11.537132,11.1393,11.135871,11.650309,12.655178,13.954991,14.332246,14.30481,14.321958,14.421415,14.243076,14.057879,14.356253,15.45715,17.103354,18.468328,17.840714,17.243965,16.609491,16.242527,16.846134,17.504614,17.367432,16.475739,15.182784,14.167625,12.836946,13.193623,14.13676,14.942713,15.261664,15.827546,15.762384,15.909856,16.79469,18.650097,19.997925,22.151705,23.598991,23.44809,21.407484,21.133118,21.019941,20.37518,19.582945,20.087093,21.150267,21.184563,20.433481,19.185112,17.799559,15.916716,13.591455,12.38424,12.377381,12.161317,12.308789,13.238208,13.96185,13.965281,13.21763,11.441104,9.928656,9.253027,9.235879,8.964942,8.769455,8.378482,8.097256,8.014946,7.997798,8.107545,8.464222,8.752307,8.940934,9.277034,9.0369625,8.64256,8.522525,8.868914,9.654288,9.884071,9.770895,9.493098,9.403929,10.041832,8.868914,7.963502,7.716572,7.9086285,7.6857057,7.7371492,7.5725293,7.4353456,6.776865,4.2595477,4.0434837,4.0606318,4.3658648,4.962613,5.802862,6.5127864,7.394191,8.004657,8.299602,8.618553,0.2469303,0.22635277,0.20920484,0.216064,0.24350071,0.25721905,0.26407823,0.22978236,0.216064,0.216064,0.15776102,0.17147937,0.15433143,0.14404267,0.14061308,0.12346515,0.106317215,0.09945804,0.11317638,0.1371835,0.17833854,0.15776102,0.16804978,0.17490897,0.17147937,0.17833854,0.21263443,0.216064,0.22292319,0.2469303,0.274367,0.36353627,0.45613512,0.5178677,0.5453044,0.5453044,0.4938606,0.52815646,0.59674823,0.66876954,0.7407909,0.7476501,0.7133542,0.70306545,0.7339317,0.7579388,0.90198153,1.039165,1.1900668,1.3752645,1.6290541,1.8725548,2.3286898,2.6407824,2.8259802,3.2889743,3.8445675,3.7931237,3.806842,3.9680326,3.7725463,3.532475,3.542764,3.8274195,4.2869844,4.6848164,5.2506986,5.675967,7.133542,9.242738,10.048691,3.6387923,1.1146159,1.3581166,2.3835633,1.3409687,0.432128,0.26064864,0.274367,0.432128,1.2003556,0.99801,0.4629943,0.14747226,0.14404267,0.08916927,0.5761707,1.0082988,1.0151579,0.70306545,0.6379033,0.69963586,0.4389872,0.216064,0.1371835,0.041155048,0.10288762,0.24350071,0.25378948,0.116605975,0.010288762,0.17833854,0.08916927,0.006859175,0.034295876,0.10288762,0.20577525,0.12689474,0.037725464,0.006859175,0.010288762,0.048014224,0.030866288,0.01371835,0.010288762,0.01371835,0.08916927,0.22978236,0.22635277,0.1097468,0.1371835,0.2469303,0.29494452,0.32238123,0.40126175,0.6379033,0.5693115,0.6036074,0.823101,1.1043272,1.1214751,1.2998136,1.2758065,1.2895249,1.3958421,1.4541451,1.0563129,0.6756287,0.38754338,0.22292319,0.17147937,0.3018037,0.37039545,0.32924038,0.23321195,0.26750782,0.4046913,0.51100856,0.47328308,0.4424168,0.8162418,0.77508676,0.90198153,1.0871792,1.1660597,0.9294182,1.0528834,0.88826317,0.65505123,0.47671264,0.36696586,0.37382504,0.28465575,0.2503599,0.2777966,0.23664154,0.23664154,0.20234565,0.19891608,0.2469303,0.31552204,0.3018037,0.31209245,0.31552204,0.32238123,0.37382504,0.42869842,0.44927597,0.4081209,0.33266997,0.30866286,0.34638834,0.4081209,0.39783216,0.32581082,0.31209245,0.4389872,0.47328308,0.6344737,0.88826317,0.94656616,1.0425946,1.0563129,1.1763484,1.3615463,1.3512574,1.4369972,1.6393428,1.7525192,1.8039631,2.0406046,2.1503513,2.2360911,2.352697,2.5378947,2.7985435,2.819121,2.510458,2.218943,2.1194851,2.2566686,2.287535,2.5756202,2.7916842,2.8877127,3.1106358,3.1380725,3.5359046,3.9268777,4.256118,4.787704,5.4599032,6.2041235,6.6053853,6.615674,6.550512,6.6876955,6.6225333,6.5950966,6.81802,7.5107965,7.4456344,7.9429245,8.22758,8.207003,8.450503,9.205012,9.80519,10.323058,10.690024,10.703742,10.782623,10.933525,11.218181,11.684605,12.38424,13.625751,14.678635,15.398848,16.016174,17.151367,17.549198,17.947031,18.12537,17.947031,17.38115,17.082775,17.315987,17.754974,18.214539,18.660385,18.516342,18.581505,18.742695,18.87302,18.828436,19.263992,19.634388,20.21399,21.006224,21.723007,22.117409,22.638706,23.314335,24.134007,25.070284,24.881657,24.374079,24.260902,24.418663,23.893936,25.293207,25.557285,27.203487,32.43018,43.085907,32.292995,27.51901,22.288889,14.373401,5.785714,5.120374,4.3521466,4.125794,4.650521,5.7136927,6.866034,8.4264965,9.853205,10.573419,9.938945,10.302481,11.345076,12.586586,13.906977,15.570327,17.185663,18.787281,19.792149,20.186552,20.505503,20.522652,20.61868,20.546658,20.056227,18.86959,19.456049,20.049368,20.53637,20.989075,21.661274,22.220297,22.46037,22.556396,22.648996,22.830763,23.533829,24.744474,25.571005,25.646456,25.135447,24.380938,23.890507,23.681301,23.839062,24.51469,23.808197,23.852781,24.682741,24.36036,18.969048,13.574307,12.576297,13.540011,14.712931,15.001016,13.001566,12.569438,12.500846,12.548861,13.38225,12.655178,12.823228,12.754636,12.487128,13.207341,11.283342,9.959522,8.934075,8.299602,8.529384,7.599966,6.9963584,6.9689217,6.9860697,5.7274113,4.3692946,3.666229,3.2203827,2.9048605,2.836269,4.5030484,6.111525,7.3221693,7.8434668,7.459353,7.7440085,7.881192,7.7680154,7.4284863,6.9963584,7.157549,7.671987,8.086967,8.193284,8.011517,7.7885933,7.3084507,6.4819202,5.5730796,5.209543,4.839148,4.5270553,4.040054,3.4981792,3.3781435,3.1243541,2.369845,1.8142518,1.6153357,1.3924125,1.1146159,1.1797781,1.2106444,1.0837497,0.9362774,1.0871792,1.2689474,1.430138,1.605047,1.9171394,2.5824795,3.2821152,4.091498,4.914599,5.4667625,7.010077,7.377043,7.051232,6.461343,5.977771,5.7308407,5.5387836,5.4084597,5.381023,5.5147767,5.857735,6.258997,6.475061,6.4373355,6.279575,5.9434752,5.4976287,5.086078,4.722542,4.280125,4.4104495,4.3349986,4.15323,4.1360826,4.7431192,4.8117113,5.0929375,5.2781353,5.3432975,5.535354,6.0497923,6.56766,7.0889573,7.5931067,8.045813,8.81747,9.80862,10.295622,10.39165,11.039842,11.441104,11.97269,12.555719,13.073587,13.361672,13.522863,13.601744,13.522863,13.128461,12.168177,12.80608,13.625751,14.164196,14.188204,13.680624,13.011855,12.624311,12.644889,12.932974,13.070158,13.289652,14.249936,15.584045,16.925014,17.902447,18.924463,19.819586,20.320305,20.21056,19.308577,20.512363,21.462358,20.913624,17.672665,10.583707,6.245279,5.5593615,5.302142,4.8837323,6.3618846,8.848335,11.756626,14.503725,15.930434,14.291091,13.855534,14.496866,17.2131,21.153696,23.636717,22.213438,21.747015,21.249723,20.574095,20.392326,19.929333,20.464348,21.225718,21.815605,22.216867,22.062536,21.472647,20.930773,20.244854,18.547209,18.598652,18.248835,18.163095,18.468328,18.759844,17.943602,17.802988,17.130789,16.170506,16.602633,10.967821,6.324159,3.4913201,2.6064866,3.1277838,4.616225,6.186976,6.276145,4.996909,4.149801,5.7925735,5.586798,5.429037,6.0703697,7.130112,8.073249,7.881192,8.525954,9.379922,7.205563,8.011517,5.528495,3.3987212,4.262977,9.764035,8.553391,3.8171308,1.4644338,2.510458,3.07634,3.683377,4.996909,5.48734,5.2164025,5.8371577,6.4819202,6.0703697,6.3893213,7.431916,7.394191,7.116394,6.677407,6.7219915,7.1232533,6.9826403,7.7748747,8.56025,8.745448,8.443645,8.488229,7.9463544,7.6925645,7.8126,8.035523,7.7371492,8.958082,9.997248,10.851214,11.4754,11.763485,12.133881,12.644889,12.699762,12.127021,11.207891,10.926665,10.991828,11.454823,12.253916,13.227919,13.694343,13.738928,13.910407,14.356253,14.79524,14.55174,14.311668,14.71636,15.861842,17.322845,16.79126,16.667795,16.667795,16.894148,17.861292,18.307138,17.823566,16.46888,14.682064,13.293081,12.459691,12.655178,13.807519,15.343974,16.204802,16.599203,16.047039,15.844694,16.510035,17.772121,19.102802,21.133118,23.081123,23.907654,22.336903,21.218857,20.217419,19.058218,17.995045,17.813278,18.6158,18.886738,18.605513,17.998474,17.508043,15.889278,13.738928,12.603734,12.665466,12.734058,12.617453,13.05301,13.152468,12.710052,12.195613,11.430815,10.179015,9.458802,9.39707,9.211872,8.995808,8.371623,8.018375,7.966932,7.596536,7.613684,8.008087,8.549961,9.167287,9.925226,9.602845,9.084977,8.772884,9.009526,10.089847,10.449953,10.30934,9.935514,9.709162,10.096705,8.669997,8.093826,8.093826,8.2481575,8.014946,8.279024,8.2310095,7.394191,5.844017,4.2252517,4.1120753,4.245829,4.6779575,5.3330083,6.001778,6.773435,7.473071,8.155559,8.858624,9.582268,0.2469303,0.21263443,0.1920569,0.20234565,0.2469303,0.28808534,0.32238123,0.33952916,0.31895164,0.26407823,0.18862732,0.2194936,0.20920484,0.18862732,0.16804978,0.14061308,0.12346515,0.13032432,0.15090185,0.17833854,0.21263443,0.16804978,0.18519773,0.20577525,0.21263443,0.22635277,0.25721905,0.28465575,0.30866286,0.33952916,0.39783216,0.47671264,0.5693115,0.6036074,0.5727411,0.5418748,0.5041494,0.5521636,0.6756287,0.8162418,0.864256,0.86082643,0.83681935,0.84367853,0.90541106,1.0014396,1.1180456,1.2483698,1.3032433,1.3752645,1.7216529,2.07833,2.4555845,2.8465576,3.292404,3.882293,4.15666,3.9886103,3.9028704,3.9474552,3.6696587,3.457024,3.6216443,4.0434837,4.6882463,5.6005163,6.6122446,6.7048435,6.7459984,7.058091,7.414768,2.534465,0.75450927,1.0185875,1.7422304,0.7956643,0.33609957,0.31552204,0.35324752,0.4424168,0.9259886,0.84367853,0.37382504,0.0548734,0.024007112,0.01371835,0.39783216,0.8779744,1.0631721,0.96371406,1.0117283,1.2792361,0.9534253,0.490431,0.15776102,0.041155048,0.28808534,0.21263443,0.17147937,0.22978236,0.13032432,0.030866288,0.0034295875,0.01371835,0.048014224,0.09602845,0.1920569,0.12346515,0.037725464,0.010288762,0.044584636,0.10288762,0.1371835,0.14404267,0.14061308,0.16119061,0.216064,0.25378948,0.18519773,0.11317638,0.31552204,0.36010668,0.31552204,0.3018037,0.3566771,0.42526886,0.42869842,0.548734,0.5418748,0.53844523,1.0254467,1.2415106,1.1729189,1.196926,1.3855534,1.5124481,0.97057325,0.58645946,0.34981793,0.26750782,0.36696586,0.5144381,0.47328308,0.3566771,0.28465575,0.39783216,0.4938606,0.4115505,0.42183927,0.5796003,0.7305021,0.66191036,0.9294182,1.1523414,1.1523414,0.94656616,0.91912943,0.8471081,0.6927767,0.52472687,0.53844523,0.44584638,0.34638834,0.3018037,0.3018037,0.26750782,0.26407823,0.20920484,0.18862732,0.22978236,0.2777966,0.2709374,0.30866286,0.30523327,0.28465575,0.37725464,0.41498008,0.432128,0.39783216,0.31895164,0.26064864,0.29494452,0.20920484,0.17147937,0.21263443,0.2503599,0.32924038,0.32238123,0.4115505,0.5624523,0.5418748,0.77851635,0.922559,1.1077567,1.2929544,1.2792361,1.3889829,1.4987297,1.5810398,1.7730967,2.3835633,2.633923,2.7813954,2.9322972,3.0420442,2.9151495,2.9151495,2.620205,2.335549,2.2258022,2.335549,2.311542,2.4247184,2.5378947,2.6750782,3.018037,3.210094,3.457024,3.6936657,4.0263357,4.7088237,5.6348124,6.3035817,6.7631464,7.0478024,7.181556,6.9792104,6.9792104,6.7665763,6.591667,7.3393173,7.6959944,8.464222,8.97866,9.050681,8.961512,9.331907,9.578837,9.80519,10.031544,10.182446,10.38479,10.700313,11.06042,11.55771,12.425395,13.505715,14.452282,15.440002,16.554619,17.7927,18.310568,18.639809,18.728977,18.53692,18.03963,17.422304,17.62122,18.20425,18.886738,19.52807,19.648108,19.757853,19.661825,19.342873,18.962189,19.514353,20.145397,20.875898,21.801888,23.087982,23.420652,23.719027,24.03455,24.487255,25.241764,25.320644,24.974257,24.970827,25.111439,24.206028,25.557285,26.644464,28.791388,33.904903,44.47832,30.845709,25.162884,21.942501,16.95931,7.239859,5.429037,4.3658648,4.046913,4.4516044,5.528495,6.375603,7.81603,9.242738,9.952662,9.146709,9.266746,10.158438,11.413667,12.854094,14.5585985,15.933864,18.224829,19.692692,20.04251,20.430052,20.78673,21.187992,21.352612,20.917053,19.435472,19.363451,19.836735,20.388897,20.879328,21.465788,22.494663,22.93708,23.094843,23.149715,23.19087,24.336353,26.092302,26.929121,26.730206,26.7645,26.35295,26.064865,25.787067,25.667032,26.133457,26.287788,26.665043,27.285797,25.495554,15.9613,10.628291,9.56512,10.412228,11.369082,11.183885,8.567109,7.3255987,7.3564653,8.1041155,8.567109,9.781183,11.067279,11.993267,12.236768,11.561139,10.045261,9.122703,7.9463544,6.866034,7.442205,6.9654922,6.5299344,6.701414,7.034084,6.077229,4.5339146,3.9028704,3.357566,3.000889,3.8548563,4.6779575,6.7631464,7.81603,7.2775846,6.310441,7.0718093,7.4696417,7.394191,7.0203657,6.8145905,6.728851,6.8900414,6.8454566,6.5059276,6.1492505,5.909179,5.65539,5.271276,4.856296,4.746549,4.40702,3.8308492,3.2992632,2.9631636,2.8294096,2.393852,1.6667795,1.1660597,1.0220171,0.939707,0.7922347,0.8196714,0.83338976,0.7476501,0.58302987,1.0151579,1.1008976,1.2277923,1.546744,1.9514352,2.7128036,3.9851806,4.98662,5.579939,6.2898636,6.9552035,6.941485,6.601956,6.121814,5.5250654,5.1238036,4.9660425,4.8768735,4.8425775,4.996909,5.5147767,5.874883,5.9640527,5.7891436,5.48734,5.302142,4.9488945,4.6573796,4.40702,3.9097297,4.1155047,3.8925817,3.508468,3.4810312,4.5647807,4.7774153,5.0312047,5.295283,5.4941993,5.4804807,6.0875177,6.5059276,7.058091,7.7371492,8.176137,8.601405,9.3593445,9.9698105,10.494537,11.5645685,12.020704,12.644889,13.29994,13.814379,14.013294,14.023583,13.663476,13.365103,13.073587,12.271064,13.3033695,13.896688,14.191633,14.325387,14.438563,13.786942,13.358243,13.320518,13.560589,13.670336,13.653188,14.184773,15.388559,16.969599,18.224829,19.390888,20.361462,21.078245,21.294308,20.577524,20.845032,21.805317,21.585823,18.70497,12.048141,8.220721,6.40304,5.2266912,4.7019644,6.186976,7.8949103,9.568549,12.061859,14.366542,13.6086035,13.848674,15.117621,18.416885,22.60441,24.391226,23.314335,22.70044,22.817045,23.537258,24.298628,24.151155,25.368658,26.250063,26.256922,26.01342,25.385807,23.911083,22.683292,21.575535,19.21255,19.068506,18.104792,17.765263,18.149376,18.022482,18.54378,20.426622,20.875898,21.397196,27.796806,16.060759,7.431916,2.74367,1.3752645,1.2346514,3.8205605,5.453044,6.094377,5.6142344,3.789694,3.4055803,3.4844608,4.5099077,6.279575,7.905199,10.024684,9.194724,9.482809,10.624862,8.028665,7.301592,4.5819287,2.8054025,3.765687,8.107545,5.3878818,2.3252604,1.6359133,3.2135234,4.1326528,4.650521,5.381023,6.262427,7.0786686,7.466212,8.31675,8.141841,8.584257,9.740028,10.1652975,9.678296,9.211872,9.205012,9.4862385,9.301042,9.983529,10.611144,10.734609,10.494537,10.621432,9.448513,8.958082,8.937505,9.071259,8.961512,9.901219,11.039842,11.784062,12.055,12.30193,12.212761,12.812939,13.245067,12.9981365,11.897239,11.146159,11.379372,12.103014,12.7272,12.562579,12.507706,12.768354,13.272504,13.972139,14.836395,14.589465,13.903547,13.841815,14.610043,15.532601,14.915276,14.925565,15.309678,16.101913,17.600643,18.097933,17.566347,16.21852,14.387119,12.531713,12.593445,12.511135,13.293081,14.832966,15.906426,16.70552,16.431154,16.088194,16.307688,17.37429,18.86959,20.169403,21.860191,23.314335,22.690151,21.736725,20.172834,18.691252,17.669235,17.171944,16.973028,16.674654,16.204802,15.810398,16.03675,15.693792,14.531162,13.529722,13.039291,12.785502,11.845795,11.396519,11.177026,11.050131,10.998687,11.46854,10.703742,9.860064,9.3936405,9.071259,9.153569,8.697433,8.2653055,8.069819,7.956643,8.110974,8.457363,9.006097,9.702303,10.456812,10.347065,9.9801,9.647429,9.712592,10.607714,10.950673,10.600855,10.045261,9.688584,9.866923,8.536243,8.272165,8.577398,8.841476,8.320179,8.423067,8.385342,7.174697,5.1855364,4.2423997,4.2286816,4.5922174,5.127233,5.7239814,6.3447366,7.1541195,7.3564653,7.8366075,8.831187,9.935514,0.22978236,0.21263443,0.216064,0.24007112,0.2777966,0.33609957,0.36010668,0.42183927,0.3841138,0.25721905,0.20577525,0.2503599,0.24350071,0.22292319,0.19891608,0.15433143,0.1371835,0.15776102,0.18176813,0.18862732,0.1920569,0.17147937,0.20234565,0.23664154,0.26064864,0.28465575,0.28808534,0.32581082,0.37382504,0.42183927,0.490431,0.50757897,0.58645946,0.61046654,0.5761707,0.5693115,0.59331864,0.66533995,0.7888051,0.90884066,0.90198153,0.864256,0.8745448,0.9259886,1.0323058,1.2380811,1.3649758,1.371835,1.3101025,1.3684053,1.8313997,2.2498093,2.6304936,3.1586502,3.7485392,4.064061,4.2423997,4.0846386,3.8308492,3.5564823,3.1895163,3.1449318,3.4227283,3.9440255,4.7808447,6.1629686,7.7028537,7.675417,5.9743414,3.5873485,2.5961976,0.78537554,0.28122616,0.2469303,0.216064,0.1097468,0.072021335,0.17833854,0.2709374,0.24007112,0.037725464,0.006859175,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.15776102,0.4389872,0.7990939,1.1454822,1.5433143,1.313532,0.8162418,0.33266997,0.058302987,0.3841138,0.19548649,0.12346515,0.28122616,0.2503599,0.06516216,0.020577524,0.034295876,0.058302987,0.07888051,0.1097468,0.072021335,0.024007112,0.01371835,0.07545093,0.14061308,0.24007112,0.3018037,0.32924038,0.4081209,0.32238123,0.18519773,0.14061308,0.25721905,0.5418748,0.47328308,0.33266997,0.274367,0.30866286,0.28465575,0.607037,0.8848336,0.84367853,0.7613684,1.4541451,1.6221949,1.4335675,1.2723769,1.2723769,1.2895249,0.85739684,0.6790583,0.548734,0.45956472,0.59674823,0.6001778,0.45270553,0.39440256,0.4698535,0.51100856,0.31895164,0.2503599,0.4355576,0.7133542,0.6241849,0.52472687,0.8779744,1.1111864,1.0460242,0.88826317,0.85739684,0.7956643,0.7339317,0.7133542,0.78537554,0.5041494,0.39097297,0.34981793,0.32581082,0.30523327,0.25721905,0.22635277,0.19548649,0.16804978,0.16804978,0.23664154,0.274367,0.3018037,0.32238123,0.34638834,0.29151493,0.35324752,0.3841138,0.33952916,0.28122616,0.25721905,0.18519773,0.17147937,0.2194936,0.23664154,0.24350071,0.21263443,0.20577525,0.25721905,0.3806842,0.99801,1.0666018,1.097468,1.2380811,1.2792361,1.4232788,1.4027013,1.488441,1.8519772,2.5790498,2.9563043,3.2443898,3.4638834,3.5118976,3.1586502,3.0866287,2.8225505,2.5721905,2.4247184,2.3561265,2.3252604,2.3767042,2.4007113,2.4624438,2.784825,3.2409601,3.4398763,3.5050385,3.7622573,4.73969,6.046363,6.1904054,6.773435,7.8434668,7.915488,7.380472,7.4765005,7.2158523,6.7631464,7.425057,8.429926,9.108984,9.5205345,9.705732,9.674867,9.825768,9.695444,9.578837,9.616563,9.80519,9.938945,10.456812,11.067279,11.732618,12.686044,13.461131,14.376831,15.5085945,16.726099,17.71382,18.293419,18.3723,18.338005,18.37573,18.45804,18.187103,18.567787,19.219408,19.86417,20.344313,20.347742,20.28601,19.895037,19.288,18.934752,19.558937,20.351171,21.136547,22.021381,23.393215,23.34863,23.574984,23.873358,24.19231,24.641586,24.963966,24.94339,25.224615,25.59501,24.977686,26.510712,27.278938,27.76937,30.657082,40.82924,30.074053,24.233465,20.543228,16.228807,8.491658,5.7925735,4.5339146,4.166949,4.4550343,5.470192,6.5196457,7.997798,9.445084,10.131001,9.016385,8.81061,9.355915,10.521975,12.260776,14.640909,15.978448,18.060207,19.270851,19.486916,20.056227,20.817596,21.242865,21.53438,21.589252,21.002794,20.131678,20.382038,21.225718,22.096832,22.398636,23.35549,23.849352,24.168303,24.339783,24.137436,25.35837,27.004572,27.025148,25.725336,25.780209,25.896814,26.627317,26.929121,26.709627,26.819374,28.890844,28.585611,27.467566,24.137436,14.273943,10.583707,9.887501,9.510246,8.23444,6.3001523,6.0086374,5.212973,5.23698,6.135532,6.7048435,7.4799304,8.172707,9.55826,10.580277,8.351046,8.738589,8.189855,6.924337,6.0223556,7.4181976,7.373613,7.191845,6.8626046,6.3653145,5.669108,5.3261495,4.9008803,4.4927597,4.5339146,5.802862,4.73969,6.591667,6.9792104,5.312431,4.804852,6.1321025,6.800872,6.8728933,6.5127864,5.994919,6.121814,5.9571934,5.501058,4.8940215,4.3933015,4.07435,3.9440255,3.9646032,4.029765,3.9440255,3.5187566,3.0660512,2.6750782,2.3458378,2.020027,1.2517995,0.8676856,0.6859175,0.6241849,0.67219913,0.5796003,0.59674823,0.6310441,0.6241849,0.53844523,1.1146159,1.0048691,1.0460242,1.4610043,1.8691251,2.836269,4.605936,5.861165,6.375603,7.040943,6.509357,6.2212715,6.15268,6.046363,5.422178,4.7534084,4.383013,4.122364,3.9954693,4.2526884,4.73969,4.9077396,4.9420357,4.976331,5.1169443,5.1409516,4.715683,4.331569,4.15323,4.029765,4.173808,3.9886103,3.5290456,3.2889743,4.2046742,4.6265135,4.7328305,5.0449233,5.4496145,5.209543,5.593657,5.994919,6.7459984,7.706283,8.285883,8.738589,9.3079,9.914937,10.659158,11.845795,12.109874,12.878101,13.725209,14.335675,14.503725,14.527733,13.886399,13.289652,12.867812,12.140739,13.29994,13.71492,13.951562,14.321958,14.891269,14.647768,14.325387,14.116182,14.05102,13.999576,13.612033,14.078457,15.333686,17.04162,18.602083,19.486916,20.382038,21.02337,21.335464,21.45207,21.081675,21.126259,21.311457,20.4472,16.434584,12.22305,7.888051,5.0003386,4.437886,6.385892,7.016936,7.596536,9.379922,12.113303,14.057879,15.611482,17.398296,20.755863,24.696459,25.924252,25.886526,26.69591,28.92514,31.805994,33.208694,32.683968,33.50364,33.788296,33.061222,32.23812,30.447878,27.748793,25.838512,24.43924,21.297739,20.639257,18.927893,18.084215,17.881868,15.930434,17.20967,21.150267,23.869928,27.1006,38.17817,21.03023,8.594546,2.3149714,0.96714365,0.65848076,2.5310357,4.4859004,5.5319247,5.435896,4.722542,3.957744,4.8940215,6.6053853,8.292743,9.290752,11.640019,11.115293,11.324498,12.22648,10.13786,7.8537555,4.887162,2.7642474,2.7813954,6.0086374,2.4212887,1.5193073,2.6990852,4.8082814,6.138962,5.6039457,6.3001523,7.764586,9.033533,8.669997,10.683165,11.046701,11.101575,11.567999,12.566009,12.13731,11.46854,11.173596,11.273054,11.177026,11.170166,11.375941,11.574858,11.742908,12.044711,10.652299,10.323058,10.360784,10.398509,10.39165,10.89237,12.089295,12.754636,12.586586,12.229909,12.603734,13.443983,14.13333,14.2362175,13.516005,12.027563,12.085866,12.9638405,13.605173,12.614022,11.790922,11.938394,12.545431,13.289652,14.044161,13.869251,13.162757,13.039291,13.618892,13.992717,13.330807,13.176475,13.605173,14.613472,16.115631,17.055338,16.780972,15.848124,14.390549,12.147599,12.590015,12.236768,12.425395,13.37882,14.184773,15.621771,16.386568,16.2974,16.187653,17.892159,19.757853,20.53637,21.28402,21.976797,21.510372,21.232576,19.747564,18.512913,18.005335,17.700102,16.849564,15.913286,14.874121,14.085316,14.280802,15.488017,15.402277,14.507155,13.317088,12.397959,10.55284,9.465661,9.455373,10.131001,10.374502,11.135871,10.854645,10.110424,9.355915,8.906639,9.314759,8.961512,8.31675,8.004657,8.803751,9.256456,9.445084,9.781183,10.275044,10.5597,10.786053,10.748327,10.521975,10.364213,10.707172,11.183885,10.820349,10.161868,9.6645775,9.671436,8.546532,8.436785,8.927217,9.328478,8.669997,8.282454,8.06296,6.8900414,5.0826488,4.40359,4.65395,5.3090014,5.885172,6.3173003,6.9517736,7.5416627,7.2775846,7.455923,8.39563,9.465661,0.22978236,0.33952916,0.37382504,0.36353627,0.32238123,0.274367,0.2503599,0.22635277,0.20920484,0.20577525,0.22978236,0.216064,0.18519773,0.15433143,0.13032432,0.106317215,0.106317215,0.13375391,0.15090185,0.14404267,0.106317215,0.15433143,0.22292319,0.2777966,0.29494452,0.26064864,0.33266997,0.38754338,0.44927597,0.5041494,0.5041494,0.58988905,0.64819205,0.65162164,0.6310441,0.65505123,0.764798,0.84024894,0.9259886,0.9842916,0.90198153,0.8162418,0.85739684,0.91227025,0.97057325,1.1283343,1.1763484,1.2003556,1.2963841,1.4781522,1.6496316,2.0749004,2.877424,3.5873485,3.9303071,3.8445675,4.383013,4.1429415,3.6696587,3.2855449,3.0660512,2.603057,2.651071,3.1586502,4.098357,5.4770513,7.613684,7.1232533,4.57164,1.5124481,0.47328308,0.20577525,0.06516216,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.030866288,0.1920569,0.65505123,0.84024894,0.85739684,0.7407909,0.51100856,0.16804978,0.044584636,0.05144381,0.082310095,0.07888051,0.030866288,0.030866288,0.07545093,0.09602845,0.09259886,0.15090185,0.116605975,0.05144381,0.010288762,0.0034295875,0.01371835,0.05144381,0.06859175,0.15090185,0.31209245,0.5178677,0.28808534,0.12689474,0.18862732,0.34638834,0.19891608,0.6379033,0.53844523,0.30523327,0.17490897,0.19891608,0.15090185,0.28465575,0.69963586,1.2209331,1.4027013,1.3306799,1.3203912,1.1797781,0.97400284,1.0220171,0.99801,1.0837497,1.1214751,0.94999576,0.4115505,0.1920569,0.34638834,0.47671264,0.41498008,0.24350071,0.20920484,0.34638834,0.4424168,0.45613512,0.5041494,0.6756287,0.85396725,0.78194594,0.59674823,0.84024894,1.0220171,0.84024894,0.77851635,0.84367853,0.5658819,0.42869842,0.37039545,0.36353627,0.36696586,0.30523327,0.25721905,0.26407823,0.25721905,0.216064,0.16804978,0.216064,0.22978236,0.30866286,0.4046913,0.31895164,0.19891608,0.28808534,0.29151493,0.18176813,0.18176813,0.15776102,0.18862732,0.19548649,0.16119061,0.1371835,0.18519773,0.25378948,0.33266997,0.490431,0.8711152,1.1626302,1.0425946,1.0734608,1.3272504,1.3889829,1.2312219,1.1351935,1.2929544,1.6633499,1.9685832,2.7368107,3.2409601,3.3369887,3.0729103,2.6716487,2.7573884,2.3835633,2.1263442,2.1229146,2.0749004,2.3561265,2.7642474,2.867135,2.7230926,2.867135,3.2958336,3.724532,3.8342788,3.8102717,4.3487167,4.9214582,5.223262,6.8557453,8.954653,8.1487,6.8900414,6.9071894,7.0958166,7.267296,8.131552,9.156999,9.424506,9.410788,9.417647,9.551401,10.065839,10.045261,9.97324,10.062409,10.268185,10.4533825,10.837497,11.588576,12.528283,13.138749,13.540011,14.291091,15.306249,16.45859,17.593784,17.995045,17.758404,17.658945,18.067066,18.921034,19.421753,20.076805,20.639257,21.064526,21.53095,21.592682,20.773012,19.925903,19.44576,19.288,19.836735,20.467777,20.827885,20.903336,21.0268,20.550089,20.632399,20.992504,21.53095,22.323185,22.895926,22.758743,22.830763,23.012531,22.172283,24.161444,25.793928,27.021719,29.659073,37.39965,27.474424,21.424633,16.448301,11.862943,9.078118,5.5387836,4.9934793,5.3844523,5.871454,6.835168,7.2158523,8.279024,10.086417,11.8115,11.749766,11.063849,11.067279,11.7086115,13.210771,16.067617,17.933313,18.962189,19.356592,19.70298,20.934202,21.62012,22.04539,22.161995,22.076254,22.062536,21.369759,22.035099,23.201159,24.168303,24.415234,24.548986,24.216316,23.808197,23.502962,23.26975,25.087433,26.421541,26.075153,24.76848,25.145735,24.987974,26.075153,26.514141,26.136887,26.490133,30.296976,25.464687,19.984205,17.082775,15.21365,9.657719,8.30646,7.2021337,4.7259717,1.587899,1.845118,2.4761622,3.8377085,5.593657,6.728851,6.0703697,6.3447366,7.3564653,8.460793,8.546532,7.5553813,6.4304767,6.0154963,6.540223,7.613684,7.822889,7.3873315,6.8214493,6.6465406,7.414768,7.64798,6.3790326,6.2864337,7.682276,8.498518,7.0478024,7.2775846,7.0889573,5.7925735,4.1189346,4.413879,4.6779575,4.9831905,5.1512403,4.7602673,5.003768,5.1100855,4.866585,4.3590055,3.9680326,3.5393343,3.2135234,3.0077481,2.9185789,2.9288676,2.7093742,2.4727325,2.1194851,1.6770682,1.313532,0.64133286,0.39097297,0.29837412,0.23321195,0.18176813,0.17147937,0.17833854,0.18176813,0.23321195,0.42869842,0.37725464,0.5041494,0.8025235,1.2723769,1.9068506,3.1655092,4.7979927,5.744559,6.001778,6.636252,6.3310184,6.245279,6.111525,5.7891436,5.2644167,4.4104495,3.765687,3.1860867,2.8465576,3.2512488,3.2992632,3.6593697,4.0606318,4.4447455,4.9591837,5.178677,5.051782,4.6608095,4.249259,4.2115335,3.5290456,3.642222,3.707384,3.4981792,3.3884325,3.875434,4.0537724,4.633373,5.381023,5.1100855,4.976331,5.3844523,6.3721733,7.7714453,9.201583,9.702303,10.13786,10.333347,10.652299,11.993267,12.175035,12.926115,13.72178,14.249936,14.417986,14.7369375,14.678635,14.195063,13.4474125,12.785502,12.7272,13.560589,14.472859,15.014734,15.138199,14.843254,14.661487,14.2533655,13.900118,14.510585,14.195063,14.654627,15.601193,16.719238,17.686382,18.015623,19.013634,20.28258,21.242865,21.133118,20.803877,20.70442,21.232576,22.172283,22.659285,17.237106,13.375391,9.798331,6.725421,5.857735,4.822,8.213862,11.2593355,13.008426,16.341984,19.514353,22.175713,25.430391,28.733084,29.892284,30.293547,36.309044,43.63464,49.320896,51.78677,47.99022,44.358284,41.954144,40.537724,38.57257,35.376194,32.78,31.164661,29.158352,23.667583,23.300617,20.344313,18.578075,17.79613,13.7938,17.017612,21.016512,20.821026,19.795578,29.631636,17.974468,8.258447,2.8568463,1.3924125,0.7339317,0.52472687,2.4144297,6.0566516,8.872343,6.025785,7.822889,9.551401,11.509696,13.358243,14.112752,15.409137,14.935853,13.145609,10.834066,9.126132,7.1849856,5.5902276,4.3452873,3.7382503,4.3487167,3.309552,4.40702,6.2075534,7.798882,8.790032,7.5690994,7.291303,8.327039,9.952662,10.329918,13.505715,12.878101,11.876661,12.127021,13.457702,13.848674,12.528283,11.478829,11.334786,11.382801,11.211322,11.286773,11.526843,11.619442,11.032983,11.05699,11.509696,11.701753,11.379372,10.7586155,11.646879,13.059869,14.112752,14.476289,14.404267,14.599753,15.683503,15.999025,15.309678,14.784951,13.248496,12.452832,12.360233,12.771784,13.320518,13.063298,11.993267,11.561139,11.993267,12.298501,12.360233,12.449403,12.55229,12.953552,14.2362175,13.663476,13.646329,14.208781,15.066177,15.638919,16.95931,16.691803,15.906426,14.723219,12.329367,11.718901,11.327928,11.670886,12.487128,12.758065,13.841815,15.553179,16.259674,16.341984,18.173384,20.663265,22.330044,22.52553,21.215427,18.982767,18.578075,18.423744,18.28999,17.991615,17.394867,17.54234,17.175373,16.077906,14.668345,14.023583,14.057879,14.116182,13.560589,12.4802685,11.688034,9.942374,9.22216,9.246168,9.544542,9.462232,9.496528,9.825768,9.72288,9.225591,9.139851,9.458802,8.621983,7.9875093,8.351046,9.962952,10.367643,10.302481,10.511685,10.960961,10.864933,10.875222,11.036412,10.81006,10.233889,9.904649,10.916377,11.170166,10.669447,9.757176,9.108984,8.512236,8.378482,8.423067,8.47451,8.498518,8.217292,8.1212635,6.941485,5.171818,5.051782,5.90575,6.7048435,7.222711,7.4284863,7.4765005,7.2947326,7.284444,7.630832,8.210432,8.573969,0.20577525,0.2469303,0.2503599,0.24007112,0.23321195,0.26407823,0.23664154,0.1920569,0.16462019,0.16462019,0.16804978,0.15433143,0.14061308,0.1371835,0.14747226,0.14404267,0.12346515,0.12346515,0.1371835,0.15776102,0.17833854,0.24007112,0.30866286,0.34295875,0.34981793,0.3806842,0.39440256,0.4081209,0.45956472,0.5590228,0.6859175,0.65505123,0.72021335,0.75450927,0.75450927,0.8265306,0.94656616,0.9328478,0.94656616,0.96714365,0.8162418,0.83681935,0.980862,1.0700313,1.0597426,1.0425946,1.1317638,1.2517995,1.3821237,1.5364552,1.7593783,2.2841053,2.9322972,3.457024,3.758828,3.9200184,4.3281393,3.5942078,2.976882,2.8705647,2.7985435,2.2669573,2.4658735,2.8396983,3.1860867,3.6456516,5.2164025,5.0586414,3.4604537,1.3649758,0.37382504,0.16462019,0.06859175,0.024007112,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.006859175,0.08916927,0.38754338,0.89169276,1.1454822,1.138623,0.85739684,0.3018037,0.10288762,0.116605975,0.14747226,0.106317215,0.017147938,0.0274367,0.041155048,0.037725464,0.034295876,0.0548734,0.037725464,0.024007112,0.024007112,0.034295876,0.0274367,0.06516216,0.12003556,0.18519773,0.22978236,0.20234565,0.14404267,0.22978236,0.37725464,0.5624523,0.7956643,0.6001778,0.5178677,0.32581082,0.07545093,0.08916927,0.1097468,0.28808534,0.4629943,0.6001778,0.7922347,0.7099246,0.5727411,0.66191036,0.9328478,1.0220171,0.8025235,0.86082643,0.805953,0.6036074,0.59674823,0.48357183,0.4972902,0.4389872,0.30866286,0.29151493,0.3841138,0.37725464,0.30866286,0.274367,0.42869842,0.4355576,0.48014224,0.4938606,0.5178677,0.70649505,0.8196714,0.823101,0.9602845,1.1146159,0.83338976,0.805953,0.5590228,0.42183927,0.42526886,0.30523327,0.35324752,0.37039545,0.35324752,0.31552204,0.2777966,0.33609957,0.41840968,0.44584638,0.4046913,0.30866286,0.29494452,0.34295875,0.31552204,0.20920484,0.17147937,0.15776102,0.14404267,0.216064,0.3018037,0.19891608,0.34638834,0.41498008,0.4046913,0.4355576,0.7339317,0.65848076,0.6962063,0.764798,0.8676856,1.0940384,1.3649758,1.4678634,1.4507155,1.5330256,2.1023371,2.3629858,2.7711067,3.0077481,2.9494452,2.633923,2.6613598,2.4727325,2.3424082,2.270387,1.978872,2.277246,2.6407824,2.7402403,2.7059445,3.1243541,3.3850029,3.3678548,3.3678548,3.566771,4.0434837,4.32471,4.887162,6.7631464,8.539673,6.3790326,5.130663,5.5593615,6.427047,7.0889573,7.4970784,8.865483,9.472521,9.825768,10.079557,10.028113,10.031544,10.069269,10.028113,9.9869585,10.233889,10.971251,11.4754,12.024134,12.72034,13.46799,13.841815,14.400838,15.155347,16.067617,17.055338,17.391438,17.676094,18.077356,18.653526,19.37374,20.028791,20.563807,20.759293,20.697561,20.762722,20.86218,20.52951,19.908754,19.281141,19.054789,19.672113,20.28601,20.646116,20.724997,20.721567,20.382038,20.073376,19.833303,19.847023,20.457489,20.86218,20.930773,21.191422,21.349182,20.29287,21.246294,22.552967,24.919382,30.523329,43.03789,27.666483,19.87789,16.554619,14.688923,11.396519,6.5882373,5.7411294,5.3330083,4.537344,5.1992545,6.5470824,7.3839016,8.477941,9.650859,9.784613,10.155008,10.984968,11.996697,13.275933,15.261664,16.650646,17.394867,17.933313,18.550638,19.37374,19.908754,21.20171,21.232576,20.124819,20.124819,20.989075,21.699,22.580404,23.28347,22.765602,22.46037,22.333473,22.261452,22.587263,24.11343,25.121729,26.274069,25.76992,24.154585,24.329493,23.554407,24.247183,25.255482,26.219196,27.549875,28.009441,21.760733,19.54522,20.02193,9.757176,5.4907694,4.2938433,3.789694,3.0077481,2.3801336,1.7079345,1.9171394,2.8019729,3.8034124,4.033195,5.40503,5.4770513,5.5593615,6.0635104,6.468202,8.64599,9.239308,9.407358,9.39021,8.529384,7.915488,7.1678376,6.7048435,6.5539417,6.3653145,7.6342616,7.466212,7.579388,8.889491,11.513125,11.417097,9.880642,7.6445503,6.101236,7.2707253,7.377043,5.8817425,4.7019644,4.372724,4.040054,3.8342788,3.9337368,3.8205605,3.3644254,2.8088322,2.4487255,2.1983654,2.1229146,2.1503513,2.0749004,1.9445761,1.7696671,1.4918705,1.0837497,0.5796003,0.2709374,0.16804978,0.14061308,0.12003556,0.1097468,0.09602845,0.08916927,0.08916927,0.106317215,0.14747226,0.15776102,0.216064,0.45613512,1.039165,2.1640697,2.9803114,4.554492,5.6485305,5.809721,5.381023,5.329579,5.137522,5.0243454,5.007198,4.911169,4.125794,3.2992632,2.5961976,2.1846473,2.2360911,2.4418662,2.6373527,3.0283258,3.590778,4.057202,4.4721823,4.8014226,4.8837323,4.804852,4.8940215,3.566771,2.9254382,2.8396983,2.9460156,2.6304936,2.7470996,3.1895163,4.0057583,4.787704,4.6848164,4.9591837,5.521636,6.327589,7.442205,9.006097,10.189304,10.912948,11.022695,10.854645,11.249047,12.1921835,13.13532,13.869251,14.318527,14.517444,14.658057,14.747226,14.527733,14.078457,13.80066,13.797231,14.291091,15.038741,15.604623,15.343974,15.3817,15.618341,15.227368,14.390549,14.328816,14.246507,14.472859,15.100473,16.012743,16.88043,17.168514,18.166525,19.94305,21.987085,23.19773,21.987085,20.69413,20.097382,20.306587,20.755863,19.54522,18.608942,14.321958,8.4093485,7.922347,6.111525,8.961512,11.530273,13.015285,16.756964,17.449741,20.100813,24.548986,29.278389,31.404732,33.42819,44.64637,58.2001,69.130196,74.370605,70.231094,64.50711,59.547928,55.09975,48.292023,43.939873,40.705772,38.716614,36.442795,30.684519,23.842491,17.058767,14.068168,14.13676,12.037852,11.276484,16.13278,18.008764,17.514904,24.494114,15.29596,8.018375,3.5016088,2.1674993,4.029765,1.8176813,1.7662375,5.219832,9.609704,8.443645,6.56766,5.9571934,8.038953,11.369082,11.650309,14.349394,15.9921665,15.374841,12.250486,7.3290286,6.2864337,4.7362604,3.5221863,3.2786856,4.434457,5.6039457,6.4819202,6.2658563,5.5422134,6.2864337,7.010077,7.73029,9.304471,11.231899,11.660598,14.277372,13.906977,13.433694,13.972139,14.860402,14.922135,14.658057,14.188204,13.481709,12.360233,12.30536,12.610593,13.173045,13.502286,12.6929035,12.120162,11.986408,12.404818,13.149038,13.649758,13.251926,14.424845,15.601193,16.228807,16.760393,16.770683,17.432592,18.04306,18.183672,17.727537,16.071047,14.417986,13.275933,12.874671,13.149038,13.059869,11.9040985,11.30735,11.588576,11.787492,11.681175,11.660598,12.092726,13.070158,14.417986,14.421415,14.417986,15.0250225,15.776102,15.127911,14.483148,14.143619,13.684054,12.97413,12.181894,11.766914,11.537132,11.585147,11.917816,12.452832,12.833516,13.855534,15.086755,16.269962,17.319416,20.052797,21.3629,21.239435,20.19684,19.250275,19.05136,19.263992,19.384027,18.982767,17.71382,17.576635,17.21996,16.321407,15.059319,14.109323,13.3033695,13.155897,13.337666,13.1421795,11.46854,9.97667,9.825768,10.31277,10.566559,9.534253,9.187865,9.527394,9.72631,9.445084,8.824328,8.964942,7.857185,7.822889,9.208443,10.377932,10.72432,10.690024,10.823778,11.091286,10.875222,10.926665,11.06042,10.796341,10.192734,9.8429165,10.590566,11.180455,10.89237,9.777754,8.669997,8.375052,8.772884,9.14328,9.105555,8.632272,8.419638,8.128122,7.1952744,5.9400454,5.562791,6.4579134,7.0752387,7.6033955,8.011517,8.049242,7.857185,7.7885933,8.086967,8.618553,8.855195,0.216064,0.26407823,0.26407823,0.26750782,0.2709374,0.23321195,0.216064,0.21263443,0.22292319,0.22978236,0.216064,0.19548649,0.17833854,0.16462019,0.16804978,0.18862732,0.18519773,0.19548649,0.22635277,0.26750782,0.29151493,0.32238123,0.33952916,0.3566771,0.37039545,0.37382504,0.39097297,0.44927597,0.50757897,0.5796003,0.72364295,0.6859175,0.6962063,0.75450927,0.84367853,0.9534253,1.0597426,0.9774324,0.89169276,0.881404,0.922559,1.0220171,1.0597426,1.0666018,1.0563129,1.0323058,1.1351935,1.2586586,1.3821237,1.546744,1.8588364,2.2326615,2.6819375,3.1106358,3.5290456,4.064061,4.266407,3.4981792,2.8877127,2.7402403,2.5207467,2.1332035,2.3835633,2.877424,3.1483612,2.6476414,3.4844608,3.6456516,2.7539587,1.2860953,0.5796003,0.23664154,0.08916927,0.0274367,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.010288762,0.020577524,0.072021335,0.2194936,0.71678376,0.9294182,0.8676856,0.6001778,0.26407823,0.14404267,0.13375391,0.14404267,0.116605975,0.034295876,0.030866288,0.048014224,0.05144381,0.041155048,0.041155048,0.0274367,0.058302987,0.061732575,0.030866288,0.01371835,0.0274367,0.09602845,0.16119061,0.17490897,0.11317638,0.15090185,0.1920569,0.31209245,0.59674823,1.1489118,0.5521636,0.31895164,0.16804978,0.037725464,0.06859175,0.1371835,0.25721905,0.35324752,0.39440256,0.42183927,0.4664239,0.4972902,0.6824879,0.9534253,0.9774324,0.8093826,0.77165717,0.71678376,0.61389613,0.5693115,0.53501564,0.50757897,0.4115505,0.30523327,0.38754338,0.33952916,0.30523327,0.26407823,0.2469303,0.31209245,0.31209245,0.32581082,0.38754338,0.52472687,0.75450927,0.9602845,0.9294182,0.939707,1.0048691,0.89169276,0.9774324,0.6379033,0.42869842,0.490431,0.5144381,0.47328308,0.44927597,0.47671264,0.50757897,0.4424168,0.4081209,0.38754338,0.33952916,0.274367,0.24007112,0.26750782,0.2469303,0.24007112,0.26064864,0.24007112,0.25721905,0.30866286,0.42526886,0.51100856,0.34981793,0.50757897,0.50757897,0.50757897,0.5590228,0.6276145,0.6036074,0.67219913,0.77165717,0.8676856,0.96714365,1.2277923,1.3443983,1.3443983,1.3958421,1.7971039,1.879414,2.2978237,2.6956558,2.8294096,2.5790498,2.627064,2.5653315,2.486451,2.393852,2.2086544,2.4795918,2.8705647,3.1380725,3.3438478,3.8479972,3.7759757,3.5290456,3.415869,3.6525106,4.3795834,4.4859004,4.73969,6.385892,7.8777623,4.8905916,3.4947495,4.266407,5.645101,6.691125,7.1026754,8.824328,9.547972,9.925226,10.203023,10.203023,10.336777,10.261326,10.213311,10.240748,10.206452,10.782623,11.303921,12.05157,12.932974,13.485138,14.225929,14.778092,15.271953,15.734947,16.081335,16.520323,17.333136,18.015623,18.502625,19.154245,19.888178,20.19341,20.258574,20.19684,20.028791,19.61724,19.576086,19.562366,19.469769,19.401176,20.028791,20.351171,20.436913,20.388897,20.351171,19.987637,19.555508,19.222837,19.171394,19.630959,20.028791,20.347742,20.423193,20.299728,20.207129,21.602972,23.69502,24.76505,26.243204,32.694256,26.503853,21.404055,18.320856,15.9921665,10.971251,7.0306544,6.2487082,5.9331865,5.144381,4.6916757,6.351596,6.9071894,7.281014,7.857185,8.488229,9.283894,10.463672,11.688034,12.682614,13.265644,14.147048,15.13134,15.916716,16.681513,18.067066,18.530062,19.589804,19.747564,19.188541,19.775002,20.899906,21.393766,21.969936,22.570116,22.354052,22.53925,22.422644,22.426073,22.961088,24.404943,24.624437,24.888515,24.007113,22.690151,23.5304,23.334913,24.621008,26.260351,28.023159,30.571342,33.380177,26.088871,23.78076,25.063425,12.082437,4.8734436,2.4452958,1.9823016,2.0817597,2.760818,3.8205605,3.1517909,3.2786856,4.232111,3.5599117,5.7377,5.7308407,4.887162,4.6436615,6.509357,8.011517,9.22902,9.736599,9.661148,9.702303,11.358793,10.666017,10.041832,9.753747,7.936065,8.495089,8.604835,9.098696,10.281903,11.938394,12.079007,10.151579,7.675417,6.166398,7.133542,6.6225333,5.2026844,4.262977,3.9097297,2.952875,2.1743584,2.0680413,2.020027,1.8108221,1.5947582,1.2963841,1.0837497,1.0117283,1.0220171,0.9568549,0.90541106,0.7682276,0.59331864,0.40126175,0.18519773,0.09259886,0.06516216,0.0548734,0.044584636,0.044584636,0.041155048,0.037725464,0.037725464,0.041155048,0.048014224,0.072021335,0.116605975,0.41840968,1.0254467,1.786815,2.2463799,3.9303071,5.055212,5.0312047,4.4516044,4.2595477,4.122364,4.040054,4.064061,4.307562,3.5461934,2.7470996,2.0886188,1.7182233,1.7182233,1.8656956,1.9891608,2.4041407,3.0317552,3.4192986,3.758828,4.3521466,4.804852,5.0312047,5.284994,3.350707,2.6716487,2.8328393,3.1655092,2.7711067,2.7299516,2.976882,3.4638834,3.9371665,3.9200184,4.554492,5.3090014,6.1972647,7.4044795,9.304471,10.858074,11.5645685,11.46854,11.046701,11.228469,12.679185,13.694343,14.280802,14.510585,14.55174,14.671775,14.839825,14.675205,14.092175,13.3033695,13.828096,14.514014,15.138199,15.505165,15.46058,15.734947,15.9613,15.570327,14.764374,14.510585,14.260224,14.891269,15.673215,16.324837,17.04505,17.799559,18.475187,19.86417,21.764162,22.978235,22.343761,21.143406,20.388897,20.385468,20.745575,21.503513,22.295748,19.161106,12.915827,9.170717,7.205563,8.80718,11.135871,12.994707,14.808959,15.234227,17.055338,21.1194,26.040857,28.204927,29.885426,39.289352,52.69561,66.44826,76.94965,79.98484,79.6213,76.66843,70.81069,60.60767,52.729908,46.676685,43.281395,41.213352,36.981243,28.280378,17.583494,11.2421875,10.343636,10.717461,7.267296,11.094715,14.260224,15.697222,21.211998,13.677195,7.222711,3.275256,3.3678548,9.153569,5.470192,3.4124396,5.271276,9.3764925,10.110424,6.427047,5.5593615,8.152129,11.842365,11.2250395,15.148488,17.566347,17.137648,13.1593275,5.5730796,4.8288593,4.3109913,3.858286,3.8137012,5.003768,5.267846,5.4084597,5.0414934,4.4584637,4.636802,5.645101,6.5059276,7.874333,9.740028,11.417097,13.564018,13.001566,12.778643,13.759505,14.637479,13.491997,13.927555,14.544881,14.565458,13.831526,14.157337,14.5243025,14.750656,14.644339,14.013294,13.982429,13.828096,14.102464,14.699212,14.850114,14.980438,16.280252,17.343424,17.813278,18.403166,17.861292,18.005335,18.838724,19.812727,19.826445,18.434032,15.892709,14.112752,13.670336,13.80409,13.797231,12.833516,11.989838,11.71547,11.80464,11.46854,11.423956,11.907528,12.929544,14.280802,14.311668,14.116182,14.517444,15.282242,15.138199,13.831526,12.977559,12.483699,12.322508,12.538571,11.910957,11.712041,11.780633,11.907528,11.852654,11.80464,12.247057,13.437123,15.021593,16.04361,17.71039,17.412016,16.684942,16.609491,17.826996,18.917604,19.46291,19.733847,19.582945,18.440891,18.087645,17.61436,16.678083,15.436573,14.55174,13.543441,13.227919,13.413116,13.330807,11.605724,10.316199,10.408798,10.864933,10.751757,9.194724,8.783174,8.971801,9.146709,9.006097,8.549961,8.635701,8.412778,8.632272,9.5205345,10.765475,10.943813,10.666017,10.703742,11.022695,10.816919,10.55284,10.467101,10.1481495,9.623423,9.342196,9.818909,10.569988,10.535692,9.674867,8.944365,8.834618,9.249598,9.5033865,9.201583,8.237869,7.98408,7.6925645,7.0752387,6.2830043,5.90232,6.893471,7.3187394,7.891481,8.621983,8.834618,8.309891,8.207003,8.282454,8.405919,8.577398,0.36353627,0.37039545,0.33609957,0.32238123,0.31552204,0.23664154,0.2469303,0.3018037,0.33266997,0.31552204,0.29151493,0.26407823,0.25721905,0.2503599,0.2503599,0.26750782,0.28122616,0.29837412,0.31552204,0.32924038,0.31895164,0.36696586,0.3806842,0.39440256,0.4046913,0.39440256,0.4424168,0.51100856,0.5555932,0.58302987,0.6379033,0.6344737,0.6756287,0.77851635,0.89855194,0.9534253,1.0254467,0.939707,0.8711152,0.91569984,1.0734608,1.1249046,1.0837497,1.0460242,1.039165,1.0254467,1.1249046,1.2620882,1.4027013,1.5673214,1.821111,2.1572106,2.534465,3.0214665,3.6182148,4.2286816,4.197815,3.5221863,2.9974594,2.7813954,2.4041407,2.0886188,2.1812177,2.5173173,2.760818,2.3732746,3.1860867,2.760818,1.7902447,0.881404,0.5693115,0.32238123,0.13375391,0.037725464,0.024007112,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.037725464,0.061732575,0.106317215,0.14061308,0.41840968,0.6824879,0.6893471,0.4698535,0.31895164,0.28808534,0.21263443,0.15433143,0.116605975,0.034295876,0.020577524,0.037725464,0.06859175,0.08573969,0.06859175,0.19548649,0.16119061,0.08573969,0.034295876,0.017147938,0.006859175,0.06859175,0.11317638,0.116605975,0.106317215,0.18862732,0.18519773,0.37725464,0.77165717,1.1180456,0.53158605,0.23664154,0.106317215,0.058302987,0.082310095,0.20234565,0.28122616,0.34295875,0.38754338,0.36010668,0.4389872,0.51100856,0.6859175,0.922559,1.0563129,0.83681935,0.72364295,0.66191036,0.6207553,0.5727411,0.65505123,0.607037,0.45613512,0.33952916,0.4972902,0.28465575,0.2777966,0.28808534,0.24350071,0.18176813,0.23664154,0.274367,0.4115505,0.6241849,0.7476501,0.97400284,0.89512235,0.7888051,0.77165717,0.78194594,0.864256,0.70306545,0.607037,0.6310441,0.59674823,0.5418748,0.5418748,0.5521636,0.53158605,0.4424168,0.4081209,0.31209245,0.23664154,0.20234565,0.17490897,0.20234565,0.20920484,0.23321195,0.29151493,0.36353627,0.45270553,0.5041494,0.5796003,0.64133286,0.5761707,0.607037,0.5521636,0.5212973,0.52815646,0.4938606,0.59331864,0.65162164,0.7682276,0.90541106,0.881404,1.0666018,1.1454822,1.2312219,1.3478279,1.4267083,1.5536032,1.9102802,2.3458378,2.6407824,2.5310357,2.668219,2.5961976,2.4384367,2.3321195,2.435007,2.5378947,2.9940298,3.4364467,3.7725463,4.1772375,3.9337368,3.74168,3.6559403,3.8548563,4.6402316,4.6573796,4.698535,5.8337283,6.914048,4.5613513,3.0454736,3.74168,4.9420357,5.909179,6.869464,8.635701,9.4862385,9.870353,10.124143,10.484249,10.501397,10.343636,10.288762,10.353925,10.295622,10.64201,11.074138,11.845795,12.744347,13.107883,14.068168,14.623761,15.151917,15.772673,16.359133,16.750105,17.655516,18.28999,18.54378,18.996485,19.78872,19.726988,19.586374,19.582945,19.356592,18.996485,18.921034,19.089085,19.349733,19.442331,19.836735,19.833303,19.644676,19.500635,19.651537,19.233126,18.934752,18.732407,18.71526,19.075365,19.54179,20.217419,20.330595,20.11453,20.821026,22.148275,24.319204,24.898806,23.773901,23.129137,28.551315,27.17605,23.149715,18.183672,11.550851,7.140401,6.012067,6.591667,6.992929,5.0140567,6.0875177,6.3824625,6.2967224,6.310441,6.9723516,8.014946,8.958082,10.034973,11.043272,11.345076,11.921246,12.826657,13.742357,14.850114,16.822126,17.573206,18.766703,19.524641,19.78872,20.323736,20.635828,21.04395,21.85676,22.8582,23.331484,23.931662,23.36921,22.8582,23.002243,23.811626,23.77733,23.931662,23.228596,22.44322,24.158014,23.797907,24.552416,25.471546,26.737064,29.683079,34.25129,30.533617,29.370987,28.84969,14.29795,5.079219,1.7936742,1.1797781,1.3992717,2.0406046,3.74168,3.059192,3.5873485,5.2335505,4.2115335,5.3570156,5.7479887,5.0174866,4.389872,6.711703,7.1952744,9.119273,9.633711,8.937505,10.257896,12.397959,12.830087,13.063298,12.764925,9.753747,9.935514,9.0644,9.033533,10.031544,10.535692,11.897239,9.595985,6.835168,5.4633327,5.953764,6.077229,5.909179,5.6073756,4.863155,2.8980014,1.3238207,0.8505377,0.77851635,0.72364295,0.6276145,0.45270553,0.32581082,0.26407823,0.2503599,0.216064,0.20920484,0.1371835,0.06516216,0.030866288,0.0274367,0.020577524,0.017147938,0.01371835,0.010288762,0.010288762,0.01371835,0.010288762,0.010288762,0.010288762,0.017147938,0.034295876,0.058302987,0.2777966,0.66876954,1.0014396,1.3512574,2.6167753,3.4776018,3.6044965,3.6696587,3.1655092,3.0626216,3.083199,3.199805,3.6319332,2.8739944,2.0989075,1.5810398,1.3924125,1.3992717,1.4918705,1.704505,2.170929,2.74367,3.0283258,3.3678548,4.0023284,4.57507,4.9008803,4.9694724,3.069481,2.5893385,2.8911421,3.2855449,3.0283258,2.952875,3.0248961,3.1415021,3.2821152,3.5153272,4.400161,5.5319247,6.6636887,7.874333,9.568549,11.111863,11.72233,11.574858,11.218181,11.567999,13.107883,13.934414,14.164196,14.1299,14.38026,14.527733,14.788382,14.730078,14.205351,13.368532,13.845244,14.579176,15.049029,15.21365,15.5085945,15.885849,15.820687,15.484588,15.073037,14.79867,14.575747,15.481158,16.331696,16.828985,17.525192,18.907316,19.270851,20.015072,21.266872,21.85676,21.956219,21.428062,21.033659,21.016512,21.088533,21.733295,23.238884,21.417774,15.87213,9.983529,8.748878,9.657719,11.348505,12.902108,13.845244,15.05246,16.05733,19.246845,23.869928,26.037428,26.051146,29.59048,37.15272,47.444912,57.390717,62.236725,64.4248,64.147,61.262722,55.28152,50.109703,46.155388,43.98103,42.544033,39.179607,29.724234,17.593784,9.280463,7.490219,11.125582,6.924337,7.9600725,10.425946,12.751206,15.587475,10.028113,5.127233,2.4830213,3.5702004,9.72288,6.6053853,5.73427,6.591667,8.368194,9.97667,7.442205,6.4819202,8.515666,12.006986,12.456262,17.412016,19.21255,17.53548,12.655178,5.4324665,5.645101,5.4907694,4.897451,4.4756117,5.504488,4.664239,4.307562,4.2423997,4.3109913,4.386442,5.3227196,6.125243,7.301592,8.779744,9.908078,11.88352,11.30049,11.077567,12.157887,13.512574,12.836946,13.354814,13.732068,13.684054,13.996146,14.599753,15.193072,15.354263,15.097044,14.850114,15.453721,15.46401,15.199932,14.788382,14.153908,15.597764,17.195951,18.293419,18.811287,19.267422,18.20082,17.861292,18.691252,20.237995,21.170843,20.100813,17.144508,15.093615,14.664916,14.517444,14.078457,13.437123,12.744347,12.147599,11.797781,10.8958,10.957532,11.650309,12.607163,13.4474125,13.841815,13.824667,14.321958,15.323397,15.875561,14.421415,13.046151,12.109874,11.777204,12.037852,11.873232,11.746337,11.777204,11.766914,11.204462,11.166737,11.159878,11.88352,13.169616,13.975569,13.951562,13.351384,12.9809885,13.443983,15.110763,17.665806,18.691252,19.099373,19.181683,18.612371,18.101362,17.494326,16.403717,15.100473,14.527733,13.656617,13.118172,12.854094,12.487128,11.317638,10.47396,10.357354,10.323058,9.856634,8.584257,8.385342,8.577398,8.862054,8.98209,8.721441,8.769455,9.187865,9.407358,9.657719,10.9541025,11.262765,10.81006,10.593996,10.714031,10.364213,10.175586,9.938945,9.582268,9.218731,9.156999,9.177576,9.911508,10.233889,9.849775,9.304471,9.139851,9.331907,9.325048,8.882631,8.083538,7.675417,7.394191,7.051232,6.667118,6.4990683,7.281014,7.613684,8.309891,9.273604,9.499957,8.632272,8.357904,8.261876,8.172707,8.158989,0.52472687,0.47328308,0.4046913,0.37039545,0.37725464,0.3841138,0.39783216,0.42183927,0.4081209,0.37039545,0.37725464,0.34638834,0.34638834,0.36696586,0.37382504,0.33952916,0.33952916,0.35324752,0.3566771,0.34638834,0.33266997,0.42183927,0.44927597,0.44927597,0.45613512,0.490431,0.5521636,0.5555932,0.5624523,0.5761707,0.548734,0.5624523,0.6859175,0.8162418,0.8848336,0.84367853,0.864256,0.864256,0.91912943,1.0357354,1.1489118,1.0940384,1.0700313,1.0528834,1.0288762,0.9945804,1.1523414,1.313532,1.4815818,1.6359133,1.7182233,2.153781,2.5824795,3.1895163,3.8857226,4.290414,4.0263357,3.433017,3.0351849,2.8705647,2.5001693,2.1297739,2.020027,2.0508933,2.201795,2.5447538,3.4227283,2.0097382,0.66191036,0.26750782,0.274367,0.31552204,0.15776102,0.05144381,0.058302987,0.05144381,0.01371835,0.0034295875,0.0034295875,0.0,0.0034295875,0.01371835,0.017147938,0.01371835,0.017147938,0.048014224,0.13032432,0.1371835,0.13032432,0.13032432,0.09945804,0.13032432,0.5178677,0.69963586,0.5693115,0.48014224,0.5144381,0.36010668,0.19891608,0.10288762,0.01371835,0.0034295875,0.006859175,0.05144381,0.1097468,0.10288762,0.39097297,0.26407823,0.10288762,0.058302987,0.0548734,0.030866288,0.0548734,0.058302987,0.05144381,0.116605975,0.17833854,0.20920484,0.5212973,0.9328478,0.77165717,0.48014224,0.2777966,0.15090185,0.09259886,0.07545093,0.25721905,0.3018037,0.34981793,0.42869842,0.4389872,0.5727411,0.58988905,0.69963586,0.9259886,1.1214751,0.78194594,0.6927767,0.66191036,0.6310441,0.6927767,0.7990939,0.764798,0.5624523,0.34638834,0.47328308,0.29151493,0.29151493,0.28465575,0.20920484,0.12346515,0.2194936,0.28808534,0.50757897,0.77165717,0.6927767,0.7476501,0.6824879,0.61389613,0.59674823,0.6001778,0.607037,0.7922347,0.881404,0.77165717,0.5178677,0.5693115,0.6173257,0.5624523,0.42183927,0.32238123,0.37382504,0.30866286,0.2503599,0.23664154,0.18519773,0.17490897,0.29151493,0.33609957,0.32581082,0.490431,0.6001778,0.5761707,0.5796003,0.66533995,0.77165717,0.6379033,0.58645946,0.5041494,0.4081209,0.432128,0.5178677,0.5418748,0.65848076,0.823101,0.77508676,0.90198153,0.9774324,1.1283343,1.2758065,1.1351935,1.4198492,1.704505,2.1023371,2.4967396,2.5413244,2.7642474,2.6304936,2.3972816,2.3081124,2.5996273,2.5378947,2.9940298,3.508468,3.865145,4.108646,3.875434,4.0366244,4.170378,4.2766957,4.763697,4.7362604,4.870014,5.4907694,6.0635104,5.1992545,4.0777793,4.3349986,4.695105,5.06893,6.574519,7.905199,8.8929205,9.493098,9.932085,10.707172,10.367643,10.220171,10.103564,10.038403,10.185875,10.566559,10.88551,11.458252,12.181894,12.528283,13.37882,13.828096,14.596324,15.87213,17.315987,17.590355,18.252264,18.684393,18.855871,19.301718,19.939621,19.555508,19.106232,18.948471,18.862732,19.263992,18.87645,18.516342,18.495766,18.62609,18.61923,18.392878,18.097933,17.947031,18.193962,17.971039,18.04649,18.056778,18.022482,18.331144,18.910746,19.86417,20.351171,20.502073,21.421204,22.155134,23.341772,24.569565,24.631298,21.52066,32.317,34.042084,29.700228,22.161995,14.171056,7.706283,5.638242,6.8145905,8.237869,5.0826488,5.254128,5.435896,5.3090014,5.0277753,5.223262,6.358455,6.7665763,7.438775,8.570539,9.544542,10.034973,10.604284,11.736049,13.457702,15.340545,16.94902,18.910746,20.37518,21.013083,21.04395,20.484926,21.016512,22.354052,23.900795,24.747904,25.543568,24.490685,23.376068,22.95423,22.967947,23.238884,23.890507,23.647005,23.424082,26.335802,24.950249,23.389786,22.19286,22.02824,23.715597,27.772799,29.707087,31.565924,29.467016,13.591455,4.846007,1.6736387,0.9602845,0.8676856,0.84024894,1.611906,1.7182233,3.316411,5.6039457,4.787704,4.712253,5.381023,5.3878818,5.127233,6.7802944,6.9826403,9.349055,9.571979,7.9120584,9.211872,9.880642,11.814929,13.413116,13.227919,9.97667,10.261326,8.110974,7.157549,7.98408,8.117833,10.748327,8.381912,5.6965446,5.1580997,7.0203657,7.3358874,7.747438,7.332458,5.7274113,3.1277838,1.2003556,0.5212973,0.39440256,0.33952916,0.09259886,0.061732575,0.041155048,0.030866288,0.030866288,0.020577524,0.017147938,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.01371835,0.07545093,0.22292319,0.5727411,1.1111864,1.6084765,2.0680413,2.7299516,2.1434922,1.9754424,2.0714707,2.3321195,2.719663,2.054323,1.3992717,1.0871792,1.1008976,1.1077567,1.2483698,1.6393428,2.0817597,2.4555845,2.719663,3.2135234,3.7211025,4.1943855,4.4687524,4.249259,3.0626216,2.6853669,2.8328393,3.1277838,3.0866287,3.0523329,3.100347,3.0900583,3.1826572,3.858286,4.945465,6.3138704,7.4765005,8.368194,9.338767,10.751757,11.375941,11.478829,11.502836,12.05843,13.248496,13.622321,13.38568,13.118172,13.776653,14.140189,14.555169,14.699212,14.544881,14.359683,14.339106,14.839825,15.069608,15.0456,15.6252,15.940722,15.587475,15.343974,15.3817,15.254805,15.398848,16.20137,16.88043,17.329706,18.118511,19.761284,19.932762,20.169403,20.776442,20.855322,21.308027,21.304598,21.239435,21.256582,21.222288,21.04395,22.508383,21.626978,17.192522,10.7757635,10.374502,11.694893,12.542002,12.775213,14.325387,16.383139,17.254255,19.871029,24.171732,27.124607,26.047716,23.451519,22.964518,25.416672,28.832542,28.757092,28.678211,29.487593,31.373867,33.81573,35.307602,37.269325,38.644592,38.630875,36.652,27.954567,16.942162,8.399059,5.8988905,11.80121,8.704293,7.1095347,7.822889,9.788043,10.069269,5.439326,2.4830213,1.471293,2.5310357,5.6348124,4.99005,7.3427467,9.030104,9.253027,10.065839,10.192734,9.033533,9.873782,13.207341,16.777542,21.318316,21.061096,17.247395,11.8869505,7.740579,8.580828,7.6274023,6.0635104,5.0312047,5.6176643,4.650521,4.331569,4.5167665,4.955754,5.3158607,6.3207297,6.910619,8.193284,9.527394,8.536243,10.065839,9.671436,9.424506,10.347065,12.394529,13.522863,13.581166,12.826657,12.236768,13.519434,14.030442,14.870691,15.282242,15.230798,15.426285,16.475739,16.636929,15.820687,14.421415,13.310229,15.117621,16.654078,17.95389,18.897026,19.188541,17.95389,17.425734,17.95046,19.325726,20.807306,20.313446,18.025911,16.29397,15.683503,14.970149,13.749216,13.327377,13.008426,12.428825,11.526843,10.302481,10.508256,11.444533,12.38424,12.562579,13.529722,13.786942,14.483148,15.721229,16.561478,15.29253,13.684054,12.13731,11.080997,10.978109,11.718901,11.770344,11.674315,11.516555,10.926665,11.245617,11.043272,11.153018,11.585147,11.533703,10.652299,11.513125,12.418536,12.682614,12.644889,15.728088,17.151367,17.648657,17.772121,17.87501,17.37429,16.564907,15.340545,14.123041,13.865822,13.310229,12.569438,11.753197,11.036412,10.659158,10.38479,9.938945,9.3936405,8.786603,8.1487,8.172707,8.56368,9.095266,9.410788,9.0369625,9.0644,9.47938,9.6645775,9.770895,10.731179,11.379372,11.153018,10.816919,10.583707,10.089847,10.100135,9.777754,9.462232,9.373062,9.592556,9.122703,9.623423,10.240748,10.343636,9.537683,9.1981535,9.071259,8.838047,8.484799,8.296172,7.8263187,7.5416627,7.3358874,7.2158523,7.274155,7.6376915,8.035523,8.868914,9.822338,9.853205,8.721441,8.176137,7.98408,7.932636,7.840037,0.36696586,0.40126175,0.42869842,0.48014224,0.59331864,0.823101,0.7373613,0.4972902,0.36353627,0.41498008,0.548734,0.48700142,0.44584638,0.4389872,0.42526886,0.29151493,0.24007112,0.26407823,0.3566771,0.48014224,0.5658819,0.6241849,0.51100856,0.4389872,0.490431,0.6241849,0.58988905,0.52472687,0.50757897,0.5624523,0.67219913,0.64819205,0.6859175,0.7305021,0.7476501,0.7476501,0.69963586,0.8779744,0.9842916,0.96714365,1.0528834,1.0666018,1.0597426,1.0220171,0.97057325,0.94656616,1.3992717,1.4815818,1.5673214,1.7422304,1.8142518,2.194936,2.5996273,3.1243541,3.6936657,4.057202,3.5599117,3.07634,2.867135,2.877424,2.7299516,2.3389788,2.4624438,2.8156912,3.0454736,2.7162333,1.6290541,0.75450927,0.22978236,0.0548734,0.09259886,0.10288762,0.06859175,0.044584636,0.041155048,0.01371835,0.0274367,0.020577524,0.010288762,0.0034295875,0.01371835,0.07545093,0.082310095,0.06516216,0.072021335,0.18176813,0.45270553,0.40126175,0.22292319,0.06516216,0.01371835,0.01371835,0.19891608,0.32581082,0.37039545,0.5041494,0.6756287,0.48700142,0.23321195,0.061732575,0.0,0.0,0.0,0.006859175,0.030866288,0.09259886,0.20234565,0.22978236,0.18519773,0.116605975,0.09259886,0.06859175,0.024007112,0.0,0.030866288,0.15090185,0.06859175,0.09259886,0.26407823,0.45613512,0.3806842,0.2469303,0.14061308,0.072021335,0.041155048,0.01371835,0.23664154,0.13375391,0.21263443,0.4389872,0.24350071,0.90198153,1.2517995,1.3546871,1.2037852,0.71678376,0.6310441,0.7373613,0.922559,1.0220171,0.84024894,0.53501564,0.7133542,0.64819205,0.24007112,0.044584636,0.31552204,0.20920484,0.09602845,0.1371835,0.26064864,0.33266997,0.4046913,0.6001778,0.84024894,0.84024894,0.5212973,0.48700142,0.548734,0.5761707,0.5041494,0.58988905,0.8676856,0.89855194,0.66533995,0.5796003,0.64133286,0.5727411,0.5178677,0.4938606,0.39783216,0.4081209,0.44927597,0.39440256,0.29494452,0.3806842,0.2709374,0.40126175,0.48014224,0.4664239,0.5658819,0.42869842,0.39783216,0.48700142,0.65162164,0.7476501,0.66191036,0.65848076,0.66533995,0.66533995,0.70306545,0.59331864,0.5007198,0.5727411,0.72707254,0.64133286,0.5418748,0.66533995,0.805953,0.8676856,0.85396725,1.3066728,1.786815,2.2806756,2.6647894,2.6990852,2.884283,2.867135,2.867135,2.9288676,2.9288676,3.0523329,3.2821152,3.7279615,4.2526884,4.4859004,4.15666,4.9420357,5.4496145,5.336438,5.3261495,5.24041,5.5559316,6.0223556,6.2144127,5.552502,6.090947,6.0223556,5.4496145,5.0003386,5.830299,6.23156,7.130112,8.327039,9.489669,10.1481495,10.110424,9.956093,9.606275,9.211872,9.126132,9.856634,10.196163,10.813489,11.7086115,12.22305,12.8197975,12.932974,13.697772,15.117621,16.081335,16.729528,17.394867,17.95046,18.656956,20.155685,19.973917,19.709839,19.085653,18.44775,18.752985,19.840164,19.058218,17.689812,16.695232,16.70895,16.489456,16.221949,16.047039,15.875561,15.412566,16.05733,16.722668,16.997036,16.976458,17.257685,18.001905,18.718689,19.593233,20.62554,21.650986,23.27661,23.489244,23.917942,24.888515,25.450968,30.26268,34.50165,33.860317,27.320093,17.151367,10.010965,6.8591747,6.2144127,5.888602,3.0214665,3.3747141,3.8034124,4.1017866,4.184097,4.07435,4.770556,5.055212,5.446185,6.0806584,6.715132,7.1061053,8.052671,10.124143,12.545431,13.227919,16.37971,18.821575,20.104242,20.53294,21.177702,21.496655,22.12427,23.225166,24.367218,24.552416,26.040857,25.505842,25.053137,24.919382,23.468666,24.140865,24.079134,23.249174,23.564695,28.901134,27.337242,22.46037,19.078794,18.03963,16.221949,20.395756,20.762722,24.175161,26.421541,12.236768,4.3521466,1.7319417,1.0906088,0.84024894,1.0837497,2.170929,2.3972816,3.316411,4.5922174,3.981751,6.4373355,5.693115,5.219832,6.3035817,8.086967,7.380472,8.100685,7.8674736,6.3893213,5.4633327,7.257007,8.988949,10.134431,9.914937,7.2775846,6.3618846,5.0174866,4.839148,5.6656785,5.5559316,5.528495,5.3330083,5.720552,8.131552,14.661487,9.633711,6.941485,4.695105,2.3595562,0.7476501,0.34638834,0.20920484,0.15090185,0.09259886,0.030866288,0.030866288,0.030866288,0.037725464,0.044584636,0.044584636,0.020577524,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.07545093,0.06516216,0.70306545,1.3375391,1.5570327,1.1900668,1.3478279,1.0597426,0.91912943,1.0460242,1.0837497,0.77851635,0.7305021,0.71678376,0.6927767,0.77851635,1.0940384,1.5124481,1.6496316,1.646202,2.1812177,2.8054025,3.1449318,3.4844608,3.882293,4.149801,3.7965534,3.2512488,3.0660512,3.2203827,3.0969174,3.1826572,3.1140654,3.2718265,3.882293,5.003768,6.433906,7.1095347,7.4353456,7.7268605,8.241299,9.9869585,10.899229,11.5645685,12.1921835,12.617453,13.155897,12.9707,12.445972,12.065289,12.421966,13.557159,14.21564,14.527733,14.675205,14.908417,15.247946,15.673215,15.515453,15.162207,16.0539,16.112202,15.916716,15.728088,15.7795315,16.280252,16.80498,17.432592,17.895588,18.28999,19.058218,19.901896,19.908754,19.884748,20.172834,20.659836,21.260014,20.930773,20.522652,20.62554,21.575535,22.44322,23.465237,23.753323,21.102251,12.006986,10.690024,13.365103,14.195063,12.713481,13.824667,16.009314,17.936743,20.759293,24.915953,30.149504,31.751122,27.326952,22.889067,20.79016,19.716698,18.115082,17.223389,16.897577,17.418875,19.469769,18.44775,20.807306,23.787619,26.812515,31.524769,29.401854,19.678972,9.849775,5.147811,8.529384,7.589677,7.2432885,8.23444,10.621432,13.7938,5.188966,1.5536032,0.6241849,1.1900668,3.083199,5.0346346,7.0718093,11.9040985,17.182234,15.488017,15.817257,15.707511,17.062197,20.917053,27.43327,27.618467,23.818485,18.509483,14.027013,12.572867,10.484249,8.23444,6.6705475,5.8988905,5.2644167,4.5819287,4.6848164,5.453044,6.355026,6.4407654,7.366754,7.023795,8.519095,11.026124,9.781183,9.266746,8.700864,8.824328,10.024684,12.343085,13.406258,12.88496,12.816368,13.910407,15.532601,15.398848,15.896138,15.995596,15.755525,16.341984,18.12537,18.423744,17.813278,16.835844,16.005884,14.79867,15.0456,16.37628,17.833855,17.881868,17.12736,17.082775,17.017612,16.767254,16.753534,17.802988,17.96418,17.63494,16.849564,15.275383,13.725209,13.032433,12.521424,11.856084,11.063849,11.183885,11.324498,11.8869505,12.754636,13.306799,13.903547,13.430264,13.461131,14.390549,15.426285,15.134769,13.697772,11.89038,10.696883,11.30735,11.842365,12.144169,12.123591,11.866373,11.595435,12.267634,12.3911,12.127021,11.410237,9.932085,11.238758,13.718349,15.433144,15.306249,13.121602,14.466,15.570327,15.96816,15.933864,16.496315,16.386568,15.093615,13.927555,13.365103,13.063298,12.9638405,12.281353,11.249047,10.39165,10.511685,10.401938,10.2921915,10.072699,9.589127,8.635701,8.416207,8.964942,9.424506,9.304471,8.498518,8.584257,8.971801,9.455373,9.815479,9.825768,10.436234,11.204462,11.581717,11.516555,11.444533,10.515115,9.908078,9.829198,10.1652975,10.484249,9.993818,9.962952,10.4533825,10.844356,9.8429165,9.571979,9.057541,8.697433,8.549961,8.330468,8.330468,8.1487,7.9086285,7.7131424,7.630832,7.936065,8.543102,9.342196,9.97667,9.8429165,8.378482,7.7268605,7.3255987,7.143831,7.706283,0.4629943,0.4698535,0.5212973,0.5796003,0.6173257,0.6036074,0.6276145,0.6241849,0.64476246,0.66876954,0.59674823,0.5178677,0.490431,0.47671264,0.45270553,0.4355576,0.48357183,0.5693115,0.6276145,0.6344737,0.6001778,0.6344737,0.6379033,0.65505123,0.67219913,0.6001778,0.5555932,0.5624523,0.59331864,0.6379033,0.70649505,0.8093826,0.823101,0.8025235,0.7956643,0.84367853,0.805953,0.84367853,0.939707,1.0734608,1.2003556,1.2517995,1.1077567,1.0323058,1.1900668,1.6530612,1.6084765,1.6633499,1.8313997,2.0131679,1.9994495,2.1126258,2.4315774,3.1620796,4.012617,4.1943855,3.3712845,3.2992632,3.3850029,3.3987212,3.4776018,3.0077481,3.2135234,3.9337368,4.2423997,2.4487255,1.1283343,0.5144381,0.25721905,0.18519773,0.31209245,0.25378948,0.33609957,0.26750782,0.06516216,0.05144381,0.0548734,0.037725464,0.041155048,0.09602845,0.23664154,0.36353627,0.21263443,0.12003556,0.216064,0.41498008,0.25378948,0.15433143,0.07888051,0.024007112,0.01371835,0.034295876,0.16462019,0.28122616,0.32581082,0.28465575,0.34638834,0.32581082,0.24007112,0.12346515,0.01371835,0.0034295875,0.0,0.006859175,0.020577524,0.041155048,0.08573969,0.14747226,0.18176813,0.16804978,0.10288762,0.05144381,0.020577524,0.017147938,0.044584636,0.12689474,0.30523327,0.4629943,0.48700142,0.38754338,0.29494452,0.17147937,0.082310095,0.034295876,0.030866288,0.06516216,0.1371835,0.25721905,0.58302987,0.8848336,0.52472687,1.3101025,1.3615463,1.155771,1.0048691,1.0357354,0.70649505,0.64133286,0.6379033,0.66191036,0.8505377,0.5761707,0.432128,0.37039545,0.31895164,0.1920569,0.18862732,0.17490897,0.22292319,0.31209245,0.30866286,0.274367,0.45270553,0.64819205,0.7407909,0.6790583,0.6276145,0.7922347,0.89169276,0.84367853,0.7613684,0.84367853,0.82996017,0.7339317,0.607037,0.53158605,0.44584638,0.4355576,0.490431,0.52472687,0.4081209,0.40126175,0.33952916,0.35324752,0.44584638,0.5041494,0.37382504,0.490431,0.5727411,0.5590228,0.58988905,0.5144381,0.5453044,0.59331864,0.6241849,0.6756287,0.77508676,0.70649505,0.66876954,0.6893471,0.6276145,0.5178677,0.52815646,0.6036074,0.7339317,0.97057325,1.1077567,1.0528834,0.97400284,0.980862,1.1351935,1.3821237,1.8108221,2.411,2.9665933,3.0420442,3.4295874,3.8137012,4.2046742,4.461893,4.297273,4.331569,4.461893,4.557922,4.6676683,4.98662,4.7945633,4.98662,5.254128,5.4736214,5.717122,5.40503,6.0395036,6.574519,6.5710897,6.2247014,6.478491,6.3721733,6.5059276,6.852316,6.7459984,6.355026,6.5642304,7.233,8.210432,9.328478,9.750318,9.650859,9.211872,8.738589,8.673427,8.937505,9.561689,10.525404,11.633161,12.5145645,12.878101,12.919256,13.344524,14.243076,15.069608,15.707511,16.221949,16.95931,18.080786,19.582945,19.634388,19.469769,18.931322,18.324286,18.423744,18.787281,18.259123,17.2131,16.074476,15.306249,15.337115,15.409137,15.532601,15.515453,14.935853,15.542891,15.978448,15.930434,15.645778,15.927004,16.770683,17.04162,17.604073,18.746124,20.21056,22.302607,23.19087,24.072275,25.60873,27.916842,31.768269,38.373653,35.75002,24.363789,17.113642,13.029003,9.009526,5.857735,3.8445675,2.702515,2.726522,2.9974594,3.4947495,4.029765,4.232111,4.420738,4.554492,4.448175,4.256118,4.479041,5.435896,6.608815,8.536243,10.97468,12.898679,14.898128,17.734396,19.236557,19.586374,21.325174,21.846472,21.980227,22.408924,23.280039,24.185452,24.247183,23.43094,23.166862,23.550978,23.358921,24.11686,24.487255,24.206028,24.706749,29.130917,28.798246,23.60928,18.238546,15.45715,16.108772,16.194511,16.856422,20.755863,23.338343,12.836946,5.096367,1.9480057,0.8779744,0.5727411,0.9259886,1.5124481,1.488441,2.054323,3.2786856,4.105216,6.3618846,4.972902,4.3692946,5.501058,5.830299,4.9077396,4.787704,4.962613,5.346727,6.3035817,5.5490727,6.5779486,7.3290286,7.3187394,7.630832,6.4819202,5.5113473,5.4153185,5.953764,5.9331865,9.424506,10.244178,10.868362,11.698323,11.050131,11.71547,11.958971,8.964942,3.724532,1.039165,0.4424168,0.23321195,0.20920484,0.20234565,0.09259886,0.061732575,0.0548734,0.06516216,0.07888051,0.06859175,0.044584636,0.024007112,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.19891608,0.5418748,0.78537554,0.8196714,0.6790583,0.7888051,0.6036074,0.44584638,0.41840968,0.38754338,0.36696586,0.36696586,0.40126175,0.4938606,0.66876954,0.7407909,1.0837497,1.3341095,1.4438564,1.670209,2.3424082,2.6613598,2.959734,3.2581081,3.2718265,3.2512488,3.0660512,2.7745364,2.534465,2.5961976,2.8396983,2.8294096,3.100347,4.0537724,5.967482,6.742569,7.39762,7.970361,8.639131,9.729739,11.201033,11.921246,12.319078,12.6757555,13.13189,13.423406,13.097594,12.459691,11.979549,12.284782,12.922686,13.598314,14.040731,14.212211,14.29795,14.668345,15.2033615,15.601193,15.899568,16.479168,16.815268,16.585485,16.424294,16.582056,16.914726,17.63494,17.95732,18.320856,18.852442,19.387459,20.073376,20.093952,20.080235,20.241425,20.36832,20.663265,20.584383,20.241425,20.145397,21.184563,22.28546,23.184011,23.084553,20.296299,12.21619,10.731179,14.500296,16.160215,14.706071,15.484588,16.743246,17.494326,19.11652,22.127699,26.171183,29.635065,28.613049,26.130028,23.753323,21.592682,20.814167,20.148827,18.746124,17.501184,19.044498,16.269962,17.336565,17.929884,19.346302,28.51016,30.252392,19.9602,8.676856,2.7985435,4.0503426,6.478491,9.328478,10.439664,9.434795,7.716572,5.689686,2.9700227,2.2463799,3.275256,2.8637056,5.9983487,7.267296,9.6988735,13.924125,18.183672,21.77788,25.368658,30.711956,37.49911,43.363705,41.31967,33.58938,25.313786,19.819586,18.591793,13.457702,9.89436,8.862054,9.595985,9.595985,6.9037595,7.140401,6.7802944,5.720552,7.281014,8.999237,10.031544,10.100135,9.510246,9.132992,9.9869585,10.81006,11.976119,13.063298,12.843805,13.4474125,12.9809885,12.55229,12.908967,14.435134,15.597764,16.897577,17.497755,17.463459,17.758404,18.945042,19.36688,19.45262,19.301718,18.667244,17.117071,16.393429,16.516893,17.178804,17.737827,17.78927,18.30028,18.890167,19.442331,20.12139,19.658396,19.075365,18.37573,17.449741,16.081335,15.29939,14.085316,12.665466,11.492548,11.245617,11.046701,11.646879,12.336226,13.011855,14.184773,15.3302555,14.79524,14.0750265,13.745787,13.485138,12.442543,11.393089,11.002116,11.269625,11.537132,12.699762,12.768354,12.548861,12.3911,12.181894,12.600305,12.696333,12.164746,11.4205265,11.592006,11.862943,13.101024,14.3974085,14.891269,13.7697935,14.760944,15.395418,15.6526375,15.690363,15.858413,15.29939,14.688923,13.96185,13.296511,13.097594,12.9809885,12.144169,11.231899,10.72432,10.964391,11.214751,11.153018,10.786053,10.065839,8.879202,8.388771,8.412778,8.594546,8.608265,8.182996,8.597976,8.711152,9.115844,9.80519,10.168727,9.880642,10.017825,10.549411,11.14273,11.177026,10.686595,10.196163,10.1652975,10.556271,10.823778,10.580277,10.508256,10.666017,10.748327,10.096705,9.205012,8.848335,8.56025,8.1487,7.6857057,7.421627,7.675417,7.891481,7.8846216,7.8503256,7.9086285,8.433355,9.2153015,9.80862,9.537683,8.453933,8.351046,8.285883,8.152129,8.694004,0.4698535,0.45613512,0.5178677,0.59331864,0.6276145,0.5761707,0.5590228,0.5624523,0.5796003,0.5796003,0.5007198,0.47328308,0.5007198,0.52472687,0.5453044,0.61046654,0.61046654,0.6173257,0.6173257,0.6036074,0.5658819,0.6824879,0.66876954,0.64133286,0.6276145,0.58645946,0.65505123,0.6927767,0.71678376,0.7305021,0.72707254,0.8093826,0.82996017,0.7956643,0.7613684,0.8162418,0.8676856,0.89855194,0.9602845,1.0220171,0.9877212,1.0117283,0.9911508,1.0597426,1.2758065,1.6221949,1.5536032,1.6496316,1.8348293,1.9857311,1.9239986,2.061182,2.719663,3.6147852,4.2869844,4.108646,3.542764,3.6182148,3.9303071,4.3109913,4.8322887,3.8479972,3.981751,4.773986,5.192395,3.6147852,1.3375391,1.8931323,1.8999915,0.66533995,0.20920484,0.13032432,0.19548649,0.22292319,0.16804978,0.09602845,0.07545093,0.041155048,0.030866288,0.07888051,0.19891608,0.21263443,0.13032432,0.18519773,0.37382504,0.45613512,0.20920484,0.07888051,0.0274367,0.01371835,0.006859175,0.044584636,0.25378948,0.47328308,0.53844523,0.25721905,0.29151493,0.28465575,0.21263443,0.09945804,0.006859175,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.037725464,0.07545093,0.1097468,0.13032432,0.106317215,0.07545093,0.037725464,0.020577524,0.037725464,0.058302987,0.25721905,0.5796003,0.65162164,0.47328308,0.42183927,0.16804978,0.082310095,0.10288762,0.18862732,0.33266997,0.31895164,0.4115505,0.58988905,0.764798,0.7888051,1.5330256,1.4164196,1.155771,1.0014396,0.764798,0.47671264,0.47328308,0.45270553,0.40126175,0.5693115,0.44927597,0.3018037,0.25721905,0.3018037,0.25721905,0.2709374,0.23664154,0.26407823,0.33952916,0.31209245,0.31552204,0.5144381,0.64476246,0.66533995,0.7613684,0.91912943,0.85739684,0.8162418,0.89169276,1.0357354,1.0597426,0.8711152,0.6962063,0.6001778,0.48357183,0.47671264,0.42526886,0.38754338,0.39097297,0.42869842,0.30866286,0.31552204,0.3841138,0.4389872,0.41498008,0.59674823,0.66533995,0.65162164,0.6036074,0.58645946,0.607037,0.59674823,0.5693115,0.5555932,0.6379033,0.7922347,0.6962063,0.6790583,0.7613684,0.64819205,0.58988905,0.65848076,0.7373613,0.7888051,0.8779744,1.08032,1.0528834,1.0357354,1.1420527,1.3512574,1.3855534,1.7936742,2.4590142,3.0900583,3.210094,3.642222,4.091498,4.4756117,4.65395,4.4447455,4.6127954,5.0140567,5.302142,5.3844523,5.40503,5.144381,5.07236,5.096367,5.2609873,5.7479887,5.470192,5.9812007,6.3173003,6.293293,6.495639,6.7871537,6.7665763,6.931196,7.1781263,6.807731,6.451054,6.711703,7.140401,7.6171136,8.375052,8.690575,8.796892,8.738589,8.608265,8.56025,8.721441,9.31133,10.055551,10.72432,11.115293,12.0138445,12.4974165,13.029003,13.732068,14.387119,14.750656,15.172495,15.858413,16.938732,18.468328,19.188541,19.524641,19.143957,18.197392,17.353712,16.942162,16.355703,15.844694,15.45715,15.035312,15.470869,15.889278,16.21166,16.29054,15.906426,15.902997,16.009314,15.608052,14.904987,14.935853,15.361122,16.050468,17.141079,18.44432,19.44919,20.882757,21.421204,22.072824,23.554407,26.26378,29.840841,34.210136,31.133795,21.7916,16.80155,15.834405,12.538571,7.6788464,3.2683969,2.5619018,2.3904223,2.5070283,2.8122618,3.1963756,3.5118976,3.6559403,3.8548563,3.882293,3.74168,3.666229,4.5956473,5.65539,7.425057,9.884071,12.397959,14.411126,16.743246,17.569777,17.192522,18.04992,18.849012,19.915615,21.417774,22.974806,23.671013,23.489244,22.666143,22.19972,22.131128,21.572105,22.707298,23.996824,24.816494,25.745913,28.575323,27.659622,23.883648,18.71526,14.79867,15.971589,15.830976,17.885298,20.21399,19.229696,9.6988735,4.098357,1.728512,0.82996017,0.5007198,0.66533995,1.1934965,1.1214751,1.5776103,2.4898806,2.568761,4.40702,3.8034124,3.192946,3.3438478,3.3609958,3.1312134,2.9906003,3.0214665,3.4913201,4.8768735,4.746549,5.4941993,5.7411294,5.8405876,7.8949103,6.8111606,6.468202,6.9346256,7.3598948,5.9914894,11.135871,14.201921,14.970149,14.249936,13.88297,16.650646,15.824117,10.782623,4.0023284,1.039165,0.5041494,0.2709374,0.24350071,0.274367,0.17833854,0.106317215,0.06516216,0.05144381,0.0548734,0.058302987,0.041155048,0.024007112,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15090185,0.29494452,0.37382504,0.37725464,0.36696586,0.36010668,0.28122616,0.22978236,0.20920484,0.12346515,0.15776102,0.1920569,0.29151493,0.4355576,0.51100856,0.6859175,0.939707,1.2277923,1.4438564,1.4232788,1.7902447,1.9925903,2.3732746,2.8637056,2.959734,2.9185789,2.5961976,2.1503513,1.8554068,2.1057668,2.3561265,2.585909,3.2066643,4.5099077,6.64997,7.298162,7.874333,8.81404,10.021255,10.88894,12.349944,12.895248,12.891819,12.871242,13.526293,14.225929,13.728639,12.936404,12.538571,12.984418,13.279363,13.718349,13.975569,14.064738,14.356253,15.035312,15.494876,15.944152,16.503176,17.20967,17.436022,17.137648,16.822126,16.753534,16.938732,17.55263,17.806417,17.998474,18.296848,18.739265,19.384027,19.54179,19.53836,19.579515,19.716698,19.425184,19.552078,19.510923,19.576086,20.886189,21.908205,22.237446,22.258022,20.61182,14.198492,12.593445,15.824117,17.638369,16.928444,17.71382,18.36544,18.691252,19.54522,21.349182,24.085993,28.458717,29.02117,27.985434,26.325514,23.78419,22.765602,21.928782,20.159115,18.163095,18.451181,15.2033615,15.594335,15.776102,16.863281,24.898806,26.76107,17.312557,7.3358874,3.7313912,9.5205345,8.069819,14.493437,17.391438,14.325387,11.842365,9.794902,8.296172,8.241299,9.386781,10.360784,16.640358,26.809086,43.751247,60.299007,59.259842,40.22906,40.184475,46.940765,52.980267,55.44957,49.656998,41.676346,33.616817,26.548437,20.498644,16.081335,13.203912,11.355364,10.295622,10.05898,10.076128,8.755736,6.8797526,5.645101,6.64997,8.484799,10.412228,10.662587,9.424506,8.862054,9.613133,10.549411,11.821788,12.833516,12.229909,13.6086035,13.38911,12.6757555,12.449403,13.54687,15.556609,17.021042,17.652086,17.878439,18.852442,19.809298,20.817596,21.541239,21.644127,20.78673,19.634388,18.499195,17.847572,17.648657,17.353712,18.677534,19.349733,20.069946,21.061096,22.055677,21.558388,20.570665,19.250275,17.809847,16.527182,15.892709,14.805529,13.588025,12.476839,11.657167,11.664027,12.511135,13.519434,14.171056,14.112752,15.011304,14.791811,14.071597,13.197053,12.229909,11.012405,10.672876,11.156448,11.993267,12.291641,13.543441,13.992717,13.519434,12.600305,12.312219,13.896688,14.160767,13.320518,12.21619,12.312219,12.476839,13.21763,14.345964,15.340545,15.350834,15.806969,15.978448,15.79325,15.234227,14.318527,14.160767,14.099034,13.728639,13.179905,13.125031,12.600305,11.55428,10.97468,11.067279,11.2593355,11.478829,11.574858,11.211322,10.419086,9.626852,8.862054,8.625413,8.584257,8.618553,8.81747,8.862054,8.848335,9.235879,10.010965,10.676306,10.031544,10.038403,10.364213,10.655728,10.549411,10.360784,10.134431,10.172156,10.39508,10.350495,10.477389,10.504827,10.545981,10.528833,10.172156,9.458802,8.934075,8.416207,7.949784,7.805741,7.534804,7.7028537,8.076678,8.464222,8.718011,8.200144,8.340756,8.862054,9.355915,9.321619,8.985519,8.899779,8.862054,8.875772,9.14328,0.6276145,0.6344737,0.6859175,0.69963586,0.66191036,0.6241849,0.5555932,0.5144381,0.5144381,0.53844523,0.53844523,0.6173257,0.6859175,0.7133542,0.71678376,0.7442205,0.6756287,0.6241849,0.6344737,0.6756287,0.6379033,0.7133542,0.67219913,0.6207553,0.607037,0.6276145,0.6927767,0.70306545,0.69963586,0.7099246,0.7373613,0.7613684,0.8025235,0.78537554,0.72707254,0.72364295,0.78537554,0.84367853,0.89169276,0.88826317,0.77508676,0.77851635,0.8848336,1.0768905,1.2758065,1.3512574,1.5261664,1.6633499,1.7525192,1.8176813,1.9239986,2.2635276,3.1517909,3.981751,4.3624353,4.1189346,3.9543142,4.232111,4.7088237,5.3227196,6.200694,5.0826488,5.0106273,4.928317,4.5167665,4.197815,1.8588364,2.609916,2.7951138,1.7765263,1.9445761,0.432128,0.116605975,0.1920569,0.22978236,0.17833854,0.09259886,0.058302987,0.072021335,0.10288762,0.09945804,0.058302987,0.0548734,0.1920569,0.39783216,0.45613512,0.22635277,0.07888051,0.01371835,0.010288762,0.01371835,0.030866288,0.2777966,0.53158605,0.58988905,0.25721905,0.26750782,0.26750782,0.18862732,0.058302987,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.030866288,0.030866288,0.044584636,0.06859175,0.06859175,0.08573969,0.05144381,0.024007112,0.017147938,0.010288762,0.11317638,0.47328308,0.6276145,0.53501564,0.5727411,0.216064,0.14747226,0.21263443,0.33609957,0.5041494,0.65162164,0.6207553,0.66533995,0.7956643,0.7922347,1.3341095,1.3203912,1.1489118,0.9259886,0.48014224,0.32924038,0.30523327,0.26407823,0.20234565,0.28465575,0.26407823,0.25378948,0.2777966,0.30866286,0.25721905,0.4355576,0.4046913,0.4698535,0.607037,0.4389872,0.42869842,0.53501564,0.61046654,0.69963586,1.0357354,1.0460242,0.7579388,0.7476501,1.0528834,1.1489118,1.0117283,0.89169276,0.7442205,0.5796003,0.48700142,0.47328308,0.4629943,0.3841138,0.30866286,0.4355576,0.34981793,0.4424168,0.53844523,0.53844523,0.42183927,0.72021335,0.7510797,0.7133542,0.6859175,0.6344737,0.65848076,0.59674823,0.52815646,0.51100856,0.5761707,0.8025235,0.6824879,0.65162164,0.78194594,0.7442205,0.66533995,0.6824879,0.7990939,0.939707,0.9568549,1.1351935,1.1592005,1.1454822,1.2003556,1.4198492,1.4232788,1.7936742,2.3321195,2.8294096,3.0900583,3.4707425,3.8342788,4.1463714,4.341858,4.3007026,4.2252517,4.7808447,5.4804807,5.9297566,5.8062916,5.381023,5.2266912,5.055212,4.99005,5.597087,5.5387836,5.744559,5.861165,5.9983487,6.7459984,6.914048,6.6396813,6.584808,6.824879,6.8557453,6.4236174,6.8111606,7.099246,7.133542,7.5245147,7.888051,8.224151,8.491658,8.676856,8.81747,9.054111,9.599416,10.216741,10.63858,10.566559,11.547421,12.130451,12.881531,13.865822,14.671775,14.767803,15.13134,15.6526375,16.37628,17.487467,18.20425,18.807858,18.849012,18.221397,17.158226,16.088194,15.29253,14.870691,14.784951,14.846684,15.834405,16.540901,17.021042,17.243965,17.089634,16.647217,16.311117,15.680074,15.018164,15.265094,15.29596,16.084764,17.237106,18.413456,19.322296,20.083664,19.77843,19.764713,20.875898,23.420652,26.713057,30.667372,28.287237,20.759293,17.487467,16.846134,14.181344,8.920357,3.2821152,2.2909644,2.0920484,2.136633,2.1846473,2.2566686,2.609916,2.6545007,2.983741,3.2649672,3.4021509,3.532475,4.139512,4.7534084,6.1972647,8.508806,10.957532,13.2862215,15.062748,15.4914465,15.079896,15.611482,16.180794,18.115082,20.35803,21.93221,21.956219,22.144846,21.602972,21.232576,21.074816,20.28601,21.589252,23.304047,24.7822,26.229485,28.712505,28.311245,25.039417,19.95677,15.512024,15.539461,14.54831,16.750105,17.754974,14.740367,6.4579134,2.7916842,1.4815818,1.0357354,0.7442205,0.6962063,1.1489118,1.0597426,1.313532,1.7936742,1.4027013,2.386993,2.4658735,2.0577524,1.605047,1.5673214,1.8554068,2.0749004,2.2292318,2.633923,3.9063,4.5990767,5.312431,5.429037,5.5593615,7.5279446,6.5470824,6.5710897,7.2604365,7.970361,7.7542973,11.89038,14.730078,15.841265,15.9578705,16.990177,19.353163,16.585485,10.213311,3.415869,1.0117283,0.72364295,0.40126175,0.26407823,0.3018037,0.3018037,0.29837412,0.18176813,0.12346515,0.14404267,0.11317638,0.06516216,0.037725464,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.12689474,0.15433143,0.15433143,0.14747226,0.14747226,0.11317638,0.1371835,0.17490897,0.18176813,0.1097468,0.106317215,0.15090185,0.25378948,0.37039545,0.3841138,0.64476246,0.77851635,0.9602845,1.1351935,1.0254467,1.1592005,1.4198492,1.8039631,2.2292318,2.4967396,2.4487255,2.1126258,1.7388009,1.5433143,1.7147937,2.0646117,2.4727325,3.3301294,4.6882463,6.258997,7.1987042,7.6376915,8.745448,10.347065,10.926665,12.55915,13.265644,13.38225,13.505715,14.472859,15.12448,14.339106,13.495427,13.334236,13.9309845,14.404267,14.685493,14.743796,14.771234,15.1862135,15.834405,16.269962,16.88386,17.669235,18.228258,18.231688,17.737827,17.250826,17.069057,17.28512,17.847572,18.097933,18.190533,18.255693,18.406595,18.45804,18.595222,18.629519,18.571217,18.636377,18.331144,18.643238,18.890167,19.239986,20.738716,21.599543,21.383478,21.462358,20.457489,14.243076,13.622321,16.842705,18.917604,18.982767,20.299728,21.016512,21.04395,20.995934,21.263443,21.987085,26.833092,28.67135,28.75023,27.789948,26.01342,24.4461,23.122278,21.572105,19.967058,19.147387,15.971589,16.108772,16.37971,17.525192,24.209457,22.213438,13.1421795,5.521636,5.2609873,15.673215,12.418536,21.935642,25.498983,20.930773,22.580404,20.392326,19.397747,21.44178,26.35295,31.939749,40.42798,64.699165,107.38039,147.21848,139.10063,75.05652,60.319584,63.01181,64.95639,61.657124,51.766193,43.830128,38.606865,33.68884,23.506393,22.011093,18.183672,13.978998,11.194174,11.499407,10.967821,8.371623,6.1732574,5.3878818,5.5559316,6.8797526,8.841476,9.668007,9.054111,8.165848,9.160428,10.244178,11.197603,11.945253,12.576297,13.622321,13.245067,12.860953,13.279363,14.699212,16.636929,17.487467,17.566347,17.682953,19.147387,20.35803,21.44864,22.096832,22.175713,21.747015,20.872469,19.977346,19.21255,18.550638,17.785841,19.102802,19.69955,20.258574,21.04052,21.897917,21.668133,20.886189,19.298288,17.463459,16.746675,16.21166,15.409137,14.287662,13.138749,12.562579,13.025573,13.9481325,14.935853,15.419425,14.661487,14.723219,14.507155,14.006435,13.107883,11.585147,10.683165,10.662587,11.5645685,12.932974,13.831526,15.395418,16.252815,15.477728,13.666906,12.926115,14.79524,15.21022,14.479718,13.310229,12.80608,13.491997,14.078457,14.901558,15.827546,16.273392,16.561478,16.846134,16.273392,14.695783,12.672326,13.341095,13.673765,13.485138,12.912396,12.428825,11.900668,11.166737,10.964391,11.345076,11.650309,11.664027,11.787492,11.447963,10.628291,9.866923,9.421077,9.383351,9.47938,9.6988735,10.2921915,9.674867,9.599416,9.938945,10.501397,11.036412,10.299051,10.134431,10.233889,10.2921915,10.024684,9.860064,9.925226,10.113853,10.192734,9.832627,10.100135,10.175586,10.254466,10.30934,10.096705,9.5033865,8.875772,8.361334,8.093826,8.186425,7.966932,7.915488,8.30646,9.006097,9.469091,8.628842,8.361334,8.570539,9.016385,9.297611,9.537683,9.342196,9.119273,9.105555,9.3764925,0.8196714,0.89512235,0.9259886,0.84367853,0.6962063,0.65505123,0.58302987,0.53844523,0.53844523,0.5796003,0.64476246,0.8162418,0.881404,0.864256,0.7990939,0.7373613,0.66876954,0.6344737,0.6962063,0.7888051,0.7442205,0.6790583,0.65162164,0.64476246,0.65162164,0.65505123,0.61046654,0.58302987,0.5693115,0.59674823,0.7133542,0.6962063,0.7373613,0.7476501,0.6962063,0.6241849,0.6207553,0.6859175,0.7476501,0.7510797,0.6859175,0.71678376,0.84367853,1.0494537,1.2243627,1.1592005,1.605047,1.7147937,1.6804979,1.728512,2.1194851,2.651071,3.5016088,4.170378,4.4516044,4.4550343,4.623084,5.2815647,5.909179,6.3790326,6.9723516,6.992929,6.3173003,4.4996185,2.6373527,3.3678548,1.9514352,1.8382589,2.1640697,2.7059445,3.8788633,0.8848336,0.20920484,0.31209245,0.3806842,0.32581082,0.13032432,0.106317215,0.17490897,0.2194936,0.072021335,0.08916927,0.08573969,0.15433143,0.29151493,0.40126175,0.21263443,0.072021335,0.024007112,0.037725464,0.0274367,0.006859175,0.18519773,0.34295875,0.3566771,0.18862732,0.17147937,0.20234565,0.15090185,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.030866288,0.017147938,0.01371835,0.024007112,0.01371835,0.06516216,0.058302987,0.037725464,0.034295876,0.06516216,0.01371835,0.25378948,0.45613512,0.53844523,0.66533995,0.28808534,0.26064864,0.33952916,0.4115505,0.48357183,0.980862,0.83338976,0.823101,0.9842916,0.6036074,0.9294182,1.2003556,1.1351935,0.7476501,0.34638834,0.28808534,0.16462019,0.08573969,0.08573969,0.13032432,0.17833854,0.26750782,0.36010668,0.39783216,0.3018037,0.5624523,0.59331864,0.7579388,0.9534253,0.6344737,0.5624523,0.548734,0.6276145,0.8505377,1.2620882,0.9568549,0.6173257,0.77851635,1.2106444,0.9568549,0.764798,0.82996017,0.77165717,0.5761707,0.61046654,0.48700142,0.5521636,0.5144381,0.3841138,0.4664239,0.53158605,0.67219913,0.764798,0.7510797,0.6379033,0.7099246,0.72707254,0.7579388,0.78194594,0.6790583,0.64819205,0.6207553,0.5796003,0.5418748,0.5693115,0.7922347,0.65848076,0.5761707,0.6756287,0.7956643,0.66191036,0.6173257,0.8093826,1.1454822,1.2758065,1.4164196,1.4369972,1.3101025,1.1832076,1.4061309,1.5055889,1.8108221,2.0508933,2.218943,2.5790498,2.9048605,3.234101,3.6113555,3.957744,4.1017866,3.765687,4.149801,5.0106273,5.8405876,5.8508763,5.435896,5.2609873,4.972902,4.7431192,5.267846,5.6142344,5.6656785,5.6313825,5.861165,6.848886,6.9860697,6.025785,5.562791,6.094377,7.0375133,6.2830043,6.6293926,6.8283086,6.677407,7.0203657,7.6342616,8.110974,8.450503,8.700864,8.961512,9.441654,10.151579,10.902658,11.430815,11.410237,11.873232,12.024134,12.730629,14.05102,15.223939,15.391989,15.806969,16.245956,16.657507,17.175373,17.072487,17.442883,17.929884,18.173384,17.813278,16.46888,15.494876,14.747226,14.291091,14.404267,15.666355,16.503176,17.168514,17.648657,17.679523,17.38115,16.671225,15.902997,15.594335,16.438013,16.486027,16.945591,17.442883,18.056778,19.318867,20.03222,19.047928,18.259123,18.814716,21.139977,24.19231,30.900583,29.820263,21.750444,19.733847,16.187653,13.049581,8.546532,3.6353626,2.0131679,1.6770682,1.6907866,1.6153357,1.488441,1.821111,1.7353712,2.085189,2.4590142,2.8122618,3.4638834,3.799983,3.998899,4.9591837,6.7494283,8.611694,10.971251,12.459691,13.121602,13.526293,14.771234,14.990726,17.113642,19.11309,20.004784,19.857311,20.69413,20.131678,19.929333,20.364891,20.227707,21.390337,22.878778,24.302057,26.10602,29.573332,30.811415,26.496992,20.971928,16.921585,15.402277,12.2093315,13.166186,13.498857,10.72432,4.6127954,1.9171394,1.2689474,1.1832076,0.9945804,0.83681935,1.1351935,0.9945804,0.94656616,1.1283343,1.2998136,1.3649758,1.4678634,1.4335675,1.2483698,1.0906088,1.3101025,1.7696671,2.4384367,3.2066643,3.8788633,4.98662,6.036074,6.3653145,6.2144127,6.728851,5.8200097,5.7891436,6.252138,7.56224,10.792912,12.000127,12.099585,13.581166,16.520323,18.571217,19.161106,14.970149,8.525954,2.867135,1.5090185,1.255229,0.6790583,0.31552204,0.29151493,0.35324752,0.44584638,0.34295875,0.33952916,0.41840968,0.24350071,0.13032432,0.072021335,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.09602845,0.14747226,0.12346515,0.082310095,0.048014224,0.0,0.020577524,0.106317215,0.16119061,0.15776102,0.15090185,0.1097468,0.14061308,0.19548649,0.2469303,0.28465575,0.47328308,0.5212973,0.5555932,0.6001778,0.5521636,0.70649505,1.0871792,1.2998136,1.3615463,1.7319417,1.8073926,1.6942163,1.5501735,1.4472859,1.3889829,1.9342873,2.4487255,3.3541365,4.48933,5.0929375,6.680836,7.0546613,7.932636,9.424506,10.007536,11.729189,12.80265,13.498857,14.208781,15.419425,15.539461,14.4145565,13.677195,13.910407,14.675205,15.731518,15.9921665,16.023033,16.19794,16.702091,16.911295,17.309128,18.193962,19.150816,19.047928,18.886738,18.190533,17.62122,17.549198,18.060207,18.691252,18.999914,19.20569,19.257133,18.831865,17.988186,17.936743,17.905876,17.669235,17.528622,17.813278,18.358582,18.814716,19.322296,20.498644,21.222288,20.899906,21.054237,20.28944,14.308239,15.127911,18.37916,20.244854,20.488356,22.436361,23.722456,23.664154,23.03311,22.041958,20.351171,24.572994,27.18634,27.930561,27.368109,26.870817,25.156025,23.664154,22.70044,21.959648,20.539799,17.724108,17.854433,17.823566,18.578075,25.10801,17.802988,8.913498,3.6147852,5.2987127,15.549749,14.959861,26.260351,29.861418,25.306927,31.277838,30.211235,28.695358,33.60653,45.016766,56.166355,63.51596,93.78207,150.26395,204.78067,197.71915,104.73274,76.79875,74.14768,72.49805,63.049538,50.840206,42.382843,39.615166,38.57943,29.425861,28.832542,21.78474,15.035312,12.168177,13.605173,9.253027,6.701414,5.4667625,5.127233,5.329579,5.9571934,7.010077,7.9120584,8.241299,7.706283,9.321619,10.580277,11.091286,11.516555,13.557159,13.29994,12.812939,13.22106,14.764374,16.780972,18.231688,18.238546,17.847572,17.88873,18.962189,20.128248,20.738716,20.906765,20.978786,21.53095,20.670124,20.385468,19.895037,19.11995,18.674105,18.996485,19.387459,19.689262,19.980776,20.574095,20.423193,20.004784,18.423744,16.46545,16.568336,16.595774,16.191082,14.997586,13.786942,14.452282,15.354263,16.149927,16.719238,16.846134,16.21852,15.3817,14.743796,14.201921,13.344524,11.458252,10.813489,10.786053,11.842365,13.666906,15.179354,17.106783,18.44432,17.923023,15.927004,14.476289,15.021593,15.450292,15.302819,14.613472,13.893259,15.042171,15.4914465,15.762384,16.108772,16.499744,16.822126,17.364002,16.575195,14.232788,11.430815,12.782072,13.371962,13.22106,12.428825,11.166737,11.105004,11.173596,11.31078,11.561139,12.068718,11.996697,11.938394,11.537132,10.690024,9.544542,9.8429165,10.254466,10.779194,11.423956,12.181894,10.923236,10.690024,10.899229,11.14273,11.204462,10.542552,10.021255,9.887501,9.966381,9.674867,9.568549,9.750318,10.069269,10.2236,9.750318,9.801761,9.784613,9.89093,10.034973,9.846346,9.136421,8.680285,8.457363,8.378482,8.292743,8.275595,8.182996,8.529384,9.277034,9.856634,9.06097,8.515666,8.447074,8.81404,9.280463,9.815479,9.623423,9.23245,9.105555,9.637141,0.5658819,0.7476501,0.77508676,0.72021335,0.64476246,0.59674823,0.5693115,0.5453044,0.47328308,0.38754338,0.4115505,0.53501564,0.53844523,0.5007198,0.4698535,0.45613512,0.4938606,0.5041494,0.51100856,0.52472687,0.548734,0.5624523,0.5453044,0.5693115,0.59674823,0.47328308,0.48357183,0.5144381,0.5521636,0.5796003,0.5796003,0.53158605,0.53844523,0.5624523,0.5761707,0.5658819,0.58988905,0.64133286,0.6962063,0.7099246,0.6241849,0.72364295,0.7922347,0.9534253,1.1489118,1.1592005,1.6221949,1.5844694,1.6324836,1.9720128,2.411,2.8739944,3.6593697,4.506478,5.137522,5.2472687,5.689686,6.831738,7.699424,7.682276,6.5470824,9.914937,7.682276,4.1155047,1.7799559,1.5124481,0.5453044,0.22292319,0.7956643,1.5090185,0.59674823,0.216064,0.19548649,0.59331864,1.0117283,0.59674823,0.25378948,0.17833854,0.28122616,0.37725464,0.18176813,0.26750782,0.20920484,0.18176813,0.20577525,0.106317215,0.044584636,0.01371835,0.07888051,0.16119061,0.01371835,0.01371835,0.041155048,0.048014224,0.030866288,0.030866288,0.041155048,0.037725464,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.017147938,0.024007112,0.01371835,0.01371835,0.0274367,0.030866288,0.072021335,0.17490897,0.31895164,0.06516216,0.09945804,0.33266997,0.6036074,0.70306545,0.33609957,0.39097297,0.4938606,0.48357183,0.4115505,1.1317638,0.94656616,0.67219913,0.6173257,0.5796003,0.9842916,1.4129901,1.3101025,0.6859175,0.1371835,0.05144381,0.030866288,0.072021335,0.13032432,0.106317215,0.38754338,0.37382504,0.40126175,0.53501564,0.59674823,0.53501564,0.6379033,0.71678376,0.6962063,0.61046654,0.64819205,0.70306545,0.86082643,1.0425946,1.0082988,0.8848336,0.6173257,0.65162164,0.823101,0.33609957,0.6893471,0.65162164,0.59674823,0.6962063,0.91569984,0.89169276,0.77508676,0.65848076,0.6001778,0.6241849,0.65162164,0.8471081,0.89855194,0.8196714,0.9911508,0.72364295,0.7579388,0.8162418,0.7510797,0.5178677,0.5693115,0.77165717,0.8025235,0.6893471,0.823101,0.6276145,0.5418748,0.45613512,0.4046913,0.5658819,0.52815646,0.7099246,0.9911508,1.2517995,1.371835,1.5330256,1.5158776,1.3889829,1.3101025,1.5398848,1.5536032,1.786815,1.7593783,1.5158776,1.6016173,1.9548649,2.5653315,3.1723683,3.5290456,3.4192986,4.0880685,4.064061,4.2252517,4.6779575,4.7774153,4.996909,4.7774153,4.482471,4.3761535,4.6093655,5.610805,6.0532217,5.90575,5.627953,6.1629686,7.3358874,5.5593615,4.2183924,4.7808447,6.8043017,6.108095,6.48535,6.7219915,6.6396813,7.0786686,7.5690994,7.9909387,8.268735,8.303031,8.011517,9.0369625,10.271614,11.115293,11.55771,12.1921835,12.459691,12.116733,12.109874,12.80608,13.975569,14.96672,15.724659,16.427725,17.161655,17.943602,16.993607,16.753534,17.010754,17.446312,17.655516,16.80155,15.88242,15.093615,14.514014,14.099034,14.503725,15.196502,16.11906,16.983316,17.288551,17.799559,17.168514,16.13278,15.570327,16.510035,17.243965,17.902447,17.826996,17.487467,18.4649,19.891607,19.1954,17.95046,17.71039,20.004784,23.653864,32.567364,32.67711,24.555847,23.406935,15.693792,10.597425,7.2158523,4.698535,2.2566686,1.1111864,0.980862,0.96714365,0.84367853,1.0528834,1.3581166,1.4164196,1.6736387,2.2566686,2.976882,3.4878905,4.0091877,4.5339146,5.1821065,6.193835,8.025234,9.280463,10.299051,11.375941,12.758065,13.903547,15.820687,17.339994,18.406595,20.066517,21.712719,19.644676,18.516342,19.579515,20.6907,21.668133,22.95423,24.089422,25.752771,29.76882,30.880005,25.3618,20.310017,18.221397,17.014183,13.3033695,13.673765,12.4974165,8.251588,3.5393343,1.5261664,0.78537554,0.58988905,0.4938606,0.33609957,0.7613684,0.5212973,0.41840968,0.8128122,1.6187652,1.6427724,1.546744,1.8759843,2.4452958,2.335549,2.1743584,2.1640697,3.1415021,4.2698364,3.0351849,5.892031,8.090397,8.412778,7.2158523,6.4236174,5.693115,5.3878818,5.754848,7.582818,12.22305,10.878652,9.318189,10.573419,15.193072,21.208569,19.853882,14.369971,8.186425,3.9268777,3.4021509,2.2292318,1.1317638,0.47328308,0.25721905,0.12346515,0.037725464,0.30866286,0.6927767,0.85396725,0.36696586,0.19548649,0.106317215,0.06859175,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.072021335,0.030866288,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.034295876,0.06516216,0.09945804,0.1371835,0.15090185,0.30866286,0.4424168,0.5041494,0.5658819,0.9431366,1.0014396,0.85396725,0.7579388,1.097468,1.2689474,1.2106444,1.0460242,0.91227025,0.9602845,1.5947582,2.3492675,3.3129816,4.2389703,4.530485,7.0958166,7.764586,7.939495,8.39563,9.263316,10.556271,11.592006,12.545431,13.529722,14.603184,14.750656,13.457702,12.939834,13.773223,14.908417,16.324837,16.513464,16.746675,17.532051,18.629519,18.44775,18.45804,19.099373,19.744135,18.708399,18.53692,17.96418,17.4566,17.487467,18.523201,19.147387,19.713268,20.399187,20.724997,19.576086,18.722118,18.574646,18.132229,17.38115,17.271402,17.96761,18.893597,19.613811,19.87446,19.60695,20.207129,20.62211,21.578964,22.61127,22.048819,22.378057,22.570116,21.849901,21.067955,22.703869,24.401514,25.26577,25.814505,25.368658,22.048819,22.683292,23.68473,24.264332,24.19917,23.818485,23.002243,22.834194,22.552967,21.674994,20.004784,18.025911,18.217968,17.243965,16.355703,21.407484,12.617453,6.1561093,2.719663,2.3664153,4.5030484,6.478491,17.494326,24.250612,23.94195,24.247183,21.7916,19.137098,25.396095,40.211914,53.78622,54.729355,60.741425,78.37979,102.1777,114.67512,82.29638,71.513756,73.50635,76.109406,63.780037,54.10174,46.23427,40.112453,36.432507,36.652,28.071173,17.86815,11.290202,9.760606,10.8958,7.390761,6.351596,5.967482,5.9640527,7.599966,8.210432,7.630832,7.507367,8.364764,9.595985,10.4533825,10.573419,10.64201,11.149589,12.421966,12.555719,13.512574,14.342535,14.87755,15.731518,17.758404,17.909306,18.574646,19.829874,19.438902,18.574646,19.006773,19.555508,19.932762,20.735287,20.20027,20.220848,19.62753,18.516342,18.235117,18.917604,18.996485,19.143957,19.682402,20.598103,20.526081,19.473198,17.415445,15.395418,15.518884,16.969599,17.545769,17.171944,16.736387,18.067066,19.102802,19.46291,19.651537,19.46634,17.991615,17.062197,16.016174,14.747226,13.279363,11.763485,10.299051,10.748327,11.993267,13.262215,14.1299,15.374841,17.936743,19.414894,18.883308,16.907866,15.3817,15.649208,16.21852,16.434584,16.492886,16.95931,17.03819,16.715809,16.523752,17.562918,17.21996,16.722668,15.806969,14.044161,10.834066,11.96926,12.747777,12.655178,11.691463,10.360784,10.593996,11.317638,11.739478,11.787492,12.130451,12.449403,12.106443,11.447963,10.621432,9.582268,10.096705,10.580277,11.410237,12.586586,13.732068,12.072148,11.338216,11.331357,11.592006,11.399949,11.067279,10.271614,9.599416,9.283894,9.184435,9.932085,9.760606,9.942374,10.518545,10.299051,9.873782,9.609704,9.506817,9.469091,9.321619,8.796892,8.803751,8.711152,8.268735,7.582818,8.279024,8.536243,8.766026,9.259886,10.161868,9.403929,8.759167,8.405919,8.4264965,8.803751,9.671436,9.657719,9.513676,9.637141,10.100135,0.39440256,0.42869842,0.48014224,0.50757897,0.5007198,0.45956472,0.47671264,0.45956472,0.4355576,0.45613512,0.607037,0.64133286,0.64476246,0.59674823,0.548734,0.6036074,0.59331864,0.5521636,0.5521636,0.5796003,0.53844523,0.5590228,0.53158605,0.5178677,0.53844523,0.58302987,0.64476246,0.6207553,0.5727411,0.52815646,0.4698535,0.52815646,0.48700142,0.45956472,0.48014224,0.5144381,0.5212973,0.61046654,0.66533995,0.64819205,0.6001778,0.8162418,0.84367853,1.0288762,1.3786942,1.5364552,1.611906,1.7079345,1.8588364,2.0817597,2.3732746,2.935727,4.190956,4.887162,5.0277753,5.871454,6.1458206,8.052671,10.556271,11.499407,7.6205435,5.892031,5.446185,4.479041,2.6887965,1.2655178,0.4081209,0.106317215,0.17147937,0.31895164,0.15433143,0.08916927,0.3806842,1.1454822,1.8656956,1.4129901,0.8162418,0.34638834,0.12346515,0.11317638,0.12346515,0.19891608,0.15776102,0.16119061,0.216064,0.16804978,0.07888051,0.13032432,0.2777966,0.33609957,0.01371835,0.17147937,0.26064864,0.216064,0.09259886,0.0548734,0.07545093,0.07888051,0.058302987,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.010288762,0.030866288,0.044584636,0.01371835,0.06516216,0.05144381,0.037725464,0.106317215,0.31895164,0.2194936,0.11317638,0.14404267,0.3841138,0.823101,0.9568549,0.9602845,0.980862,1.0940384,1.313532,0.823101,0.5555932,0.5727411,0.88826317,1.4472859,1.430138,1.138623,0.85396725,0.65848076,0.4424168,0.26064864,0.4046913,0.3841138,0.22978236,0.51100856,0.4664239,0.5007198,0.4938606,0.5007198,0.7305021,0.7373613,0.71678376,0.7579388,0.9259886,1.2689474,0.90541106,0.89855194,1.0700313,1.1146159,0.5796003,0.96714365,0.91912943,0.91227025,0.9568549,0.6036074,0.58645946,0.52815646,0.5624523,0.65505123,0.6241849,0.5590228,0.5727411,0.6036074,0.65162164,0.77165717,0.52472687,0.6241849,0.6379033,0.5212973,0.61389613,0.5693115,0.58645946,0.66533995,0.77508676,0.83681935,0.77851635,0.83681935,0.7888051,0.71678376,1.0082988,0.548734,0.48357183,0.5453044,0.6173257,0.7339317,0.66876954,0.72707254,0.90541106,1.1763484,1.4815818,1.6427724,1.5741806,1.4953002,1.4850113,1.4918705,1.6599203,1.961724,2.0817597,1.978872,1.8691251,2.0577524,2.393852,2.4795918,2.4384367,2.9048605,3.234101,3.690236,4.1017866,4.383013,4.5201964,5.2164025,5.302142,5.1169443,4.945465,5.0106273,5.2506986,5.627953,5.562791,5.3913116,6.3481665,7.1198235,6.108095,4.911169,4.5270553,5.353586,4.6676683,5.3432975,6.1286726,6.6739774,7.5450926,8.179566,8.450503,8.937505,9.547972,9.499957,9.606275,9.938945,10.323058,10.569988,10.484249,10.535692,10.717461,11.125582,11.917816,13.293081,14.273943,14.987297,15.676644,16.341984,16.722668,16.37628,16.12249,16.005884,16.13278,16.654078,16.071047,15.347404,14.983868,15.014734,14.990726,14.904987,15.083325,15.62863,16.259674,16.300829,16.80155,16.571766,16.256245,16.156786,16.228807,16.20137,17.189093,17.861292,18.091074,18.938183,20.20027,20.759293,18.488907,16.328266,22.275171,20.03565,25.807646,27.84825,23.554407,19.476627,12.144169,10.882081,10.569988,8.4093485,3.9543142,1.8108221,1.0357354,0.980862,1.0597426,0.7613684,1.0734608,1.3546871,1.7730967,2.3595562,3.0111778,3.6799474,4.262977,4.482471,4.4275975,4.57164,6.012067,7.599966,9.273604,10.799771,11.766914,13.101024,14.55174,16.03675,17.62808,19.552078,19.003344,18.231688,18.694681,19.857311,19.202261,22.384918,23.396646,24.645016,27.378397,31.685959,26.870817,22.220297,17.806417,14.30481,12.9981365,13.505715,11.183885,8.2310095,5.422178,2.0886188,1.2243627,0.8025235,0.64476246,0.5761707,0.39783216,0.47328308,0.45270553,0.6927767,1.1626302,1.4232788,2.1297739,2.411,2.644212,2.867135,2.784825,3.340418,4.1155047,5.164959,5.970912,5.442755,6.111525,5.909179,5.90575,6.759717,8.718011,8.251588,8.700864,10.508256,13.817808,18.495766,15.738377,15.62863,15.577187,15.501736,17.826996,17.422304,13.090735,8.06296,4.8905916,5.429037,3.690236,1.762808,0.78537554,0.82996017,0.89169276,0.5041494,0.45613512,0.94999576,1.6153357,1.5364552,0.8093826,0.31209245,0.07888051,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.020577524,0.020577524,0.024007112,0.041155048,0.041155048,0.08916927,0.25721905,0.42183927,0.26064864,0.490431,0.548734,0.5453044,0.5555932,0.6344737,1.1283343,1.1729189,1.0906088,1.1008976,1.3169615,2.0474637,2.585909,3.2375305,4.064061,4.8734436,6.23499,6.8969,7.082098,7.0203657,6.931196,8.14527,9.170717,10.213311,11.345076,12.5145645,12.123591,11.701753,12.151029,13.505715,14.946142,16.420864,17.384579,17.463459,17.28512,18.471758,18.945042,19.123379,19.027351,18.663815,18.0362,17.775553,17.672665,17.559488,17.497755,17.744686,18.502625,19.353163,19.826445,19.871029,19.857311,18.427174,17.672665,17.04162,16.681513,17.432592,18.20425,18.54035,19.092514,19.984205,20.827885,21.397196,22.998814,24.473536,25.60187,27.1006,27.735073,27.731644,27.230925,26.723345,27.049156,25.60187,24.727325,24.696459,24.569565,22.196291,21.647556,22.508383,23.28347,23.674442,24.576424,24.871368,24.579853,23.653864,22.131128,20.124819,19.428614,19.12681,19.174824,20.015072,22.580404,14.514014,7.346176,3.649081,3.1483612,2.7059445,2.2909644,4.972902,8.663138,11.8115,13.395968,11.115293,10.39508,13.176475,19.504065,27.532728,32.50563,37.24875,43.14764,50.305187,57.52104,50.38064,47.931915,49.516384,50.943092,44.48518,34.793163,29.034887,27.230925,27.663052,26.836521,24.243753,17.87158,12.13731,9.160428,8.783174,6.989499,5.9812007,5.7822843,6.574519,8.711152,10.501397,11.190743,11.454823,11.677745,11.952112,10.912948,10.854645,11.286773,11.862943,12.360233,12.6586075,12.833516,13.341095,13.9138365,13.54687,14.754086,14.874121,15.196502,16.108772,17.096493,17.549198,18.632948,18.941612,18.677534,19.637817,20.018501,20.385468,19.833303,18.530062,17.720678,19.167965,19.480057,19.79901,20.440342,20.917053,21.03023,20.258574,18.663815,16.811838,15.762384,15.409137,17.017612,18.842154,19.761284,19.274282,19.346302,19.281141,19.147387,18.643238,17.099922,17.566347,17.302269,16.19794,14.599753,13.289652,11.561139,11.688034,12.8197975,13.694343,12.617453,13.138749,14.973578,17.014183,18.303709,18.005335,16.743246,16.842705,17.576635,18.324286,18.581505,18.019053,17.096493,16.359133,16.184223,16.780972,16.811838,17.007324,16.62664,15.3302555,13.166186,12.346515,12.4974165,12.079007,10.840926,9.81205,10.443094,11.667457,12.751206,13.317088,13.327377,12.843805,12.651748,12.188754,11.502836,11.255906,11.406808,11.80121,12.295071,12.878101,13.684054,11.965831,10.899229,10.81006,11.228469,10.899229,10.88894,10.563129,9.935514,9.273604,9.088407,9.668007,9.89436,10.268185,10.604284,10.041832,9.97667,9.836057,9.671436,9.482809,9.187865,8.937505,9.098696,8.999237,8.488229,7.963502,8.56025,9.208443,9.630281,9.904649,10.456812,9.386781,8.697433,8.618553,8.903209,8.851766,9.095266,9.146709,9.366203,9.853205,10.443094,0.33266997,0.37725464,0.41498008,0.4698535,0.5178677,0.48357183,0.5212973,0.53844523,0.58988905,0.6893471,0.82996017,0.67219913,0.6893471,0.67219913,0.58645946,0.5590228,0.59331864,0.548734,0.53844523,0.5521636,0.45956472,0.48357183,0.5212973,0.5658819,0.6001778,0.59331864,0.607037,0.5658819,0.52815646,0.51100856,0.48700142,0.4938606,0.48014224,0.4664239,0.4698535,0.51100856,0.490431,0.53158605,0.59331864,0.6310441,0.59674823,0.84024894,0.94656616,1.1729189,1.4953002,1.6221949,1.7525192,1.7902447,1.9480057,2.287535,2.7128036,3.5393343,4.7499785,5.312431,5.4496145,6.6225333,8.038953,11.430815,14.754086,14.925565,7.8331776,4.6916757,4.166949,3.8788633,2.843128,1.471293,0.764798,0.42183927,0.31895164,0.3841138,0.5761707,0.7510797,0.6036074,0.9431366,1.5364552,1.1214751,0.8505377,0.6962063,0.44927597,0.15090185,0.07888051,0.116605975,0.22292319,0.33266997,0.40126175,0.4389872,0.4664239,0.70649505,0.94999576,0.9294182,0.29837412,0.28122616,0.28465575,0.26407823,0.19548649,0.05144381,0.06859175,0.06859175,0.048014224,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.06859175,0.32924038,0.6207553,0.29837412,0.17833854,0.08916927,0.037725464,0.061732575,0.22978236,0.14747226,0.19891608,0.39097297,0.67219913,0.96371406,1.3821237,1.3375391,1.1797781,1.0700313,0.97400284,0.61389613,0.7442205,0.9877212,1.2586586,1.7559488,1.4918705,1.0837497,0.7990939,0.66533995,0.42869842,0.35324752,0.47671264,0.5658819,0.5555932,0.5658819,0.4355576,0.44927597,0.48700142,0.52815646,0.64476246,0.66876954,0.71678376,0.805953,0.9259886,1.039165,0.8471081,0.91227025,0.9602845,0.8505377,0.5727411,0.881404,0.823101,0.7305021,0.7373613,0.77165717,0.52472687,0.51100856,0.65162164,0.764798,0.59674823,0.50757897,0.5555932,0.58645946,0.61046654,0.8093826,0.5796003,0.6241849,0.6276145,0.5727411,0.72021335,0.607037,0.6344737,0.64476246,0.6344737,0.7339317,0.6756287,0.72021335,0.77508676,0.8471081,1.0082988,0.58302987,0.5624523,0.6379033,0.6824879,0.7407909,0.6756287,0.7373613,0.8676856,1.0425946,1.2620882,1.5158776,1.4850113,1.4850113,1.546744,1.3889829,1.7353712,1.9823016,2.16064,2.2738166,2.311542,2.510458,2.301253,2.1915064,2.3595562,2.6476414,2.9151495,3.3472774,3.7451096,4.0434837,4.3007026,5.0826488,5.171818,5.038064,4.9351764,4.9008803,4.547633,4.695105,5.0106273,5.6485305,7.281014,8.694004,7.0443726,4.8288593,3.6696587,4.338428,4.1189346,4.979761,5.8474464,6.4887795,7.531374,8.06296,8.501947,9.026674,9.589127,9.908078,9.904649,9.914937,10.034973,10.1481495,9.908078,9.932085,10.155008,10.662587,11.530273,12.8197975,13.862392,14.637479,15.169065,15.549749,15.923574,15.88242,15.656067,15.415996,15.29939,15.405707,15.121051,14.678635,14.555169,14.685493,14.479718,14.318527,14.479718,14.805529,15.114192,15.227368,15.642348,15.844694,16.149927,16.561478,16.780972,16.80498,17.319416,17.785841,18.221397,19.21255,20.207129,20.519222,18.574646,17.21996,23.722456,20.697561,22.484375,24.843931,23.821915,15.748666,10.645439,12.600305,13.828096,10.991828,5.192395,2.3321195,1.0871792,0.8711152,1.0323058,0.823101,0.96714365,1.196926,1.5810398,2.1194851,2.7573884,3.1483612,3.4638834,3.6113555,3.6936657,4.0091877,4.897451,6.574519,8.224151,9.496528,10.494537,12.408247,13.272504,14.411126,16.115631,17.63151,16.78783,17.024471,17.62122,18.344864,19.442331,22.100262,23.132568,26.208908,30.50275,30.68109,24.94682,20.663265,16.095055,12.041282,11.845795,11.982979,9.277034,5.8200097,3.0523329,1.7593783,1.3478279,1.0117283,0.7407909,0.53844523,0.42183927,0.47328308,0.53158605,0.7476501,1.0940384,1.3649758,2.1194851,2.8259802,3.6044965,4.4413157,5.195825,5.6073756,5.7994323,6.2830043,7.0032177,7.3530354,6.8145905,5.5902276,5.7274113,7.658269,10.189304,9.743458,10.175586,11.982979,14.88098,17.802988,16.352274,16.091625,15.223939,13.989287,14.675205,13.862392,10.593996,6.8283086,4.3658648,4.863155,3.0660512,1.6084765,1.138623,1.3821237,1.1489118,0.6379033,0.44927597,0.7133542,1.3272504,1.9239986,1.6256244,0.7442205,0.15090185,0.0548734,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.010288762,0.0034295875,0.006859175,0.034295876,0.034295876,0.14061308,0.22635277,0.26064864,0.31895164,0.28122616,0.32924038,0.36353627,0.34981793,0.31895164,0.7682276,0.7990939,0.8093826,0.96714365,1.2312219,2.2292318,2.7333813,3.1346428,3.7794054,4.9694724,5.48734,6.0497923,6.4887795,6.701414,6.660259,7.2021337,8.008087,9.22216,10.587136,11.417097,10.9369545,11.231899,12.017275,13.121602,14.496866,16.108772,17.343424,17.63494,17.69667,19.514353,20.045938,19.757853,18.828436,17.761833,17.38115,16.976458,16.859852,17.034761,17.278261,17.134218,17.878439,18.523201,18.653526,18.54378,19.140528,18.231688,17.55263,17.315987,17.55263,18.12194,18.636377,18.866161,19.390888,20.217419,20.78673,21.500084,23.20802,25.087433,26.953129,29.254381,29.326403,29.34012,30.067194,30.51647,27.909983,24.957108,23.86307,23.821915,23.835632,22.727877,21.421204,21.548098,22.347193,23.266321,23.959099,25.406384,25.903673,25.27949,23.801336,22.19972,21.630407,21.551527,21.678423,21.421204,19.898466,12.648318,7.6651278,4.7534084,3.3678548,2.5961976,2.2498093,1.879414,2.9254382,5.2575574,7.1369715,7.3358874,8.40249,10.0041065,12.298501,15.96816,19.929333,22.967947,25.042849,26.548437,28.3524,28.071173,28.455288,29.247522,28.92857,24.734184,17.556059,17.573206,18.12194,18.108221,22.03167,19.994495,15.37827,10.72775,7.606825,6.5710897,6.3447366,5.4599032,5.0174866,5.9880595,9.1981535,11.4376745,12.044711,11.609154,11.135871,12.020704,12.542002,12.977559,12.737488,12.103014,12.178465,12.500846,12.253916,12.596875,13.46799,13.594885,13.9138365,14.13333,14.634049,15.590904,16.95931,18.070496,19.28457,19.744135,19.305147,18.547209,19.078794,19.377169,19.095943,18.389448,17.895588,18.506054,18.752985,19.435472,20.327166,20.179693,19.630959,19.21255,18.53692,17.62122,16.88386,15.741806,17.240536,19.315437,20.488356,19.871029,19.853882,20.165974,19.836735,18.71183,17.442883,18.656956,18.499195,17.29541,15.618341,14.30481,13.169616,13.114742,13.406258,13.334236,12.21962,12.061859,12.991278,14.740367,16.592344,17.364002,17.178804,17.53891,18.183672,18.917604,19.6241,18.279701,17.062197,16.431154,16.276823,15.909856,15.745236,15.587475,15.37827,14.634049,12.428825,11.218181,11.399949,10.912948,9.668007,9.571979,10.6145735,11.849225,12.80265,13.101024,12.47341,12.0309925,12.085866,11.705182,11.046701,11.372512,11.197603,11.341646,11.8115,12.445972,12.895248,11.578287,10.88551,10.333347,9.949233,10.288762,10.830637,11.094715,10.998687,10.508256,9.602845,9.736599,9.918367,10.30591,10.683165,10.491108,10.089847,9.89436,9.6817255,9.270175,8.522525,8.580828,9.095266,9.39707,9.249598,8.872343,9.057541,9.585697,10.158438,10.604284,10.88551,9.561689,8.704293,8.652849,9.256456,9.880642,9.321619,9.31133,9.671436,10.14472,10.408798,0.40126175,0.47671264,0.44927597,0.45613512,0.5041494,0.45270553,0.4698535,0.52472687,0.61046654,0.70649505,0.7922347,0.6173257,0.6173257,0.6036074,0.52815646,0.47328308,0.5521636,0.53158605,0.5178677,0.5212973,0.45956472,0.490431,0.5453044,0.59331864,0.61046654,0.58645946,0.61389613,0.5761707,0.548734,0.5521636,0.5178677,0.45956472,0.47671264,0.48357183,0.47328308,0.4938606,0.490431,0.50757897,0.5761707,0.65162164,0.61389613,0.83681935,1.039165,1.3169615,1.5673214,1.5090185,1.7525192,1.7730967,1.9480057,2.411,3.0557625,3.9543142,5.1238036,5.994919,6.601956,7.5690994,9.856634,14.997586,18.814716,17.62808,8.261876,4.5784993,3.223812,2.6956558,2.1983654,1.6221949,1.0254467,0.6859175,0.5796003,0.67219913,0.91227025,1.2517995,0.7476501,0.6173257,0.94656616,0.6962063,0.6310441,0.7476501,0.61046654,0.2469303,0.15090185,0.12003556,0.25721905,0.39440256,0.45956472,0.45613512,0.48014224,0.82996017,1.3101025,1.4953002,0.7613684,0.432128,0.28465575,0.26407823,0.26750782,0.12003556,0.072021335,0.048014224,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.09945804,0.22292319,0.5761707,0.97057325,0.84367853,0.52472687,0.26407823,0.09602845,0.048014224,0.13032432,0.11317638,0.37725464,0.65848076,0.85739684,1.0185875,1.4164196,1.646202,1.471293,0.9842916,0.6001778,0.78194594,0.97057325,1.1283343,1.2655178,1.4507155,1.2175035,0.91227025,0.7407909,0.67219913,0.44584638,0.41840968,0.53501564,0.61389613,0.6036074,0.5658819,0.47328308,0.50757897,0.53844523,0.52472687,0.5041494,0.5521636,0.70306545,0.7682276,0.7442205,0.8162418,0.7922347,0.8711152,0.8505377,0.7407909,0.77508676,0.823101,0.7682276,0.7373613,0.77851635,0.8265306,0.5624523,0.58645946,0.6962063,0.77165717,0.7476501,0.7133542,0.6893471,0.6379033,0.59674823,0.6927767,0.5555932,0.607037,0.70306545,0.77165717,0.83681935,0.66876954,0.6824879,0.66191036,0.58645946,0.6173257,0.61046654,0.66191036,0.7373613,0.7922347,0.7613684,0.6824879,0.7305021,0.7442205,0.70649505,0.75450927,0.7133542,0.7442205,0.823101,0.89855194,0.89855194,1.1454822,1.1180456,1.2003556,1.4027013,1.371835,1.9068506,2.3321195,2.5961976,2.750529,2.935727,3.07634,2.5927682,2.3561265,2.486451,2.369845,2.668219,3.0523329,3.5393343,3.99204,4.1155047,4.756838,4.7671266,4.7088237,4.746549,4.6436615,4.184097,4.372724,4.9591837,5.953764,7.6033955,9.304471,6.944915,4.2698364,3.2375305,4.016047,4.0880685,4.955754,5.720552,6.2864337,7.349606,7.747438,8.364764,8.824328,9.156999,9.798331,10.179015,10.100135,10.14129,10.377932,10.374502,10.329918,10.532263,11.080997,11.962401,13.029003,13.762935,14.263655,14.500296,14.586036,14.802099,14.754086,14.678635,14.599753,14.441993,14.003006,14.020154,13.828096,13.759505,13.7526455,13.334236,13.227919,13.536582,13.80409,13.941273,14.225929,14.345964,14.726648,15.261664,15.851553,16.396858,17.014183,17.247395,17.758404,18.588364,19.157675,19.52807,19.473198,18.588364,18.605513,23.403505,21.719578,24.428951,25.876238,22.546108,13.080446,10.521975,14.356253,16.03675,12.5145645,6.245279,2.8499873,1.2277923,0.78537554,0.8848336,0.8779744,0.90198153,0.97400284,1.2003556,1.611906,2.1332035,2.3321195,2.5721905,2.8705647,3.2718265,3.875434,4.173808,5.5319247,6.8900414,7.9463544,9.139851,11.039842,11.499407,12.531713,14.239647,14.839825,14.846684,16.225378,16.993607,17.54234,20.639257,21.819035,23.122278,27.083452,31.126936,27.594461,21.94593,19.181683,16.005884,12.401388,11.616013,10.117283,7.4353456,4.3349986,2.136633,2.7059445,2.3732746,3.0146074,2.4795918,0.922559,0.8128122,0.9842916,1.1797781,1.4507155,1.8245405,2.3149714,2.942586,4.0023284,4.9591837,5.7411294,6.759717,6.944915,6.276145,6.276145,7.1095347,7.5725293,7.531374,6.444195,6.509357,8.179566,10.189304,9.952662,10.281903,11.201033,12.734058,14.88098,15.357693,14.856973,14.05102,13.306799,12.703192,10.799771,8.172707,5.689686,4.190956,4.479041,3.2032347,2.6407824,2.2669573,1.9239986,1.8313997,1.1832076,1.0460242,1.1283343,1.5433143,2.8328393,2.1812177,0.9294182,0.14747226,0.058302987,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.01371835,0.044584636,0.041155048,0.17833854,0.21263443,0.15776102,0.29494452,0.15776102,0.18519773,0.20920484,0.17833854,0.14747226,0.41840968,0.47328308,0.59674823,0.864256,1.1077567,2.194936,2.7985435,3.0900583,3.4947495,4.6882463,4.7842746,5.3844523,6.121814,6.660259,6.708273,6.842027,7.6033955,8.999237,10.491108,10.995257,11.067279,11.917816,12.80265,13.543441,14.531162,15.638919,16.636929,17.442883,18.440891,20.478067,20.224277,19.164536,17.717249,16.499744,16.352274,16.434584,16.513464,16.70552,16.901007,16.746675,17.233677,17.62465,17.778982,17.833855,18.20768,18.176813,18.063637,18.533491,19.312008,19.157675,19.294859,19.6241,20.141968,20.807306,21.578964,22.563255,24.209457,26.095732,28.074602,30.296976,30.59192,31.17152,31.878016,31.240112,26.469557,24.562706,24.120289,23.86307,23.345201,22.957659,21.62012,20.934202,21.328604,22.36434,22.721018,24.281479,25.416672,25.52985,24.634727,23.328054,22.817045,23.578413,23.550978,20.906765,14.05102,9.160428,6.186976,4.2526884,3.0111778,2.633923,2.5173173,1.8176813,1.9548649,3.3678548,5.5079174,6.7357097,8.340756,10.0041065,11.640019,13.402828,15.086755,16.681513,17.53891,17.29198,15.834405,17.065628,18.588364,19.342873,18.653526,16.225378,13.937843,16.002455,16.739817,16.143068,19.857311,15.6252,11.55428,8.443645,6.461343,5.130663,5.360445,4.931747,4.791134,5.744559,8.440215,10.902658,11.444533,11.012405,10.803201,12.271064,13.80066,14.363112,14.054449,13.38225,13.258785,13.166186,12.830087,12.782072,13.087306,13.368532,13.63261,14.105893,14.688923,15.560039,17.165085,18.725548,20.03222,20.539799,19.987637,18.403166,18.742695,18.893597,18.728977,18.440891,18.516342,18.451181,18.499195,18.931322,19.500635,19.442331,18.54035,18.097933,17.720678,17.312557,17.079346,16.503176,17.79613,19.277712,20.12139,20.334024,20.697561,21.074816,20.556948,19.281141,18.434032,19.829874,19.504065,17.95389,15.920145,14.359683,14.023583,14.068168,13.999576,13.522863,12.548861,11.499407,11.770344,12.88496,14.421415,16.009314,16.575195,17.240536,18.008764,18.752985,19.222837,18.03963,17.264544,17.12393,17.117071,16.005884,15.391989,14.3974085,13.958421,13.512574,10.988399,10.388221,10.7586155,10.247607,9.102125,9.647429,11.249047,12.418536,13.022143,12.826657,11.509696,11.451392,11.492548,11.218181,10.782623,10.88894,10.676306,10.587136,10.988399,11.760056,12.271064,11.297061,10.80663,9.97324,9.14328,9.836057,10.64201,11.317638,11.633161,11.379372,10.374502,10.076128,10.079557,10.39165,10.844356,11.070708,10.155008,9.860064,9.613133,9.081548,8.193284,8.354475,9.002667,9.613133,9.89093,9.764035,9.595985,9.72288,10.216741,10.88551,11.2593355,9.650859,8.4264965,8.327039,9.301042,10.497967,9.654288,9.554831,9.815479,10.14129,10.30591,0.51100856,0.59674823,0.5041494,0.44927597,0.4664239,0.40126175,0.37039545,0.44584638,0.5041494,0.5212973,0.5521636,0.5178677,0.48700142,0.44927597,0.41840968,0.4389872,0.5144381,0.53158605,0.53501564,0.5453044,0.5624523,0.5761707,0.5727411,0.5590228,0.5590228,0.6344737,0.7133542,0.6824879,0.6379033,0.59674823,0.51100856,0.4389872,0.4629943,0.48014224,0.4629943,0.4664239,0.5212973,0.5555932,0.61389613,0.6790583,0.6790583,0.8745448,1.1214751,1.4198492,1.605047,1.3443983,1.5913286,1.7079345,1.9823016,2.5207467,3.2581081,4.029765,5.212973,6.677407,8.021805,8.594546,10.786053,16.921585,20.666695,18.245405,8.443645,4.2286816,2.3081124,1.5090185,1.2380811,1.4815818,0.9911508,0.7888051,0.71678376,0.71678376,0.83338976,1.2517995,0.77165717,0.4389872,0.52472687,0.51100856,0.36696586,0.4424168,0.4115505,0.26407823,0.30866286,0.26407823,0.26407823,0.29837412,0.31209245,0.18862732,0.09602845,0.40126175,1.039165,1.5638919,1.138623,0.6207553,0.37039545,0.30866286,0.31895164,0.2469303,0.12346515,0.072021335,0.05144381,0.030866288,0.010288762,0.0034295875,0.0,0.0034295875,0.024007112,0.08916927,0.116605975,0.32581082,0.53844523,0.7613684,1.1934965,0.8848336,0.4629943,0.16119061,0.058302987,0.072021335,0.16462019,0.5521636,0.823101,0.91912943,1.1489118,1.2175035,1.7456601,1.6770682,0.97400284,0.58988905,1.2175035,1.0734608,0.96714365,1.0528834,0.84367853,0.89169276,0.71678376,0.6379033,0.6859175,0.6241849,0.5555932,0.64133286,0.5624523,0.39783216,0.65162164,0.58302987,0.65848076,0.6379033,0.5144381,0.5144381,0.6001778,0.72021335,0.6893471,0.59331864,0.78194594,0.7579388,0.7442205,0.7579388,0.805953,0.91227025,0.82996017,0.8505377,1.0048691,1.1214751,0.82996017,0.7099246,0.70306545,0.6927767,0.7373613,1.0597426,1.0734608,0.9328478,0.77165717,0.65162164,0.53844523,0.4972902,0.66533995,0.85739684,0.9259886,0.7476501,0.6962063,0.71678376,0.72364295,0.70649505,0.72364295,0.6927767,0.7442205,0.77165717,0.7099246,0.5178677,0.84024894,0.9431366,0.85396725,0.7133542,0.7888051,0.764798,0.7476501,0.7888051,0.8025235,0.58988905,0.7339317,0.6893471,0.864256,1.2792361,1.5433143,2.1915064,2.8499873,3.2443898,3.3712845,3.5221863,3.4981792,3.117495,2.8088322,2.603057,2.136633,2.5138876,2.9391565,3.5221863,4.0503426,3.9851806,4.465323,4.40702,4.4104495,4.5853586,4.5442033,4.3795834,4.7842746,5.336438,5.967482,6.975781,8.131552,5.761707,3.7519686,3.5461934,4.166949,4.3281393,4.979761,5.579939,6.1149545,7.0786686,7.486789,8.217292,8.652849,8.848335,9.530824,10.319629,10.251037,10.371073,10.868362,11.080997,11.050131,11.341646,11.907528,12.668896,13.505715,13.708061,13.735497,13.677195,13.6086035,13.605173,13.430264,13.471419,13.612033,13.574307,12.895248,13.001566,12.785502,12.55229,12.346515,11.955542,11.989838,12.466551,12.833516,13.004995,13.368532,13.090735,13.310229,13.701202,14.191633,14.946142,16.20137,16.650646,17.689812,19.03078,18.694681,18.62266,18.739265,18.78042,19.390888,22.10712,20.392326,27.803665,28.757092,20.28258,12.037852,12.984418,16.37971,16.71238,12.610593,6.835168,3.2032347,1.3581166,0.7099246,0.70649505,0.8162418,0.823101,0.7442205,0.77851635,0.9911508,1.2929544,1.5433143,1.9068506,2.3801336,2.9631636,3.642222,3.590778,4.4859004,5.521636,6.5230756,7.905199,9.205012,9.647429,10.851214,12.432255,12.000127,13.46799,15.769243,17.333136,18.478617,21.404055,21.345753,24.806206,28.472435,28.921711,22.62156,16.602633,16.595774,16.167076,13.238208,10.072699,7.5210853,5.007198,3.0317552,2.5721905,5.099797,4.1463714,6.042933,5.5833683,2.5413244,1.6736387,1.8588364,2.352697,3.4810312,4.5819287,4.0229063,4.6848164,5.7891436,6.15268,5.8680243,6.276145,6.0703697,5.06893,5.0929375,6.159539,6.4990683,8.179566,8.008087,7.630832,7.936065,9.043822,9.314759,9.647429,9.863494,10.456812,12.590015,14.644339,14.441993,14.267084,14.212211,12.175035,9.0644,6.6705475,5.127233,4.5167665,4.8905916,4.9008803,4.8940215,3.9954693,2.6167753,2.452155,1.9891608,2.085189,2.0131679,2.0886188,3.666229,2.2395205,0.7990939,0.07545093,0.06516216,0.041155048,0.006859175,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.0274367,0.030866288,0.041155048,0.030866288,0.1097468,0.16804978,0.16462019,0.1097468,0.06516216,0.061732575,0.06859175,0.07545093,0.08916927,0.216064,0.32924038,0.5693115,0.91227025,1.1626302,2.0063086,2.644212,2.942586,3.1723683,4.029765,4.173808,5.096367,6.101236,6.715132,6.694555,6.7871537,7.6033955,8.999237,10.456812,11.118723,12.024134,13.258785,14.105893,14.507155,15.059319,15.536031,15.995596,17.12393,18.866161,20.430052,19.143957,17.53891,16.002455,15.0250225,15.196502,16.235666,16.955881,17.003895,16.63007,16.681513,16.715809,17.027903,17.63151,18.231688,18.224829,18.924463,19.263992,20.11453,21.050808,20.361462,20.28258,20.711279,21.236006,22.069395,24.051697,25.084003,26.737064,28.318104,29.583622,30.75997,31.83686,33.09209,32.766277,29.964306,24.645016,24.404943,24.127148,23.225166,22.131128,22.295748,21.77445,20.728426,20.515793,21.19828,21.558388,22.26831,23.35549,23.890507,23.571554,22.714157,22.44665,23.787619,23.629858,19.294859,8.543102,6.111525,4.201245,3.1552205,2.819121,2.534465,2.5756202,2.4247184,2.884283,4.32471,6.680836,7.3427467,8.330468,10.333347,13.022143,15.049029,15.762384,16.595774,16.859852,15.985307,13.519434,16.571766,18.183672,18.879879,18.986197,18.602083,20.570665,20.60839,21.187992,21.740154,18.684393,12.253916,8.158989,6.385892,5.9812007,5.0826488,4.3281393,4.530485,5.2438393,6.1629686,7.1061053,9.8429165,10.940384,11.492548,12.253916,13.656617,14.7026415,14.946142,15.285671,15.704081,15.258235,14.935853,14.7026415,14.13676,13.395968,13.190193,13.732068,14.267084,14.647768,15.3302555,17.38115,19.277712,20.632399,20.94449,20.265432,19.21255,19.315437,19.301718,19.003344,18.728977,19.260563,19.19197,18.87302,18.578075,18.61923,19.353163,18.732407,17.95389,17.178804,16.70895,16.990177,17.652086,18.749556,19.46291,19.826445,20.752434,21.825895,21.95279,21.421204,20.587814,19.87446,20.872469,20.29287,18.259123,15.584045,13.756075,13.7938,13.9138365,14.112752,14.030442,12.9707,11.05699,11.080997,11.677745,12.521424,14.335675,15.21022,16.242527,17.487467,18.434032,18.008764,17.590355,17.508043,17.857862,18.087645,16.969599,15.700651,14.177915,13.529722,13.111313,10.494537,10.535692,10.830637,10.295622,9.383351,10.117283,12.154458,13.203912,13.529722,13.090735,11.537132,11.63659,11.595435,11.55428,11.341646,10.4705305,10.357354,10.251037,10.467101,11.063849,11.852654,11.094715,10.508256,9.777754,9.177576,9.592556,10.30934,10.933525,11.170166,11.036412,10.864933,10.583707,10.422516,10.518545,10.851214,11.2421875,10.240748,9.815479,9.513676,9.091836,8.484799,8.546532,8.98209,9.56512,10.055551,10.209882,9.925226,9.630281,9.870353,10.6145735,11.245617,9.465661,8.080108,8.018375,9.136421,10.230459,9.513676,9.702303,9.89436,9.873782,10.106995,0.48700142,0.5727411,0.5693115,0.58645946,0.6344737,0.61046654,0.548734,0.6173257,0.6241849,0.53844523,0.5041494,0.48014224,0.4629943,0.44584638,0.4389872,0.48700142,0.52472687,0.58988905,0.6310441,0.64819205,0.67219913,0.59674823,0.5144381,0.51100856,0.61046654,0.7922347,0.7442205,0.7407909,0.65505123,0.51100856,0.48700142,0.41498008,0.45956472,0.490431,0.48014224,0.5041494,0.5761707,0.58645946,0.61046654,0.6893471,0.823101,1.0323058,1.2655178,1.4610043,1.529596,1.3581166,1.5055889,1.7593783,2.2738166,2.942586,3.4192986,4.197815,5.0277753,6.625963,8.594546,9.400499,10.741467,15.498305,17.62465,14.390549,6.392751,2.74367,1.4541451,1.1008976,0.96714365,1.0528834,0.85739684,0.9911508,0.91912943,0.6241849,0.6241849,1.0151579,0.70306545,0.31209245,0.18176813,0.36696586,0.2194936,0.12689474,0.09602845,0.16119061,0.3806842,0.5521636,0.42869842,0.24007112,0.10288762,0.030866288,0.006859175,0.09945804,0.31895164,0.6379033,0.9911508,0.7476501,0.59674823,0.5041494,0.42869842,0.31895164,0.23664154,0.19548649,0.15776102,0.106317215,0.044584636,0.010288762,0.0,0.01371835,0.041155048,0.07545093,0.01371835,0.06516216,0.07545093,0.12003556,0.47328308,0.6310441,0.34295875,0.1097468,0.08573969,0.061732575,0.13375391,0.5453044,1.0357354,1.4541451,1.786815,1.2963841,1.2312219,1.0666018,0.7099246,0.5041494,1.3958421,1.2620882,1.2346514,1.371835,0.6241849,1.0528834,1.0048691,0.8196714,0.7339317,0.85396725,0.8676856,0.65162164,0.45956472,0.48014224,0.8093826,0.5658819,0.5761707,0.59674823,0.6241849,0.9294182,1.0151579,0.7888051,0.7613684,0.85396725,0.42869842,0.45270553,0.3566771,0.4115505,0.607037,0.65505123,0.77851635,0.83681935,1.0494537,1.2586586,0.91569984,0.90198153,0.7888051,0.7888051,1.0357354,1.5707511,1.3992717,1.2209331,0.9842916,0.7339317,0.6241849,0.7476501,1.2003556,1.2655178,0.85739684,0.5041494,0.7339317,0.922559,0.9328478,0.881404,1.1146159,0.8196714,0.89512235,1.1077567,1.1900668,0.823101,1.1043272,1.155771,0.9568549,0.6790583,0.71678376,0.64476246,0.75450927,0.8505377,0.8093826,0.5658819,0.69963586,0.7339317,1.1043272,1.728512,1.9823016,2.4830213,2.7573884,3.2066643,3.7176728,3.6319332,3.5221863,3.2649672,3.1792276,3.100347,2.3801336,2.942586,3.2478194,3.3815732,3.5221863,3.9371665,4.4859004,4.3487167,4.245829,4.4584637,4.835718,4.897451,5.086078,5.2506986,5.4736214,6.0737996,6.279575,4.839148,3.9851806,4.1772375,4.105216,4.7259717,4.928317,5.2472687,5.857735,6.591667,7.250148,8.220721,8.886061,9.115844,9.263316,9.836057,9.9801,10.30934,10.751757,10.542552,11.019264,11.46854,11.842365,12.250486,12.9707,13.1421795,13.183334,13.111313,13.118172,13.581166,13.543441,13.2862215,13.197053,13.227919,12.908967,12.456262,11.612583,10.878652,10.491108,10.405369,10.81006,11.578287,12.171606,12.442543,12.648318,12.185325,12.041282,12.243628,12.843805,13.9309845,15.138199,15.927004,17.21996,18.499195,17.7927,18.79414,19.53836,19.263992,19.154245,22.340332,15.234227,23.10856,26.915403,20.96164,12.895248,21.133118,20.52951,15.87213,10.47396,6.1629686,2.8945718,1.1592005,0.51100856,0.5212973,0.77851635,0.7305021,0.58988905,0.4972902,0.5144381,0.61046654,0.9774324,1.1420527,1.4644338,2.07833,2.884283,3.175798,4.1120753,4.863155,5.501058,6.989499,8.124693,9.030104,10.237319,11.180455,10.192734,13.440554,15.313108,17.981327,20.683842,19.744135,19.305147,30.0912,34.50851,27.258362,15.319967,9.55826,12.037852,12.9707,9.301042,4.698535,2.0028791,1.2175035,1.3443983,3.1449318,9.139851,5.892031,6.958633,7.8777623,6.468202,2.8088322,2.6133456,3.525616,7.3084507,10.63858,5.096367,6.169828,6.64997,5.885172,4.4550343,4.149801,2.4418662,2.177788,2.8259802,4.1326528,6.135532,9.0644,10.014396,9.235879,7.8846216,8.056101,8.923786,9.057541,10.333347,12.247057,11.917816,15.361122,15.717799,15.748666,15.566897,12.648318,8.683716,6.526505,4.90431,3.8137012,4.547633,6.9037595,6.4579134,5.23698,3.7691166,1.0837497,2.0474637,2.4624438,1.8828435,1.0528834,1.9068506,1.8108221,0.72364295,0.05144381,0.12346515,0.19891608,0.041155048,0.06516216,0.06516216,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.061732575,0.072021335,0.07545093,0.01371835,0.0274367,0.020577524,0.12346515,0.24350071,0.061732575,0.037725464,0.020577524,0.034295876,0.06516216,0.07545093,0.17490897,0.2709374,0.5453044,0.9911508,1.4198492,1.7250825,2.0097382,2.2978237,2.6407824,3.1277838,3.8479972,5.4187484,6.701414,7.3050213,7.599966,7.366754,7.8126,8.7283,10.041832,11.825217,12.936404,14.376831,14.853543,14.54831,15.121051,16.62321,16.640358,16.95931,17.988186,18.770132,17.669235,16.462019,15.100473,14.160767,14.832966,16.259674,17.851004,17.95046,16.911295,17.1205,16.657507,17.072487,18.187103,19.61724,20.752434,21.753874,21.434921,21.294308,21.630407,21.544668,21.78817,22.151705,22.841053,24.418663,27.786518,28.0163,29.274958,30.705097,31.294985,29.892284,30.207806,31.041197,31.435598,30.039757,25.084003,22.36434,19.685833,18.03277,18.084215,20.234566,21.332033,20.954779,20.62211,20.838173,21.1194,21.20514,21.592682,21.218857,20.567236,21.650986,21.236006,21.253153,20.7833,17.905876,9.688584,5.501058,5.223262,5.267846,4.307562,3.2821152,5.2335505,5.3570156,5.06893,5.3981705,6.9723516,8.913498,9.455373,11.194174,14.400838,17.014183,19.404606,20.361462,21.95279,23.163433,19.8676,23.321196,21.421204,19.346302,19.092514,19.469769,19.140528,19.847023,23.68473,26.448978,17.62465,11.825217,7.548522,5.360445,5.288424,6.790583,3.957744,4.3933015,5.5490727,6.334448,7.140401,10.278474,12.363663,13.656617,14.5585985,15.608052,16.842705,17.168514,17.473747,17.55263,16.112202,17.28512,17.103354,16.503176,16.105343,16.204802,15.498305,15.165636,15.278812,16.245956,18.79757,20.652975,21.53781,21.606401,21.04395,20.080235,20.056227,19.62753,19.133669,18.989626,19.69955,19.600092,18.506054,18.077356,18.842154,20.172834,19.939621,19.075365,18.1288,17.95389,19.69955,20.577524,20.659836,20.62211,20.728426,20.814167,23.060547,23.722456,23.825344,23.499533,21.973368,21.839613,20.917053,18.44432,15.21022,13.5503,12.902108,12.346515,12.531713,13.080446,12.603734,10.600855,10.679735,11.269625,11.684605,12.099585,13.749216,15.6252,17.504614,18.61923,17.655516,17.226818,17.075916,17.29884,17.655516,17.532051,15.189643,14.466,14.520873,14.171056,11.8869505,11.204462,10.858074,10.371073,10.079557,11.153018,12.80265,13.306799,13.4474125,13.416546,12.816368,12.205902,12.778643,13.13189,12.449403,10.484249,10.055551,10.377932,10.508256,10.374502,10.803201,10.535692,10.1652975,9.750318,9.421077,9.383351,10.041832,9.870353,9.441654,9.386781,10.374502,11.122152,10.820349,10.326488,10.155008,10.497967,10.569988,9.846346,9.403929,9.400499,9.095266,9.105555,9.174147,9.3764925,9.674867,9.918367,9.709162,9.266746,9.369633,10.014396,10.39165,8.913498,8.453933,8.656279,9.14328,9.5205345,8.436785,9.993818,10.690024,9.815479,9.458802,0.42869842,0.4938606,0.607037,0.64819205,0.59674823,0.52472687,0.51100856,0.53501564,0.5555932,0.548734,0.5041494,0.490431,0.45270553,0.44584638,0.4629943,0.4629943,0.4424168,0.5144381,0.5658819,0.5761707,0.61046654,0.7510797,0.77508676,0.7407909,0.6859175,0.6344737,0.5178677,0.48357183,0.45270553,0.39783216,0.35324752,0.33952916,0.42869842,0.52472687,0.5796003,0.61389613,0.66876954,0.6790583,0.7476501,0.881404,1.0082988,1.1866373,1.2826657,1.2209331,1.1454822,1.3958421,1.786815,2.0440342,2.411,2.8911421,3.2581081,4.4104495,5.960623,7.346176,8.673427,10.731179,10.216741,9.613133,9.2153015,7.963502,3.415869,1.7559488,1.1797781,1.0563129,1.0151579,0.9431366,0.7099246,0.7510797,0.78194594,0.72707254,0.7476501,0.8745448,0.5521636,0.2469303,0.22292319,0.5727411,0.37725464,0.274367,0.24007112,0.37039545,0.881404,1.0734608,0.77851635,0.42526886,0.18519773,0.006859175,0.0,0.020577524,0.08916927,0.22635277,0.45613512,0.5144381,0.5453044,0.6207553,0.65848076,0.42869842,0.30523327,0.19891608,0.14061308,0.1371835,0.14404267,0.048014224,0.017147938,0.010288762,0.006859175,0.01371835,0.0034295875,0.01371835,0.1097468,0.216064,0.13032432,0.16462019,0.14061308,0.106317215,0.08916927,0.13375391,0.30523327,0.29494452,1.0323058,2.0063086,1.2620882,0.52815646,0.41498008,0.58302987,0.7099246,0.5041494,1.0323058,1.3443983,1.1317638,0.71678376,1.0151579,1.4129901,2.486451,2.435007,1.3238207,1.0734608,0.91227025,1.3375391,1.313532,0.823101,0.8711152,0.86082643,0.6173257,0.61389613,0.7956643,0.5658819,0.7373613,0.70306545,0.7956643,0.922559,0.5727411,0.8505377,0.75450927,0.77508676,1.0151579,1.1797781,1.0288762,0.9534253,0.8505377,0.7922347,1.0254467,0.85739684,0.7407909,1.0768905,1.5433143,1.0837497,1.0014396,0.9431366,0.9842916,1.039165,0.8711152,1.0700313,0.9568549,0.7990939,0.6824879,0.5041494,0.6859175,0.8745448,0.9362774,0.9328478,1.1249046,0.764798,0.84367853,0.89512235,0.84367853,0.9945804,0.69963586,0.75450927,0.77851635,0.70306545,0.77851635,0.65505123,0.8711152,0.96714365,0.86082643,0.8196714,0.77851635,0.8196714,1.1763484,1.6804979,1.7525192,2.3801336,2.784825,3.2615378,3.7451096,3.8274195,3.3369887,3.2992632,3.1346428,2.7711067,2.6373527,2.9254382,3.309552,3.7313912,3.9851806,3.7176728,4.2286816,4.5201964,4.664239,4.671098,4.482471,4.6608095,4.746549,4.976331,5.4907694,6.355026,6.3653145,6.0052075,5.0312047,3.7931237,3.199805,4.5853586,4.846007,4.822,5.0174866,5.6039457,6.691125,7.425057,7.8949103,8.30646,8.98209,9.280463,9.709162,10.278474,10.72432,10.508256,10.583707,10.871792,11.4205265,12.027563,12.250486,12.010415,12.082437,12.308789,12.607163,12.9809885,12.878101,12.397959,12.048141,11.893809,11.5645685,11.105004,10.63858,10.072699,9.561689,9.517105,9.626852,10.357354,11.008976,11.266195,11.22161,11.283342,11.303921,11.698323,12.607163,13.858963,15.350834,15.923574,16.904436,18.434032,19.46291,19.459478,19.60695,19.593233,20.083664,22.741594,22.168854,27.340672,26.545008,18.663815,13.162757,17.556059,17.446312,14.04759,9.325048,5.994919,2.7916842,1.1694894,0.72364295,0.89855194,1.0117283,0.8745448,0.65848076,0.490431,0.41498008,0.41498008,0.6344737,0.90884066,1.1146159,1.3169615,1.7593783,2.0817597,2.6133456,3.3712845,4.3178506,5.377593,7.3701835,8.999237,10.357354,11.252477,11.180455,15.093615,16.657507,16.54433,15.364552,13.642899,16.942162,27.951138,30.718815,21.335464,7.922347,4.4275975,5.579939,5.8817425,3.758828,1.587899,0.6173257,0.41840968,0.71678376,1.7010754,4.012617,4.5853586,9.084977,11.859513,9.616563,1.4541451,1.7662375,2.5413244,3.7039545,4.262977,2.3252604,2.901431,3.5290456,4.033195,4.5201964,5.346727,3.0111778,3.9200184,4.245829,3.923448,6.660259,9.335337,9.784613,10.158438,11.129011,11.876661,12.411677,12.682614,13.924125,16.074476,17.775553,18.69811,18.163095,16.856422,14.754086,11.122152,8.875772,6.492209,4.602506,3.875434,5.0003386,6.632822,5.7582774,5.2815647,4.9660425,1.4129901,1.4610043,1.7490896,1.8279701,1.4541451,0.58988905,2.719663,1.3546871,0.09602845,0.1097468,0.11317638,0.024007112,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.0034295875,0.006859175,0.0034295875,0.030866288,0.06516216,0.048014224,0.12346515,0.16804978,0.22292319,0.2777966,0.26064864,0.26064864,0.25378948,0.33266997,0.5418748,0.881404,1.2758065,1.4815818,1.762808,2.0989075,2.1880767,3.542764,4.3658648,5.2918534,6.0978065,5.7068334,5.768566,6.4407654,7.7920227,9.513676,10.933525,12.298501,13.365103,13.687484,13.529722,13.838386,15.323397,15.54632,15.704081,16.269962,17.010754,17.072487,15.981877,15.162207,15.258235,16.12592,17.250826,17.991615,18.094503,17.504614,16.362562,16.369421,17.28169,18.279701,19.178253,20.423193,21.891056,22.299177,22.597551,22.906214,22.498095,23.729315,25.378946,26.448978,27.251501,29.408712,30.355278,31.929459,33.308155,33.76772,32.67368,33.383606,33.352737,32.625664,30.255821,24.305487,18.807858,15.594335,16.942162,21.513802,24.346642,21.822466,19.823015,18.825006,18.800999,19.239986,20.145397,21.03023,20.848463,19.980776,20.237995,21.44178,21.644127,20.910194,18.499195,12.864383,8.3922,6.8866115,5.826869,5.0483527,6.7459984,8.532814,7.2021337,6.8557453,8.107545,8.05953,11.036412,12.977559,14.071597,16.45516,24.202599,23.334913,22.762173,21.52066,20.388897,21.918493,21.582394,18.71183,18.252264,20.152256,19.349733,19.222837,19.768143,20.711279,20.406046,15.817257,10.6145735,7.582818,7.8846216,9.081548,5.1409516,4.928317,5.2472687,5.8165803,6.756287,8.604835,10.912948,12.181894,12.850664,13.63261,15.512024,15.563468,15.704081,15.566897,15.241087,15.29596,16.448301,17.12393,17.737827,18.396307,18.914175,19.239986,18.612371,18.28656,18.886738,20.37175,21.174273,21.808746,22.408924,22.87192,22.865059,23.091412,22.398636,21.20171,20.018501,19.46634,19.397747,18.800999,18.0362,17.4566,17.388008,18.4649,19.401176,19.562366,19.171394,19.294859,19.198832,19.565796,19.644676,19.805868,21.53438,23.78076,24.425522,24.085993,23.043398,21.253153,20.248285,19.476627,17.971039,15.645778,13.293081,12.665466,12.144169,11.766914,11.585147,11.677745,11.609154,11.543991,11.495977,11.664027,12.442543,14.342535,15.999025,17.394867,18.341434,18.46147,18.766703,18.516342,18.571217,18.893597,18.54378,13.622321,12.672326,13.474849,13.807519,11.447963,10.998687,10.659158,10.422516,10.501397,11.362224,12.415107,12.439114,12.253916,12.315649,12.730629,13.155897,13.042721,12.778643,12.154458,10.323058,10.093276,10.127572,10.124143,9.959522,9.692014,10.545981,10.494537,9.925226,9.290752,9.126132,9.006097,9.201583,9.325048,9.410788,9.901219,10.576848,10.940384,10.662587,9.860064,9.119273,10.364213,10.518545,10.230459,9.956093,9.97324,9.331907,9.373062,9.544542,9.568549,9.441654,8.923786,8.567109,8.738589,9.4862385,10.549411,9.757176,8.930646,8.800322,9.06097,8.385342,8.344186,10.14472,11.2250395,10.943813,10.5597,0.4938606,0.6276145,0.64133286,0.61389613,0.59331864,0.59674823,0.6241849,0.6241849,0.6207553,0.6241849,0.64133286,0.6207553,0.5693115,0.5555932,0.58988905,0.61389613,0.6344737,0.6859175,0.70649505,0.69963586,0.7133542,0.77851635,0.7510797,0.67219913,0.5796003,0.48357183,0.432128,0.41498008,0.41498008,0.41840968,0.42183927,0.39783216,0.4389872,0.53844523,0.65162164,0.6859175,0.85396725,0.91569984,0.94999576,1.0220171,1.1797781,1.2346514,1.3546871,1.3443983,1.3512574,1.8416885,1.8999915,2.253239,2.9151495,3.6113555,3.7691166,5.336438,7.0203657,9.023245,11.396519,14.054449,10.947243,7.1232533,4.7259717,3.758828,2.0920484,1.3581166,1.1523414,1.196926,1.3066728,1.4095604,1.0425946,0.88826317,0.82996017,0.78194594,0.70649505,0.6790583,0.45956472,0.25378948,0.19548649,0.36010668,0.22635277,0.15776102,0.14404267,0.25378948,0.65162164,1.1592005,1.0631721,0.72021335,0.37039545,0.12003556,0.044584636,0.034295876,0.048014224,0.10288762,0.2469303,0.30866286,0.5178677,0.7373613,0.8128122,0.58645946,0.4355576,0.29151493,0.18519773,0.14061308,0.15776102,0.072021335,0.024007112,0.0034295875,0.0,0.0,0.006859175,0.024007112,0.08573969,0.15090185,0.09945804,0.25378948,0.18519773,0.13032432,0.16462019,0.17833854,0.6756287,0.5144381,0.91227025,1.6256244,0.96371406,0.4424168,0.70306545,1.0494537,1.0631721,0.61389613,0.9294182,1.1523414,0.9294182,0.5453044,0.9294182,1.8485477,2.7299516,2.6922262,1.8759843,1.4404267,1.4438564,1.5055889,1.3478279,1.1317638,1.4541451,1.2517995,0.99801,0.7922347,0.6824879,0.6379033,0.8265306,0.77508676,0.864256,1.0117283,0.6756287,0.89855194,0.89855194,0.9294182,1.0494537,1.1283343,0.8128122,0.77508676,0.72364295,0.64476246,0.7956643,0.6859175,0.70649505,0.91569984,1.097468,0.7682276,1.0734608,0.90541106,0.82996017,0.96371406,0.9842916,1.2792361,1.0288762,0.90541106,1.0563129,1.1249046,0.88826317,0.83681935,0.8162418,0.85396725,1.1489118,0.90198153,0.9362774,0.8745448,0.7442205,0.9842916,0.77165717,0.67219913,0.72364295,0.84024894,0.84024894,0.7922347,0.9362774,1.0254467,0.99801,0.9568549,0.7990939,0.83338976,1.2483698,1.8005334,1.8313997,2.386993,2.9494452,3.5187566,3.9337368,3.858286,3.5290456,3.3781435,3.100347,2.8122618,3.0660512,3.192946,3.5770597,3.9337368,4.0263357,3.6525106,3.82399,4.262977,4.5167665,4.434457,4.1463714,4.297273,4.431027,4.506478,4.7088237,5.442755,5.802862,5.73427,4.770556,3.4981792,3.5702004,4.2595477,4.7671266,5.0826488,5.2987127,5.6210938,6.6705475,7.1232533,7.425057,7.932636,8.8929205,9.218731,9.647429,10.134431,10.545981,10.672876,11.063849,11.447963,11.859513,12.181894,12.123591,11.585147,11.519984,11.718901,11.965831,12.055,12.048141,11.413667,10.772334,10.367643,10.05898,10.131001,10.048691,9.846346,9.602845,9.448513,9.287323,9.956093,10.521975,10.666017,10.679735,10.89237,11.293632,12.130451,13.255356,14.13333,15.9578705,16.96617,18.097933,19.476627,20.412905,23.341772,20.793589,18.962189,19.922474,21.644127,25.76649,28.218645,26.126596,20.649546,17.000465,17.53891,15.995596,12.655178,8.580828,5.593657,2.6064866,1.0768905,0.6824879,0.8779744,0.9294182,0.8093826,0.6310441,0.47671264,0.39440256,0.3841138,0.42869842,0.5590228,0.6927767,0.8676856,1.2517995,1.704505,2.3595562,3.1312134,3.9268777,4.6436615,6.4819202,7.98065,9.695444,11.22161,11.180455,13.749216,15.151917,15.951012,15.666355,12.747777,16.602633,22.182571,21.232576,12.929544,3.8925817,1.9102802,2.2600982,2.3424082,1.4404267,0.72707254,0.29837412,0.28465575,0.6379033,1.2483698,1.9445761,3.0146074,5.2987127,6.3721733,5.1238036,1.7353712,2.7093742,3.0866287,3.2958336,3.8479972,5.329579,9.541112,11.4033785,12.535142,13.440554,13.526293,7.7783046,6.451054,6.40304,6.701414,8.594546,9.054111,10.062409,11.996697,14.273943,15.367981,15.313108,14.915276,16.643787,19.651537,19.78186,21.167414,19.36688,15.803539,11.732618,8.213862,6.5950966,4.6436615,3.4776018,3.5290456,4.554492,5.895461,5.645101,5.878313,5.926327,2.3732746,1.8554068,1.3992717,1.0940384,0.8779744,0.5521636,1.8108221,0.9294182,0.09602845,0.041155048,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.07888051,0.09259886,0.11317638,0.14404267,0.14061308,0.17490897,0.36010668,0.48700142,0.5453044,0.6927767,0.8505377,0.96714365,1.2929544,1.7765263,2.0714707,2.7230926,3.2821152,4.1429415,4.9591837,4.6848164,5.2644167,5.809721,6.619104,7.7885933,9.201583,10.923236,12.38767,13.179905,13.567448,14.507155,15.71437,15.505165,15.193072,15.278812,15.453721,15.755525,15.680074,15.415996,15.343974,16.009314,17.71039,18.224829,18.193962,17.813278,16.832415,17.679523,18.499195,19.137098,19.661825,20.36832,21.301168,22.234016,23.427511,24.61415,25.005123,25.94826,27.639046,28.92857,30.039757,32.553646,34.885765,35.59226,35.365906,34.693707,33.90147,34.31988,33.640823,30.845709,26.959988,25.042849,19.857311,17.717249,17.851004,19.363451,21.236006,20.334024,19.473198,19.586374,20.011642,18.512913,24.411804,20.659836,16.307688,15.069608,15.333686,16.249386,16.173935,16.585485,16.12935,10.607714,9.246168,7.380472,7.1061053,10.192734,18.087645,15.570327,10.47396,8.22758,9.438225,9.887501,14.5585985,15.566897,15.854982,17.665806,22.53239,22.69358,22.679861,22.041958,21.908205,25.001692,22.957659,20.347742,20.601532,22.059107,17.971039,18.241976,17.669235,16.743246,15.402277,13.039291,9.633711,8.954653,9.22902,8.879202,6.4887795,5.9160385,6.0669403,6.783724,8.131552,10.39165,11.2593355,11.506266,11.622872,12.103014,13.437123,14.057879,15.302819,15.697222,15.165636,15.035312,15.618341,15.854982,16.016174,16.424294,17.449741,19.236557,20.810738,21.633839,21.832754,22.196291,22.021381,21.935642,22.391777,23.211449,23.568125,23.904224,23.304047,22.244305,21.153696,20.426622,19.493774,18.807858,18.084215,17.364002,17.021042,18.132229,18.897026,19.027351,18.87302,19.404606,19.70298,19.747564,19.480057,19.558937,21.36633,23.705309,25.286348,25.142305,23.304047,20.79016,19.349733,18.567787,17.658945,16.047039,13.365103,12.679185,12.507706,12.38424,12.041282,11.406808,11.506266,11.523414,11.962401,12.850664,13.718349,14.54831,15.357693,16.105343,16.828985,17.63494,18.307138,18.663815,19.065077,19.493774,19.569225,14.147048,12.706621,12.9638405,12.939834,10.926665,11.537132,11.701753,11.393089,11.067279,11.660598,12.1921835,11.797781,11.38966,11.348505,11.5645685,12.243628,11.924676,11.334786,10.837497,10.449953,10.113853,10.048691,9.750318,9.39021,9.798331,10.738038,10.693454,10.151579,9.523964,9.136421,8.700864,9.081548,9.355915,9.362774,9.709162,10.089847,10.340206,10.031544,9.23245,8.525954,9.517105,10.045261,10.1481495,10.021255,10.010965,9.297611,9.239308,9.277034,9.1810055,9.047252,8.567109,8.279024,8.519095,9.146709,9.582268,8.776315,8.385342,8.207003,8.093826,7.963502,9.050681,10.360784,11.348505,11.71547,11.427385,0.58645946,0.7339317,0.66876954,0.6310441,0.70306545,0.8025235,0.7442205,0.71678376,0.6893471,0.65505123,0.65848076,0.6310441,0.6001778,0.61046654,0.65505123,0.69963586,0.7305021,0.72021335,0.6927767,0.67219913,0.67219913,0.6379033,0.59331864,0.53501564,0.48014224,0.4664239,0.4424168,0.4389872,0.44584638,0.45613512,0.48700142,0.4698535,0.490431,0.5761707,0.7099246,0.8093826,1.0082988,1.0631721,1.0768905,1.1146159,1.2037852,1.2483698,1.4335675,1.5364552,1.6187652,2.0097382,1.9925903,2.627064,3.426158,4.166949,4.897451,6.728851,8.220721,10.501397,13.491997,15.906426,12.538571,7.425057,3.5976372,2.0234566,1.605047,1.2792361,1.2792361,1.3752645,1.4610043,1.5673214,1.2620882,1.0940384,0.980862,0.8745448,0.7407909,0.6859175,0.58302987,0.4389872,0.30866286,0.28808534,0.18176813,0.13032432,0.1097468,0.16462019,0.38754338,0.96714365,1.0734608,0.82996017,0.4389872,0.17490897,0.1097468,0.106317215,0.116605975,0.17833854,0.42526886,0.42526886,0.607037,0.7682276,0.7888051,0.6036074,0.48014224,0.34295875,0.216064,0.1371835,0.15776102,0.12346515,0.06859175,0.024007112,0.0034295875,0.0,0.01371835,0.030866288,0.06516216,0.10288762,0.14404267,0.6001778,0.548734,0.37039545,0.274367,0.2709374,0.65848076,0.66876954,1.1694894,1.9582944,1.7696671,1.4472859,1.5673214,1.5673214,1.255229,0.8265306,0.84367853,0.8196714,0.6824879,0.5693115,0.8025235,2.1057668,2.6613598,2.5310357,2.0714707,1.9171394,1.6427724,1.3101025,1.1454822,1.2277923,1.488441,1.0460242,1.0940384,1.0220171,0.8025235,1.0151579,1.0185875,0.9362774,1.0117283,1.1249046,0.7956643,1.0151579,0.9945804,0.97400284,1.0082988,0.9568549,0.75450927,0.7922347,0.7613684,0.66876954,0.8196714,0.6824879,0.7888051,0.83338976,0.77508676,0.84367853,1.1420527,1.0151579,0.89169276,0.980862,1.2655178,1.2963841,1.1214751,1.138623,1.3855534,1.5364552,1.1832076,1.0048691,0.8848336,0.84367853,1.0494537,0.91227025,0.91227025,0.8196714,0.70306545,0.922559,0.89855194,0.70306545,0.7099246,0.90884066,0.89855194,0.8093826,0.8676856,0.9534253,1.0151579,1.0666018,0.939707,0.9362774,1.2415106,1.6736387,1.6976458,2.3424082,2.884283,3.3266997,3.5564823,3.3644254,3.1689389,3.0660512,2.9700227,2.9494452,3.2375305,3.3129816,3.666229,3.9714622,4.029765,3.7622573,3.6216443,3.9268777,4.0777793,3.9337368,3.8171308,3.8548563,4.081209,4.184097,4.2698364,4.8768735,5.7479887,6.3378778,5.545643,3.9851806,3.9680326,4.3521466,4.945465,5.3673043,5.562791,5.761707,6.385892,6.742569,7.0752387,7.579388,8.399059,9.170717,9.602845,10.031544,10.539123,10.947243,11.015835,11.207891,11.334786,11.324498,11.235329,10.957532,10.926665,11.015835,11.091286,11.012405,10.991828,10.501397,9.9698105,9.599416,9.345626,9.585697,9.595985,9.595985,9.637141,9.595985,9.3079,9.9698105,10.521975,10.72432,11.1393,11.201033,11.653738,12.744347,14.195063,15.169065,17.278261,18.519772,19.558937,20.334024,20.03565,22.93708,20.834743,20.61182,22.309467,19.099373,25.927681,27.27208,25.715046,22.62156,18.159666,16.774113,15.395418,12.696333,8.697433,4.763697,2.218943,0.94656616,0.6241849,0.764798,0.7305021,0.67219913,0.607037,0.53844523,0.4698535,0.41498008,0.39097297,0.42526886,0.548734,0.77508676,1.097468,1.5364552,2.270387,2.9631636,3.4878905,3.9131594,5.3981705,6.5470824,8.553391,10.854645,11.149589,12.871242,14.7369375,15.971589,15.837835,13.656617,15.501736,16.287111,13.37882,7.421627,2.3252604,1.0048691,0.9294182,0.939707,0.66533995,0.5178677,0.25721905,0.28122616,0.5727411,1.0768905,1.7010754,3.0729103,3.450165,3.5942078,3.799983,3.8891523,4.7088237,4.557922,4.3761535,5.079219,7.548522,12.991278,15.662926,17.03819,18.327715,20.498644,15.079896,12.120162,10.820349,10.707172,11.633161,11.646879,12.874671,14.726648,16.252815,16.13621,14.856973,14.273943,16.39,19.384027,17.604073,18.54378,16.047039,11.938394,7.956643,5.754848,4.3007026,3.0866287,2.6887965,3.07634,3.6010668,4.8082814,5.662249,6.3893213,6.0566516,2.5824795,2.0680413,1.2380811,0.5590228,0.33952916,0.71678376,1.0768905,1.3752645,0.9259886,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.010288762,0.006859175,0.020577524,0.037725464,0.13032432,0.33266997,0.4664239,0.52472687,0.66876954,0.5693115,0.6859175,1.0288762,1.5021594,1.8897027,2.201795,2.7368107,3.4398763,4.1017866,4.372724,5.1752477,5.5387836,5.90575,6.636252,8.018375,9.918367,11.533703,12.524854,13.179905,14.428274,16.019604,15.772673,14.891269,14.198492,14.147048,14.764374,15.484588,15.734947,15.752095,16.582056,18.259123,18.488907,18.293419,18.084215,17.652086,18.567787,19.185112,19.709839,20.29287,21.033659,21.342323,22.395206,24.092852,25.958548,27.124607,27.896265,29.364128,30.657082,31.716825,33.280716,35.81518,36.0141,35.208145,34.49822,34.72114,34.74515,33.83631,30.667372,26.486704,25.114868,21.45207,20.543228,19.6241,18.756414,20.814167,21.167414,21.0268,21.335464,21.3629,18.718689,27.412693,18.996485,10.621432,8.652849,8.635701,9.458802,9.033533,11.005547,13.138749,7.3118806,7.517656,6.1149545,9.56512,18.214539,26.298077,18.255693,11.211322,8.176137,9.023245,10.48082,14.87755,17.086205,17.096493,16.016174,16.091625,17.463459,18.578075,19.281141,20.237995,22.94051,21.45893,20.841602,21.52066,21.476076,16.225378,15.433144,14.781522,14.325387,14.157337,14.4317045,12.665466,11.962401,10.443094,8.1487,7.0375133,5.6656785,6.169828,7.610255,9.379922,11.177026,11.286773,10.868362,10.64201,11.002116,12.05157,13.951562,15.488017,15.851553,15.254805,14.946142,15.028452,14.658057,14.38026,14.678635,15.971589,18.595222,21.465788,23.26975,23.708738,23.506393,23.437801,23.34863,23.811626,24.627867,24.837072,25.132017,24.264332,23.386356,22.882208,22.354052,21.143406,20.207129,19.239986,18.344864,18.04306,18.732407,18.61923,18.399736,18.602083,19.552078,19.963629,19.750994,19.630959,20.045938,21.170843,23.019392,24.833643,24.963966,23.139427,20.488356,18.547209,17.528622,16.753534,15.638919,13.690913,13.1421795,13.3033695,13.495427,13.203912,12.079007,11.646879,11.766914,12.586586,13.786942,14.586036,14.033872,14.448852,15.234227,16.091625,17.024471,18.413456,19.257133,19.648108,19.634388,19.219408,14.953001,13.615462,13.025573,12.202472,11.365653,12.699762,12.758065,12.044711,11.362224,11.787492,12.151029,11.509696,11.087856,11.163307,11.084427,11.180455,10.573419,10.014396,9.846346,10.0041065,9.897789,9.928656,9.619993,9.22902,9.781183,10.672876,10.789482,10.38479,9.705732,8.954653,8.567109,8.886061,9.14328,9.15014,9.280463,9.410788,9.335337,9.06097,8.690575,8.423067,8.800322,9.482809,9.921797,9.956093,9.801761,9.23245,9.0644,8.971801,8.868914,8.927217,8.519095,8.179566,8.275595,8.618553,8.471081,7.6171136,7.548522,7.606825,7.689135,8.241299,9.283894,10.189304,11.201033,12.044711,11.948683,0.6036074,0.72021335,0.69963586,0.72364295,0.8505377,0.9945804,0.7956643,0.7407909,0.70649505,0.64819205,0.607037,0.59331864,0.607037,0.6379033,0.67219913,0.6824879,0.67219913,0.59674823,0.53844523,0.5212973,0.52472687,0.4698535,0.4938606,0.4938606,0.47328308,0.5453044,0.4938606,0.48700142,0.48014224,0.48014224,0.5144381,0.53158605,0.6036074,0.69963586,0.8162418,0.9945804,1.0768905,1.0563129,1.0666018,1.1283343,1.1214751,1.3169615,1.4987297,1.6599203,1.7902447,1.879414,2.1983654,3.083199,3.6799474,4.3521466,6.6876955,8.045813,9.156999,11.022695,13.474849,15.169065,15.398848,11.063849,5.9331865,2.393852,1.4541451,1.3272504,1.3546871,1.3924125,1.3649758,1.2860953,1.2106444,1.1832076,1.1008976,0.9568549,0.85396725,0.86082643,0.84367853,0.7373613,0.5796003,0.52472687,0.39783216,0.29151493,0.20577525,0.18176813,0.31895164,0.66191036,0.7990939,0.66876954,0.3806842,0.20920484,0.22978236,0.23664154,0.2194936,0.29151493,0.6859175,0.77851635,0.8162418,0.78194594,0.66876954,0.50757897,0.432128,0.33609957,0.23664154,0.16462019,0.16804978,0.18519773,0.12689474,0.0548734,0.010288762,0.0034295875,0.010288762,0.020577524,0.06859175,0.1371835,0.15090185,0.7613684,0.83681935,0.59674823,0.31552204,0.32581082,0.32581082,0.7888051,1.903421,3.0660512,2.8980014,2.5893385,2.1846473,1.7079345,1.2758065,1.0906088,0.72707254,0.5521636,0.5418748,0.65505123,0.8265306,1.9342873,2.4967396,2.3286898,1.862266,2.1469216,1.3409687,1.1077567,1.1008976,1.0906088,0.97400284,0.61389613,0.97400284,1.1660597,1.0837497,1.4198492,1.1180456,1.039165,1.0906088,1.1214751,0.91569984,1.2826657,1.08032,0.9431366,1.0254467,0.9945804,0.9568549,1.0528834,0.96371406,0.77851635,1.0117283,0.86082643,0.9259886,0.9328478,0.88826317,1.0940384,1.0082988,1.0940384,1.1008976,1.0871792,1.4232788,1.0666018,1.0528834,1.2072148,1.3924125,1.5021594,1.4129901,1.3238207,1.1420527,0.9259886,0.8711152,0.72707254,0.72707254,0.71678376,0.69963586,0.82996017,0.8265306,0.70649505,0.71678376,0.8505377,0.8779744,0.6893471,0.70649505,0.78194594,0.8779744,1.0837497,1.0323058,1.039165,1.1283343,1.2655178,1.3409687,2.1915064,2.4555845,2.5584722,2.633923,2.5378947,2.3081124,2.4007113,2.5927682,2.767677,2.9322972,3.0660512,3.3987212,3.7279615,3.9268777,3.9371665,3.6353626,3.7485392,3.7862647,3.6559403,3.666229,3.6456516,3.882293,4.190956,4.588788,5.295283,6.560801,7.8606143,7.2604365,5.0655007,3.82399,4.57164,4.9420357,5.178677,5.453044,5.861165,5.967482,6.3961806,6.8454566,7.233,7.7097125,9.043822,9.517105,9.904649,10.460241,10.930096,10.251037,10.093276,10.007536,9.856634,9.818909,10.031544,10.113853,10.14129,10.14472,10.089847,9.959522,9.860064,9.794902,9.702303,9.455373,9.47938,9.407358,9.342196,9.373062,9.568549,9.362774,10.000677,10.624862,11.087856,11.952112,11.934964,12.130451,13.121602,14.812388,16.441442,18.608942,19.730417,20.395756,20.467777,19.106232,18.708399,19.973917,23.338343,24.922812,16.558048,24.223177,26.040857,25.862518,23.794477,16.191082,14.623761,15.333686,13.886399,9.2153015,3.6353626,1.6873571,0.84024894,0.6893471,0.77851635,0.58988905,0.58645946,0.66191036,0.6893471,0.64476246,0.607037,0.53158605,0.59331864,0.7407909,0.94999576,1.214074,1.5124481,2.1880767,2.7470996,3.0283258,3.2032347,4.4584637,5.4016004,7.473071,10.271614,11.571428,13.756075,15.947581,15.748666,13.958421,14.562028,13.687484,12.154458,9.321619,5.5147767,1.99602,0.8128122,0.5693115,0.5418748,0.42183927,0.31209245,0.23664154,0.34638834,0.59331864,1.214074,2.7573884,5.638242,6.5059276,6.7391396,6.8043017,6.279575,6.4579134,5.785714,5.31929,5.5662203,6.4887795,9.163857,11.194174,12.346515,14.325387,20.773012,19.524641,17.53891,15.258235,13.656617,14.229359,15.608052,16.029892,16.077906,15.536031,13.399398,11.303921,11.207891,13.05301,14.750656,12.199042,11.30735,9.177576,6.6293926,4.5956473,4.1360826,2.8739944,2.2978237,2.2360911,2.4041407,2.411,3.5461934,5.288424,6.276145,5.4599032,2.095478,1.7799559,1.1592005,0.548734,0.25378948,0.5761707,0.980862,2.1674993,1.7799559,0.08573969,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.041155048,0.14061308,0.14747226,0.24007112,0.44584638,0.65848076,0.48014224,0.7133542,1.0254467,1.2723769,1.4815818,2.0817597,2.5961976,3.0523329,3.5804894,4.40702,5.003768,5.2609873,5.6656785,6.48535,7.7577267,9.561689,10.851214,11.705182,12.346515,13.128461,15.189643,15.532601,14.544881,13.29994,13.5503,14.695783,15.6526375,16.29397,16.904436,18.180243,18.79071,18.36544,18.063637,18.183672,18.156237,18.37573,19.188541,20.059656,20.923914,22.175713,22.350622,23.338343,24.902235,26.630747,27.9237,29.172071,30.657082,31.76141,32.176388,31.884874,33.465916,33.74028,33.620247,33.863747,35.08468,34.83775,34.182697,32.653103,29.861418,25.495554,23.01596,22.251163,21.500084,21.263443,24.240324,23.832203,23.36921,22.748453,21.908205,20.817596,26.846811,16.6335,6.7871537,3.5530527,2.8088322,4.1326528,3.649081,6.7391396,10.971251,6.077229,5.1821065,4.5339146,12.154458,24.398085,25.94826,15.151917,8.81404,6.543653,7.226141,9.019815,11.290202,16.510035,17.007324,12.339656,9.287323,11.108434,12.792361,14.147048,15.22051,16.311117,16.698662,18.485476,19.555508,18.574646,14.983868,13.087306,13.2862215,14.239647,15.717799,18.584934,17.78927,14.928994,11.351934,8.213862,6.468202,5.2506986,6.135532,8.038953,9.914937,10.7586155,11.149589,10.816919,10.6317215,11.0981455,12.377381,14.839825,15.700651,15.614912,15.251375,15.29253,14.836395,14.085316,14.013294,14.925565,16.479168,18.694681,20.61182,22.295748,23.568125,23.993395,24.833643,25.51956,26.26721,26.83995,26.541578,26.675331,25.478405,24.730755,24.682741,24.065414,23.228596,22.20315,20.992504,19.984205,19.939621,20.097382,19.318867,18.986197,19.469769,20.097382,19.905325,19.6241,19.977346,20.855322,21.318316,22.059107,22.8582,22.967947,22.048819,20.183123,17.830425,16.37285,15.343974,14.503725,13.817808,13.457702,13.7526455,14.057879,13.934414,13.149038,12.569438,12.723769,13.138749,13.570878,14.027013,12.984418,13.855534,15.278812,16.510035,17.442883,19.44919,20.37518,20.37518,19.5315,17.830425,15.237658,14.483148,13.457702,12.1921835,12.843805,13.742357,12.9707,11.808069,11.218181,11.842365,12.432255,11.694893,11.362224,11.681175,11.427385,10.521975,9.623423,9.445084,9.757176,9.386781,9.80862,10.065839,10.017825,9.743458,9.537683,10.4533825,10.765475,10.504827,9.770895,8.707723,8.388771,8.405919,8.64599,8.855195,8.64256,8.604835,8.340756,8.224151,8.357904,8.597976,8.690575,9.331907,9.81205,9.884071,9.753747,9.342196,9.0644,8.81747,8.690575,8.97523,8.707723,8.224151,7.939495,7.8983397,7.764586,7.0443726,6.852316,7.267296,8.086967,8.824328,9.074688,9.925226,11.094715,12.055,12.037852,0.45613512,0.64133286,0.7682276,0.805953,0.7990939,0.8848336,0.7613684,0.70649505,0.6790583,0.70649505,0.84024894,0.91227025,0.90198153,0.8676856,0.8162418,0.7339317,0.72021335,0.65162164,0.6276145,0.65848076,0.67219913,0.59674823,0.6893471,0.6824879,0.5590228,0.53501564,0.5212973,0.5007198,0.5007198,0.53844523,0.6241849,0.66191036,0.8265306,0.980862,1.08032,1.1900668,1.0666018,1.0014396,0.96371406,0.9842916,1.1454822,1.546744,1.5741806,1.7388009,2.0749004,2.136633,2.6476414,3.2272418,3.525616,4.6745276,9.277034,8.433355,9.012956,10.213311,11.605724,13.107883,20.749004,19.737276,12.46312,3.8720043,1.4815818,1.371835,1.0666018,1.0082988,1.1866373,1.1763484,1.138623,1.1008976,1.0048691,0.8676856,0.7922347,0.8779744,0.90884066,0.8848336,0.84367853,0.85396725,0.7579388,0.5041494,0.26407823,0.14747226,0.18176813,0.4389872,0.4389872,0.37382504,0.37039545,0.5041494,0.5041494,0.42869842,0.29494452,0.20920484,0.3806842,0.881404,1.0631721,0.9774324,0.7373613,0.5178677,0.432128,0.36696586,0.32924038,0.29151493,0.16804978,0.15433143,0.09602845,0.037725464,0.0034295875,0.01371835,0.0034295875,0.037725464,0.10288762,0.16462019,0.15090185,0.16462019,0.18519773,0.16119061,0.106317215,0.106317215,0.40126175,1.471293,2.8088322,3.4364467,1.9239986,1.5433143,1.4232788,1.5124481,1.6016173,1.2963841,0.69963586,0.65162164,0.7476501,0.8265306,0.9602845,1.0837497,1.728512,1.8862731,1.4987297,1.4507155,1.0460242,1.4404267,1.3992717,0.864256,0.9602845,1.4129901,1.3992717,1.08032,0.8711152,1.4198492,0.9911508,0.85739684,0.77165717,0.72021335,0.91569984,1.4267083,1.0082988,0.7888051,1.0940384,1.4335675,0.9945804,1.1694894,1.2312219,0.9534253,0.61046654,0.91569984,0.90198153,0.91227025,0.9945804,0.8848336,0.7510797,0.85396725,0.91569984,0.8128122,0.5796003,0.5555932,0.77851635,0.96714365,1.097468,1.4027013,1.4027013,1.4678634,1.2963841,0.9431366,0.8093826,0.52815646,0.5693115,0.7613684,0.8779744,0.61046654,0.45270553,0.6241849,0.78194594,0.7682276,0.61046654,0.6344737,0.6036074,0.6344737,0.7305021,0.77851635,0.5693115,0.7922347,0.90198153,0.88826317,1.2655178,2.0097382,1.7593783,1.6290541,1.9274281,2.136633,1.9651536,1.903421,1.7833855,1.7250825,2.1503513,2.4315774,2.7779658,2.983741,3.2032347,3.9371665,3.5461934,3.841138,4.2526884,4.386442,4.0434837,4.2389703,4.2526884,4.5510626,5.31929,6.4544835,7.795452,8.076678,7.346176,5.693115,3.2512488,3.7142432,3.6559403,4.180667,5.411889,6.48535,6.4716315,6.8728933,7.133542,7.2707253,7.8434668,9.15014,9.47595,9.451943,9.513676,9.904649,9.829198,9.959522,10.041832,9.966381,9.736599,9.517105,9.277034,9.3079,9.541112,9.551401,9.541112,9.719451,9.928656,9.942374,9.489669,9.760606,9.990388,9.740028,9.201583,9.201583,9.297611,9.661148,10.240748,10.964391,11.732618,12.319078,12.586586,13.197053,14.486577,16.46545,18.221397,19.44919,20.059656,20.107672,19.792149,19.11995,20.982216,21.45893,19.490345,16.877,23.907654,26.078583,27.628757,26.918833,16.434584,14.126471,15.9750185,14.664916,8.748878,2.6716487,1.2415106,0.82996017,0.9328478,1.0528834,0.6859175,0.6756287,0.83681935,0.90198153,0.9259886,1.2655178,0.84024894,0.8779744,1.0117283,1.1900668,1.6770682,1.99602,2.8808534,3.4295874,3.450165,3.450165,4.400161,5.3707337,7.2432885,9.949233,12.449403,15.563468,15.875561,13.780083,11.938394,15.258235,14.05102,10.069269,6.0532217,3.2409601,1.371835,0.53158605,0.29151493,0.30523327,0.36010668,0.39783216,0.5178677,0.89855194,1.3615463,2.428148,5.3090014,10.569988,12.528283,10.048691,5.6348124,5.4016004,6.0978065,5.0346346,4.5784993,4.852866,3.7553983,2.9734523,2.411,2.4590142,4.636802,11.581717,11.986408,13.560589,13.728639,12.730629,13.594885,14.476289,13.111313,11.485688,10.103564,7.98065,7.956643,8.1041155,8.508806,8.327039,5.813151,4.629943,3.9954693,3.2855449,2.510458,2.3046827,1.6084765,1.1214751,0.9328478,0.9945804,1.1283343,2.3629858,3.9165888,5.0757895,4.9420357,2.4247184,1.5227368,1.1592005,0.84367853,0.4424168,0.19891608,0.45613512,0.35324752,0.18862732,0.08573969,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.020577524,0.30866286,0.70649505,0.548734,0.5727411,0.9842916,1.2312219,1.2517995,1.4335675,1.7388009,2.0268862,2.527606,3.2958336,4.2115335,4.4550343,4.616225,5.2575574,6.451054,7.781734,9.283894,10.374502,11.519984,12.493987,12.360233,12.895248,13.893259,14.208781,13.965281,14.527733,15.71094,16.767254,17.583494,18.313997,19.363451,18.471758,17.113642,16.828985,17.604073,17.899017,17.826996,19.730417,21.335464,22.03167,22.87192,23.643576,24.998262,26.133457,26.836521,27.495003,29.545897,31.305275,32.118088,32.25184,32.896603,34.25129,34.141544,33.8123,33.76772,33.76772,33.205265,33.222412,33.363026,32.797146,30.317553,27.436699,24.741043,23.11199,22.895926,23.911083,23.043398,23.146286,22.755312,22.868488,26.946268,24.713608,16.263103,7.7611566,2.6133456,1.4644338,2.5756202,2.6887965,5.7479887,10.14129,8.711152,6.7357097,6.1321025,12.319078,20.810738,17.195951,11.458252,6.0326443,4.0057583,5.1409516,5.861165,7.006647,11.907528,13.471419,10.323058,6.8214493,10.556271,11.526843,12.703192,14.040731,12.466551,13.906977,15.364552,16.664366,17.034761,15.107333,16.558048,16.300829,15.505165,15.46058,17.549198,17.37772,14.167625,10.569988,8.261876,7.9189177,8.090397,7.822889,8.40249,9.671436,10.024684,11.207891,11.917816,12.394529,12.915827,13.7938,14.280802,15.265094,16.156786,16.70895,17.014183,15.121051,13.852104,14.2190695,16.21166,18.79757,19.188541,18.61923,18.962189,20.86904,23.773901,24.799347,25.93454,26.702768,26.737064,25.77335,25.711617,25.44068,25.334362,25.029129,23.406935,22.247734,21.500084,21.287449,21.685282,22.734735,22.11398,21.44521,21.524092,22.172283,22.247734,21.479506,20.920483,20.779871,21.088533,21.699,21.342323,20.402617,20.018501,20.159115,19.6241,17.768692,15.810398,14.38369,13.574307,12.939834,12.205902,12.418536,12.867812,13.173045,13.258785,14.016724,14.13333,13.248496,11.866373,11.351934,12.096155,13.996146,15.638919,16.846134,18.677534,19.579515,20.409475,20.464348,19.442331,17.439453,15.22051,14.417986,13.834956,13.46799,14.479718,13.310229,11.835506,10.762046,10.717461,12.267634,13.2690735,12.476839,12.000127,12.089295,11.122152,9.657719,9.201583,9.654288,10.388221,10.254466,10.803201,11.2593355,11.314209,10.902658,10.206452,10.696883,10.563129,10.319629,9.9869585,9.108984,8.303031,7.8537555,8.1487,8.738589,8.361334,8.032094,7.8846216,7.8503256,8.073249,8.927217,9.352485,9.544542,9.599416,9.692014,10.069269,9.815479,9.355915,8.783174,8.412778,8.803751,9.132992,8.556821,7.795452,7.3598948,7.5690994,6.944915,6.4407654,6.9792104,8.296172,8.958082,9.72631,10.604284,11.519984,12.099585,11.674315,0.4698535,0.50757897,0.64819205,0.91569984,1.1694894,1.1180456,0.9842916,0.939707,0.89169276,0.8505377,0.9259886,1.0185875,1.0220171,0.9945804,0.97400284,0.9774324,1.0323058,0.9534253,0.8128122,0.72021335,0.82996017,0.7579388,0.6790583,0.607037,0.53844523,0.48357183,0.5418748,0.6241849,0.72364295,0.7956643,0.78537554,0.78194594,0.84024894,0.90541106,0.97057325,1.08032,0.99801,0.9774324,0.9774324,1.0254467,1.1934965,1.5776103,1.6942163,1.9239986,2.2326615,2.1983654,2.6887965,3.350707,4.2218223,5.861165,9.349055,7.1712675,8.467651,10.230459,11.653738,14.13333,28.637054,26.490133,16.441442,6.090947,1.8828435,1.646202,1.3272504,1.1626302,1.2346514,1.4678634,1.529596,1.3101025,1.097468,0.9774324,0.8676856,0.97057325,1.0288762,0.97057325,0.864256,0.91569984,0.8471081,0.6001778,0.3566771,0.24007112,0.30523327,0.45270553,0.5144381,0.47328308,0.4972902,0.9431366,1.0700313,0.86082643,0.5590228,0.36010668,0.39440256,0.61046654,0.9911508,1.08032,0.7990939,0.432128,0.39783216,0.37725464,0.33609957,0.25721905,0.14404267,0.15090185,0.13375391,0.08916927,0.030866288,0.01371835,0.0034295875,0.006859175,0.020577524,0.034295876,0.041155048,0.07545093,0.09259886,0.09259886,0.082310095,0.082310095,0.4355576,1.4918705,2.2498093,2.3835633,2.2292318,2.5996273,2.4555845,1.8931323,1.1934965,0.8196714,0.8471081,0.764798,0.7613684,0.7407909,0.33952916,1.4267083,2.1812177,2.1263442,1.5158776,1.3409687,0.89855194,1.1146159,1.1008976,0.7956643,0.9602845,1.5776103,1.1866373,0.7956643,0.82996017,1.1249046,0.922559,0.8745448,1.0837497,1.3546871,1.2072148,1.2037852,1.0700313,0.9774324,1.0151579,1.1900668,0.9259886,0.9534253,1.0460242,0.9842916,0.5727411,0.7922347,0.7888051,0.7476501,0.7956643,1.0185875,1.08032,0.881404,0.7956643,0.82996017,0.6173257,0.6207553,0.70649505,0.96371406,1.3203912,1.5364552,0.8745448,0.96371406,1.0254467,0.85396725,0.7956643,0.8196714,0.8025235,0.90541106,0.9774324,0.5624523,0.71678376,0.6207553,0.5796003,0.5796003,0.29151493,0.5521636,0.6241849,0.69963586,0.7922347,0.75450927,0.66191036,0.7407909,0.8676856,0.94999576,0.88826317,1.214074,1.2277923,1.2895249,1.4987297,1.6976458,1.5741806,1.4232788,1.2998136,1.2415106,1.2483698,1.7147937,2.4212887,3.0283258,3.4227283,3.7039545,3.0317552,3.3815732,4.0537724,4.540774,4.5201964,4.8014226,4.8151407,5.192395,6.0497923,6.9792104,6.992929,7.250148,7.3187394,6.3173003,2.9082901,3.1586502,3.57363,4.2355404,5.055212,5.7754254,6.5367937,6.7185616,6.684266,6.694555,6.914048,8.357904,9.259886,9.56512,9.541112,9.80519,9.623423,9.527394,9.403929,9.3079,9.465661,9.959522,9.613133,9.338767,9.273604,8.80718,8.676856,8.961512,9.441654,9.853205,9.870353,9.9801,9.846346,9.585697,9.369633,9.407358,9.3593445,9.760606,10.343636,10.906088,11.293632,11.842365,12.120162,12.665466,13.526293,14.243076,15.415996,16.530611,17.405157,17.902447,17.936743,18.231688,19.017063,18.166525,15.834405,14.472859,17.62465,23.44809,27.85511,26.833092,16.434584,17.926455,17.545769,13.265644,6.48535,2.037175,1.0940384,1.0323058,1.2449403,1.2277923,0.58988905,0.59674823,0.6824879,0.75450927,0.85739684,1.1797781,1.1454822,1.0906088,1.2758065,1.8005334,2.6304936,2.4212887,2.983741,3.1655092,3.1312134,4.3521466,4.396731,5.1992545,6.831738,9.301042,12.535142,12.857523,11.290202,12.360233,16.359133,19.346302,15.618341,9.506817,4.5442033,2.0165975,0.97057325,0.34295875,0.14404267,0.12689474,0.15776102,0.21263443,0.42526886,0.85396725,1.4678634,2.9494452,6.6876955,11.88352,12.055,8.347616,3.9611735,4.170378,3.8685746,3.333559,2.8808534,2.8328393,3.5221863,3.0317552,3.234101,3.4913201,4.1463714,6.492209,6.543653,6.725421,6.5539417,6.3138704,7.0546613,7.394191,7.7783046,7.599966,7.058091,7.15069,7.233,7.5416627,8.608265,8.872343,4.6779575,2.8396983,2.0406046,1.6427724,1.3786942,1.3752645,1.1900668,0.9842916,1.1351935,1.6530612,2.177788,2.8465576,4.0537724,4.914599,4.8940215,3.806842,2.2463799,1.5158776,1.1146159,0.764798,0.39440256,0.2777966,0.20920484,0.12346515,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.16462019,0.31895164,0.3018037,0.1371835,0.0,0.037725464,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.06516216,0.06859175,0.2777966,0.6001778,0.59674823,0.66191036,0.9328478,1.097468,1.1351935,1.3375391,1.5844694,1.9514352,2.411,3.0797696,4.197815,4.3761535,4.8425775,5.813151,7.2364297,8.783174,9.170717,10.093276,11.132441,12.037852,12.713481,12.517994,12.672326,13.265644,14.184773,15.086755,16.153357,17.394867,18.139088,18.389448,18.814716,17.943602,16.602633,16.074476,16.417435,16.496315,17.223389,19.613811,22.11055,24.085993,25.828222,25.999702,26.407824,26.860529,27.316664,27.885975,29.967735,31.065203,32.131805,33.42133,34.49822,35.14984,34.227283,32.567364,31.027477,30.458166,29.439579,28.856548,28.678211,29.01431,30.111778,29.652214,27.573883,25.10115,23.386356,23.533829,23.44809,24.669024,25.128588,24.250612,22.967947,17.45317,13.039291,7.8503256,7.7440085,26.291218,7.997798,4.2423997,7.2775846,11.2421875,12.168177,10.89237,11.63659,14.064738,16.63007,16.561478,11.050131,6.478491,5.0757895,6.341307,7.0306544,9.818909,12.55915,14.784951,15.861842,14.973578,11.856084,12.795791,13.96871,13.944703,13.687484,15.038741,14.198492,13.536582,13.392539,12.079007,15.484588,14.623761,12.421966,11.129011,12.298501,11.063849,10.340206,11.036412,12.524854,12.63117,11.862943,11.331357,11.036412,11.06042,11.550851,12.05157,13.37882,14.503725,14.908417,14.586036,14.363112,14.404267,14.822677,15.364552,15.415996,15.29939,15.302819,15.892709,16.976458,17.895588,18.842154,19.421753,20.320305,21.37662,21.575535,22.035099,23.533829,24.346642,24.398085,25.258911,26.28093,26.589592,26.215767,25.059996,22.868488,21.153696,20.817596,21.290878,22.014523,22.429502,21.565247,21.033659,21.174273,21.829325,22.333473,22.20658,22.072824,22.247734,22.384918,21.503513,20.749004,19.569225,19.20569,19.552078,19.171394,18.262554,16.80155,15.199932,13.96871,13.684054,13.46799,13.581166,13.584596,13.646329,14.555169,15.614912,16.221949,15.683503,14.171056,12.730629,13.457702,14.733508,15.786391,16.568336,17.785841,18.231688,19.281141,19.901896,19.45262,17.686382,14.839825,13.485138,13.152468,13.430264,13.954991,13.166186,11.859513,11.47197,12.247057,13.231348,13.88297,13.29994,12.096155,10.751757,9.623423,8.868914,9.112414,9.997248,10.861504,10.717461,11.434244,11.331357,10.868362,10.545981,10.916377,10.456812,10.532263,10.347065,9.6645775,8.803751,9.054111,8.597976,8.508806,8.899779,8.923786,8.124693,8.176137,8.40249,8.604835,9.047252,9.455373,9.595985,9.489669,9.431366,9.9869585,10.069269,9.626852,8.9100685,8.289313,8.2310095,8.707723,7.9772205,7.407909,7.3598948,7.164408,7.0032177,6.6293926,6.7357097,7.431916,8.2481575,10.347065,11.739478,12.319078,12.085866,11.159878,0.42869842,0.39783216,0.53158605,0.7888051,1.0357354,1.039165,0.99801,1.0014396,0.96714365,0.89855194,0.8711152,0.9774324,0.96371406,0.89855194,0.84367853,0.85396725,0.8471081,0.805953,0.7476501,0.7133542,0.7613684,0.6790583,0.67219913,0.70649505,0.7305021,0.6824879,0.6241849,0.70306545,0.805953,0.86082643,0.83338976,0.8128122,0.82996017,0.9362774,1.0906088,1.1351935,1.1489118,1.097468,1.1454822,1.3032433,1.4164196,1.6187652,1.7525192,1.9548649,2.1743584,2.1846473,2.9220085,3.724532,4.8734436,6.4304767,8.241299,7.64798,9.822338,11.334786,12.46998,17.237106,29.453297,27.395544,17.36057,6.341307,2.0303159,1.5330256,1.1317638,1.0254467,1.2312219,1.5673214,1.3684053,1.0768905,0.9328478,0.97057325,1.0323058,1.1489118,1.2586586,1.1832076,0.9945804,1.0048691,0.922559,0.6379033,0.37382504,0.2469303,0.29151493,0.4938606,0.52472687,0.432128,0.40126175,0.7510797,1.2689474,1.1729189,0.7990939,0.48357183,0.5796003,0.64476246,0.85739684,0.96371406,0.8711152,0.65162164,0.64819205,0.59331864,0.4664239,0.3018037,0.1920569,0.20577525,0.20920484,0.15090185,0.0548734,0.024007112,0.020577524,0.058302987,0.08916927,0.12003556,0.18862732,0.15090185,0.1371835,0.12689474,0.12003556,0.10288762,0.432128,1.5741806,2.2841053,2.4247184,2.9734523,3.2272418,2.6579304,1.978872,1.5090185,1.1694894,1.0940384,1.2517995,1.1900668,1.0254467,1.4472859,2.0303159,1.8554068,1.6084765,1.4781522,1.138623,0.7613684,0.88826317,0.9431366,0.881404,1.1797781,0.96714365,0.91227025,0.980862,1.0563129,0.9431366,1.0323058,0.96371406,1.1214751,1.4267083,1.3272504,1.2517995,1.1900668,1.0837497,0.9328478,0.7888051,0.90198153,0.91227025,0.89512235,0.8711152,0.84024894,0.7407909,0.7476501,0.7888051,0.83338976,0.88826317,0.7579388,0.6962063,0.64476246,0.58302987,0.5418748,0.548734,0.6379033,0.82996017,1.0151579,0.96714365,0.7099246,0.881404,0.922559,0.805953,1.039165,1.1660597,0.96714365,0.94656616,1.0425946,0.65162164,0.8745448,0.6790583,0.5624523,0.61046654,0.50757897,0.50757897,0.5555932,0.66876954,0.8162418,0.90198153,0.805953,0.9294182,1.0425946,0.9945804,0.7305021,1.08032,1.2072148,1.3992717,1.6564908,1.6976458,1.5433143,1.605047,1.5707511,1.3546871,1.1043272,1.5604624,2.4384367,3.3884325,4.1017866,4.32471,3.4535947,3.4844608,4.125794,4.852866,4.9214582,5.3878818,5.4016004,5.6142344,6.2075534,6.910619,7.5725293,8.196714,8.275595,6.917478,2.8122618,2.8465576,3.683377,4.623084,5.5662203,6.999788,7.226141,6.9380555,6.8797526,7.284444,7.874333,9.438225,10.281903,10.621432,10.6488695,10.511685,10.0041065,9.630281,9.23245,8.988949,9.39021,9.616563,9.692014,9.523964,9.067829,8.320179,7.98408,8.244728,8.803751,9.355915,9.571979,9.1981535,9.06097,9.054111,9.0644,8.964942,9.012956,9.301042,9.822338,10.405369,10.72775,11.2421875,11.533703,11.965831,12.596875,13.183334,13.982429,14.706071,15.638919,16.561478,16.756964,17.082775,16.938732,15.902997,14.411126,13.742357,17.405157,22.741594,23.513252,19.37031,15.858413,21.650986,18.989626,11.924676,4.664239,1.546744,0.97057325,1.1283343,1.3203912,1.1660597,0.5727411,0.607037,0.6927767,0.7579388,0.8196714,0.9774324,1.1694894,1.2620882,1.4953002,2.301253,4.32471,3.3026927,3.5153272,3.875434,3.8857226,3.625074,4.139512,5.785714,7.507367,8.940934,10.432805,13.63604,13.402828,13.649758,14.781522,13.687484,9.644,5.4941993,2.784825,1.7113642,1.1249046,0.5521636,0.25378948,0.13032432,0.1097468,0.15090185,0.31552204,0.53158605,0.8265306,1.6667795,3.957744,5.778855,5.6313825,4.6436615,3.6456516,3.1655092,3.875434,2.7916842,1.6942163,1.4541451,2.0646117,2.3149714,2.702515,2.5996273,2.3801336,3.415869,3.2306714,4.0194764,4.73969,5.0003386,5.051782,5.192395,5.3330083,5.669108,6.169828,6.5779486,6.5779486,6.2658563,7.016936,7.9189177,5.7479887,3.309552,2.0577524,1.4815818,1.2106444,1.0254467,1.4027013,1.4404267,1.4678634,1.7250825,2.3424082,3.07634,4.081209,4.3521466,3.782835,3.1517909,2.4041407,1.8588364,1.4610043,1.1729189,0.94656616,0.85396725,0.9774324,0.65848076,0.0274367,0.010288762,0.0034295875,0.0,0.0,0.024007112,0.12689474,0.39440256,0.39097297,0.24007112,0.082310095,0.072021335,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.09602845,0.2194936,0.4355576,0.764798,0.53844523,0.9259886,1.0734608,0.922559,1.2037852,1.3101025,1.5673214,2.085189,2.8911421,3.9303071,3.9851806,4.448175,5.3330083,6.6122446,8.22758,8.213862,9.335337,10.127572,10.484249,11.650309,11.842365,12.271064,13.083877,14.112752,14.88098,14.445422,15.433144,16.674654,17.37429,17.137648,16.901007,16.026463,16.21166,17.367432,17.61779,19.497204,21.53438,23.808197,25.999702,27.381826,26.18833,25.814505,26.418112,27.642475,28.626766,29.607628,30.643364,31.809423,33.122955,34.539375,35.455074,33.829453,31.994621,30.783978,29.542467,28.932,28.054026,26.980564,26.641035,28.815393,29.539038,29.888855,29.367558,27.916842,25.917393,26.8571,25.663603,25.546997,26.315224,24.37065,16.695232,10.532263,8.604835,11.447963,17.405157,9.575408,9.441654,11.362224,12.905538,14.843254,13.481709,13.176475,13.903547,15.103903,15.680074,14.339106,11.712041,9.095266,7.8777623,9.55826,12.926115,14.057879,15.758954,18.173384,18.79757,17.436022,17.830425,18.30028,18.516342,19.510923,16.925014,13.426835,12.80608,14.4145565,13.1421795,15.038741,14.150477,12.9707,12.504276,12.295071,11.958971,12.22648,13.1421795,14.21564,14.4145565,13.594885,12.092726,11.187314,11.4754,12.867812,14.030442,15.409137,16.04018,15.923574,16.002455,16.245956,16.434584,16.732958,17.055338,17.055338,17.343424,17.343424,16.815268,16.239098,16.828985,18.015623,18.451181,19.215979,20.649546,22.36434,22.196291,22.117409,22.484375,23.61957,25.817934,27.721355,28.887415,28.719366,26.990854,23.852781,23.256033,22.069395,21.476076,21.657845,21.767591,20.12139,19.099373,19.654966,21.431492,22.77589,23.647005,24.058556,23.818485,22.834194,21.11597,19.9602,18.547209,17.504614,16.925014,16.359133,17.21653,17.436022,16.427725,14.980438,15.251375,15.066177,14.500296,13.80066,13.5503,14.675205,15.920145,16.520323,16.012743,14.644339,13.38911,13.749216,14.568888,15.680074,16.756964,17.29884,16.79126,17.806417,18.756414,18.718689,17.425734,15.505165,14.544881,14.171056,14.009865,13.660047,12.435684,11.842365,11.862943,12.199042,12.264205,11.187314,11.578287,11.784062,11.063849,9.585697,9.239308,9.448513,10.350495,11.286773,10.796341,10.600855,10.419086,10.30591,10.443094,11.129011,10.63858,10.429376,10.031544,9.349055,8.656279,9.174147,8.553391,8.272165,8.748878,9.349055,8.577398,8.495089,8.594546,8.772884,9.325048,9.3936405,9.626852,9.72288,9.661148,9.72631,9.705732,9.623423,9.253027,8.663138,8.207003,8.412778,8.261876,8.049242,7.8777623,7.6857057,7.5519514,7.2295704,7.1369715,7.5862474,8.820899,11.492548,13.279363,13.756075,12.843805,10.813489,0.48357183,0.4424168,0.58302987,0.7682276,0.922559,1.0117283,1.0323058,1.0117283,0.9877212,0.97057325,0.9294182,1.0117283,0.96714365,0.86082643,0.764798,0.7510797,0.66876954,0.67219913,0.7099246,0.7407909,0.72364295,0.6962063,0.6927767,0.72364295,0.7579388,0.72707254,0.6824879,0.77508676,0.8676856,0.90884066,0.91227025,0.90884066,0.91912943,1.0357354,1.1934965,1.1900668,1.3032433,1.2998136,1.3478279,1.4747226,1.5673214,1.6530612,1.8485477,2.020027,2.1400626,2.287535,3.100347,3.875434,5.394741,7.349606,8.364764,9.191295,10.645439,11.516555,13.673765,22.059107,28.503302,24.789059,15.395418,5.844017,2.719663,1.6530612,1.08032,0.97400284,1.1729189,1.4027013,1.1317638,0.9259886,0.9259886,1.097468,1.2209331,1.2483698,1.2895249,1.1934965,1.0151579,1.0048691,0.89169276,0.6207553,0.36010668,0.22635277,0.2709374,0.44927597,0.4938606,0.4355576,0.42526886,0.72021335,1.3889829,1.2895249,0.84024894,0.4389872,0.4698535,0.5212973,0.61389613,0.72364295,0.823101,0.8745448,0.9328478,0.8025235,0.58988905,0.37725464,0.2469303,0.29494452,0.32581082,0.24350071,0.08916927,0.037725464,0.041155048,0.08916927,0.15433143,0.30866286,0.70306545,0.490431,0.3566771,0.29494452,0.25378948,0.15090185,0.6379033,1.9925903,2.8328393,3.0386145,3.758828,3.4878905,2.6373527,1.937717,1.6770682,1.7113642,1.4918705,1.704505,1.8348293,1.8142518,2.0337453,1.9754424,1.587899,1.3992717,1.4198492,1.138623,0.7407909,0.89855194,1.0151579,1.0220171,1.3512574,0.7305021,0.8093826,1.097468,1.2312219,0.9842916,1.2895249,1.1832076,1.1660597,1.2929544,1.1763484,1.255229,1.1866373,1.0220171,0.8025235,0.5693115,0.7682276,0.7922347,0.78194594,0.8128122,0.89512235,0.8505377,0.823101,0.805953,0.7956643,0.77165717,0.6344737,0.59331864,0.61046654,0.6173257,0.50757897,0.5418748,0.607037,0.72364295,0.7990939,0.6241849,0.64476246,0.7990939,0.764798,0.66191036,1.0460242,1.0357354,0.90541106,0.864256,0.881404,0.6927767,0.83338976,0.6927767,0.64819205,0.7373613,0.67219913,0.51100856,0.5693115,0.66191036,0.77508676,1.0871792,0.881404,0.9294182,0.99801,0.9842916,0.91227025,1.3478279,1.5124481,1.6873571,1.8485477,1.6907866,1.6427724,1.7422304,1.8416885,1.8279701,1.605047,1.8005334,2.4075704,3.3061223,4.2218223,4.722542,4.091498,3.8137012,4.184097,4.866585,4.90431,5.3398676,5.5422134,5.9228973,6.5230756,7.006647,8.056101,8.488229,8.124693,6.5470824,3.1072063,3.532475,4.57164,5.360445,6.012067,7.641121,7.5725293,7.2295704,7.380472,8.086967,8.704293,10.175586,10.864933,11.183885,11.269625,10.988399,10.39508,9.925226,9.647429,9.602845,9.81205,9.273604,9.369633,9.129561,8.385342,7.7714453,7.490219,7.7748747,8.182996,8.40249,8.275595,7.8949103,7.9429245,8.268735,8.591117,8.525954,8.783174,9.088407,9.47595,9.880642,10.103564,10.264755,10.573419,11.039842,11.732618,12.758065,13.238208,13.612033,14.359683,15.254805,15.364552,15.806969,15.481158,15.114192,15.155347,15.762384,20.426622,23.581844,20.94792,15.662926,18.293419,24.068846,18.735836,10.206452,3.6627994,1.546744,1.3169615,1.4644338,1.5090185,1.2106444,0.5624523,0.5555932,0.65505123,0.7579388,0.823101,0.86082643,1.1180456,1.3581166,1.6427724,2.3904223,4.372724,3.2478194,3.9337368,4.972902,5.267846,4.0846386,4.90431,7.5039372,9.156999,10.017825,13.118172,15.254805,13.975569,11.825217,9.640571,6.557371,3.799983,2.1126258,1.529596,1.5638919,1.2003556,0.8128122,0.4664239,0.2777966,0.22978236,0.1920569,0.28465575,0.34638834,0.39097297,0.6001778,1.2860953,0.9774324,0.9362774,1.6153357,2.49331,2.0714707,3.0111778,2.0714707,1.155771,0.96714365,0.9842916,1.5570327,1.6976458,1.4061309,1.1626302,1.920569,1.8108221,2.9494452,4.671098,6.0806584,6.0566516,5.562791,5.1992545,5.6485305,6.5985265,6.711703,6.619104,5.8988905,5.809721,6.2864337,5.950334,4.3692946,2.867135,1.9582944,1.6633499,1.5124481,2.0337453,2.054323,1.862266,1.8897027,2.6956558,3.2855449,3.981751,3.758828,2.719663,2.085189,1.8588364,1.587899,1.3512574,1.214074,1.2277923,1.3066728,1.3032433,0.8093826,0.072021335,0.010288762,0.0034295875,0.0,0.0,0.024007112,0.12689474,0.31209245,0.23664154,0.15776102,0.15090185,0.14061308,0.17833854,0.106317215,0.030866288,0.010288762,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.07888051,0.15776102,0.31895164,0.764798,0.59674823,0.8711152,0.96714365,0.85739684,1.1214751,1.0631721,1.3066728,1.8519772,2.6133456,3.4192986,3.5976372,3.7759757,4.2595477,5.2506986,6.835168,7.284444,8.375052,9.177576,9.695444,10.837497,11.327928,12.2093315,13.13532,13.992717,14.898128,14.181344,14.682064,15.700651,16.619781,16.907866,16.558048,16.396858,16.986746,18.152807,18.965618,21.548098,23.170294,24.826784,26.521,27.27208,26.246634,26.099161,26.716486,27.728214,28.51016,28.637054,29.388136,30.948597,32.82801,33.887753,34.024937,32.19011,30.622786,29.779108,28.3524,27.649334,27.17605,26.455837,26.332373,28.956007,30.10492,31.805994,32.16953,30.67423,28.17749,30.221525,26.812515,29.484163,35.461933,27.6802,18.238546,11.9040985,15.402277,21.013083,6.5642304,9.781183,10.782623,11.1393,12.089295,14.544881,13.88983,12.662037,12.243628,12.864383,13.581166,14.7026415,13.88983,11.893809,10.504827,12.535142,14.493437,14.654627,16.064188,18.852442,20.237995,20.718138,21.11597,20.793589,20.066517,20.21056,16.307688,11.910957,11.550851,14.249936,13.522863,14.63062,14.71636,14.788382,15.011304,14.688923,14.496866,14.393978,14.212211,14.05102,14.30481,13.179905,11.537132,11.084427,12.21962,14.044161,15.29253,16.45173,16.86671,16.901007,17.933313,18.71183,19.490345,19.552078,18.986197,18.71526,19.226267,18.842154,17.823566,17.12393,18.37573,18.61923,18.276272,18.557497,20.066517,22.796469,22.77589,22.230585,22.515242,23.911083,25.636166,27.121178,28.42785,28.75023,27.481285,24.212887,24.013971,22.576975,20.800447,19.45262,19.19197,17.806417,17.03819,17.919594,20.097382,21.829325,23.653864,24.494114,24.048267,22.494663,20.484926,19.44919,17.943602,16.496315,15.481158,15.107333,16.355703,17.024471,16.410576,15.326826,16.095055,15.786391,14.572317,13.361672,12.984418,14.181344,15.237658,15.87213,15.721229,15.035312,14.692352,15.001016,15.244516,15.549749,15.865272,15.944152,15.954441,17.103354,17.748116,17.408587,16.743246,16.20137,15.642348,15.107333,14.490007,13.543441,11.701753,11.427385,11.533703,11.334786,10.652299,9.22216,10.264755,11.794352,12.154458,10.031544,9.445084,9.73317,10.628291,11.321068,10.456812,9.482809,9.47938,9.788043,10.185875,10.89237,10.693454,10.398509,9.97324,9.414218,8.745448,8.80718,8.251588,8.049242,8.512236,9.294182,8.855195,8.601405,8.519095,8.673427,9.205012,9.22216,9.465661,9.688584,9.72288,9.513676,9.253027,9.47595,9.4862385,9.126132,8.772884,8.711152,8.865483,8.841476,8.570539,8.296172,8.23444,8.241299,8.484799,9.146709,10.415657,12.411677,13.745787,13.975569,12.984418,10.9541025,0.6207553,0.6001778,0.7373613,0.8676856,0.939707,1.039165,1.0631721,0.9877212,0.9774324,1.0528834,1.08032,1.1180456,1.0597426,0.94999576,0.84367853,0.8162418,0.70649505,0.7099246,0.75450927,0.78537554,0.764798,0.8196714,0.72707254,0.65848076,0.65848076,0.66191036,0.75450927,0.8745448,0.94999576,0.980862,1.039165,1.0563129,1.08032,1.1592005,1.2415106,1.2037852,1.3889829,1.4781522,1.471293,1.4610043,1.605047,1.6770682,1.9239986,2.054323,2.1229146,2.5447538,3.0626216,3.74168,5.826869,8.64942,9.609704,10.960961,10.494537,10.81006,14.71636,25.234905,26.10602,19.490345,11.032983,4.7945633,3.2375305,1.8519772,1.2415106,1.0631721,1.0734608,1.1283343,1.0768905,1.0700313,1.1832076,1.3443983,1.3375391,1.2175035,1.1043272,0.9945804,0.922559,0.9568549,0.8128122,0.58645946,0.36696586,0.23664154,0.26407823,0.29837412,0.39097297,0.45270553,0.5658819,0.9911508,1.5124481,1.2826657,0.78537554,0.36353627,0.1920569,0.25721905,0.34981793,0.4629943,0.6207553,0.8745448,1.0117283,0.8471081,0.61389613,0.42183927,0.28465575,0.3566771,0.39097297,0.29494452,0.12003556,0.0548734,0.0548734,0.06859175,0.14061308,0.39440256,1.0563129,0.7922347,0.61046654,0.5658819,0.607037,0.5761707,1.2483698,2.5138876,3.2855449,3.4467354,3.8479972,3.210094,2.4761622,1.8108221,1.4953002,1.9445761,1.8039631,1.8554068,2.2738166,2.5481834,1.4850113,1.4335675,1.5501735,1.5364552,1.3786942,1.3306799,0.8128122,1.0734608,1.1866373,1.0597426,1.4335675,1.0323058,0.9362774,1.0906088,1.3032433,1.2449403,1.4644338,1.3375391,1.2003556,1.1214751,0.89512235,1.1420527,1.0288762,0.8505377,0.72707254,0.6276145,0.6173257,0.64133286,0.7339317,0.84024894,0.8265306,1.1283343,1.0734608,0.8779744,0.7476501,0.8471081,0.8471081,0.6310441,0.6962063,0.9362774,0.61046654,0.6790583,0.66191036,0.7339317,0.84367853,0.70649505,0.6036074,0.6173257,0.5590228,0.4938606,0.764798,0.5521636,0.66876954,0.6824879,0.5590228,0.64819205,0.71678376,0.6859175,0.78537554,0.9294182,0.7305021,0.65505123,0.7613684,0.78194594,0.77508676,1.1489118,0.90198153,0.8128122,0.8711152,1.0220171,1.2003556,1.5913286,1.786815,1.8382589,1.7525192,1.5055889,1.6633499,1.6667795,1.8862731,2.2463799,2.253239,2.0680413,2.1023371,2.6236343,3.5461934,4.4104495,4.3624353,4.046913,4.170378,4.6608095,4.695105,4.852866,5.4324665,6.23499,7.0135064,7.449064,8.086967,7.9017696,7.010077,5.645101,4.1772375,5.2747054,6.2830043,6.540223,6.39961,7.226141,7.2707253,7.2535777,7.579388,8.158989,8.40249,9.530824,10.106995,10.484249,10.731179,10.621432,10.30934,10.1481495,10.364213,10.714031,10.460241,9.3593445,8.97523,8.405919,7.596536,7.346176,7.164408,7.459353,7.599966,7.31531,6.7048435,6.8557453,7.0923867,7.623973,8.268735,8.453933,8.838047,9.242738,9.47595,9.561689,9.746887,9.438225,9.668007,10.192734,11.050131,12.555719,12.929544,13.118172,13.560589,14.092175,13.9481325,15.014734,15.066177,15.529172,16.925014,18.866161,23.266321,25.241764,22.542679,18.62609,22.642136,23.914513,16.29054,8.134981,3.5118976,2.1640697,2.1674993,2.0989075,1.903421,1.4541451,0.5624523,0.45956472,0.5418748,0.6790583,0.77851635,0.7990939,1.0082988,1.3203912,1.6907866,2.1915064,3.0317552,2.6613598,4.033195,5.6313825,6.5196457,6.310441,7.1026754,9.530824,10.518545,11.4033785,17.95732,15.086755,10.55284,6.5813785,3.998899,2.253239,1.3272504,0.9431366,1.0563129,1.313532,1.0597426,0.922559,0.64476246,0.47328308,0.4355576,0.31895164,0.32924038,0.37039545,0.4046913,0.39783216,0.32238123,0.19891608,0.2194936,0.3566771,0.61046654,1.0357354,1.08032,1.0700313,1.0768905,1.039165,0.7476501,1.0563129,0.91227025,0.8093826,0.9602845,1.3032433,1.3992717,2.0097382,3.8788633,6.2864337,7.0752387,6.3310184,6.0154963,6.307011,6.9037595,7.0135064,7.0786686,6.447624,5.562791,4.979761,5.363875,5.271276,4.07435,3.100347,2.7951138,2.726522,2.8705647,2.651071,2.3972816,2.609916,3.9508848,4.338428,4.4859004,3.6765177,2.194936,1.3169615,0.94999576,0.922559,0.9568549,0.9602845,1.0494537,1.2346514,0.88826317,0.4355576,0.116605975,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.15090185,0.30866286,0.16119061,0.3566771,0.25378948,0.12689474,0.09945804,0.15090185,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.044584636,0.12346515,0.28122616,0.6036074,0.7613684,0.75450927,0.805953,0.9534253,1.0254467,0.89169276,1.2380811,1.7422304,2.253239,2.7745364,3.1415021,3.0626216,3.1586502,3.841138,5.295283,6.6465406,7.5759587,8.597976,9.794902,10.820349,11.30735,12.404818,13.29994,14.05102,15.601193,15.916716,15.772673,15.851553,16.55119,17.977898,17.075916,17.69667,18.303709,18.680964,19.94305,22.175713,23.674442,24.881657,25.793928,25.955118,26.579304,27.577312,28.105469,28.153484,28.565035,28.52731,28.791388,30.547335,32.817722,32.491913,31.363577,30.296976,29.974594,30.046616,29.120626,27.611609,27.409264,27.577312,28.393555,31.343,32.1661,33.60996,33.513927,31.91917,31.109787,33.49678,29.35384,36.41536,47.45863,30.290117,18.886738,14.438563,22.44665,30.029469,5.895461,10.175586,7.922347,6.917478,9.431366,12.195613,12.435684,11.598865,10.532263,10.127572,11.30049,12.363663,12.6929035,13.149038,14.0750265,15.285671,14.38026,15.769243,18.11165,20.179693,20.855322,20.176264,21.184563,20.899906,18.70154,16.321407,13.066729,10.899229,10.782623,12.0138445,12.233338,13.96185,15.179354,15.683503,15.8138275,16.45173,15.553179,14.5414505,13.622321,13.042721,13.070158,11.38623,10.652299,11.38966,13.1593275,14.582606,15.261664,16.235666,16.945591,17.597214,19.161106,20.19341,21.37319,21.102251,19.576086,18.787281,19.342873,18.95533,18.828436,19.589804,21.287449,20.189981,19.19197,18.948471,19.802439,21.77445,22.799898,23.496103,24.161444,24.69303,24.583282,24.744474,25.10115,25.584723,25.461258,23.321196,22.61127,21.764162,19.648108,16.942162,16.143068,15.827546,15.659496,16.311117,17.727537,19.11995,21.414345,22.453508,22.2786,21.11597,19.384027,18.9519,17.717249,16.54433,15.995596,16.324837,16.393429,15.906426,15.12448,14.668345,15.536031,15.371411,14.352823,13.258785,12.860953,13.9138365,14.339106,15.059319,15.477728,15.614912,16.13621,16.719238,15.916716,14.448852,13.313659,13.814379,15.3302555,16.585485,16.513464,15.590904,15.820687,16.314548,15.995596,15.498305,14.778092,13.094165,11.032983,10.635151,10.669447,10.374502,9.445084,9.119273,10.028113,11.852654,13.004995,10.618003,9.448513,10.000677,10.882081,11.074138,9.928656,8.793462,8.999237,9.493098,9.860064,10.316199,10.425946,10.429376,10.230459,9.753747,8.954653,8.320179,7.98065,7.9875093,8.30646,8.81061,8.721441,8.440215,8.292743,8.39563,8.666568,8.927217,9.098696,9.31133,9.496528,9.403929,9.098696,9.400499,9.554831,9.451943,9.616563,9.469091,9.400499,9.355915,9.205012,8.759167,9.006097,9.4862385,10.213311,11.0981455,11.945253,12.63803,12.79922,12.644889,12.199042,11.290202,0.65505123,0.65505123,0.7099246,0.764798,0.78194594,0.7339317,0.8162418,0.85739684,0.9294182,1.0323058,1.0666018,1.0666018,1.0597426,1.0117283,0.9534253,0.9774324,0.85396725,0.7613684,0.71678376,0.71678376,0.71678376,0.7407909,0.7373613,0.77508676,0.8711152,0.9911508,1.0151579,1.0220171,1.0117283,1.0151579,1.1146159,1.0906088,1.1214751,1.2620882,1.3992717,1.2517995,1.4953002,1.4747226,1.4061309,1.4472859,1.6770682,1.6907866,1.786815,1.7490896,1.8485477,2.8396983,2.7402403,3.6696587,6.358455,9.427936,9.352485,11.952112,10.926665,11.283342,14.870691,20.402617,17.569777,10.792912,5.086078,2.3458378,1.3581166,1.2106444,1.1489118,1.039165,0.94656616,1.1283343,1.2517995,1.4267083,1.5090185,1.4335675,1.2517995,1.0940384,0.9602845,0.90198153,0.9328478,1.0666018,0.8848336,0.6207553,0.42526886,0.31209245,0.15090185,0.09259886,0.12346515,0.23321195,0.490431,1.0528834,1.5055889,1.3889829,1.039165,0.6927767,0.47328308,0.36353627,0.30866286,0.28465575,0.31552204,0.47328308,0.65505123,0.6001778,0.48014224,0.3806842,0.31895164,0.29494452,0.22635277,0.15776102,0.116605975,0.09259886,0.041155048,0.030866288,0.037725464,0.0548734,0.09259886,0.3841138,0.5761707,0.864256,1.3581166,2.0920484,2.4212887,2.4212887,2.49331,2.5790498,2.1503513,1.9823016,1.7182233,1.5090185,1.430138,1.4815818,1.5055889,1.5844694,1.8691251,1.9514352,0.84024894,1.646202,1.2517995,1.0734608,1.4027013,1.4027013,0.8162418,1.1489118,1.1043272,0.77508676,1.6187652,1.08032,1.1763484,1.3821237,1.488441,1.587899,1.1214751,0.980862,0.9294182,0.881404,0.8711152,1.0768905,0.8162418,0.77508676,0.9842916,0.823101,0.77508676,0.8162418,0.78194594,0.8025235,1.3272504,1.5227368,1.5638919,1.3786942,1.1283343,1.1900668,0.7990939,0.6379033,0.75450927,0.9774324,0.91569984,0.91569984,0.88826317,0.881404,0.85396725,0.67219913,0.6824879,0.5693115,0.53158605,0.59674823,0.59674823,0.51100856,0.52472687,0.47671264,0.41498008,0.61046654,0.85396725,0.7956643,0.94999576,1.2655178,1.1454822,1.1077567,1.1523414,1.1523414,1.0631721,0.91569984,1.0014396,1.1489118,1.3341095,1.3821237,0.9911508,1.2346514,1.4987297,1.4815818,1.2483698,1.2346514,1.3958421,1.7730967,2.0063086,2.0440342,2.1674993,1.7765263,1.4953002,1.7936742,2.6407824,3.4947495,3.8377085,3.8857226,4.245829,4.8768735,5.096367,4.962613,5.9434752,6.6705475,6.9620624,7.8263187,8.4264965,8.40249,7.3255987,6.046363,6.667118,7.4627824,8.299602,8.344186,7.6788464,7.3255987,6.715132,6.6431108,6.6122446,6.5813785,6.9723516,7.6342616,7.881192,8.453933,9.22902,9.2153015,9.362774,10.086417,10.690024,10.827208,10.497967,9.911508,9.297611,8.601405,7.966932,7.7371492,6.931196,6.893471,6.931196,6.776865,6.6053853,7.1678376,7.380472,7.7920227,8.429926,8.820899,8.97866,9.211872,9.325048,9.489669,10.2236,10.089847,9.945804,10.086417,10.786053,12.298501,13.251926,13.334236,13.63261,14.140189,13.762935,15.789821,15.803539,16.163645,17.487467,18.646667,21.894485,26.641035,26.733635,22.971376,23.11542,19.905325,12.247057,6.2212715,3.8960114,3.309552,3.1415021,2.784825,2.3389788,1.7216529,0.67219913,0.5007198,0.4938606,0.51100856,0.50757897,0.5178677,0.6893471,1.08032,1.605047,2.2738166,3.1895163,3.7382503,3.940596,4.8117113,6.5779486,8.666568,10.278474,9.866923,9.184435,9.716022,12.696333,10.545981,6.468202,3.1277838,1.5433143,1.0666018,1.0323058,1.0666018,1.1420527,1.1797781,1.0837497,0.84024894,0.65848076,0.5693115,0.53844523,0.48700142,0.35324752,0.36696586,0.39097297,0.34638834,0.21263443,0.17833854,0.28808534,0.34638834,0.38754338,0.65505123,0.7888051,0.9259886,0.91227025,0.77165717,0.6859175,0.6756287,0.83681935,0.9534253,0.88826317,0.59674823,0.4972902,0.6927767,1.039165,1.8005334,3.6319332,5.439326,5.6348124,5.212973,5.0586414,5.950334,6.7700057,6.2967224,5.360445,5.1580997,7.233,6.169828,6.060081,5.802862,5.0449233,4.166949,3.724532,3.3129816,3.2958336,4.1463714,6.4544835,7.7611566,7.0889573,4.8254294,2.0749004,0.67219913,0.48700142,0.881404,1.138623,1.0014396,0.67219913,0.72021335,0.48357183,0.24007112,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07888051,0.18519773,0.1371835,0.1371835,0.2194936,0.34295875,0.4046913,0.26064864,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06859175,0.15090185,0.28808534,0.5796003,0.4938606,0.6276145,0.8676856,0.9877212,0.67219913,0.7339317,1.0666018,1.5193073,1.9445761,2.2120838,2.201795,2.4624438,2.702515,3.0866287,4.256118,5.9297566,7.4113383,8.344186,9.15014,11.015835,11.979549,13.193623,13.852104,14.476289,16.907866,17.175373,16.19794,15.88242,16.660936,17.501184,17.576635,18.903887,20.227707,21.054237,21.650986,22.079683,23.650434,25.001692,25.368658,24.61415,25.979126,28.006012,29.367558,30.18723,32.042637,32.056355,32.478195,32.797146,32.16267,29.405283,29.624777,30.876575,34.57024,38.92582,38.98412,36.898933,34.765728,33.09895,32.78343,35.08125,34.347317,35.719154,37.132145,37.99297,39.2139,39.628883,35.07439,39.84152,47.417477,30.485603,16.434584,9.537683,12.771784,18.386019,7.874333,11.399949,7.6685576,6.1972647,9.253027,11.842365,10.364213,11.101575,11.266195,10.703742,11.8869505,14.4145565,15.364552,16.383139,17.545769,17.350283,14.140189,21.997374,27.042297,25.128588,21.819035,19.342873,20.62554,22.432932,22.326614,18.677534,10.216741,14.006435,15.446862,11.784062,12.099585,13.015285,13.4474125,13.629181,13.838386,14.390549,14.438563,13.471419,12.816368,12.4974165,11.214751,9.873782,9.993818,11.207891,12.737488,13.395968,14.654627,15.755525,16.324837,16.585485,17.38115,18.770132,19.5315,19.37374,18.434032,17.271402,16.492886,17.147938,18.807858,20.406046,20.248285,19.895037,19.219408,18.663815,18.821575,20.430052,22.823904,24.593573,25.4544,25.303495,24.216316,24.007113,22.594122,21.860191,22.11398,22.065966,21.980227,21.143406,19.836735,18.36544,17.058767,16.595774,15.196502,14.5585985,15.028452,15.638919,17.446312,18.475187,18.646667,18.139088,17.394867,17.480608,17.171944,16.80155,16.835844,17.899017,17.021042,15.46401,14.157337,13.584596,13.780083,14.5243025,15.570327,15.642348,14.915276,15.001016,14.486577,14.805529,15.107333,15.145059,15.306249,15.87899,13.155897,10.251037,9.482809,12.373952,13.461131,13.972139,13.591455,13.22106,14.953001,15.673215,15.971589,16.204802,15.415996,11.338216,10.007536,9.856634,10.034973,9.983529,9.445084,9.078118,9.2153015,10.679735,12.449403,11.64345,10.484249,10.789482,11.286773,11.0981455,9.719451,8.793462,8.98209,9.616563,10.034973,9.582268,9.9869585,10.343636,10.2921915,9.760606,8.940934,8.320179,7.805741,7.764586,8.114404,8.347616,8.237869,8.172707,8.069819,8.008087,8.241299,8.4093485,8.663138,9.06097,9.414218,9.294182,9.4862385,9.692014,9.661148,9.578837,10.055551,9.959522,9.668007,9.582268,9.661148,9.431366,10.124143,10.63858,10.88894,11.039842,11.506266,11.993267,11.245617,10.933525,11.255906,10.926665,0.864256,0.980862,0.96371406,0.9842916,1.0597426,1.0494537,1.1043272,1.08032,1.0940384,1.1592005,1.1660597,1.0871792,1.1111864,1.155771,1.155771,1.0734608,1.0014396,0.9328478,0.89512235,0.8848336,0.864256,0.8779744,0.94656616,1.0082988,1.0254467,0.9911508,0.9877212,1.0425946,1.08032,1.0906088,1.138623,1.2003556,1.2826657,1.3066728,1.3238207,1.5193073,1.3238207,1.2826657,1.3615463,1.4404267,1.2998136,1.4404267,1.6839274,1.7696671,1.9651536,3.083199,3.1895163,4.7602673,7.56224,10.360784,10.9541025,17.106783,16.671225,13.591455,10.947243,10.930096,8.954653,5.5730796,2.8225505,1.4541451,0.89512235,0.8162418,0.78537554,0.8779744,1.1317638,1.5193073,1.5536032,1.5330256,1.4987297,1.4472859,1.313532,1.1146159,1.155771,1.196926,1.1729189,1.1900668,0.94999576,0.7407909,0.61046654,0.4938606,0.23664154,0.1371835,0.12346515,0.14061308,0.25378948,0.65162164,1.3272504,1.4781522,1.2620882,0.90884066,0.7305021,0.6207553,0.47671264,0.39440256,0.4081209,0.51100856,0.61389613,0.66533995,0.64476246,0.58302987,0.5521636,0.53844523,0.48357183,0.34981793,0.17147937,0.07888051,0.06859175,0.06859175,0.058302987,0.048014224,0.0548734,0.12346515,0.16462019,0.2469303,0.44584638,0.85739684,0.6893471,0.77851635,0.939707,1.1146159,1.371835,1.1489118,1.0288762,1.0597426,1.2243627,1.4198492,1.5981878,1.6153357,1.9137098,2.2155135,1.5364552,1.587899,1.5570327,1.7696671,1.9102802,1.0117283,1.0906088,1.0460242,1.1866373,1.4987297,1.6187652,1.196926,1.2346514,1.3101025,1.2483698,1.1214751,0.89512235,1.0151579,1.2758065,1.3066728,0.5521636,1.1592005,1.1900668,1.2072148,1.255229,0.86082643,1.0082988,1.2586586,1.4678634,1.4507155,1.0117283,1.1180456,1.1351935,1.1729189,1.1592005,0.86082643,0.8711152,0.8745448,0.7990939,0.7339317,0.91569984,1.08032,0.72364295,0.45613512,0.51100856,0.72021335,0.5178677,0.3841138,0.39097297,0.5178677,0.64476246,0.5796003,0.6207553,0.70649505,0.78537554,0.7922347,0.823101,0.78537554,0.97057325,1.3375391,1.4987297,1.3341095,1.6256244,1.5981878,1.2209331,1.2209331,1.4027013,1.1180456,1.1249046,1.3478279,0.8711152,1.2517995,1.371835,1.3684053,1.3375391,1.3341095,1.7182233,1.9754424,1.9685832,1.8554068,2.0920484,2.0234566,1.9582944,2.2120838,2.8156912,3.4947495,4.108646,4.461893,4.835718,5.3673043,6.036074,6.3790326,6.9037595,6.9723516,6.90033,7.963502,8.100685,9.242738,11.705182,12.761495,6.6568294,5.8680243,6.444195,6.7391396,6.3207297,5.9571934,6.1458206,6.5059276,6.56766,6.293293,6.0703697,6.7665763,7.39762,8.320179,9.095266,8.508806,9.513676,9.784613,9.990388,10.31277,10.460241,10.30591,9.8429165,9.177576,8.515666,8.176137,7.9086285,7.720001,7.442205,7.2535777,7.6685576,8.162418,7.7577267,7.8023114,8.429926,8.587687,8.940934,9.544542,9.935514,10.172156,10.844356,10.251037,10.542552,11.156448,11.797781,12.432255,12.915827,13.262215,14.102464,15.076467,14.826107,16.657507,15.323397,16.071047,19.421753,21.184563,27.52587,30.670801,27.786518,20.906765,16.904436,14.994157,9.89093,5.7822843,4.190956,3.9954693,3.7553983,3.4947495,2.9563043,2.1057668,1.1214751,0.7373613,0.58988905,0.5453044,0.52472687,0.50757897,0.70649505,1.0254467,1.5090185,2.2429502,3.3369887,3.0351849,3.07634,4.2595477,5.9228973,5.919468,7.599966,8.251588,11.842365,15.837835,11.231899,6.5024977,3.4638834,1.6873571,1.097468,1.9582944,1.3169615,0.9602845,0.8093826,0.7682276,0.7305021,0.59331864,0.58645946,0.53844523,0.4629943,0.548734,0.33609957,0.26407823,0.25378948,0.31209245,0.53158605,0.39783216,0.34295875,0.30523327,0.2709374,0.26407823,0.3806842,0.6276145,0.823101,0.8779744,0.77165717,0.7510797,1.1866373,1.5021594,1.5638919,1.6804979,2.2669573,1.9685832,2.2360911,3.5187566,5.2438393,6.7459984,8.124693,9.856634,11.194174,10.161868,8.001227,7.0546613,6.7357097,6.8111606,7.4044795,6.3790326,6.0154963,5.7102633,5.267846,4.897451,4.341858,4.5682106,5.518206,7.1541195,9.431366,10.97468,9.136421,5.9743414,2.952875,0.9534253,0.37725464,0.45613512,0.84367853,1.214074,1.2449403,0.6790583,0.274367,0.06859175,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.037725464,0.0274367,0.0274367,0.10288762,0.12689474,0.082310095,0.05144381,0.010288762,0.072021335,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.0274367,0.058302987,0.13032432,0.28808534,0.5144381,0.881404,1.0117283,0.8779744,0.7922347,0.922559,1.1729189,1.4541451,1.7422304,2.0920484,2.3218307,2.726522,3.0900583,3.4604537,4.122364,5.178677,6.3447366,7.8263187,9.427936,10.55284,12.641459,13.906977,14.832966,15.71437,16.650646,16.87014,16.050468,16.016174,17.079346,18.03963,18.571217,19.53836,20.21399,20.673553,21.798458,21.4555,22.679861,23.821915,24.487255,25.51613,26.863958,28.637054,29.854559,30.797695,32.99606,34.776016,37.5094,38.792065,38.171307,37.128716,35.26988,34.99208,38.06499,42.351974,41.81696,41.868404,41.14133,40.050724,39.265347,39.707764,38.884663,39.24134,39.59802,39.72834,40.362816,43.922726,48.295452,51.62215,48.528664,30.132355,15.086755,12.003556,15.3302555,18.056778,11.705182,11.026124,8.8929205,8.98209,10.4533825,7.936065,5.7068334,6.989499,7.720001,7.56224,9.897789,11.05699,11.434244,13.481709,15.87899,13.516005,21.417774,23.478956,23.60585,22.94737,19.905325,19.682402,19.421753,20.11796,20.601532,17.518333,12.542002,11.667457,10.9369545,9.73317,10.782623,10.261326,10.158438,10.618003,11.393089,11.825217,11.30735,11.070708,10.8958,10.679735,10.432805,10.799771,11.231899,11.718901,12.363663,13.38568,14.7026415,16.45516,17.977898,18.948471,19.37031,20.378609,20.186552,18.931322,17.161655,15.844694,16.70552,17.470318,18.694681,19.70641,18.602083,18.804428,18.310568,18.44432,19.071936,18.612371,19.932762,21.688711,23.256033,23.749893,22.017952,21.28402,20.382038,19.54179,18.722118,17.607502,17.484037,17.597214,17.322845,16.263103,14.263655,14.081886,13.876111,13.972139,14.46943,15.223939,15.920145,16.595774,17.20624,17.837284,18.71183,17.508043,16.849564,16.606062,16.575195,16.496315,15.937293,15.062748,14.46943,14.4317045,14.901558,15.148488,16.12249,16.194511,15.13134,14.085316,13.406258,13.516005,13.965281,14.29452,14.023583,13.814379,12.531713,10.851214,10.028113,11.8869505,11.616013,12.123591,13.594885,15.45715,16.369421,16.798119,16.911295,15.954441,13.917266,11.55771,10.597425,10.912948,11.262765,11.331357,11.739478,11.499407,10.672876,10.878652,11.931535,11.838936,10.511685,10.079557,10.072699,10.124143,9.97667,9.448513,9.716022,10.14129,10.419086,10.569988,10.329918,10.38479,10.446524,10.161868,9.15014,8.193284,7.8777623,7.747438,7.7097125,8.028665,8.220721,8.06639,7.857185,7.874333,8.351046,8.7145815,8.848335,8.889491,8.971801,9.218731,9.1810055,9.040393,9.146709,9.602845,10.275044,9.757176,9.97667,10.381361,10.587136,10.39508,10.532263,10.789482,10.923236,10.991828,11.358793,11.592006,11.382801,11.47197,11.4205265,9.606275,0.6241849,0.7407909,0.7613684,0.8093826,0.90884066,0.9842916,1.0597426,1.08032,1.0666018,1.0220171,0.9328478,0.8711152,0.90198153,0.9877212,1.0768905,1.097468,1.138623,1.0940384,1.0597426,1.0734608,1.1008976,1.0700313,1.1008976,1.1454822,1.1626302,1.1214751,1.138623,1.2243627,1.3101025,1.3546871,1.3443983,1.4232788,1.4335675,1.3752645,1.3101025,1.3581166,1.2792361,1.2723769,1.2860953,1.2449403,1.0494537,1.3306799,1.5227368,1.6770682,2.095478,3.3438478,3.525616,5.8234396,8.961512,12.22648,15.481158,23.321196,21.050808,14.006435,7.2947326,5.796003,5.079219,3.5221863,2.0474637,1.1763484,1.0151579,1.2175035,1.3546871,1.3821237,1.3752645,1.4987297,1.4438564,1.3649758,1.255229,1.2312219,1.5090185,1.4198492,1.3546871,1.255229,1.1694894,1.2312219,1.0323058,0.78194594,0.64133286,0.61389613,0.5624523,0.37725464,0.24350071,0.16462019,0.20577525,0.48357183,0.9534253,1.155771,1.1351935,0.9945804,0.91227025,0.64819205,0.41840968,0.31552204,0.35324752,0.44584638,0.45613512,0.4938606,0.61389613,0.8025235,0.9774324,0.85396725,1.0185875,0.8779744,0.4081209,0.15776102,0.13032432,0.106317215,0.07888051,0.05144381,0.037725464,0.048014224,0.05144381,0.06859175,0.12689474,0.26407823,0.15433143,0.274367,0.3806842,0.4424168,0.6344737,0.83338976,0.72021335,0.9842916,1.4507155,1.0837497,1.4438564,1.6736387,1.961724,2.1915064,1.9548649,1.8073926,1.670209,1.6942163,1.762808,1.4747226,1.4335675,1.4953002,1.7147937,1.8965619,1.6187652,1.2483698,1.2106444,1.1592005,0.9602845,0.66876954,0.77508676,0.9259886,1.0700313,1.0151579,0.42869842,1.1729189,1.2449403,1.3478279,1.488441,1.0082988,1.0425946,1.0871792,1.2037852,1.255229,0.89512235,1.097468,1.1111864,1.0425946,0.99801,1.0906088,0.9877212,1.0666018,0.96714365,0.7305021,0.805953,0.6756287,0.53501564,0.48357183,0.52815646,0.58645946,0.44584638,0.4046913,0.41840968,0.5041494,0.7305021,0.53501564,0.6173257,0.69963586,0.6893471,0.6824879,0.7476501,0.70649505,0.90198153,1.2655178,1.3306799,1.2895249,1.6633499,1.7422304,1.4575747,1.4061309,1.4987297,1.4678634,1.529596,1.5947582,1.2792361,1.255229,1.2895249,1.4027013,1.5673214,1.704505,1.5673214,1.821111,2.061182,2.1297739,2.1194851,2.5721905,2.9700227,2.9631636,2.8534167,3.566771,4.2938433,4.7979927,5.2609873,5.754848,6.23499,6.5813785,6.8283086,6.6396813,6.4098988,7.2638664,7.205563,9.081548,11.705182,12.778643,8.89635,4.729401,4.846007,5.528495,5.4736214,5.7891436,6.7802944,6.9723516,6.8591747,6.6431108,6.217842,7.431916,8.241299,8.964942,9.386781,8.735159,9.31133,9.702303,9.863494,9.774324,9.472521,9.239308,8.995808,8.484799,7.922347,8.001227,8.182996,8.385342,8.2310095,7.9463544,8.381912,8.601405,8.128122,8.032094,8.354475,8.107545,9.191295,9.788043,9.97324,10.034973,10.497967,10.172156,10.518545,11.327928,12.322508,13.162757,13.207341,13.605173,14.534592,15.433144,14.96329,16.561478,16.592344,18.79071,22.26831,21.527521,29.655643,33.157253,28.136335,18.056778,13.749216,13.070158,10.038403,6.495639,4.0606318,4.139512,4.290414,4.249259,3.6559403,2.6476414,1.8691251,1.3546871,1.0425946,0.8848336,0.8093826,0.7407909,0.84024894,1.1111864,1.5913286,2.1880767,2.6853669,2.452155,2.4761622,3.8137012,5.7651367,5.892031,6.944915,6.012067,8.371623,12.260776,8.868914,4.105216,2.0028791,1.3649758,1.4027013,1.7422304,1.2655178,0.94999576,0.86082643,0.8745448,0.65848076,0.53501564,0.53501564,0.5007198,0.4115505,0.3806842,0.2503599,0.26064864,0.2777966,0.30866286,0.48357183,0.4629943,0.42526886,0.41840968,0.4355576,0.4046913,0.47328308,0.78537554,1.2723769,1.7010754,1.6736387,1.978872,2.170929,2.277246,2.3801336,2.620205,3.1963756,3.7519686,5.4941993,8.080108,9.637141,12.003556,12.127021,12.435684,13.399398,13.540011,11.1393,9.0644,8.268735,8.423067,7.905199,6.9723516,5.960623,4.931747,4.0537724,3.5873485,3.3678548,3.82399,5.0312047,6.8626046,8.97866,8.827758,6.9209075,4.6402316,2.6236343,0.78537554,0.48700142,0.7579388,0.89512235,0.7133542,0.5658819,0.37039545,0.17490897,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.030866288,0.0,0.0,0.0,0.037725464,0.037725464,0.034295876,0.16462019,0.15090185,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.0548734,0.106317215,0.16462019,0.2503599,0.72364295,0.9877212,0.97400284,0.8265306,0.89855194,1.0425946,1.1626302,1.2449403,1.3889829,1.821111,2.335549,2.9494452,3.4055803,3.6353626,3.7691166,4.5990767,5.6176643,6.6739774,7.7783046,9.091836,11.30735,12.984418,14.164196,15.175924,16.660936,17.271402,17.017612,17.243965,18.067066,18.37573,18.142517,18.903887,19.514353,19.901896,21.057667,21.033659,21.832754,22.813616,23.928232,25.704758,26.579304,28.033447,29.000591,29.384705,30.056904,32.601658,37.00182,41.22707,45.15052,50.55212,56.914005,62.53853,66.48941,67.04157,61.68799,56.492165,50.70988,45.88102,43.48031,44.88987,44.876152,44.018757,43.260815,43.38771,45.023624,52.20518,54.26293,50.631,40.294224,21.78817,20.141968,16.667795,13.3033695,10.422516,6.842027,8.008087,8.440215,9.095266,9.530824,7.9017696,8.639131,7.658269,7.4799304,9.568549,14.325387,15.700651,14.949572,14.71636,15.642348,16.37628,19.6241,20.128248,19.092514,18.166525,19.45262,18.965618,15.656067,13.094165,11.924676,9.877212,10.13786,10.703742,10.792912,10.693454,11.780633,11.4205265,11.478829,11.845795,12.082437,11.396519,10.377932,9.925226,9.688584,9.630281,10.045261,11.029553,11.465111,11.917816,12.895248,14.856973,17.182234,19.435472,20.954779,21.62012,21.86362,23.297188,22.77932,20.86218,18.307138,16.074476,15.577187,15.62863,16.503176,17.370861,16.283682,16.619781,15.978448,15.927004,16.664366,17.051908,18.019053,18.924463,20.015072,20.954779,20.817596,19.613811,18.629519,17.689812,16.767254,15.981877,16.074476,16.63007,16.582056,15.594335,14.057879,12.96727,12.161317,11.900668,12.13731,12.511135,13.711491,14.661487,15.96816,17.669235,19.243416,18.670673,18.296848,18.416885,18.62609,17.820137,16.54433,15.940722,15.758954,15.789821,15.885849,15.422854,15.803539,15.645778,14.572317,13.203912,12.703192,12.075578,12.614022,13.978998,14.188204,13.505715,11.989838,10.751757,10.72432,12.662037,12.672326,13.522863,15.443433,17.532051,17.748116,16.695232,16.492886,15.673215,14.061309,12.747777,11.286773,11.571428,11.996697,11.852654,11.345076,10.220171,9.637141,9.89436,10.600855,10.679735,9.822338,9.829198,9.705732,9.386781,9.719451,9.836057,9.932085,9.962952,9.932085,9.89436,9.863494,10.028113,10.082987,9.839486,9.201583,8.368194,7.9875093,7.8194594,7.706283,7.56567,7.373613,7.4353456,7.641121,7.922347,8.241299,8.522525,8.539673,8.659708,9.0644,9.750318,9.345626,9.057541,9.383351,10.14129,10.504827,9.918367,10.213311,10.796341,11.1393,10.81006,10.422516,10.659158,11.166737,11.561139,11.451392,11.159878,11.495977,11.862943,11.430815,9.122703,0.4938606,0.59331864,0.607037,0.6241849,0.6824879,0.78194594,0.88826317,0.97057325,1.0014396,0.9568549,0.823101,0.7922347,0.864256,0.97400284,1.0734608,1.1214751,1.3615463,1.3924125,1.3581166,1.3375391,1.3443983,1.3443983,1.3409687,1.3238207,1.2963841,1.2895249,1.4610043,1.4061309,1.3546871,1.371835,1.3581166,1.3375391,1.3066728,1.2415106,1.1592005,1.1146159,1.1489118,1.1283343,1.0871792,1.0597426,1.08032,1.3546871,1.5158776,1.8999915,2.6716487,3.8137012,4.029765,6.910619,10.106995,13.598314,19.70641,27.062874,22.652426,13.375391,5.346727,3.9165888,4.602506,3.7005248,2.1915064,0.9945804,0.94999576,1.3238207,1.6427724,1.6290541,1.3786942,1.371835,1.3169615,1.2689474,1.1729189,1.1351935,1.3992717,1.471293,1.2998136,1.1660597,1.155771,1.138623,1.039165,0.7990939,0.6276145,0.59674823,0.64133286,0.4081209,0.2709374,0.19548649,0.23321195,0.51100856,0.9945804,1.1729189,1.1626302,1.0631721,0.9842916,0.6790583,0.4115505,0.274367,0.28122616,0.35324752,0.36010668,0.42869842,0.61389613,0.9294182,1.3443983,1.138623,1.1729189,0.9294182,0.41840968,0.16462019,0.15433143,0.14404267,0.1097468,0.058302987,0.024007112,0.061732575,0.0548734,0.048014224,0.05144381,0.06516216,0.08573969,0.20234565,0.24350071,0.20234565,0.24350071,0.6241849,0.548734,0.77165717,1.1797781,0.77851635,1.0940384,1.5433143,1.9857311,2.1915064,1.8348293,1.920569,1.6084765,1.4164196,1.5604624,1.9857311,1.9171394,1.879414,1.8382589,1.7833855,1.728512,1.4369972,1.3032433,1.1489118,0.9328478,0.7407909,0.94999576,0.8848336,0.7510797,0.6824879,0.72021335,1.2106444,1.214074,1.2620882,1.3786942,1.0666018,0.94656616,0.97400284,0.96714365,0.90198153,0.9362774,0.89169276,0.9911508,0.91569984,0.7922347,1.2106444,0.9877212,1.0151579,0.9602845,0.764798,0.66533995,0.45613512,0.4664239,0.53501564,0.5624523,0.51100856,0.66191036,0.6001778,0.5693115,0.6379033,0.70649505,0.51100856,0.6207553,0.6859175,0.6241849,0.58645946,0.69963586,0.6927767,0.89512235,1.2243627,1.1832076,1.3752645,1.587899,1.7250825,1.6839274,1.371835,1.4027013,1.5707511,1.7079345,1.6976458,1.4507155,1.3272504,1.3306799,1.4404267,1.6084765,1.7593783,1.6221949,1.9754424,2.3904223,2.6064866,2.5481834,2.8739944,3.2786856,3.3644254,3.3026927,3.8377085,4.5784993,5.1066556,5.518206,5.778855,5.751418,6.001778,6.2041235,6.0737996,5.919468,6.6465406,6.701414,8.848335,11.146159,11.900668,9.647429,4.4859004,4.341858,5.24041,5.5490727,5.970912,7.267296,7.3255987,7.3084507,7.5279446,7.459353,8.553391,9.3593445,9.798331,9.897789,9.801761,9.856634,10.089847,10.209882,10.014396,9.369633,8.591117,8.258447,7.864044,7.5862474,8.299602,8.721441,9.1981535,9.174147,8.800322,8.913498,8.81747,8.529384,8.64942,9.043822,8.865483,9.753747,9.897789,9.822338,9.921797,10.467101,10.39508,10.8958,11.670886,12.562579,13.55373,13.924125,14.325387,15.031882,15.642348,15.097044,16.86671,17.415445,19.658396,22.645567,21.558388,31.768269,36.32619,29.611057,16.386568,11.787492,12.521424,10.13786,6.5642304,3.7965534,3.923448,4.307562,4.280125,3.7108135,2.8396983,2.2566686,1.7833855,1.4369972,1.2209331,1.1111864,1.0220171,1.1454822,1.2860953,1.6770682,2.1263442,2.037175,2.0817597,2.5207467,3.9165888,5.802862,6.691125,6.601956,5.2575574,5.9743414,8.220721,7.630832,3.6387923,2.1057668,1.821111,1.7936742,1.2860953,1.1934965,1.1008976,1.0700313,1.0494537,0.8779744,0.70649505,0.59674823,0.4972902,0.38754338,0.30866286,0.22292319,0.2777966,0.32924038,0.34981793,0.44584638,0.53501564,0.53501564,0.548734,0.64476246,0.84024894,0.9842916,1.2346514,1.605047,1.9925903,2.1983654,2.6647894,2.6476414,2.8465576,3.340418,3.5976372,3.4878905,4.0606318,5.586798,7.6205435,9.023245,11.190743,12.065289,12.977559,14.085316,14.363112,13.203912,11.434244,10.847785,11.170166,10.069269,8.086967,6.5299344,5.2301207,4.187526,3.5530527,3.2203827,3.4844608,4.3933015,5.888602,7.8263187,6.807731,5.120374,3.4433057,2.1263442,1.1626302,1.2106444,1.4438564,1.1351935,0.36353627,0.034295876,0.13375391,0.09602845,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.16462019,0.15090185,0.058302987,0.06516216,0.12689474,0.0,0.072021335,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.1097468,0.1371835,0.16804978,0.28465575,0.41840968,0.34295875,0.91227025,1.0666018,1.0048691,0.9362774,1.0563129,1.1523414,1.138623,1.1420527,1.3101025,1.8108221,2.194936,2.6853669,3.0557625,3.2649672,3.4398763,4.2595477,4.880303,5.4941993,6.310441,7.5416627,9.575408,11.372512,12.788932,14.321958,17.130789,18.437462,18.413456,18.667244,19.387459,19.315437,18.12537,18.502625,19.260563,19.895037,20.604961,20.752434,21.45207,22.210009,23.074265,24.638157,25.447538,26.51757,26.881107,26.61703,26.83995,28.76395,32.478195,37.16987,42.90757,50.620712,63.817764,79.88195,94.317085,102.34232,98.9093,91.343636,77.78304,63.91379,54.043438,51.11114,49.38263,47.438053,46.368023,45.89131,44.354855,48.099964,44.80756,38.195316,30.317553,21.585823,28.208357,22.594122,15.385129,10.700313,6.108095,6.461343,7.157549,9.801761,13.004995,12.397959,11.777204,8.543102,7.829748,11.348505,17.394867,18.413456,17.593784,15.518884,14.232788,17.21996,16.352274,15.971589,15.45715,15.525743,18.238546,17.302269,13.337666,9.499957,7.157549,5.895461,8.176137,10.364213,11.430815,11.502836,11.852654,11.410237,11.63659,11.96926,11.9040985,11.012405,9.993818,9.644,9.674867,9.983529,10.669447,11.866373,12.46998,13.13532,14.565458,17.518333,19.672113,21.500084,22.480946,22.597551,22.333473,23.475527,22.504953,20.330595,17.751545,15.443433,13.978998,13.807519,14.143619,14.291091,13.646329,14.044161,13.557159,13.485138,14.229359,15.278812,15.752095,15.981877,16.55119,17.532051,18.512913,17.933313,17.494326,16.674654,15.512024,14.603184,15.05246,15.577187,15.412566,14.496866,13.454271,11.938394,10.597425,10.079557,10.329918,10.590566,12.0309925,13.145609,14.685493,16.691803,18.512913,19.37031,19.329155,19.572655,19.980776,19.137098,16.417435,16.108772,16.403717,16.414005,16.173935,15.343974,15.083325,14.531162,13.536582,12.662037,11.828648,11.094715,11.653738,13.255356,14.205351,13.1593275,12.253916,11.691463,11.592006,11.989838,12.836946,13.982429,15.604623,17.161655,17.384579,16.221949,15.9578705,15.601193,14.7369375,13.54687,12.247057,12.908967,13.275933,12.445972,10.868362,10.179015,9.89436,9.9698105,10.189304,10.189304,9.72631,10.007536,9.918367,9.455373,9.757176,10.052121,9.72288,9.294182,9.047252,9.026674,9.355915,9.513676,9.541112,9.451943,9.242738,8.766026,8.244728,8.049242,8.018375,7.442205,7.0203657,7.226141,7.630832,7.9086285,7.8606143,7.915488,8.014946,8.320179,8.855195,9.530824,9.407358,9.379922,9.791472,10.446524,10.600855,10.285333,10.5597,11.087856,11.441104,11.122152,10.244178,10.275044,10.72089,10.988399,10.381361,10.326488,11.080997,11.578287,11.163307,9.578837,0.5693115,0.6344737,0.59331864,0.5418748,0.53501564,0.58988905,0.70306545,0.7956643,0.89169276,0.9534253,0.881404,0.85396725,0.980862,1.1111864,1.1626302,1.1351935,1.4850113,1.6256244,1.6084765,1.5124481,1.4644338,1.4953002,1.4953002,1.4541451,1.3958421,1.3786942,1.646202,1.4164196,1.1626302,1.097468,1.1489118,1.0048691,0.9911508,0.96371406,0.90884066,0.94656616,0.9294182,0.8711152,0.8745448,1.0082988,1.2895249,1.5124481,1.8073926,2.5241764,3.5290456,4.2081037,4.8734436,8.028665,10.762046,13.872682,21.843042,26.740494,21.163984,12.185325,5.1992545,3.9200184,5.353586,4.530485,2.5824795,0.7922347,0.5658819,0.91569984,1.3032433,1.371835,1.1866373,1.2517995,1.2826657,1.3066728,1.2998136,1.2346514,1.0666018,1.1934965,1.0220171,1.0151579,1.155771,0.96371406,0.96714365,0.8093826,0.61389613,0.4664239,0.41498008,0.20920484,0.17490897,0.18176813,0.25378948,0.5727411,1.3443983,1.5398848,1.3615463,1.0631721,0.9568549,0.8128122,0.5555932,0.34295875,0.2469303,0.28808534,0.40126175,0.548734,0.7133542,0.96371406,1.471293,1.1763484,0.8025235,0.4424168,0.17490897,0.08573969,0.14061308,0.16462019,0.13032432,0.058302987,0.01371835,0.07545093,0.061732575,0.034295876,0.030866288,0.05144381,0.07545093,0.17490897,0.19548649,0.14747226,0.19548649,0.3806842,0.39097297,0.41498008,0.52472687,0.65162164,0.6927767,1.1283343,1.7010754,1.978872,1.3478279,1.7216529,1.4061309,1.2209331,1.4918705,2.054323,2.2223728,1.9891608,1.6564908,1.5124481,1.8176813,1.587899,1.3752645,1.1934965,1.0837497,1.1283343,1.1694894,0.9534253,0.7099246,0.72021335,1.3375391,1.2517995,1.2277923,1.1454822,1.0254467,1.0151579,0.91227025,1.1214751,1.0082988,0.66533995,0.91227025,0.6036074,0.7990939,0.7956643,0.6241849,1.0494537,0.864256,0.7956643,0.75450927,0.67219913,0.5178677,0.5658819,0.5178677,0.48014224,0.4972902,0.52472687,0.9294182,0.75450927,0.67219913,0.78537554,0.6241849,0.51100856,0.61389613,0.7339317,0.7476501,0.58645946,0.78537554,0.8471081,0.9945804,1.2003556,1.1832076,1.5433143,1.4267083,1.529596,1.7422304,1.1454822,1.3066728,1.4027013,1.5638919,1.7147937,1.605047,1.611906,1.5364552,1.5055889,1.5433143,1.5844694,1.9994495,2.411,2.7059445,2.884283,3.0729103,2.8499873,2.935727,3.415869,4.057202,4.280125,4.839148,5.2266912,5.4941993,5.5387836,5.1409516,5.4667625,5.802862,5.7822843,5.6965446,6.492209,6.992929,8.97523,11.317638,12.133881,8.766026,5.579939,5.4153185,6.169828,6.697984,6.8111606,7.7577267,7.864044,8.100685,8.669997,8.988949,9.352485,10.103564,10.401938,10.30591,10.789482,10.607714,10.39508,10.484249,10.679735,10.261326,9.22902,8.690575,8.330468,8.354475,9.489669,9.904649,10.261326,10.096705,9.527394,9.249598,9.050681,8.999237,9.400499,10.052121,10.237319,10.31277,10.031544,10.014396,10.460241,11.153018,10.933525,11.670886,12.30536,12.713481,13.71492,14.767803,15.179354,15.649208,16.067617,15.512024,17.669235,17.463459,18.87645,22.429502,25.159454,35.767166,39.90668,31.442457,15.824117,10.106995,11.664027,9.0369625,5.6073756,3.4947495,3.5770597,3.841138,3.6216443,3.1792276,2.7093742,2.2978237,1.99602,1.7319417,1.5330256,1.4061309,1.3341095,1.5981878,1.6016173,1.8416885,2.2052248,1.9445761,2.0989075,2.935727,4.170378,5.5319247,6.7665763,5.919468,6.0635104,6.6876955,7.4627824,8.261876,5.3981705,3.7691166,2.9254382,2.301253,1.2037852,1.3169615,1.4232788,1.3546871,1.1832076,1.2415106,0.9945804,0.7373613,0.5007198,0.34981793,0.35324752,0.26750782,0.32924038,0.3841138,0.4081209,0.51100856,0.61046654,0.61389613,0.6036074,0.7133542,1.1489118,1.488441,1.6667795,1.6770682,1.6907866,2.0680413,2.3286898,2.4007113,3.1723683,4.3624353,4.496189,3.8274195,3.5530527,3.2512488,3.223812,4.48933,5.456474,8.790032,13.018714,16.12249,15.518884,14.959861,14.503725,14.349394,14.195063,13.227919,10.031544,8.06639,6.8214493,5.977771,5.3844523,4.8425775,4.623084,4.839148,5.641671,7.2124224,6.4407654,4.835718,3.1106358,1.9480057,1.99602,2.2635276,2.1434922,1.3992717,0.38754338,0.06859175,0.082310095,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16119061,0.34295875,0.09945804,0.23664154,0.18862732,0.1371835,0.13032432,0.044584636,0.010288762,0.006859175,0.006859175,0.0,0.0,0.0,0.037725464,0.08573969,0.16804978,0.35324752,0.37039545,0.432128,0.61046654,0.77851635,0.6001778,1.0906088,1.1934965,1.1866373,1.2003556,1.2346514,1.2758065,1.2175035,1.2860953,1.5741806,2.037175,2.095478,2.2086544,2.3732746,2.6647894,3.2649672,4.180667,4.1943855,4.7259717,5.926327,6.677407,8.433355,10.007536,11.519984,13.646329,17.638369,19.517782,19.589804,19.826445,20.567236,20.491785,18.862732,18.95533,19.908754,20.889618,21.11597,21.006224,21.7916,22.343761,22.559826,23.36921,24.319204,24.922812,24.559277,23.94538,25.145735,25.814505,27.10403,29.34698,32.615376,36.724022,47.921627,68.74265,93.25734,113.36159,118.82492,116.68143,103.22715,85.32813,68.80096,58.429882,52.918533,48.768734,46.14167,43.048183,35.3419,30.869717,24.60729,20.697561,21.325174,26.699339,31.970613,27.121178,22.131128,18.763273,10.539123,7.2775846,6.1149545,10.618003,17.583494,17.024471,12.236768,8.443645,8.110974,11.441104,16.345413,15.385129,15.518884,14.068168,12.106443,14.479718,15.093615,14.778092,15.062748,16.163645,16.96617,15.059319,12.3533745,9.836057,8.1384115,7.5690994,8.447074,10.017825,10.861504,10.611144,9.945804,9.235879,9.427936,9.825768,10.021255,9.911508,9.373062,9.716022,10.515115,11.447963,12.274493,13.756075,14.699212,15.4914465,16.88043,19.9602,20.773012,21.602972,21.860191,21.335464,20.183123,20.186552,18.752985,16.828985,15.062748,13.7938,12.891819,13.066729,12.7272,11.746337,11.430815,11.777204,11.780633,12.006986,12.55229,13.049581,12.898679,12.97413,13.443983,14.2190695,14.973578,15.721229,16.352274,15.999025,14.555169,12.648318,13.2690735,13.663476,13.584596,13.029003,12.243628,11.101575,9.997248,9.613133,9.938945,10.288762,11.204462,12.507706,13.982429,15.539461,17.20624,19.215979,19.346302,19.497204,19.997925,19.60695,15.88242,15.54632,15.9613,15.954441,15.803539,15.004445,14.459141,13.732068,12.915827,12.644889,11.039842,10.816919,11.454823,12.545431,13.783512,12.55915,13.149038,13.509145,12.600305,10.388221,11.485688,12.668896,13.87954,14.994157,15.851553,16.098484,16.12249,15.985307,15.402277,13.759505,13.454271,14.682064,14.853543,13.282792,11.197603,11.945253,11.7257595,11.30049,10.984968,10.652299,10.360784,10.535692,10.600855,10.422516,10.329918,10.048691,9.06097,8.354475,8.31332,8.694004,9.030104,9.026674,9.047252,9.156999,9.112414,8.958082,8.423067,8.275595,8.40249,7.7920227,7.421627,7.610255,7.8777623,7.891481,7.4765005,7.3084507,7.579388,7.966932,8.340756,8.755736,9.283894,9.736599,10.1481495,10.494537,10.679735,10.72432,11.06042,11.38966,11.499407,11.276484,9.993818,9.6645775,9.661148,9.472521,8.704293,9.3593445,10.364213,10.840926,10.652299,10.429376,0.45613512,0.39783216,0.42869842,0.4389872,0.41840968,0.4424168,0.52815646,0.5418748,0.5761707,0.66191036,0.7476501,0.69963586,0.77851635,0.91227025,1.0254467,1.039165,1.0734608,1.2483698,1.3032433,1.2312219,1.2826657,1.097468,1.08032,1.2380811,1.4027013,1.2209331,1.0871792,1.0700313,0.9842916,0.881404,1.0528834,0.96714365,0.9362774,0.89512235,0.83681935,0.823101,0.83681935,0.85739684,0.9568549,1.1283343,1.313532,1.8005334,2.4898806,3.2889743,3.8925817,3.7691166,6.125243,9.122703,10.902658,13.251926,21.575535,22.724447,17.38115,10.573419,5.6313825,4.166949,4.2869844,3.7965534,2.4487255,0.83338976,0.3806842,0.6756287,0.85739684,1.039165,1.1763484,1.0666018,1.1763484,1.2517995,1.3169615,1.3203912,1.1146159,0.96714365,0.84024894,0.8711152,0.9774324,0.85396725,0.91569984,0.8025235,0.58302987,0.35324752,0.24350071,0.13375391,0.12346515,0.1371835,0.19548649,0.42869842,1.196926,1.5158776,1.2586586,0.77165717,0.8711152,1.0288762,0.78537554,0.4424168,0.22635277,0.274367,0.5555932,0.67219913,0.7990939,1.0082988,1.2517995,0.65162164,0.29151493,0.09602845,0.024007112,0.061732575,0.14747226,0.14061308,0.08573969,0.0274367,0.01371835,0.01371835,0.024007112,0.017147938,0.01371835,0.07545093,0.05144381,0.09945804,0.1371835,0.14747226,0.18176813,0.23321195,0.24350071,0.39783216,0.6379033,0.6859175,0.4664239,0.48357183,0.58988905,0.7613684,1.1283343,1.1900668,1.0940384,1.1214751,1.3101025,1.4815818,1.6393428,2.0268862,2.1983654,1.9891608,1.5261664,1.1489118,0.9431366,0.91227025,0.9568549,0.8848336,0.7373613,1.1146159,1.2860953,1.2758065,1.862266,1.1420527,1.3101025,1.2963841,0.9431366,0.9911508,1.2586586,1.2449403,0.8711152,0.40126175,0.4115505,1.0117283,1.0666018,0.7579388,0.48700142,0.91569984,0.7682276,0.7682276,0.6036074,0.32238123,0.33609957,0.5178677,0.5178677,0.4629943,0.42869842,0.42869842,0.59674823,0.45613512,0.4389872,0.6241849,0.7339317,0.42869842,0.48014224,0.7407909,0.91569984,0.548734,1.1592005,1.2586586,1.1420527,1.0254467,1.039165,1.2689474,0.91569984,0.9945804,1.3992717,0.90198153,1.4610043,1.5638919,1.7250825,2.1915064,2.959734,2.311542,1.9137098,1.8039631,1.8897027,1.937717,2.2566686,2.4075704,2.4144297,2.4384367,2.7916842,2.901431,3.2958336,3.8274195,4.355576,4.746549,4.647091,4.633373,4.979761,5.4839106,5.446185,6.1904054,6.697984,6.39961,5.830299,6.636252,7.932636,9.407358,10.988399,11.705182,9.705732,8.484799,8.224151,8.378482,8.800322,9.764035,9.911508,9.911508,9.80862,9.589127,9.184435,9.331907,10.220171,10.563129,10.1652975,9.932085,9.373062,9.266746,9.6645775,10.285333,10.528833,11.039842,10.8958,10.5597,10.528833,11.321068,11.530273,11.499407,10.748327,9.602845,9.201583,9.482809,9.571979,9.626852,9.650859,9.489669,10.209882,10.545981,11.218181,12.068718,12.068718,11.252477,11.797781,12.38424,12.9707,14.802099,15.326826,15.693792,16.410576,16.96617,15.854982,17.806417,18.296848,21.53781,28.76395,38.22275,41.933567,41.14819,30.26611,14.270514,8.7283,8.742019,6.9689217,4.6608095,3.0523329,3.357566,3.4192986,3.1209247,2.901431,2.836269,2.6407824,2.5070283,2.2806756,2.0646117,1.920569,1.845118,2.1023371,2.201795,2.411,2.6887965,2.6990852,2.750529,2.7882545,3.3198407,4.2526884,4.897451,5.312431,6.461343,7.394191,8.2481575,10.237319,9.702303,6.975781,4.7842746,3.642222,1.862266,1.7525192,1.862266,1.7765263,1.4987297,1.4507155,1.1454822,0.77508676,0.432128,0.2194936,0.24350071,0.29151493,0.50757897,0.53844523,0.40126175,0.48700142,0.53844523,0.5590228,0.5212973,0.5144381,0.7476501,1.2106444,1.6187652,1.8656956,1.9342873,1.9239986,1.7147937,2.1194851,3.5976372,5.2644167,4.897451,5.3741636,5.528495,5.192395,4.928317,6.025785,7.1026754,9.575408,15.587475,22.817045,24.490685,20.913624,19.826445,17.648657,14.596324,14.695783,13.251926,10.6145735,8.378482,7.239859,6.958633,7.7268605,6.9860697,6.2830043,6.307011,6.883182,5.2815647,3.6010668,2.4658735,2.0577524,2.1057668,2.668219,2.4590142,1.5124481,0.37382504,0.09259886,0.116605975,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17147937,0.4424168,0.5041494,0.45613512,0.5693115,0.6927767,0.64476246,0.22978236,0.044584636,0.037725464,0.037725464,0.0,0.0,0.0,0.18176813,0.42869842,0.6241849,0.67219913,0.5624523,0.96371406,1.1283343,1.0048691,1.2346514,1.4918705,1.4198492,1.4267083,1.5158776,1.2963841,1.4061309,1.5158776,1.6873571,1.903421,2.0749004,2.452155,2.5378947,2.5927682,2.8019729,3.2649672,4.3281393,4.0263357,4.636802,6.324159,7.140401,8.251588,9.818909,11.022695,12.6586075,17.151367,18.739265,19.95677,20.70785,20.882757,20.37175,19.198832,19.984205,21.256582,22.213438,22.751883,22.642136,23.02625,23.660725,24.27462,24.566135,24.566135,24.61415,24.085993,23.595562,24.963966,25.622448,25.715046,26.136887,26.812515,26.702768,23.883648,26.219196,32.24155,40.932125,51.749046,62.415062,74.40833,79.130875,74.81302,66.51342,59.45533,49.169994,38.795494,29.566473,20.814167,15.453721,11.204462,9.606275,11.159878,15.337115,20.207129,25.883097,25.9414,19.13024,9.352485,8.14527,6.615674,7.3050213,10.113853,12.298501,11.664027,9.537683,9.736599,12.291641,13.426835,8.923786,9.373062,11.262765,12.771784,13.749216,15.199932,20.03222,20.683842,17.610931,19.270851,12.864383,8.477941,6.941485,7.6788464,8.7283,9.362774,9.163857,8.669997,8.06639,7.1884155,7.98065,8.207003,8.450503,8.766026,8.666568,8.604835,9.513676,11.05356,12.785502,14.191633,16.276823,17.28512,17.905876,18.6158,19.654966,20.11796,20.86561,20.474638,18.756414,16.753534,16.033321,15.093615,14.167625,13.488567,13.306799,13.440554,13.337666,12.579727,11.4205265,10.772334,10.504827,10.786053,10.858074,10.5597,10.316199,10.340206,10.436234,11.022695,11.859513,12.055,13.018714,13.790371,14.30481,13.845244,11.063849,11.135871,12.024134,12.840376,13.1593275,13.001566,11.976119,11.444533,10.9541025,10.432805,10.179015,10.652299,13.179905,15.361122,16.410576,17.182234,19.023922,19.349733,19.713268,20.37518,20.27915,18.019053,16.20137,15.151917,14.949572,15.426285,14.596324,14.46257,14.479718,14.195063,13.227919,11.410237,11.111863,12.154458,13.639469,13.9309845,13.077017,13.615462,14.143619,13.670336,11.595435,11.170166,12.106443,13.38911,14.616901,16.023033,16.911295,17.364002,17.106783,16.067617,14.359683,14.675205,15.313108,15.172495,13.821238,11.489118,11.7086115,11.893809,12.037852,11.825217,10.604284,10.703742,11.276484,11.814929,11.880091,11.122152,9.623423,7.798882,7.4044795,8.378482,8.865483,8.597976,8.666568,8.721441,8.601405,8.330468,8.1487,7.956643,8.107545,8.464222,8.378482,7.7542973,7.9737906,8.279024,8.220721,7.658269,7.4524937,7.5382333,7.8434668,8.364764,9.170717,9.366203,9.956093,10.583707,11.008976,11.094715,11.129011,11.622872,11.701753,11.214751,10.72775,9.201583,8.848335,9.023245,9.191295,8.9100685,9.156999,10.323058,10.6488695,10.110424,10.4533825,0.44584638,0.4424168,0.4664239,0.48357183,0.48357183,0.48014224,0.4664239,0.490431,0.548734,0.61389613,0.65162164,0.6790583,0.72021335,0.764798,0.83681935,0.9774324,0.9259886,1.1008976,1.214074,1.1660597,1.039165,1.0700313,0.980862,0.96714365,1.039165,1.0117283,0.90884066,0.89169276,0.823101,0.71678376,0.77165717,0.83338976,0.8676856,0.922559,0.9842916,0.9842916,1.0151579,1.1008976,1.2792361,1.5433143,1.8245405,2.2841053,2.7470996,3.2478194,3.9131594,4.9523244,7.6205435,9.451943,12.411677,17.734396,25.93454,21.650986,13.762935,7.606825,4.866585,3.566771,3.0729103,2.8911421,2.1469216,0.9534253,0.39440256,0.48014224,0.58988905,0.6036074,0.5693115,0.70306545,0.84024894,1.1111864,1.214074,1.1180456,1.0768905,0.9877212,0.7956643,0.69963586,0.7407909,0.7922347,0.91227025,0.77851635,0.53844523,0.31209245,0.18176813,0.17147937,0.22978236,0.29494452,0.32924038,0.31895164,0.71678376,1.0666018,1.1146159,0.9431366,0.9911508,0.9945804,0.7407909,0.47671264,0.36696586,0.4938606,0.51100856,0.4972902,0.6173257,0.91912943,1.2998136,0.8779744,0.4664239,0.18176813,0.06516216,0.061732575,0.116605975,0.10288762,0.058302987,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.06859175,0.058302987,0.058302987,0.08916927,0.09602845,0.18519773,0.28808534,0.36696586,0.4046913,0.4046913,0.6241849,0.65162164,0.5727411,0.53844523,0.7373613,0.8676856,1.1351935,1.3889829,1.5844694,1.786815,1.9720128,2.1983654,2.1263442,1.7010754,1.1592005,1.3581166,1.2895249,1.0185875,0.83681935,1.2517995,1.0666018,1.4095604,1.3855534,0.9602845,0.97057325,0.9534253,1.430138,1.5158776,1.2037852,1.371835,1.5913286,1.3341095,0.9911508,0.8093826,0.89855194,1.4678634,1.1180456,0.64819205,0.48700142,0.67219913,0.7407909,0.72021335,0.6036074,0.490431,0.5796003,0.65505123,0.5418748,0.4629943,0.4698535,0.4389872,0.6207553,0.61389613,0.5658819,0.53501564,0.48700142,0.4664239,0.6173257,0.6859175,0.607037,0.52472687,1.1729189,1.0700313,0.89512235,1.0460242,1.6359133,1.2998136,1.3101025,1.3889829,1.3478279,1.0837497,1.587899,1.7182233,1.786815,1.9514352,2.253239,2.0749004,2.1057668,2.270387,2.4624438,2.5619018,2.603057,2.4555845,2.6613598,3.0317552,2.633923,3.2889743,3.4844608,3.5564823,3.7794054,4.355576,4.5099077,4.698535,4.7979927,4.9214582,5.411889,5.861165,6.3310184,6.8145905,7.449064,8.529384,8.241299,8.255017,9.006097,9.757176,8.594546,8.299602,8.961512,10.096705,11.324498,12.377381,11.694893,11.077567,10.864933,10.840926,10.2236,10.134431,10.209882,10.127572,9.887501,9.81205,9.798331,9.860064,10.134431,10.593996,11.05356,11.626302,12.116733,12.47341,12.610593,12.408247,12.168177,11.849225,11.166737,10.357354,10.189304,9.962952,9.89436,10.124143,10.388221,10.0041065,10.655728,11.180455,12.055,12.922686,12.569438,12.346515,12.641459,13.056439,13.917266,16.266533,15.940722,17.261114,18.6158,19.092514,18.478617,21.554956,21.94936,26.455837,34.378185,37.540264,35.616264,31.000042,22.573545,13.190193,9.6817255,8.745448,6.7631464,4.9488945,3.9611735,3.8925817,3.8857226,3.7211025,3.525616,3.3850029,3.3369887,3.1415021,3.1586502,3.316411,3.4947495,3.5187566,3.6970954,4.0194764,4.2869844,4.4104495,4.420738,3.8171308,3.5530527,3.6010668,3.9165888,4.4447455,5.302142,5.9126086,6.550512,7.366754,8.4093485,9.297611,8.333898,6.3653145,4.249259,2.8396983,2.6407824,2.603057,2.5584722,2.3321195,1.7662375,1.1283343,0.77851635,0.6036074,0.48014224,0.28122616,0.23321195,0.45613512,0.5761707,0.51100856,0.5007198,0.48014224,0.39097297,0.39097297,0.61046654,1.1249046,2.1160555,3.1037767,4.139512,4.513337,2.7539587,2.136633,3.0248961,4.180667,4.887162,4.9591837,6.478491,5.4907694,4.5201964,4.839148,6.468202,8.107545,9.815479,13.197053,17.679523,20.522652,15.512024,15.810398,17.566347,17.919594,15.001016,11.489118,8.851766,7.442205,7.2638664,7.9600725,8.512236,7.7542973,7.2467184,7.2192817,6.5642304,4.6608095,3.175798,2.4212887,2.1915064,1.7525192,2.0886188,1.605047,0.84024894,0.2777966,0.34638834,0.18519773,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.08916927,0.09945804,0.30523327,0.3841138,0.4664239,0.58645946,0.6790583,0.64476246,0.6344737,0.64819205,0.66191036,0.6241849,0.72021335,0.9259886,1.196926,1.4781522,1.7216529,1.7490896,1.8039631,1.8279701,1.8142518,1.821111,1.845118,1.786815,1.8108221,1.8862731,1.786815,1.903421,1.9582944,1.9582944,2.095478,2.7333813,2.8499873,2.8259802,3.083199,3.57363,3.7519686,4.0537724,4.081209,4.695105,6.0532217,7.6033955,8.961512,10.456812,12.349944,15.141628,19.603521,19.648108,20.550089,21.174273,20.989075,20.066517,19.041069,19.9602,21.61326,22.923363,22.923363,22.295748,23.060547,24.374079,25.488693,25.763062,24.933102,25.10115,24.60386,23.787619,25.001692,26.44212,26.037428,25.145735,24.590141,24.665592,25.145735,26.922262,27.206917,26.35638,27.868828,29.141205,32.82115,38.044415,43.41858,47.033363,53.745064,50.39436,37.896942,21.959648,13.063298,8.776315,6.684266,6.094377,6.608815,8.097256,15.2033615,24.281479,26.18147,19.263992,9.3764925,8.333898,6.6122446,6.6533995,8.1384115,7.9909387,8.244728,8.491658,10.213311,12.569438,12.415107,12.511135,13.9309845,13.522863,11.873232,13.310229,20.95135,29.058895,29.041746,21.301168,15.206791,11.355364,8.937505,8.838047,10.041832,9.606275,11.571428,12.435684,12.024134,10.1481495,6.6122446,6.773435,7.160979,7.7028537,8.368194,9.167287,9.633711,11.201033,12.836946,14.212211,15.704081,17.412016,18.338005,18.307138,17.960749,18.763273,19.305147,19.003344,18.152807,16.935303,15.412566,14.651197,13.944703,13.3033695,12.826657,12.682614,12.504276,12.037852,11.31078,10.487679,9.870353,9.530824,9.760606,10.0041065,9.901219,9.277034,9.047252,8.8929205,8.862054,9.194724,10.295622,10.878652,11.365653,11.869802,12.061859,11.173596,10.902658,11.14273,11.369082,11.444533,11.595435,10.950673,10.371073,10.30591,10.943813,12.1921835,13.203912,15.419425,16.88386,17.350283,18.255693,17.785841,17.96761,19.11309,20.659836,21.20514,18.938183,15.944152,13.488567,12.593445,14.033872,14.13333,14.390549,14.21564,13.416546,12.21619,11.245617,10.830637,11.629731,13.207341,14.030442,13.869251,14.277372,14.565458,14.009865,11.866373,10.72432,10.779194,11.149589,11.80464,13.581166,15.896138,17.034761,17.158226,16.664366,16.163645,15.367981,14.819247,13.756075,12.267634,11.293632,11.22161,11.324498,11.4033785,11.286773,10.837497,11.365653,11.7086115,12.147599,12.267634,10.964391,9.277034,8.045813,7.864044,8.539673,9.098696,8.779744,8.968371,9.088407,9.057541,9.294182,8.388771,8.05953,8.207003,8.7283,9.513676,9.1810055,8.947794,8.793462,8.488229,7.5759587,7.0752387,7.3290286,7.857185,8.361334,8.707723,8.920357,9.294182,10.1481495,11.204462,11.581717,11.47197,11.746337,11.72233,11.146159,10.179015,9.493098,9.39021,9.421077,9.287323,8.851766,9.544542,10.196163,10.590566,10.412228,9.23245,0.41498008,0.39783216,0.3841138,0.38754338,0.4081209,0.432128,0.47671264,0.5693115,0.65848076,0.7407909,0.85396725,0.86082643,0.89512235,0.922559,0.94656616,1.0151579,1.0528834,1.1866373,1.2517995,1.1866373,1.0597426,1.1077567,0.97400284,0.8848336,0.89169276,0.88826317,0.8848336,0.8711152,0.8505377,0.8505377,0.939707,0.9877212,0.9774324,1.0151579,1.1111864,1.1763484,1.2723769,1.3924125,1.5227368,1.7113642,2.0817597,2.7368107,3.199805,3.923448,5.038064,6.3378778,8.580828,11.550851,15.642348,20.361462,24.332924,19.301718,11.379372,6.1321025,4.57164,3.1517909,2.2635276,2.1640697,2.0063086,1.5227368,1.0117283,0.65162164,0.52815646,0.5212973,0.5693115,0.6824879,0.66191036,0.91912943,1.1043272,1.1146159,1.0768905,0.8711152,0.70649505,0.6036074,0.6241849,0.86082643,0.980862,0.8471081,0.58302987,0.31209245,0.15090185,0.16119061,0.26407823,0.33609957,0.33952916,0.32581082,0.4115505,0.6344737,0.91569984,1.2003556,1.471293,1.0768905,0.70306545,0.5418748,0.6756287,1.0700313,1.0425946,0.7990939,0.6241849,0.66533995,0.9294182,1.3684053,1.1626302,0.6927767,0.25721905,0.061732575,0.058302987,0.041155048,0.020577524,0.0034295875,0.0,0.0,0.006859175,0.01371835,0.024007112,0.0548734,0.048014224,0.020577524,0.0274367,0.07888051,0.16804978,0.28122616,0.36010668,0.44584638,0.5041494,0.42869842,0.6756287,0.5727411,0.5212973,0.6276145,0.70649505,0.89512235,1.2209331,1.3272504,1.2277923,1.313532,1.646202,1.5810398,1.5055889,1.4678634,1.1763484,1.1454822,1.0700313,1.0837497,1.1454822,1.0220171,0.97400284,1.3684053,1.2860953,0.8025235,0.9774324,0.980862,1.4575747,1.5330256,1.2415106,1.5021594,1.488441,1.3066728,1.155771,1.1317638,1.2312219,1.3615463,1.097468,0.9294182,0.96371406,0.89512235,0.90541106,0.78194594,0.78194594,0.86082643,0.6790583,0.6173257,0.5658819,0.61046654,0.7133542,0.7339317,0.6927767,0.6241849,0.6344737,0.66533995,0.490431,0.67219913,0.72364295,0.7407909,0.7476501,0.6824879,1.1832076,1.0254467,0.8848336,1.0528834,1.4198492,1.0460242,1.2483698,1.4027013,1.3306799,1.3203912,1.6496316,1.6324836,1.7765263,2.085189,2.0920484,2.0920484,2.5207467,2.7368107,2.651071,2.7162333,2.7059445,2.8911421,3.210094,3.3438478,2.7128036,3.4913201,3.6044965,3.5290456,3.673088,4.3761535,4.2081037,4.914599,5.528495,5.7136927,5.7479887,6.193835,6.7871537,7.5450926,8.347616,8.930646,8.333898,8.364764,8.985519,9.410788,8.114404,7.864044,8.570539,9.434795,10.237319,11.317638,11.043272,10.583707,10.487679,10.792912,11.022695,11.602294,11.567999,11.362224,11.108434,10.604284,10.179015,10.275044,10.398509,10.504827,11.002116,11.917816,12.620882,13.454271,14.016724,13.183334,12.075578,11.742908,11.561139,11.341646,11.341646,11.129011,11.111863,11.293632,11.612583,11.924676,12.737488,12.9707,13.639469,14.562028,14.369971,14.627191,14.788382,15.13134,15.9921665,17.758404,17.37429,19.408035,20.845032,21.174273,22.384918,27.484715,27.117748,30.718815,37.526546,36.56283,31.384155,26.887966,20.76958,14.099034,11.31078,10.47396,8.64256,6.9552035,5.8817425,5.209543,4.9420357,4.681387,4.4447455,4.232111,4.0229063,3.6387923,3.6285036,3.8342788,4.081209,4.166949,4.763697,5.6793966,7.2021337,8.433355,7.2878733,6.8626046,6.15268,5.528495,5.302142,5.751418,6.526505,6.6053853,6.694555,7.0375133,7.4181976,7.8366075,7.486789,6.48535,5.24041,4.465323,4.046913,3.7039545,3.3198407,2.877424,2.4590142,1.5261664,1.1626302,1.0631721,0.94656616,0.53844523,0.4115505,0.805953,1.0425946,0.9259886,0.70649505,0.6241849,0.48357183,0.4389872,0.58302987,0.9294182,2.8499873,3.7348208,4.9008803,5.9640527,4.863155,2.9734523,3.8548563,4.616225,4.619654,5.4770513,7.363324,6.4544835,5.4084597,5.5730796,6.9792104,8.615124,8.347616,9.047252,11.187314,12.867812,13.296511,13.615462,15.3302555,17.20281,15.247946,10.408798,8.440215,8.282454,8.635701,7.98065,7.1198235,6.684266,6.56766,6.2967224,5.038064,3.309552,2.270387,1.9994495,1.9925903,1.1592005,1.9102802,1.5055889,0.823101,0.39097297,0.40126175,0.1371835,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1371835,0.23664154,0.29837412,0.40126175,0.70306545,1.3032433,1.5707511,1.6393428,1.762808,2.3149714,2.452155,2.8568463,3.0420442,2.9322972,2.843128,3.117495,2.9871707,2.7813954,2.6373527,2.5070283,2.5447538,2.4967396,2.4384367,2.4487255,2.5927682,2.6133456,2.5447538,2.6407824,2.8225505,2.6716487,3.5530527,3.5564823,3.5153272,3.6868064,3.7382503,4.2218223,4.5613513,5.302142,6.6053853,8.251588,10.319629,12.161317,15.13134,18.728977,20.584383,20.879328,20.858751,20.587814,19.973917,18.78042,17.95389,19.023922,20.941061,22.384918,21.736725,21.472647,22.18943,23.406935,24.617579,25.26577,24.792488,24.254042,23.69159,23.61957,25.029129,26.788507,26.397535,25.094292,24.247183,25.382378,26.83995,27.066305,27.26522,27.289227,25.622448,23.736176,23.921373,25.93797,28.92857,31.439028,36.92294,34.961216,29.521889,22.9508,15.985307,11.705182,9.081548,7.8023114,7.781734,9.132992,11.64345,16.496315,18.149376,14.620332,7.507367,5.3501563,4.201245,4.9008803,7.0615206,9.081548,8.399059,9.256456,10.792912,12.9707,16.575195,13.6086035,14.143619,13.169616,11.372512,15.148488,26.033998,32.639385,31.970613,24.459818,13.978998,11.588576,12.130451,12.144169,10.563129,8.711152,9.5033865,11.917816,11.324498,7.953213,6.917478,6.7871537,7.442205,8.176137,8.940934,10.353925,11.530273,13.173045,14.009865,13.934414,14.003006,15.594335,16.345413,16.527182,16.492886,16.671225,16.691803,15.937293,15.148488,14.603184,14.116182,13.96871,13.155897,12.2093315,11.592006,11.677745,12.151029,11.633161,10.861504,10.158438,9.414218,9.352485,9.523964,9.496528,9.071259,8.275595,8.172707,7.706283,7.3255987,7.466212,8.546532,9.410788,9.801761,10.521975,11.30735,10.834066,10.185875,9.469091,9.527394,10.281903,10.741467,10.714031,10.089847,9.836057,10.535692,12.401388,13.821238,15.05246,15.930434,16.516893,17.106783,17.2131,17.806417,18.818146,19.795578,19.87446,18.166525,15.522313,13.594885,13.138749,13.989287,13.375391,12.867812,12.38767,11.718901,10.535692,10.48082,10.106995,10.1481495,10.930096,12.349944,13.433694,14.627191,15.138199,14.376831,11.952112,10.508256,9.839486,10.247607,11.406808,12.367092,14.805529,15.542891,15.446862,15.223939,15.443433,14.750656,13.118172,11.869802,11.561139,11.952112,11.327928,11.132441,11.149589,11.279913,11.543991,11.989838,12.771784,13.149038,12.6929035,11.283342,10.216741,9.4862385,9.273604,9.39707,9.31133,8.440215,8.4093485,8.824328,9.31133,9.499957,8.207003,7.9875093,8.381912,8.999237,9.5033865,9.283894,9.1981535,9.057541,8.790032,8.440215,7.8537555,8.128122,8.676856,9.088407,9.122703,9.129561,9.537683,10.30934,11.177026,11.657167,11.314209,11.331357,11.2593355,10.991828,10.755186,9.736599,9.211872,9.091836,9.108984,8.81747,9.585697,9.465661,9.551401,9.959522,9.832627,0.32238123,0.3018037,0.28465575,0.31209245,0.37382504,0.4081209,0.5658819,0.66191036,0.7099246,0.7510797,0.8779744,0.85396725,0.9294182,1.0117283,1.0528834,1.0768905,1.1043272,1.1214751,1.1249046,1.1214751,1.1317638,1.1214751,1.0048691,0.89512235,0.8711152,0.9568549,0.980862,0.9534253,0.9568549,1.0220171,1.1214751,1.1660597,1.2037852,1.255229,1.3272504,1.4267083,1.488441,1.6016173,1.6873571,1.8554068,2.3972816,3.333559,3.9268777,4.8597255,6.1561093,7.205563,11.945253,16.245956,18.687822,18.835295,17.240536,13.341095,8.1041155,4.8494368,3.8685746,2.4452958,1.5741806,1.6153357,2.0474637,2.3286898,1.8656956,1.1797781,0.864256,0.7613684,0.7373613,0.6790583,0.66876954,0.86082643,1.0563129,1.1489118,1.138623,0.8711152,0.65848076,0.5212973,0.5212973,0.7682276,0.805953,0.7099246,0.53158605,0.32238123,0.15090185,0.16119061,0.2469303,0.32924038,0.39783216,0.51100856,0.4046913,0.40126175,0.65848076,1.0940384,1.371835,0.88826317,0.5521636,0.4629943,0.6241849,0.96714365,1.1454822,1.2517995,1.097468,0.8128122,0.82996017,1.7422304,1.670209,1.0734608,0.39783216,0.08573969,0.030866288,0.006859175,0.0034295875,0.0034295875,0.0,0.0034295875,0.010288762,0.020577524,0.034295876,0.06859175,0.024007112,0.017147938,0.0548734,0.1371835,0.26064864,0.33609957,0.41840968,0.5178677,0.59674823,0.5693115,0.75450927,0.6310441,0.64819205,0.86082643,0.91912943,1.0837497,1.2243627,1.1763484,0.9945804,0.939707,1.371835,1.2449403,1.2277923,1.3889829,1.1660597,1.196926,1.1008976,1.1351935,1.2449403,1.0288762,0.97057325,1.2346514,1.2003556,0.939707,1.2277923,1.1694894,1.4335675,1.4472859,1.2449403,1.4781522,1.2998136,1.2106444,1.1523414,1.1420527,1.2689474,1.2723769,1.1283343,1.0940384,1.1489118,0.9911508,0.881404,0.86082643,0.8848336,0.8779744,0.70649505,0.6379033,0.66533995,0.7579388,0.84367853,0.8196714,0.72364295,0.6824879,0.70649505,0.72021335,0.5693115,0.70649505,0.67219913,0.6962063,0.78537554,0.7579388,0.91912943,1.0220171,1.0768905,1.1283343,1.2346514,1.0425946,1.0425946,1.2243627,1.4472859,1.4369972,1.6804979,1.7833855,1.978872,2.218943,2.1983654,2.469303,2.9391565,3.1380725,3.0454736,3.1072063,3.1106358,3.6285036,3.9508848,3.7862647,3.275256,3.998899,3.865145,3.8102717,4.105216,4.3349986,4.5784993,5.223262,5.826869,6.228131,6.550512,6.9654922,7.514226,8.001227,8.447074,9.0644,9.091836,9.208443,9.355915,9.15014,7.888051,7.421627,7.7028537,8.23444,8.8929205,9.914937,10.103564,10.062409,10.082987,10.398509,11.201033,12.6757555,12.648318,12.373952,12.271064,11.910957,11.351934,11.30049,11.153018,10.991828,11.55771,12.449403,13.361672,14.287662,14.79867,14.0750265,12.898679,12.833516,13.13189,13.361672,13.399398,13.3033695,13.313659,13.227919,13.334236,14.441993,14.942713,15.151917,15.830976,16.822126,17.062197,17.532051,17.658945,18.28999,19.404606,20.100813,20.395756,23.067406,24.634727,25.619019,30.557625,33.215553,34.378185,40.167328,47.074516,41.98158,34.117535,28.465576,22.134558,15.697222,13.1593275,12.109874,10.518545,8.923786,7.582818,6.495639,5.768566,5.2747054,4.9488945,4.6745276,4.2835546,3.9028704,3.82399,3.9851806,4.32471,4.7945633,5.381023,6.3721733,8.076678,9.585697,8.783174,8.388771,7.956643,7.966932,8.296172,8.224151,8.1487,8.011517,8.008087,8.134981,8.200144,8.049242,7.9017696,7.582818,7.0272245,6.2418494,5.579939,4.623084,3.9440255,3.542764,2.8259802,2.3561265,1.7422304,1.3821237,1.2415106,0.8676856,0.65505123,0.9431366,1.1660597,1.08032,0.77165717,0.71678376,0.59674823,0.53158605,0.5555932,0.6173257,2.2395205,2.8980014,3.9268777,5.1855364,5.0483527,3.234101,3.5050385,3.7005248,3.566771,4.763697,5.7891436,6.125243,6.3481665,6.6396813,6.790583,8.903209,8.045813,7.5862474,8.529384,9.513676,13.193623,13.96185,14.466,15.158776,14.280802,9.901219,8.440215,8.433355,8.405919,6.8763227,5.7239814,5.717122,5.7925735,5.2609873,3.799983,2.3389788,1.6667795,1.6290541,1.646202,0.72021335,1.5810398,1.2209331,0.7510797,0.5555932,0.30523327,0.24007112,0.1371835,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.09602845,0.14747226,0.14747226,0.058302987,0.29151493,0.53501564,0.71678376,1.0323058,1.7696671,2.2429502,2.5584722,2.8945718,3.5050385,3.7348208,4.1360826,4.3007026,4.197815,4.166949,4.557922,4.4413157,4.125794,3.875434,3.9063,3.9131594,3.8720043,3.8137012,3.8788633,4.331569,4.307562,3.8925817,3.7553983,3.8514268,3.4192986,4.523626,4.8014226,4.6676683,4.479041,4.554492,5.2335505,5.7308407,6.6533995,8.155559,9.918367,12.185325,14.586036,17.885298,21.184563,21.894485,22.261452,21.904776,20.94449,19.62067,18.324286,18.139088,18.886738,20.248285,21.493225,21.486366,21.44178,22.007662,22.597551,23.03654,23.568125,23.403505,22.933651,23.256033,24.518122,25.93111,27.330383,27.066305,25.725336,24.511261,25.224615,26.887966,26.898254,27.94085,29.467016,27.690489,26.274069,26.044287,26.301506,26.730206,27.392115,27.34753,24.398085,23.636717,24.52498,20.872469,14.904987,12.655178,11.578287,11.074138,12.483699,9.873782,10.353925,10.576848,9.160428,6.715132,3.3438478,2.620205,3.7725463,6.2727156,9.832627,8.652849,11.050131,13.807519,16.180794,19.87446,14.922135,14.575747,14.771234,14.658057,16.619781,24.202599,24.991404,22.823904,19.041069,12.504276,13.042721,14.102464,12.21962,8.217292,7.1849856,7.414768,10.683165,10.14472,6.691125,8.930646,7.932636,8.261876,8.961512,9.887501,11.71547,13.488567,15.158776,15.29596,13.965281,12.7272,13.430264,13.944703,14.46257,14.908417,14.932424,14.544881,13.807519,13.262215,13.1421795,13.358243,13.38568,12.590015,11.698323,11.132441,10.998687,11.427385,11.228469,10.7586155,10.30591,10.086417,10.103564,9.993818,9.355915,8.282454,7.366754,7.1026754,6.4373355,6.0566516,6.351596,7.4113383,8.244728,8.827758,9.613133,10.47396,10.710602,10.024684,8.796892,8.604835,9.5033865,10.034973,10.844356,10.813489,10.573419,10.792912,12.195613,14.105893,14.5414505,14.891269,15.693792,16.62321,17.065628,17.12393,17.511473,18.104792,17.96418,17.490896,15.724659,14.339106,13.900118,13.865822,12.607163,11.592006,10.950673,10.491108,9.692014,10.072699,9.626852,9.191295,9.47938,11.0981455,12.596875,13.972139,14.249936,13.238208,11.537132,9.921797,8.858624,9.153569,10.388221,10.930096,12.836946,13.615462,13.80066,13.852104,14.150477,13.478279,12.123591,11.502836,11.931535,12.617453,11.598865,11.245617,11.331357,11.773774,12.644889,13.004995,14.0750265,14.29795,13.365103,12.229909,11.780633,11.297061,10.871792,10.343636,9.318189,8.333898,8.501947,9.187865,9.856634,10.069269,8.453933,8.23444,8.724871,9.280463,9.321619,9.06097,9.126132,9.263316,9.318189,9.253027,8.522525,8.656279,9.112414,9.513676,9.671436,9.424506,9.825768,10.412228,10.930096,11.321068,10.899229,10.463672,10.155008,10.124143,10.55284,10.052121,9.561689,9.253027,9.095266,8.865483,9.170717,8.604835,8.604835,9.506817,10.545981,0.26064864,0.26407823,0.28122616,0.34981793,0.4389872,0.44584638,0.6859175,0.72364295,0.66876954,0.6310441,0.72021335,0.6824879,0.805953,0.9602845,1.0768905,1.1694894,1.0768905,0.94999576,0.9362774,1.0494537,1.1763484,1.097468,1.0117283,0.9294182,0.91227025,1.0871792,1.08032,1.0631721,1.0666018,1.1043272,1.1729189,1.2655178,1.4198492,1.5090185,1.546744,1.6770682,1.6084765,1.7250825,1.8554068,2.1091962,2.8568463,3.9783216,4.698535,5.7308407,7.1232533,8.272165,17.607502,21.836184,19.963629,13.893259,8.447074,6.334448,4.722542,3.6147852,2.7333813,1.5124481,1.0014396,1.2620882,2.037175,2.702515,2.2360911,1.6084765,1.3546871,1.1523414,0.8779744,0.59674823,0.8025235,0.9362774,1.0288762,1.1043272,1.1489118,0.9774324,0.6927767,0.4938606,0.4629943,0.5521636,0.4629943,0.432128,0.4081209,0.34638834,0.17490897,0.18519773,0.20234565,0.28465575,0.45270553,0.6824879,0.5796003,0.39440256,0.4081209,0.6036074,0.64476246,0.4389872,0.3018037,0.24007112,0.23321195,0.2469303,0.7682276,1.6256244,1.7902447,1.2758065,1.1420527,1.9925903,1.8416885,1.1489118,0.40126175,0.106317215,0.030866288,0.006859175,0.01371835,0.020577524,0.006859175,0.020577524,0.0274367,0.0274367,0.034295876,0.041155048,0.034295876,0.05144381,0.12003556,0.22292319,0.31552204,0.32581082,0.45613512,0.5521636,0.59331864,0.70649505,0.8505377,0.8711152,0.9294182,1.0597426,1.1351935,1.1900668,1.0871792,0.9911508,0.94656616,0.91912943,1.2929544,1.3238207,1.3341095,1.3272504,0.9774324,1.6084765,1.4438564,1.1592005,1.0906088,1.2620882,1.1317638,1.1660597,1.2449403,1.3409687,1.5158776,1.4781522,1.4541451,1.3169615,1.1763484,1.3649758,1.1694894,1.0768905,0.99801,0.94999576,1.0460242,1.2963841,1.1934965,1.0494537,0.9774324,0.922559,0.7476501,0.91569984,0.88826317,0.6790583,0.84024894,0.7990939,0.8162418,0.84024894,0.8265306,0.72021335,0.70649505,0.7579388,0.7407909,0.65848076,0.66876954,0.58645946,0.5212973,0.5555932,0.66533995,0.70649505,0.5693115,1.0185875,1.2655178,1.1626302,1.2209331,1.255229,0.90884066,1.039165,1.5261664,1.2792361,1.5844694,2.0714707,2.2978237,2.2395205,2.2978237,2.8945718,3.216953,3.474172,3.6936657,3.7279615,3.8171308,4.249259,4.4687524,4.341858,4.139512,4.5956473,4.245829,4.2595477,4.616225,4.0880685,5.3878818,5.2815647,5.3432975,6.125243,7.160979,7.582818,7.9429245,8.032094,8.196714,9.349055,10.086417,10.041832,9.547972,8.80718,7.888051,7.455923,7.5107965,8.141841,9.084977,9.743458,10.028113,10.326488,10.350495,10.316199,10.9369545,12.905538,12.96727,12.682614,12.737488,12.950122,12.651748,12.367092,12.079007,12.065289,12.898679,13.2862215,14.291091,15.031882,15.193072,15.014734,14.592895,14.870691,15.426285,15.79325,15.46058,15.5085945,15.587475,15.446862,15.529172,16.983316,16.818697,17.353712,18.231688,19.109661,19.682402,20.316875,20.632399,21.753874,23.280039,23.300617,24.638157,27.484715,29.408712,31.854008,40.139893,37.104706,41.23393,50.661865,57.730247,49.001945,39.33051,31.51105,23.979675,17.480608,15.059319,13.3033695,11.763485,10.199594,8.628842,7.349606,6.1801167,5.422178,4.9351764,4.540774,4.0434837,3.8137012,3.7862647,3.998899,4.523626,5.4736214,5.689686,6.3138704,7.0546613,7.8023114,8.632272,8.333898,8.844906,10.155008,11.355364,10.652299,9.678296,9.750318,10.055551,10.240748,10.381361,10.432805,10.30934,9.89093,9.050681,7.641121,6.728851,5.2335505,4.4275975,4.15323,2.819121,3.1895163,2.2360911,1.4369972,1.2449403,1.0768905,0.83681935,0.8025235,0.8848336,0.9259886,0.70306545,0.6893471,0.6344737,0.59674823,0.5624523,0.4664239,0.7613684,1.2483698,2.0165975,2.8259802,3.1072063,2.7779658,2.393852,2.3252604,2.7333813,3.5633414,3.069481,4.523626,6.420188,7.5450926,6.9792104,9.626852,9.544542,9.211872,9.770895,11.029553,12.9707,14.191633,13.975569,12.662037,11.650309,9.095266,7.9257765,7.2432885,6.5642304,5.830299,5.751418,5.8543057,5.6245236,4.7945633,3.3472774,2.1434922,1.786815,1.6804979,1.371835,0.5418748,0.99801,0.7133542,0.5693115,0.65505123,0.2709374,0.5144381,0.33952916,0.106317215,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.048014224,0.14404267,0.274367,0.39440256,0.4355576,0.274367,0.59674823,1.0082988,1.3443983,1.6770682,1.9857311,2.4555845,3.0214665,3.4878905,3.5153272,3.8445675,4.1189346,4.506478,5.007198,5.4633327,5.73427,5.768566,5.65539,5.597087,5.9126086,5.751418,5.826869,5.909179,6.1286726,6.992929,6.7700057,5.7411294,5.1340923,5.188966,5.127233,5.9983487,6.5642304,6.540223,6.245279,6.608815,6.989499,7.4524937,8.47451,10.1481495,12.185325,14.284232,17.233677,19.94305,21.942501,23.376068,23.02625,23.098272,22.326614,20.755863,19.757853,20.145397,20.03908,20.172834,20.903336,22.220297,22.011093,22.422644,22.230585,21.500084,21.561817,21.290878,21.78474,23.629858,26.088871,27.11089,27.693918,27.68363,26.627317,24.994833,24.19231,25.804216,26.750782,27.752222,28.451859,27.388685,26.836521,27.241213,28.640486,30.766829,33.030357,29.388136,25.02227,23.060547,23.561266,23.52354,16.983316,16.143068,15.63206,14.157337,14.493437,9.692014,9.0644,8.532814,7.531374,8.988949,5.147811,4.523626,5.4324665,7.174697,10.048691,9.277034,12.754636,16.88043,19.428614,19.548649,17.233677,16.331696,17.480608,18.972477,16.777542,15.662926,10.9369545,8.008087,8.443645,9.993818,12.614022,11.876661,8.385342,4.897451,6.327589,7.034084,9.249598,9.14328,7.654839,10.508256,8.851766,8.580828,9.016385,9.997248,11.849225,13.824667,15.707511,15.954441,14.5414505,12.946692,12.000127,12.2093315,12.867812,13.498857,13.838386,13.594885,13.152468,12.80608,12.7272,12.97413,12.80265,12.452832,12.21962,12.027563,11.434244,11.026124,11.269625,11.393089,11.327928,11.691463,11.245617,10.655728,9.537683,8.06296,6.9654922,6.0840883,5.295283,5.0312047,5.4907694,6.632822,7.1266828,8.045813,8.752307,9.287323,10.347065,10.096705,9.160428,8.848335,9.3936405,9.935514,11.375941,12.085866,11.96926,11.516555,11.80121,13.88983,14.081886,14.208781,15.179354,16.990177,16.839275,15.854982,15.6869335,16.400288,16.479168,17.243965,16.475739,15.1862135,14.05102,13.38911,12.22305,11.393089,10.861504,10.511685,10.151579,10.271614,9.801761,9.534253,9.935514,11.132441,11.989838,12.730629,12.308789,11.026124,10.542552,9.14328,7.9600725,7.7097125,8.357904,9.112414,10.254466,11.523414,12.542002,13.152468,13.416546,12.79922,12.754636,12.854094,12.895248,12.905538,11.646879,11.355364,11.80121,12.823228,14.30481,14.5414505,15.093615,14.695783,13.488567,13.035862,12.96727,12.583157,11.938394,10.947243,9.373062,8.834618,9.523964,10.31277,10.772334,11.153018,9.331907,8.786603,9.006097,9.3593445,9.095266,8.940934,9.033533,9.448513,9.873782,9.595985,8.992378,8.98209,9.218731,9.547972,9.9801,9.705732,10.007536,10.436234,10.731179,10.827208,10.532263,9.743458,9.218731,9.256456,9.6988735,10.295622,10.401938,10.034973,9.489669,9.3079,8.762596,8.014946,8.128122,9.263316,10.696883,0.4424168,0.4664239,0.5178677,0.5418748,0.53158605,0.5178677,0.7373613,0.764798,0.6859175,0.64819205,0.85396725,0.7579388,0.86082643,1.0117283,1.1694894,1.3889829,1.3272504,1.1832076,1.1832076,1.2998136,1.2517995,1.0940384,0.9534253,0.9294182,0.9774324,0.91569984,0.9774324,1.1111864,1.1283343,1.0734608,1.2209331,1.3443983,1.4095604,1.4232788,1.4815818,1.8005334,1.6427724,1.903421,2.177788,2.4898806,3.2958336,4.32128,4.979761,6.3481665,8.738589,11.701753,22.384918,24.10314,18.224829,9.301042,5.0655007,5.7377,4.9077396,3.450165,2.0028791,0.9774324,0.805953,1.1283343,1.4781522,1.5158776,1.0528834,1.0288762,1.3169615,1.3581166,1.0254467,0.61046654,0.90198153,0.939707,0.90198153,0.8779744,0.85396725,0.9294182,0.7990939,0.66533995,0.6001778,0.5658819,0.41840968,0.4355576,0.47328308,0.41840968,0.19891608,0.20920484,0.16804978,0.16119061,0.24350071,0.42869842,0.59674823,0.4938606,0.29837412,0.14404267,0.106317215,0.106317215,0.08916927,0.06516216,0.05144381,0.07545093,0.83338976,1.7902447,1.8999915,1.3238207,1.4335675,2.5070283,2.0714707,1.1008976,0.29151493,0.044584636,0.010288762,0.017147938,0.041155048,0.0548734,0.030866288,0.0548734,0.06859175,0.082310095,0.09259886,0.09259886,0.09259886,0.12689474,0.17833854,0.24007112,0.34981793,0.36353627,0.4938606,0.59674823,0.65848076,0.7922347,0.82996017,1.0048691,1.0906088,1.039165,0.9774324,0.90198153,0.82996017,0.6276145,0.48014224,0.8711152,0.9911508,1.0220171,1.0048691,0.9294182,0.7339317,1.8931323,1.4129901,1.0768905,1.2483698,0.8711152,1.1008976,1.2415106,1.4678634,1.7971039,2.0920484,1.8965619,1.6633499,1.1797781,0.75450927,1.2037852,1.0597426,0.91227025,0.91912943,0.9842916,0.77851635,1.0460242,1.1420527,1.1180456,1.08032,1.1900668,1.0563129,0.9774324,0.9945804,1.1214751,1.3272504,1.0357354,0.90541106,0.881404,0.91569984,0.9774324,0.70649505,0.59674823,0.6001778,0.6927767,0.84024894,0.66876954,0.48014224,0.5590228,0.805953,0.7339317,0.7682276,1.0425946,1.0734608,0.84367853,0.7922347,1.0631721,0.96371406,1.0014396,1.1214751,0.71678376,1.1214751,1.8073926,2.253239,2.2978237,2.1503513,2.651071,3.2718265,3.8137012,4.0846386,3.875434,4.266407,3.998899,4.0537724,4.540774,4.698535,4.3590055,4.4996185,4.5270553,4.2355404,3.8445675,5.3090014,4.4756117,4.756838,6.341307,6.193835,7.085528,7.4936485,7.9086285,8.556821,9.400499,9.55826,9.89093,9.9869585,9.561689,8.436785,8.669997,9.650859,10.621432,11.050131,10.635151,10.978109,11.365653,11.290202,10.899229,10.984968,12.425395,13.207341,13.245067,12.812939,12.55915,11.897239,11.561139,11.828648,12.764925,14.205351,14.033872,14.359683,15.018164,15.601193,15.443433,15.429714,15.700651,16.335125,16.606062,14.983868,15.470869,16.005884,16.911295,18.1288,19.239986,18.95876,19.613811,20.179693,20.388897,20.70442,22.02481,23.077694,24.308916,25.656744,26.534718,28.585611,30.204376,32.478195,36.305614,42.434284,38.246758,42.08104,48.07596,50.017105,41.33682,33.157253,27.909983,23.636717,19.771572,17.134218,15.182784,13.193623,11.228469,9.3764925,7.750868,6.6396813,5.7308407,4.9248877,4.190956,3.5564823,3.2375305,3.450165,3.974892,4.6436615,5.3398676,5.878313,6.7459984,7.514226,8.107545,8.803751,10.086417,11.211322,11.681175,11.509696,11.214751,10.981539,11.574858,11.794352,11.640019,12.298501,13.238208,12.713481,11.406808,9.791472,8.117833,6.8728933,5.8371577,4.887162,3.9543142,3.0523329,3.1380725,2.253239,1.4404267,1.0906088,0.9294182,0.90541106,0.83681935,0.85396725,0.922559,0.823101,0.66533995,0.66191036,0.6310441,0.5521636,0.5658819,0.5144381,0.70649505,0.9602845,1.2895249,1.862266,2.3149714,2.452155,3.508468,5.0655007,5.0655007,4.0537724,3.9646032,5.295283,7.798882,10.48082,11.80121,11.231899,10.251037,9.846346,10.528833,9.246168,8.285883,8.327039,8.755736,7.6445503,6.351596,6.0086374,5.888602,6.0497923,7.3530354,7.8537555,7.157549,5.8988905,4.506478,3.1895163,2.393852,2.6819375,2.4761622,1.430138,0.4424168,0.490431,0.84367853,0.8711152,0.6001778,0.6859175,0.7339317,0.36353627,0.06516216,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.08916927,0.08916927,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.1371835,0.2469303,0.34638834,0.42183927,0.51100856,0.71678376,1.0700313,1.0768905,1.0666018,1.2860953,1.9068506,2.0920484,2.411,2.7093742,2.819121,2.5619018,2.784825,3.340418,4.396731,5.610805,6.135532,6.0737996,6.2212715,6.800872,7.548522,7.706283,7.3530354,7.8777623,8.182996,8.405919,9.932085,8.772884,6.944915,6.4407654,7.0786686,6.5299344,8.495089,8.786603,8.371623,8.23444,9.369633,8.868914,9.191295,10.010965,11.30735,13.38225,16.21509,19.438902,21.434921,22.10712,22.889067,21.825895,22.247734,22.919933,23.27318,23.406935,22.8582,21.740154,20.989075,21.02337,21.743584,21.53781,21.630407,21.04395,20.12139,20.522652,20.241425,21.232576,23.571554,26.10945,26.490133,26.466127,27.26522,27.203487,26.229485,25.924252,26.706198,27.021719,28.211786,29.635065,28.67135,25.52299,25.310356,28.479294,33.520786,36.988102,33.41104,27.957996,23.44809,21.839613,24.230036,24.497543,22.745024,19.52807,15.981877,13.810948,10.367643,11.228469,13.437123,15.093615,15.350834,12.260776,11.993267,12.47341,13.173045,15.090185,14.308239,12.905538,12.905538,14.507155,16.081335,19.390888,17.04162,15.014734,15.398848,16.386568,7.051232,5.9228973,6.992929,7.5039372,7.98065,4.6127954,3.450165,3.8960114,5.425607,7.599966,7.548522,5.586798,6.029215,8.213862,6.5162163,6.931196,7.0786686,7.14726,7.455923,8.467651,9.993818,12.188754,13.7697935,14.092175,13.152468,10.871792,10.655728,11.365653,12.140739,12.421966,13.018714,12.912396,12.593445,12.325937,12.130451,12.593445,13.296511,13.862392,14.071597,13.838386,13.313659,13.5503,14.027013,14.13333,13.169616,11.567999,10.573419,9.938945,9.235879,7.857185,6.23499,5.1409516,4.557922,4.506478,5.0826488,5.8988905,6.927767,7.829748,8.320179,8.1487,8.711152,8.831187,9.472521,10.717461,11.780633,12.782072,12.764925,11.893809,10.738038,10.299051,11.214751,11.592006,12.346515,13.80409,15.6697855,15.755525,15.577187,15.6869335,15.9921665,15.748666,16.2974,16.80155,16.194511,14.620332,13.413116,12.71691,12.22305,12.05157,11.955542,11.321068,10.6145735,10.7586155,11.276484,11.780633,11.962401,12.048141,12.435684,11.763485,10.14129,9.139851,9.126132,7.805741,7.140401,7.5759587,8.025234,8.368194,9.074688,10.456812,12.229909,13.5503,14.575747,14.942713,14.335675,13.234778,12.895248,11.149589,10.923236,12.229909,14.575747,16.96617,16.431154,15.179354,13.087306,11.255906,12.024134,12.401388,12.349944,11.794352,10.923236,10.179015,9.932085,10.511685,11.214751,11.691463,11.948683,10.408798,9.098696,8.680285,8.800322,8.117833,8.766026,9.098696,9.496528,9.863494,9.644,10.350495,10.518545,10.316199,10.028113,10.041832,10.333347,10.652299,10.988399,11.132441,10.679735,10.569988,10.261326,10.2236,10.429376,10.347065,10.065839,10.388221,10.491108,10.347065,10.710602,9.3936405,8.038953,7.795452,8.889491,10.635151,0.34638834,0.4389872,0.5521636,0.6824879,0.8128122,0.89855194,0.864256,0.7888051,0.7339317,0.72364295,0.7442205,0.72364295,0.8848336,0.9877212,0.9945804,1.0460242,1.1043272,1.1283343,1.1317638,1.0940384,0.9568549,0.9362774,0.9328478,0.96714365,1.0014396,0.939707,0.9911508,1.2312219,1.3238207,1.2689474,1.4164196,1.488441,1.3752645,1.2758065,1.3101025,1.5193073,1.5261664,1.9685832,2.3561265,2.8739944,4.383013,4.928317,5.5422134,6.883182,9.506817,13.838386,19.812727,20.128248,15.501736,8.783174,4.9694724,4.897451,4.6436615,3.7965534,2.469303,1.3066728,0.77508676,0.72707254,0.8162418,0.864256,0.8711152,1.0700313,1.2586586,1.1317638,0.7339317,0.47671264,0.58302987,0.6036074,0.66876954,0.8196714,1.0014396,1.1146159,0.9294182,0.72707254,0.6310441,0.61389613,0.45613512,0.5761707,0.65505123,0.53844523,0.20920484,0.12346515,0.09602845,0.082310095,0.15776102,0.47671264,0.78537554,0.64819205,0.3841138,0.17833854,0.09602845,0.044584636,0.058302987,0.10288762,0.14061308,0.12346515,0.5418748,1.1351935,1.3375391,1.1694894,1.2380811,2.2841053,1.9514352,1.0837497,0.31552204,0.06859175,0.01371835,0.0034295875,0.006859175,0.01371835,0.017147938,0.024007112,0.0274367,0.034295876,0.05144381,0.09259886,0.13032432,0.1920569,0.2469303,0.274367,0.2777966,0.29837412,0.37382504,0.53844523,0.70306545,0.67219913,1.0014396,1.0494537,0.96371406,0.8505377,0.78194594,0.7682276,0.7305021,0.53501564,0.33952916,0.61389613,0.66876954,0.78194594,0.9877212,1.1626302,1.0254467,1.7559488,1.3581166,1.2380811,1.4918705,0.91912943,1.1317638,1.3032433,1.4644338,1.6427724,1.845118,1.4850113,1.4541451,1.3752645,1.155771,0.9602845,1.0700313,0.9568549,0.85396725,0.84024894,0.8265306,0.96714365,1.1283343,1.2380811,1.2620882,1.1763484,1.1523414,1.155771,1.2346514,1.3203912,1.255229,1.2243627,1.1694894,1.097468,0.9945804,0.82996017,0.58988905,0.5796003,0.607037,0.61046654,0.66876954,0.45956472,0.59674823,0.7099246,0.6893471,0.6962063,0.8196714,1.0940384,1.2037852,1.1249046,1.1351935,1.2380811,1.1351935,1.08032,1.1523414,1.2655178,1.3169615,1.4541451,1.6324836,1.9651536,2.7368107,2.6133456,3.0557625,3.4021509,3.5290456,3.8377085,4.2595477,4.1429415,4.3590055,4.822,4.4927597,5.0106273,5.40503,5.439326,5.188966,5.0414934,5.4016004,4.9008803,4.9934793,5.610805,5.1683884,6.090947,6.958633,7.610255,8.189855,9.119273,8.652849,9.084977,9.201583,8.886061,9.122703,9.72631,10.412228,10.88894,10.930096,10.377932,10.7586155,11.129011,10.971251,10.436234,10.326488,11.797781,13.426835,14.291091,14.153908,13.498857,12.830087,12.30536,12.147599,12.576297,13.80409,14.246507,14.96672,15.666355,16.084764,16.016174,16.160215,16.256245,16.564907,16.87014,16.486027,16.486027,16.846134,17.319416,17.96761,19.154245,18.962189,20.430052,21.62012,21.884197,21.829325,23.266321,24.19231,25.69104,27.546446,28.26666,30.317553,32.217545,35.729443,40.5,44.070198,47.266575,53.03857,52.266914,44.468033,37.82149,31.984333,27.17605,23.19087,20.464348,20.052797,18.001905,15.319967,12.809509,10.823778,9.290752,8.375052,7.380472,6.3893213,5.442755,4.5442033,4.098357,3.9886103,4.170378,4.664239,5.535354,6.3173003,6.783724,7.6342616,8.937505,10.110424,10.367643,11.015835,11.945253,12.826657,13.118172,13.354814,13.3033695,13.107883,13.183334,14.21564,14.754086,13.697772,11.506266,9.091836,7.798882,6.574519,5.8165803,4.996909,4.0194764,3.234101,2.4898806,2.07833,1.6736387,1.2655178,1.1763484,1.4815818,1.786815,1.8759843,1.6633499,1.214074,0.9877212,0.9294182,0.84024894,0.71678376,0.7613684,0.88826317,0.96714365,1.0460242,1.371835,2.386993,2.7779658,2.7745364,3.199805,3.8514268,3.4913201,4.098357,4.2835546,4.3692946,4.8768735,6.526505,7.613684,7.373613,7.298162,7.582818,7.133542,7.6616983,7.829748,7.7577267,7.4799304,6.9723516,6.3035817,7.3873315,8.913498,9.956093,9.942374,7.7783046,6.3173003,4.887162,3.4638834,2.6647894,2.3595562,2.4761622,2.2395205,1.4198492,0.34638834,0.29494452,0.44584638,0.4664239,0.3841138,0.5761707,1.1934965,0.64476246,0.106317215,0.0,0.0,0.0,0.0,0.010288762,0.082310095,0.30866286,0.26407823,0.22635277,0.1371835,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16462019,0.37725464,0.22292319,0.45956472,0.6790583,0.82996017,0.91569984,0.99801,1.0288762,1.2620882,1.3272504,1.2415106,1.3958421,1.6256244,1.7525192,1.978872,2.2498093,2.2463799,2.4761622,3.1963756,4.0674906,4.835718,5.3398676,6.2658563,6.728851,6.5367937,6.3207297,7.5210853,8.056101,9.434795,9.084977,7.5107965,8.272165,7.864044,6.6053853,6.48535,7.5450926,7.8846216,8.210432,8.923786,9.263316,9.091836,8.930646,9.14328,9.746887,10.950673,13.025573,16.311117,19.143957,20.714708,21.314886,21.3629,21.410915,19.569225,18.95876,19.919044,21.884197,23.393215,24.212887,23.729315,23.86307,24.593573,23.976246,21.825895,20.982216,20.78673,20.666695,20.131678,20.35803,21.647556,23.211449,24.466677,25.001692,25.296637,25.797358,26.370098,26.67876,26.167753,28.853119,29.717375,29.727665,29.84427,31.037767,29.168642,30.904013,38.66174,51.37522,64.50025,70.85528,60.8546,45.503765,34.216995,34.800022,34.062664,30.26268,24.240324,18.358582,16.520323,19.003344,19.421753,19.075365,18.37573,16.815268,14.448852,18.307138,17.329706,11.746337,13.077017,10.635151,10.353925,10.792912,11.780633,14.411126,18.20768,16.62321,13.646329,11.358793,9.956093,4.6608095,5.209543,6.7871537,7.1198235,6.492209,6.4716315,6.64997,6.958633,7.490219,8.501947,8.539673,8.117833,8.035523,8.100685,7.1266828,6.7802944,6.694555,6.7185616,6.8385973,7.1884155,8.196714,10.539123,13.090735,14.699212,14.177915,12.257345,11.423956,11.331357,11.653738,12.092726,12.620882,13.128461,13.594885,14.033872,14.46257,15.7966795,16.492886,17.20967,17.689812,16.79469,16.2974,15.7795315,15.097044,14.112752,12.679185,11.1393,10.460241,10.436234,10.381361,9.126132,7.7783046,6.4819202,5.5319247,5.103226,5.2781353,5.6656785,5.98463,6.447624,7.14726,8.049242,8.114404,8.7283,10.031544,11.701753,12.939834,12.932974,12.456262,11.660598,10.789482,10.151579,11.067279,11.290202,12.017275,13.5503,15.278812,14.428274,14.315098,14.520873,14.603184,14.088745,14.520873,15.395418,15.542891,14.740367,13.718349,13.920695,13.152468,12.723769,12.816368,12.493987,11.989838,11.746337,11.814929,12.027563,11.986408,11.986408,11.451392,10.381361,9.246168,8.968371,9.054111,7.888051,7.250148,7.905199,9.623423,8.824328,8.879202,9.853205,11.578287,13.660047,14.754086,14.55174,13.9138365,13.533153,13.944703,13.485138,13.3033695,13.697772,14.730078,16.235666,14.634049,13.056439,11.986408,11.55428,11.571428,11.4033785,11.427385,11.019264,10.196163,9.626852,9.472521,9.225591,9.5205345,10.377932,11.190743,10.679735,9.2153015,8.447074,8.601405,8.484799,8.964942,9.595985,10.113853,10.4533825,10.741467,10.765475,10.748327,10.511685,10.076128,9.637141,10.456812,10.762046,10.751757,10.504827,9.9869585,9.434795,9.438225,10.014396,10.693454,10.528833,10.532263,10.14129,10.024684,10.477389,11.4205265,10.422516,9.098696,8.203573,8.14527,8.961512,0.4664239,0.53158605,0.72707254,0.91569984,1.0597426,1.2312219,1.0151579,0.90541106,0.8505377,0.8196714,0.77165717,0.90541106,1.0185875,1.0254467,0.980862,1.0906088,1.1660597,1.2380811,1.2723769,1.255229,1.1694894,1.138623,1.138623,1.1694894,1.2106444,1.2312219,1.2860953,1.3752645,1.3752645,1.3032433,1.3169615,1.2689474,1.3032433,1.3924125,1.4781522,1.4850113,1.6530612,2.3252604,2.8328393,3.3472774,4.863155,4.822,5.442755,7.1541195,9.949233,13.38568,18.804428,18.759844,15.319967,10.316199,5.336438,4.2081037,3.474172,2.7745364,2.0474637,1.5261664,0.9774324,0.7305021,0.6379033,0.6276145,0.70649505,1.0494537,1.1934965,1.0288762,0.6859175,0.52472687,0.64476246,0.65848076,0.71678376,0.85396725,0.9911508,0.939707,0.7133542,0.5693115,0.548734,0.48014224,0.33609957,0.4115505,0.45956472,0.36353627,0.14061308,0.058302987,0.041155048,0.037725464,0.10288762,0.37039545,0.7476501,0.7613684,0.58988905,0.37039545,0.1920569,0.1097468,0.14061308,0.18862732,0.18519773,0.1097468,0.24007112,0.58645946,0.84024894,0.94999576,1.1077567,1.9548649,1.7250825,1.0220171,0.34295875,0.07545093,0.024007112,0.0034295875,0.0034295875,0.006859175,0.006859175,0.01371835,0.037725464,0.044584636,0.05144381,0.12689474,0.12689474,0.12003556,0.12003556,0.14061308,0.20577525,0.24350071,0.36696586,0.4938606,0.6001778,0.7339317,0.9877212,1.0048691,0.82996017,0.6893471,0.9602845,0.6036074,0.5796003,0.5658819,0.47328308,0.42869842,0.58302987,0.71678376,1.0460242,1.3478279,0.9602845,1.6496316,1.3684053,1.4918705,1.9480057,1.214074,1.4438564,1.2826657,1.1592005,1.2415106,1.4472859,1.1694894,1.2929544,1.3546871,1.196926,0.9842916,0.8676856,0.922559,0.94656616,0.89512235,0.89512235,1.0494537,1.0117283,1.0425946,1.1729189,1.2209331,1.4267083,1.2792361,1.1934965,1.2449403,1.1626302,1.2346514,1.0768905,0.9328478,0.864256,0.7476501,0.5453044,0.490431,0.5007198,0.5041494,0.45270553,0.42183927,0.69963586,0.77165717,0.58645946,0.5693115,0.5761707,0.8265306,1.0117283,1.0185875,0.91912943,0.9945804,0.97057325,0.88826317,0.8711152,1.1283343,1.2312219,1.2346514,1.3478279,1.5947582,1.8142518,1.9274281,2.6304936,3.0969174,3.2478194,3.782835,4.1600895,3.940596,4.057202,4.540774,4.523626,5.007198,5.5833683,5.5662203,4.996909,4.65395,4.5784993,5.329579,5.8543057,5.885172,5.919468,6.392751,6.800872,7.298162,7.8949103,8.443645,7.864044,8.152129,8.412778,8.553391,9.266746,9.880642,10.611144,11.019264,10.978109,10.672876,10.316199,10.2236,10.127572,10.134431,10.738038,11.492548,12.857523,14.243076,15.028452,14.565458,14.085316,13.577737,13.560589,14.174485,15.175924,15.481158,16.002455,16.314548,16.300829,16.149927,16.969599,17.151367,17.28512,17.63494,18.132229,18.025911,18.560926,19.36688,20.183123,20.855322,20.779871,22.264881,23.44809,23.914513,24.69303,25.10115,26.140316,27.741934,29.525318,30.814844,32.697685,34.947495,38.80921,43.775253,47.582096,55.933144,64.41108,62.247013,51.11457,45.099075,38.363365,30.458166,24.699888,22.374628,22.741594,20.073376,17.257685,14.788382,12.932974,11.742908,10.899229,9.757176,8.508806,7.39762,6.742569,5.977771,5.535354,5.442755,5.744559,6.4990683,7.208993,7.6205435,8.30646,9.345626,10.319629,10.604284,12.343085,14.2190695,15.402277,15.563468,14.476289,13.443983,12.723769,12.507706,12.936404,11.441104,9.685155,7.840037,6.293293,5.662249,6.001778,5.3981705,4.712253,4.2766957,3.8925817,3.000889,2.5413244,2.170929,1.8073926,1.646202,2.287535,2.277246,2.0508933,1.7730967,1.3409687,1.2037852,1.2346514,1.2620882,1.1900668,0.9842916,0.9259886,0.89512235,0.9534253,1.2723769,2.1332035,2.3218307,2.07833,2.1572106,2.5070283,2.2360911,3.2512488,3.8171308,4.664239,5.802862,6.5367937,8.073249,8.035523,7.596536,7.250148,6.8283086,8.303031,8.858624,8.56368,7.864044,7.5759587,7.4799304,8.405919,10.443094,12.257345,11.101575,7.932636,5.9743414,4.2183924,2.668219,2.3046827,5.56965,5.5113473,3.6182148,1.3889829,0.31895164,0.18176813,0.58988905,0.65505123,0.4424168,0.97057325,1.5227368,0.86082643,0.21263443,0.037725464,0.0,0.0,0.0,0.0034295875,0.058302987,0.23664154,0.21263443,0.16462019,0.09259886,0.0274367,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.216064,0.4972902,0.33609957,0.764798,0.85739684,0.922559,1.0117283,0.91227025,0.96714365,1.3101025,1.4027013,1.1592005,0.9568549,1.2929544,1.5090185,1.6599203,1.8759843,2.3389788,2.3389788,2.527606,2.867135,3.357566,4.033195,4.9934793,5.0346346,4.852866,4.99005,5.8371577,6.0806584,7.1198235,7.4181976,6.831738,6.6122446,6.883182,6.6465406,7.2432885,8.364764,8.076678,7.932636,8.652849,9.5205345,9.89093,9.167287,9.054111,9.887501,11.077567,12.912396,16.568336,19.099373,19.709839,20.344313,20.965069,19.54179,18.6158,17.940172,18.12537,19.411465,21.671564,22.44322,22.549538,23.52697,24.888515,24.140865,22.412354,21.53438,21.332033,21.493225,21.544668,21.253153,21.476076,21.575535,21.434921,21.45893,22.673002,23.78419,25.121729,26.119738,25.324074,27.673342,29.419,29.964306,29.463587,28.829113,30.722244,36.792614,47.60953,63.159283,82.84168,103.99881,98.58006,74.57981,48.31603,44.420017,44.258827,38.692604,31.93632,26.747353,24.411804,23.574984,22.583834,22.041958,21.393766,18.948471,18.008764,16.108772,13.011855,10.110424,10.422516,9.235879,9.211872,9.174147,9.410788,11.694893,12.442543,12.415107,11.705182,10.113853,7.174697,5.2335505,5.6245236,6.118384,6.1321025,6.7219915,7.956643,8.056101,8.165848,8.587687,8.772884,8.776315,8.601405,8.453933,8.323608,7.98408,7.5931067,7.3873315,7.1987042,7.0135064,6.9860697,7.5725293,9.14328,11.324498,13.248496,13.574307,12.277924,11.399949,10.933525,10.89237,11.341646,11.955542,12.71691,13.612033,14.627191,15.731518,17.947031,19.510923,20.838173,21.585823,20.652975,19.922474,18.588364,16.763824,14.764374,13.13532,12.055,11.71547,11.506266,11.087856,10.377932,9.551401,8.659708,7.8983397,7.2295704,6.385892,6.3618846,6.090947,5.9297566,6.1801167,7.1095347,7.3701835,7.939495,9.256456,10.998687,12.075578,12.157887,11.869802,11.2593355,10.573419,10.264755,10.782623,10.827208,11.423956,12.80608,14.4145565,14.126471,14.177915,14.198492,13.941273,13.306799,13.7526455,14.5585985,15.093615,15.0250225,14.29795,13.876111,13.145609,13.190193,13.817808,13.574307,13.121602,12.408247,12.027563,12.089295,12.202472,12.202472,11.149589,10.134431,9.637141,9.530824,8.4093485,7.531374,7.366754,8.124693,9.767465,8.851766,8.440215,8.752307,10.028113,12.524854,14.740367,14.778092,14.627191,15.073037,15.6697855,15.316538,14.836395,14.870691,15.278812,15.155347,13.454271,12.212761,12.024134,12.511135,12.346515,11.9040985,11.502836,11.111863,10.518545,9.373062,9.465661,9.205012,9.3079,9.938945,10.700313,10.082987,9.283894,8.985519,9.156999,9.043822,9.263316,9.554831,9.80519,10.010965,10.302481,10.419086,10.504827,10.515115,10.203023,9.088407,9.80519,10.072699,10.021255,9.740028,9.263316,8.903209,9.108984,9.774324,10.549411,10.858074,10.412228,9.884071,9.788043,10.360784,11.578287,11.513125,10.422516,8.745448,7.486789,8.23444,0.53501564,0.58645946,0.8162418,0.97400284,1.0528834,1.3032433,1.138623,1.0288762,0.9362774,0.8505377,0.78537554,1.0323058,1.0220171,0.9431366,0.91569984,0.9842916,1.0837497,1.2312219,1.3341095,1.3649758,1.3752645,1.2723769,1.2277923,1.2175035,1.2483698,1.371835,1.5193073,1.4987297,1.4164196,1.3512574,1.3615463,1.2723769,1.3821237,1.5158776,1.611906,1.7113642,2.0234566,2.651071,3.0797696,3.40901,4.3590055,4.448175,5.23698,7.0752387,9.925226,13.37882,19.349733,19.438902,16.026463,10.8958,5.2266912,3.666229,2.7093742,2.095478,1.670209,1.3855534,1.0597426,0.94999576,0.82996017,0.70306545,0.7956643,1.1694894,1.1249046,0.89855194,0.66533995,0.53844523,0.607037,0.65162164,0.78194594,0.9842916,1.1317638,0.864256,0.53158605,0.3841138,0.40126175,0.3018037,0.24007112,0.25378948,0.23664154,0.15776102,0.072021335,0.0274367,0.01371835,0.0274367,0.1097468,0.37382504,0.77165717,0.84367853,0.7133542,0.48700142,0.26407823,0.14404267,0.1371835,0.15433143,0.1371835,0.061732575,0.06516216,0.274367,0.5555932,0.83681935,1.1214751,1.7216529,1.6221949,1.0837497,0.4389872,0.09602845,0.0274367,0.0034295875,0.0034295875,0.006859175,0.0,0.006859175,0.030866288,0.037725464,0.041155048,0.10288762,0.08573969,0.058302987,0.037725464,0.048014224,0.11317638,0.14747226,0.26407823,0.37382504,0.45270553,0.53844523,0.764798,0.7579388,0.59331864,0.5521636,1.0940384,0.5521636,0.5007198,0.5212973,0.45956472,0.42526886,0.66191036,0.65162164,0.8779744,1.2037852,0.864256,1.2380811,1.2723769,1.4541451,1.6427724,1.0631721,1.4232788,1.1523414,0.97400284,1.097468,1.2449403,1.2072148,1.2209331,1.1832076,1.0940384,1.0563129,0.89855194,1.0837497,1.1180456,0.94999576,0.97400284,1.0631721,0.881404,0.89169276,1.1489118,1.3066728,1.5124481,1.3101025,1.1214751,1.0940384,1.0906088,1.2175035,1.1249046,1.0151579,0.91569984,0.6927767,0.5624523,0.45613512,0.4389872,0.47328308,0.432128,0.490431,0.6344737,0.61046654,0.48700142,0.64819205,0.4938606,0.72707254,0.881404,0.8162418,0.70649505,0.84367853,1.0220171,0.97057325,0.78537554,0.91569984,0.9945804,1.1043272,1.2346514,1.3684053,1.4644338,1.6667795,2.2360911,2.5824795,2.7642474,3.4776018,3.7279615,3.6936657,3.7725463,4.1292233,4.712253,4.9523244,4.979761,4.996909,4.9488945,4.5442033,4.3349986,5.7479887,6.5710897,6.416758,6.725421,7.250148,7.0718093,7.414768,8.275595,8.412778,8.841476,9.482809,9.517105,9.136421,9.5205345,9.770895,10.494537,10.827208,10.635151,10.508256,10.106995,10.017825,9.846346,9.860064,10.988399,11.458252,12.164746,13.4645605,14.867262,15.018164,15.138199,15.206791,15.230798,15.505165,16.592344,16.750105,17.099922,16.973028,16.410576,16.13278,17.480608,17.984756,18.163095,18.430603,19.12681,19.661825,20.697561,21.908205,22.751883,22.474087,22.933651,24.164873,24.905664,25.286348,26.815945,26.514141,27.94085,29.789396,31.445887,33.02007,36.0724,38.130154,41.861546,47.657547,53.61817,61.19413,67.264496,64.455666,54.715637,49.30375,41.954144,32.99606,26.76107,24.394655,23.852781,20.632399,18.077356,16.156786,14.815818,13.965281,13.88297,12.401388,10.744898,9.633711,9.31133,8.255017,7.7748747,7.7268605,8.097256,8.985519,9.163857,9.458802,10.055551,10.837497,11.372512,11.674315,13.989287,15.951012,16.345413,15.107333,12.655178,11.423956,10.545981,9.702303,9.105555,6.509357,4.7671266,3.7211025,3.234101,3.1826572,4.139512,4.0194764,3.875434,3.99204,3.8891523,3.3850029,3.0557625,2.7402403,2.386993,2.0440342,2.4418662,2.4144297,2.1812177,1.8416885,1.3889829,1.4850113,1.6084765,1.6907866,1.5810398,1.0494537,0.7990939,0.70306545,0.7922347,1.1077567,1.6942163,1.7113642,1.4027013,1.546744,2.2498093,2.9322972,4.3007026,4.5339146,5.892031,8.423067,9.966381,10.220171,10.669447,10.518545,9.606275,8.4264965,9.6645775,9.527394,8.80718,8.158989,8.073249,7.7851634,7.8263187,9.764035,12.243628,11.012405,7.8503256,5.7479887,4.057202,2.8945718,3.1140654,7.6685576,7.0306544,4.3007026,1.6427724,0.29151493,0.31552204,0.94656616,1.0425946,0.72364295,1.3478279,1.3581166,0.71678376,0.1920569,0.037725464,0.0,0.0,0.017147938,0.0274367,0.037725464,0.08916927,0.09259886,0.06516216,0.037725464,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.034295876,0.2469303,0.490431,0.30523327,0.8128122,0.8162418,0.77165717,0.84024894,0.8711152,0.939707,1.1249046,1.1454822,0.9362774,0.64476246,1.2277923,1.3855534,1.3341095,1.3375391,1.6873571,1.937717,1.8519772,1.9342873,2.3252604,2.8259802,3.5942078,3.5221863,3.5221863,3.957744,4.6608095,4.338428,4.972902,5.7479887,6.0223556,5.336438,5.5902276,6.427047,7.4181976,8.018375,7.5759587,7.332458,8.351046,9.325048,9.702303,9.668007,9.3593445,10.38479,11.667457,13.197053,16.029892,17.751545,18.975908,19.912186,20.207129,18.924463,19.03764,19.548649,19.387459,19.143957,21.061096,21.129688,20.752434,21.061096,21.908205,21.884197,21.887627,21.921923,21.94936,21.94593,21.894485,21.647556,21.397196,20.430052,19.342873,20.049368,21.815605,22.87192,24.058556,25.056566,24.401514,25.495554,26.709627,27.323523,27.158903,26.582733,35.887203,46.5395,57.582775,69.04102,81.90541,100.809296,104.25946,86.8543,59.582222,49.80447,50.87793,45.037342,38.030697,33.644253,33.705986,26.68562,23.547548,22.930222,23.053686,21.729866,18.78042,12.747777,8.793462,8.114404,7.9737906,8.4093485,8.39563,8.086967,7.936065,8.721441,7.486789,8.351046,9.163857,8.56025,5.9434752,5.5422134,5.7719955,5.744559,5.693115,6.9654922,8.22758,8.056101,8.30646,9.218731,9.414218,9.582268,9.547972,9.438225,9.335337,9.294182,9.006097,8.875772,8.56025,8.008087,7.442205,7.431916,7.915488,9.263316,10.981539,11.701753,11.077567,10.446524,9.908078,9.644,9.918367,10.597425,11.513125,12.679185,14.126471,15.913286,18.169954,19.901896,21.417774,22.288889,21.338894,20.60839,19.44919,17.730967,15.810398,14.527733,13.900118,13.7938,13.289652,12.240198,11.2593355,10.748327,10.220171,9.626852,8.762596,7.284444,6.8900414,6.276145,5.768566,5.7308407,6.5539417,7.373613,7.949784,9.105555,10.624862,11.252477,11.698323,11.362224,10.714031,10.340206,10.933525,11.05356,10.912948,11.190743,12.185325,13.814379,13.066729,13.306799,13.756075,13.780083,12.891819,13.443983,14.123041,14.603184,14.637479,14.04759,12.9809885,12.4802685,13.190193,14.476289,14.441993,14.078457,13.090735,12.38767,12.264205,12.397959,11.97269,11.084427,10.573419,10.436234,9.8429165,8.388771,7.6274023,7.466212,7.840037,8.738589,7.840037,7.1884155,7.4627824,8.992378,11.780633,14.435134,15.076467,15.251375,15.6252,15.971589,15.265094,14.376831,14.232788,14.46943,13.426835,12.421966,12.47341,13.358243,14.239647,13.690913,13.035862,12.13731,11.4754,10.940384,9.836057,9.767465,9.6817255,9.9869585,10.662587,11.266195,10.161868,9.578837,9.455373,9.513676,9.239308,9.80519,9.767465,9.554831,9.47938,9.740028,10.189304,10.415657,10.532263,10.244178,8.844906,9.019815,9.012956,9.054111,9.115844,8.920357,8.663138,8.834618,9.431366,10.353925,11.396519,10.549411,10.364213,10.336777,10.597425,11.907528,12.624311,11.324498,9.009526,7.31531,8.525954,0.5007198,0.5521636,0.7510797,0.84367853,0.86082643,1.1283343,1.1214751,1.039165,0.9362774,0.8505377,0.805953,1.0666018,0.939707,0.8196714,0.823101,0.7613684,0.9568549,1.2243627,1.3478279,1.3306799,1.3992717,1.2277923,1.1729189,1.1592005,1.2037852,1.4129901,1.6530612,1.611906,1.4953002,1.4404267,1.529596,1.5158776,1.5501735,1.5844694,1.704505,2.1263442,2.486451,2.8019729,2.935727,2.983741,3.2821152,4.1635194,5.209543,6.893471,9.877212,15.001016,20.676983,20.45406,16.067617,9.860064,4.787704,3.3987212,2.6716487,2.1743584,1.6633499,1.0734608,1.0048691,1.1626302,1.1351935,0.94999576,1.097468,1.3272504,1.0494537,0.77508676,0.66533995,0.53501564,0.52472687,0.5658819,0.78194594,1.1283343,1.3786942,0.9877212,0.5418748,0.29494452,0.2503599,0.17147937,0.21263443,0.19548649,0.13375391,0.06516216,0.044584636,0.020577524,0.017147938,0.030866288,0.12003556,0.4081209,0.71678376,0.71678376,0.58645946,0.42869842,0.28465575,0.13375391,0.048014224,0.024007112,0.034295876,0.020577524,0.08916927,0.23664154,0.47328308,0.7990939,1.1797781,1.6290541,1.704505,1.2929544,0.6001778,0.13375391,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.044584636,0.0548734,0.058302987,0.0548734,0.044584636,0.048014224,0.09602845,0.22635277,0.33266997,0.16119061,0.47328308,0.5007198,0.38754338,0.4046913,0.9294182,0.5590228,0.4424168,0.33952916,0.29837412,0.64819205,0.7682276,0.58645946,0.58988905,0.7922347,0.75450927,0.6927767,1.0254467,1.0906088,0.8093826,0.6790583,1.0837497,1.0117283,1.0425946,1.2483698,1.2209331,1.4095604,1.2243627,1.0871792,1.1283343,1.1832076,1.1523414,1.3375391,1.2758065,1.0014396,1.0323058,1.0117283,0.8128122,0.8848336,1.2209331,1.3409687,1.3169615,1.1934965,1.0666018,1.0117283,1.0700313,1.2037852,1.3203912,1.2860953,1.0631721,0.6893471,0.61389613,0.51100856,0.48014224,0.52472687,0.5796003,0.5796003,0.4355576,0.33952916,0.432128,0.7888051,0.5727411,0.7407909,0.78194594,0.64476246,0.7476501,0.86082643,1.1454822,1.1763484,0.9294182,0.7956643,0.7956643,1.0082988,1.1523414,1.2929544,1.8416885,1.8108221,1.8862731,1.9514352,2.201795,3.1312134,3.1277838,3.4844608,3.57363,3.5873485,4.5030484,4.73969,3.9851806,4.0366244,4.9351764,4.955754,4.962613,6.159539,6.8900414,6.917478,7.459353,8.30646,7.9120584,8.2310095,9.325048,9.349055,11.032983,12.072148,11.657167,10.336777,10.014396,9.887501,10.336777,10.408798,10.014396,9.952662,10.182446,10.545981,10.254466,9.750318,10.693454,11.561139,11.780633,12.545431,13.886399,14.668345,15.440002,16.304258,16.242527,15.731518,16.750105,17.171944,17.586924,17.247395,16.345413,16.023033,17.20624,18.094503,18.54378,18.770132,19.329155,20.893047,22.405495,23.660725,24.120289,22.93708,23.996824,25.053137,25.320644,25.35837,27.049156,26.877676,28.84626,31.068632,32.91375,35.029808,39.83809,41.281944,45.023624,52.424675,60.556225,62.991234,62.915783,58.584213,51.426662,46.05593,39.457405,32.99263,28.733084,26.462696,23.671013,20.436913,18.36887,16.973028,16.012743,15.501736,16.482597,14.771234,12.751206,11.598865,11.273054,10.319629,10.175586,10.467101,11.070708,12.130451,12.154458,12.151029,12.521424,13.13189,13.334236,13.2862215,14.764374,15.415996,14.188204,11.317638,8.676856,8.025234,7.414768,6.1629686,4.870014,2.7093742,1.6530612,1.2620882,1.2449403,1.4267083,1.6907866,2.1469216,2.651071,3.018037,2.9974594,3.0386145,3.1106358,3.0146074,2.7128036,2.3149714,2.1160555,2.3252604,2.3046827,1.8828435,1.3409687,1.6359133,1.7902447,1.8245405,1.6256244,0.9568549,0.69963586,0.61046654,0.70306545,0.9534253,1.2826657,1.2277923,1.1214751,1.5776103,2.7333813,4.2526884,6.540223,6.711703,8.038953,11.111863,13.824667,12.199042,13.80066,14.712931,13.38568,10.655728,9.966381,8.776315,7.936065,7.699424,7.747438,6.615674,5.994919,7.4799304,10.082987,10.251037,7.9772205,6.1492505,4.8837323,4.4516044,5.284994,7.332458,6.217842,4.07435,2.0508933,0.30523327,0.52815646,1.1489118,1.2758065,1.0357354,1.5433143,0.84367853,0.31895164,0.05144381,0.0,0.0,0.0,0.037725464,0.0548734,0.041155048,0.01371835,0.0034295875,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08916927,0.25721905,0.37725464,0.22978236,0.6824879,0.66876954,0.5658819,0.64476246,1.0528834,0.9842916,0.89855194,0.8025235,0.6927767,0.5693115,1.255229,1.1592005,0.90541106,0.7613684,0.64819205,1.4472859,1.5844694,1.7833855,2.1846473,2.3389788,2.7128036,2.8877127,3.07634,3.4913201,4.307562,3.8617156,4.3795834,4.8905916,4.955754,4.65395,4.588788,6.0806584,6.958633,6.7871537,6.8591747,6.5367937,7.905199,8.762596,8.844906,9.846346,10.209882,11.382801,12.8197975,14.2362175,15.621771,16.647217,19.075365,19.905325,19.071936,19.44919,19.682402,21.69557,22.422644,21.78474,22.673002,21.963078,20.570665,19.260563,18.588364,18.910746,20.268862,21.270302,21.801888,21.743584,20.975357,21.332033,21.369759,20.028791,18.608942,20.755863,22.61813,23.36921,24.10314,24.891945,24.792488,24.76848,24.476965,24.730755,26.785078,32.32386,55.147766,74.41176,83.64078,81.32238,70.899864,69.80239,78.23918,77.18287,63.6017,50.486958,51.687313,46.23084,39.265347,35.122406,37.3242,28.314674,23.986534,22.94394,23.468666,23.499533,16.04018,10.655728,7.431916,6.094377,5.9983487,7.3393173,7.534804,7.414768,7.2364297,6.684266,5.9743414,6.6636887,7.0889573,6.636252,5.720552,5.23698,5.675967,6.0635104,6.262427,6.9552035,7.846896,7.8846216,8.488229,9.729739,10.329918,10.786053,11.05699,10.947243,10.600855,10.494537,10.203023,10.100135,9.764035,9.023245,7.9429245,7.3050213,6.8866115,7.394191,8.553391,9.105555,9.102125,8.772884,8.351046,8.073249,8.186425,8.745448,9.647429,10.80663,12.277924,14.243076,15.659496,16.61292,17.63494,18.334574,17.394867,17.1205,17.055338,16.650646,15.971589,15.690363,15.54632,15.566897,15.062748,13.828096,12.106443,11.595435,10.912948,10.007536,8.820899,7.2707253,6.756287,6.1904054,5.778855,5.8200097,6.7391396,8.06296,8.930646,9.873782,10.772334,10.875222,11.417097,10.792912,10.031544,10.014396,11.454823,11.742908,11.646879,11.602294,12.212761,14.2362175,12.487128,12.418536,13.059869,13.365103,12.205902,12.891819,13.570878,13.814379,13.495427,12.795791,11.595435,11.489118,12.71691,14.479718,14.953001,14.644339,13.570878,12.624311,12.140739,11.859513,11.050131,10.762046,10.912948,10.9198065,9.729739,8.937505,7.9772205,7.332458,7.1232533,7.099246,6.23499,5.6313825,6.3653145,8.543102,11.297061,13.426835,14.836395,15.097044,14.620332,14.668345,13.814379,12.788932,12.562579,12.881531,12.267634,12.445972,13.797231,15.275383,15.940722,14.973578,13.978998,12.8197975,11.794352,11.015835,10.39508,10.089847,10.364213,11.0981455,12.024134,12.7272,11.461681,10.477389,9.853205,9.47938,9.047252,10.268185,10.254466,9.877212,9.678296,9.89436,10.422516,10.443094,10.264755,9.839486,8.762596,8.340756,8.025234,8.200144,8.694004,8.779744,8.453933,8.536243,9.040393,10.076128,11.828648,11.283342,11.571428,11.622872,11.516555,12.493987,13.677195,12.343085,10.000677,8.405919,9.541112,0.548734,0.51100856,0.6310441,0.77165717,0.8711152,0.94656616,0.8128122,0.77851635,0.84367853,0.96371406,1.039165,1.1729189,1.0768905,0.980862,0.97057325,1.0082988,1.4472859,1.7319417,1.6564908,1.371835,1.371835,1.2037852,1.2895249,1.4404267,1.6084765,1.8759843,1.9514352,1.7593783,1.5638919,1.4541451,1.3581166,1.430138,1.4953002,1.7216529,2.1263442,2.5790498,2.7128036,2.7745364,2.6167753,2.452155,2.8534167,4.232111,5.3844523,7.1884155,10.789482,17.576635,21.239435,18.924463,13.985858,8.903209,5.2644167,3.690236,2.719663,2.1640697,1.7696671,1.2209331,1.1111864,1.1283343,1.1523414,1.1729189,1.2826657,1.1111864,0.9294182,0.8745448,0.89855194,0.77851635,0.97400284,0.8025235,0.8162418,1.1111864,1.3443983,1.039165,0.65162164,0.34638834,0.18176813,0.12346515,0.13375391,0.1097468,0.09602845,0.09602845,0.044584636,0.010288762,0.0274367,0.0274367,0.006859175,0.030866288,0.006859175,0.0274367,0.09945804,0.20920484,0.31895164,0.19891608,0.08573969,0.017147938,0.010288762,0.044584636,0.33952916,0.39440256,0.4424168,0.6310441,1.0220171,1.546744,1.862266,1.5501735,0.7579388,0.18176813,0.048014224,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.05144381,0.05144381,0.044584636,0.058302987,0.106317215,0.06859175,0.14404267,0.23664154,0.2709374,0.19891608,0.4424168,0.7133542,0.5727411,0.19891608,0.3806842,0.3806842,0.18176813,0.106317215,0.37725464,1.097468,0.72021335,0.71678376,0.6790583,0.4972902,0.34981793,0.6790583,0.70649505,0.72021335,0.8711152,1.1900668,1.0666018,1.0940384,1.214074,1.2689474,0.9774324,1.1351935,1.2655178,1.4610043,1.646202,1.587899,1.1832076,1.2037852,1.2929544,1.2517995,1.0082988,1.1043272,0.881404,0.85739684,1.0837497,1.1454822,1.0357354,0.8505377,0.8745448,1.0837497,1.1454822,1.1317638,1.1660597,1.0014396,0.7373613,0.823101,0.64133286,0.58645946,0.5624523,0.5418748,0.5796003,0.5796003,0.33266997,0.32581082,0.53158605,0.39783216,0.34638834,0.28122616,0.28808534,0.48014224,0.9911508,0.6756287,0.4938606,0.64133286,0.8711152,0.5041494,0.89512235,0.881404,0.96714365,1.196926,1.1592005,1.2346514,1.3786942,1.6907866,2.301253,3.3884325,2.935727,3.1346428,2.9563043,2.4795918,2.867135,3.5633414,3.426158,3.1963756,3.4295874,4.5167665,5.518206,6.5539417,7.0752387,7.5690994,9.582268,9.630281,9.561689,9.8429165,10.446524,10.847785,11.701753,11.533703,11.22161,10.978109,10.329918,10.573419,10.4533825,10.1481495,9.928656,10.1481495,10.182446,10.504827,10.515115,10.240748,10.316199,11.571428,11.9040985,12.319078,13.118172,13.886399,14.435134,15.285671,15.580616,15.199932,14.784951,15.9578705,16.489456,16.324837,15.803539,15.656067,15.570327,16.527182,17.466888,18.169954,19.257133,21.160555,22.46037,23.211449,23.204588,21.973368,22.583834,23.725885,24.096281,24.044838,25.557285,25.985985,28.345541,30.725674,33.297863,38.31535,42.427425,43.723812,48.43606,57.088913,64.50025,64.280754,62.92264,57.596493,48.81675,40.465702,34.618256,31.60022,30.715385,29.580193,24.123718,21.767591,20.227707,18.351723,16.516893,16.602633,17.357141,16.245956,14.38026,12.603734,11.506266,11.578287,11.989838,12.583157,13.155897,13.474849,15.549749,15.217079,14.445422,14.188204,14.359683,13.978998,13.491997,11.698323,8.879202,6.790583,5.7891436,5.4016004,5.096367,4.602506,3.9063,2.3321195,1.6907866,1.3855534,1.1489118,1.039165,1.0871792,1.2826657,1.5433143,1.786815,1.9239986,2.0337453,2.253239,2.435007,2.5481834,2.6716487,2.5481834,2.16064,1.728512,1.3409687,0.9602845,1.1214751,1.196926,1.2449403,1.2003556,0.8711152,0.8711152,0.84367853,0.84367853,0.84367853,0.7339317,0.65848076,0.9431366,1.5158776,2.0406046,1.9068506,5.7411294,8.940934,11.382801,12.775213,12.665466,13.275933,17.034761,18.097933,15.29596,12.144169,7.130112,6.324159,6.773435,6.9071894,6.5162163,4.856296,4.8425775,5.4976287,6.8214493,9.81205,9.678296,8.580828,7.500508,7.1884155,8.179566,6.310441,6.200694,4.8322887,2.0508933,0.548734,0.30523327,0.78537554,1.039165,1.0563129,1.7388009,0.6276145,0.14061308,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12003556,0.12003556,0.09602845,0.47328308,0.88826317,0.71678376,0.6001778,0.84367853,1.4198492,1.1249046,1.1180456,0.9945804,0.77508676,0.8848336,0.90884066,0.66876954,0.58988905,0.7922347,1.097468,1.6359133,1.9994495,2.311542,2.6785078,3.2032347,2.301253,2.1400626,2.8294096,3.7211025,3.4021509,3.8171308,4.0949273,3.9200184,3.7005248,4.5922174,5.3501563,6.5196457,7.051232,6.773435,6.4098988,6.15268,6.7185616,7.8263187,8.868914,8.940934,11.149589,12.397959,13.4474125,14.5243025,15.306249,17.20967,18.581505,18.69811,18.228258,19.239986,18.166525,19.829874,22.813616,25.468117,25.893385,24.747904,23.917942,22.638706,20.803877,18.996485,18.996485,19.188541,19.963629,20.999365,21.256582,21.19485,20.649546,19.123379,17.765263,19.363451,21.647556,24.230036,26.483274,27.930561,28.2598,28.040308,27.909983,29.655643,37.389362,57.555336,103.758736,145.38707,153.64552,124.43915,78.383224,60.086372,58.141796,59.09865,56.087475,48.81332,46.419468,39.13159,33.723133,30.818274,24.871368,25.77678,24.408375,23.893936,23.962528,20.934202,12.500846,7.3255987,5.1752477,4.852866,4.180667,6.0978065,6.9792104,6.893471,6.5230756,7.1712675,7.781734,7.8983397,7.6342616,7.332458,7.5519514,6.831738,6.7802944,7.140401,7.613684,7.857185,8.796892,9.609704,10.117283,10.30591,10.329918,10.707172,10.813489,10.7586155,10.580277,10.237319,9.908078,9.22216,8.742019,8.433355,7.675417,6.931196,6.2041235,5.888602,6.0669403,6.5299344,7.0923867,6.958633,6.725421,6.7459984,7.1095347,7.233,7.5553813,8.008087,8.553391,9.201583,9.688584,9.993818,10.203023,10.268185,10.010965,10.597425,11.338216,12.096155,12.96727,14.29795,15.151917,15.302819,15.234227,14.949572,13.96185,13.365103,11.684605,9.678296,7.7714453,6.0875177,6.0395036,6.1286726,6.0840883,6.1629686,7.140401,8.447074,9.770895,10.206452,9.825768,9.705732,9.777754,9.541112,9.205012,9.184435,10.100135,11.869802,12.542002,12.620882,13.296511,16.434584,16.63007,14.819247,12.79922,11.399949,10.497967,11.2421875,12.024134,12.456262,12.271064,11.30735,10.038403,10.542552,12.0138445,13.708061,14.953001,14.342535,13.035862,11.712041,10.576848,9.369633,9.661148,9.654288,10.031544,10.511685,9.825768,8.752307,7.267296,6.557371,6.5127864,5.7068334,5.535354,5.346727,5.919468,7.380472,9.184435,10.991828,13.375391,14.016724,13.145609,13.533153,13.3033695,12.9707,12.939834,13.416546,14.404267,15.830976,16.280252,16.191082,15.889278,15.608052,13.9481325,12.977559,12.0309925,10.81006,9.369633,10.0041065,11.427385,12.312219,12.689473,13.9481325,13.529722,12.466551,11.012405,9.633711,8.988949,9.866923,10.288762,10.80663,11.31078,11.015835,10.930096,9.866923,8.903209,8.419638,8.1041155,7.613684,7.5279446,7.888051,8.327039,8.073249,8.05953,8.495089,8.776315,9.301042,11.4754,12.452832,12.740917,12.97413,13.176475,12.785502,14.5585985,15.227368,14.123041,11.910957,10.604284,0.548734,0.5041494,0.53158605,0.61389613,0.6962063,0.6893471,0.84024894,0.91912943,1.0597426,1.2998136,1.5981878,1.2929544,1.3306799,1.4232788,1.5021594,1.7147937,1.8416885,1.7971039,1.6290541,1.4438564,1.4335675,1.3306799,1.3306799,1.430138,1.6256244,1.9137098,1.9102802,1.7182233,1.5981878,1.5638919,1.4198492,1.4918705,1.6359133,1.8348293,2.085189,2.4212887,2.253239,2.1194851,2.201795,2.5138876,2.9254382,4.0537724,5.768566,8.141841,11.842365,18.152807,19.713268,15.649208,10.093276,5.703404,3.6765177,2.4452958,1.8142518,1.704505,1.7765263,1.4404267,1.1832076,1.0768905,1.1351935,1.2655178,1.2586586,1.0460242,1.0631721,1.0288762,0.84024894,0.58302987,0.7476501,0.65848076,0.72021335,1.0254467,1.3546871,1.0597426,0.6824879,0.39440256,0.25721905,0.20920484,0.22978236,0.15776102,0.106317215,0.09602845,0.044584636,0.037725464,0.048014224,0.044584636,0.030866288,0.0548734,0.05144381,0.12003556,0.15776102,0.16462019,0.23664154,0.17147937,0.08916927,0.030866288,0.017147938,0.034295876,0.14061308,0.20234565,0.26750782,0.4046913,0.66876954,1.3581166,1.862266,1.6221949,0.7888051,0.19548649,0.05144381,0.006859175,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.030866288,0.044584636,0.044584636,0.037725464,0.05144381,0.082310095,0.116605975,0.15090185,0.29494452,0.28808534,0.18176813,0.13375391,0.4046913,0.20234565,0.2777966,0.3566771,0.41498008,0.6962063,0.5727411,0.61046654,0.5796003,0.4972902,0.64476246,0.7476501,0.5796003,0.5555932,0.764798,0.9945804,0.89169276,1.0837497,1.3066728,1.3821237,1.196926,1.5193073,1.6496316,1.5124481,1.2998136,1.4541451,1.3238207,1.3203912,1.2415106,1.08032,1.0323058,1.0323058,0.90884066,0.8779744,0.9534253,0.9362774,0.91569984,1.039165,1.1180456,1.0871792,1.0220171,0.85396725,0.91569984,0.84367853,0.6241849,0.59331864,0.47671264,0.42526886,0.36696586,0.33266997,0.45613512,0.50757897,0.39783216,0.3566771,0.38754338,0.26407823,0.32238123,0.3018037,0.28465575,0.37725464,0.72364295,0.58988905,0.6276145,0.66533995,0.61046654,0.42869842,1.0357354,1.1214751,1.1317638,1.2175035,1.2209331,1.4095604,1.8588364,1.9102802,1.6736387,2.0097382,2.2395205,2.4247184,2.5138876,2.6647894,3.2718265,3.6456516,3.974892,4.105216,4.091498,4.2115335,5.3878818,6.6876955,7.56567,8.337327,10.206452,10.604284,11.324498,11.790922,12.068718,12.850664,12.5145645,12.1921835,12.411677,12.922686,12.686044,11.952112,12.151029,12.085866,11.4376745,10.7586155,10.628291,10.899229,11.228469,11.681175,12.72034,13.128461,13.275933,13.615462,14.174485,14.592895,15.258235,15.621771,15.402277,15.004445,15.518884,15.947581,15.978448,15.748666,15.354263,14.826107,15.237658,15.858413,16.160215,16.331696,17.29198,18.159666,19.298288,20.28258,20.803877,20.652975,21.733295,22.148275,22.875349,24.408375,26.791937,27.35439,29.484163,32.23469,35.599117,40.5,42.83555,46.46748,53.841095,62.075535,62.974087,65.54627,67.38796,63.317043,53.67647,44.31027,39.440254,36.360485,32.735413,27.76594,22.172283,23.544119,22.834194,19.682402,15.594335,13.951562,13.87954,13.035862,12.449403,12.30193,11.945253,12.915827,13.077017,13.179905,13.557159,14.109323,15.433144,15.138199,15.066177,15.522313,15.275383,14.064738,13.245067,11.55771,9.0369625,7.010077,6.166398,5.171818,4.139512,3.2409601,2.7230926,2.750529,2.1263442,1.5844694,1.3306799,1.0734608,1.6496316,1.3752645,1.2723769,1.5364552,1.5433143,1.6942163,1.8656956,1.9548649,2.0474637,2.4144297,1.978872,1.6084765,1.2826657,1.0357354,0.94999576,1.1180456,1.1729189,1.2723769,1.2415106,0.58988905,0.6756287,0.70649505,0.70649505,0.69963586,0.6962063,0.7305021,0.7613684,0.94999576,1.3615463,1.978872,3.059192,6.636252,10.353925,11.955542,9.259886,11.255906,14.13333,14.2362175,11.941824,11.633161,8.423067,6.5539417,5.5593615,5.0655007,4.7808447,3.8548563,5.7754254,9.441654,11.962401,8.663138,8.375052,7.8023114,7.1369715,7.016936,8.532814,5.7651367,4.098357,2.7162333,1.5055889,1.0494537,0.39440256,0.33952916,0.39097297,0.77851635,2.4487255,0.59331864,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.34638834,0.50757897,0.5624523,1.0597426,0.72364295,0.58302987,0.7613684,0.9362774,0.3566771,0.71678376,0.805953,0.7339317,0.58302987,0.4081209,0.83338976,0.8025235,0.72364295,0.8162418,1.1111864,1.3169615,1.9102802,2.1400626,1.99602,2.2292318,1.821111,1.5433143,1.8931323,2.6236343,2.7573884,3.1620796,3.450165,3.508468,3.6593697,4.6779575,5.1992545,5.754848,6.1492505,6.5024977,7.250148,7.1129646,8.025234,9.325048,10.48082,11.091286,12.459691,13.498857,14.733508,15.786391,15.37827,16.890718,18.893597,19.294859,18.307138,18.423744,18.482046,18.941612,20.27572,22.052248,22.926792,22.971376,22.055677,20.70785,19.414894,18.595222,19.267422,18.852442,18.910746,19.360022,18.471758,18.900457,18.855871,19.013634,19.980776,22.292318,22.552967,23.616138,25.135447,26.476416,26.69591,27.042297,27.539587,30.286688,38.99784,58.99576,88.407906,101.59124,93.758064,72.1791,56.217796,52.575577,53.079723,50.932804,44.684093,38.219322,35.82547,29.624777,25.989414,26.232914,26.61703,29.151493,28.777668,25.920822,21.493225,16.894148,11.125582,6.5813785,4.1292233,3.5976372,3.765687,5.212973,7.39762,8.704293,8.694004,8.100685,8.251588,8.309891,8.210432,8.213862,8.920357,7.9737906,7.1198235,6.9346256,7.363324,7.723431,8.968371,9.554831,9.884071,10.113853,10.158438,9.9698105,9.832627,9.623423,9.362774,9.177576,8.553391,7.8983397,7.4696417,7.1712675,6.550512,6.0806584,5.5833683,5.144381,4.9420357,5.2506986,5.381023,5.2575574,5.1409516,5.1512403,5.254128,5.3570156,5.2438393,5.1580997,5.223262,5.429037,5.576509,5.809721,6.042933,6.2692857,6.5813785,7.507367,8.2481575,8.81404,9.424506,10.501397,11.434244,12.336226,13.083877,13.564018,13.670336,12.922686,11.787492,10.038403,7.891481,6.001778,5.3673043,5.0106273,5.1238036,5.7994323,7.0203657,7.8674736,9.016385,9.637141,9.407358,8.532814,8.615124,7.963502,7.500508,7.7131424,8.64942,10.408798,11.122152,11.094715,11.537132,14.565458,14.273943,13.162757,11.698323,10.388221,9.777754,10.230459,10.336777,10.271614,10.182446,10.182446,9.246168,10.179015,11.523414,12.627741,13.660047,13.323947,12.545431,11.609154,10.5597,9.235879,9.712592,9.712592,9.441654,8.971801,8.241299,8.543102,7.7097125,7.1987042,7.0752387,5.9743414,6.7631464,6.6122446,6.6225333,7.2535777,8.368194,9.705732,11.314209,12.63117,13.440554,13.838386,13.334236,13.255356,13.790371,14.863832,16.13621,17.175373,15.971589,14.946142,14.983868,15.4742985,14.119612,13.461131,12.4802685,11.22161,10.796341,10.912948,11.862943,12.370522,12.363663,12.946692,13.673765,12.63117,11.279913,10.576848,10.964391,10.88551,10.923236,11.046701,11.125582,10.9198065,10.511685,9.791472,9.040393,8.56025,8.652849,8.98209,8.759167,8.4264965,8.237869,8.255017,8.378482,8.073249,8.251588,9.3079,11.122152,12.977559,13.440554,13.059869,12.22305,11.187314,12.109874,13.080446,13.05301,11.993267,10.861504,0.59674823,0.53158605,0.5796003,0.66876954,0.75450927,0.8162418,1.0871792,1.1523414,1.2723769,1.5090185,1.704505,1.7422304,1.920569,2.0714707,2.1160555,2.0577524,1.8416885,1.7662375,1.6496316,1.4850113,1.4507155,1.4815818,1.6324836,1.7456601,1.8108221,1.9514352,1.8519772,1.6393428,1.529596,1.5261664,1.4335675,1.5227368,1.6084765,1.7662375,1.9239986,1.8862731,2.037175,2.1263442,2.3081124,2.760818,3.7039545,4.6436615,7.8434668,10.583707,12.092726,13.543441,13.673765,11.406808,8.008087,4.8014226,3.1723683,2.095478,1.4781522,1.3443983,1.4541451,1.313532,1.0323058,0.9568549,1.1660597,1.471293,1.3992717,1.1043272,1.1660597,1.1454822,0.90884066,0.64476246,0.6790583,0.6824879,0.823101,1.1454822,1.5501735,1.2346514,0.78194594,0.4355576,0.28465575,0.26407823,0.30523327,0.29494452,0.24350071,0.16462019,0.072021335,0.072021335,0.082310095,0.07545093,0.07888051,0.16119061,0.33609957,0.34295875,0.23664154,0.12003556,0.12346515,0.08916927,0.041155048,0.01371835,0.006859175,0.01371835,0.037725464,0.072021335,0.12003556,0.25378948,0.6173257,1.2689474,1.7319417,1.4575747,0.6207553,0.12346515,0.030866288,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.010288762,0.030866288,0.044584636,0.048014224,0.048014224,0.041155048,0.0274367,0.030866288,0.0548734,0.09945804,0.14061308,0.12346515,0.09602845,0.12346515,0.28465575,0.16804978,0.2777966,0.32581082,0.30866286,0.4938606,0.45613512,0.45613512,0.4972902,0.5418748,0.4972902,0.64819205,0.5796003,0.6001778,0.77165717,0.90198153,0.9774324,1.2380811,1.2929544,1.1523414,1.214074,1.4061309,1.3066728,1.1420527,1.0837497,1.2620882,1.0117283,1.08032,1.0460242,0.8779744,0.9362774,0.8471081,0.7888051,0.8471081,0.939707,0.7922347,0.7407909,0.83681935,0.85739684,0.78537554,0.8265306,0.7579388,0.69963586,0.6207553,0.5041494,0.37039545,0.37382504,0.31895164,0.26407823,0.274367,0.4355576,0.33609957,0.32924038,0.30866286,0.23664154,0.1371835,0.23664154,0.2503599,0.274367,0.36353627,0.53844523,0.58302987,0.6379033,0.64476246,0.6001778,0.5693115,0.96371406,0.939707,0.9328478,1.0357354,1.0254467,1.4953002,1.611906,1.5398848,1.4781522,1.646202,2.1126258,2.2463799,2.417859,2.7951138,3.3369887,3.8274195,4.3281393,4.698535,4.8254294,4.629943,6.2692857,7.623973,8.484799,9.184435,10.590566,10.878652,11.519984,11.893809,12.127021,13.094165,12.761495,13.118172,13.522863,13.687484,13.670336,13.416546,13.272504,13.347955,13.323947,12.456262,12.21962,11.962401,12.006986,12.6586075,14.2190695,15.247946,15.45715,15.402277,15.385129,15.419425,15.721229,15.608052,15.117621,14.867262,16.05733,15.539461,15.151917,14.939283,14.949572,15.21365,15.54632,15.697222,15.570327,15.673215,17.130789,17.61436,18.344864,19.123379,19.826445,20.388897,21.218857,21.976797,23.60242,26.016851,28.126047,29.624777,32.34787,35.51338,38.936108,43.051613,45.79871,51.759335,60.539078,68.327675,67.87496,73.07079,72.89245,65.34736,53.67647,46.333725,42.64692,38.558853,33.555084,28.150053,23.869928,25.546997,24.487255,20.649546,15.837835,13.673765,12.912396,11.684605,11.012405,10.923236,10.4533825,12.05843,12.956982,12.668896,12.127021,13.690913,14.743796,14.843254,15.217079,15.762384,15.035312,13.186764,11.818358,10.082987,7.9875093,6.4064693,5.5113473,4.355576,3.2375305,2.4418662,2.253239,2.1023371,1.5433143,1.1797781,1.155771,1.155771,1.1043272,1.0117283,1.1351935,1.4095604,1.4575747,1.5947582,1.6599203,1.6290541,1.5741806,1.6633499,1.430138,1.1832076,0.91227025,0.7305021,0.8711152,1.0082988,1.0220171,1.0323058,1.0082988,0.764798,0.5761707,0.52472687,0.52472687,0.5144381,0.4664239,0.5727411,0.58645946,0.7099246,1.097468,1.8416885,2.651071,5.5113473,8.988949,11.002116,8.838047,10.960961,11.677745,11.550851,11.393089,12.264205,9.650859,6.8763227,4.8940215,4.1155047,4.420738,5.295283,5.7994323,7.082098,8.505377,7.6274023,8.117833,8.419638,7.7748747,6.5779486,6.385892,4.355576,2.510458,1.3238207,0.82996017,0.6241849,0.29494452,0.4081209,1.0700313,1.8039631,1.5536032,0.33609957,0.01371835,0.0,0.0,0.0,0.0,0.0,0.07545093,0.15433143,0.0,0.044584636,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.23321195,0.32581082,0.4115505,0.9568549,0.66876954,0.66191036,0.64133286,0.4629943,0.1371835,0.48700142,0.53501564,0.5555932,0.6036074,0.490431,0.8848336,0.7613684,0.64819205,0.75450927,1.0048691,1.3615463,1.9857311,2.2669573,2.2429502,2.5790498,2.2086544,2.061182,2.4247184,3.083199,3.2889743,2.836269,3.3266997,4.15323,4.931747,5.504488,6.0703697,6.728851,7.490219,8.351046,9.263316,9.383351,10.871792,12.120162,12.524854,12.4802685,13.485138,13.985858,14.908417,16.13621,16.513464,18.001905,19.421753,19.771572,19.167965,18.821575,19.12681,19.970488,20.749004,21.239435,21.592682,21.887627,20.508932,19.198832,18.3723,17.103354,18.478617,18.95533,19.60695,20.159115,19.003344,18.440891,18.643238,20.145397,22.456938,24.058556,23.492674,23.02968,23.623,25.303495,27.17605,26.565584,25.93454,27.398973,32.601658,42.694935,57.064907,62.18528,60.295578,55.52159,53.86167,54.13261,51.262043,45.843296,39.282494,33.781437,29.587051,25.865948,26.016851,30.293547,35.787746,35.91121,31.76141,25.063425,17.583494,11.14273,12.404818,7.6788464,4.9488945,6.0223556,6.5196457,6.3481665,7.0718093,7.5759587,8.337327,11.417097,8.824328,7.822889,7.7577267,8.110974,8.501947,7.3839016,6.6122446,6.5642304,7.130112,7.7268605,8.783174,9.256456,9.510246,9.692014,9.740028,9.39707,9.338767,9.129561,8.663138,8.179566,7.682276,6.8866115,6.3790326,6.142391,5.593657,5.329579,5.06893,4.7259717,4.4241676,4.48933,4.396731,4.2183924,4.1155047,4.1155047,4.122364,4.0880685,3.875434,3.7553983,3.8034124,3.899441,3.998899,4.266407,4.5613513,4.8940215,5.446185,6.166398,7.0135064,7.6857057,8.186425,8.820899,9.465661,10.052121,10.741467,11.345076,11.345076,11.163307,10.662587,9.290752,7.2638664,5.579939,4.7534084,4.420738,4.664239,5.4736214,6.742569,7.8194594,9.012956,9.80519,9.877212,9.108984,8.200144,7.4113383,7.191845,7.6788464,8.707723,9.599416,9.853205,9.647429,9.880642,12.195613,13.039291,12.80265,11.945253,10.789482,9.506817,9.424506,9.499957,9.301042,8.838047,8.573969,8.196714,9.719451,11.14273,11.756626,12.147599,12.243628,11.808069,11.417097,10.864933,9.126132,8.848335,8.505377,8.368194,8.31332,7.8331776,8.532814,8.049242,7.3564653,6.8900414,6.5470824,6.715132,6.495639,6.2830043,6.451054,7.349606,8.512236,9.606275,10.714031,11.739478,12.404818,13.114742,13.824667,14.747226,15.861842,16.928444,16.513464,15.038741,14.277372,14.579176,14.88441,14.123041,13.893259,13.262215,12.30193,12.116733,12.133881,12.689473,13.138749,13.173045,12.840376,13.71492,13.214201,12.30193,11.698323,11.897239,12.085866,11.921246,11.2421875,10.401938,10.264755,9.89093,9.582268,9.146709,8.920357,9.767465,10.100135,9.609704,8.964942,8.611694,8.748878,8.577398,8.536243,8.838047,9.571979,10.731179,12.569438,13.461131,13.025573,11.664027,10.539123,10.172156,10.621432,11.434244,11.986408,11.454823,0.6927767,0.6962063,0.7133542,0.764798,0.8848336,1.1043272,1.3958421,1.4438564,1.5433143,1.7388009,1.8485477,2.0337453,2.1057668,2.1469216,2.1434922,2.0097382,1.8313997,1.8519772,1.786815,1.6084765,1.5055889,1.5947582,1.845118,1.9308578,1.821111,1.7559488,1.6907866,1.5536032,1.471293,1.4507155,1.371835,1.4610043,1.4507155,1.5810398,1.7696671,1.6221949,2.194936,2.4315774,2.603057,3.1380725,4.6402316,5.7925735,9.938945,12.627741,12.363663,10.6145735,9.633711,8.800322,7.1129646,4.7979927,3.2992632,2.3218307,1.5227368,1.1351935,1.1180456,1.1523414,1.0151579,0.99801,1.2175035,1.5261664,1.4953002,1.313532,1.3889829,1.5227368,1.5158776,1.1763484,0.8676856,0.89512235,0.9877212,1.1146159,1.488441,1.2312219,0.84024894,0.53501564,0.39440256,0.3566771,0.4355576,0.4355576,0.35324752,0.22292319,0.1097468,0.14404267,0.15433143,0.13032432,0.1097468,0.1920569,0.4355576,0.42183927,0.274367,0.116605975,0.0548734,0.030866288,0.010288762,0.0,0.0,0.0,0.0,0.010288762,0.058302987,0.24007112,0.72021335,1.1180456,1.3443983,1.0425946,0.37725464,0.058302987,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.010288762,0.024007112,0.034295876,0.037725464,0.0548734,0.041155048,0.0274367,0.024007112,0.037725464,0.058302987,0.044584636,0.0548734,0.06516216,0.07545093,0.12346515,0.14061308,0.26407823,0.28808534,0.24007112,0.40126175,0.40126175,0.37039545,0.4115505,0.4938606,0.44927597,0.6001778,0.5590228,0.61389613,0.805953,0.94999576,1.0597426,1.2106444,1.2620882,1.196926,1.1420527,1.1934965,1.0151579,0.9328478,1.0048691,1.0082988,0.72021335,0.84367853,0.84367853,0.6790583,0.764798,0.6859175,0.7305021,0.805953,0.7956643,0.59331864,0.65848076,0.59674823,0.5041494,0.4698535,0.5658819,0.5796003,0.53158605,0.48014224,0.42869842,0.33952916,0.34981793,0.31209245,0.29494452,0.31895164,0.34638834,0.32238123,0.34981793,0.30866286,0.1920569,0.11317638,0.16462019,0.1920569,0.26064864,0.37725464,0.47671264,0.4629943,0.5007198,0.5144381,0.53158605,0.66533995,0.7682276,0.71678376,0.7373613,0.83338976,0.78194594,1.3443983,1.2449403,1.2277923,1.5055889,1.7662375,2.1229146,2.1332035,2.2566686,2.702515,3.415869,3.865145,4.1360826,4.4413157,4.7774153,4.9351764,6.475061,7.7131424,8.844906,9.901219,10.741467,11.231899,11.430815,11.746337,12.199042,12.397959,12.144169,12.816368,13.38568,13.522863,13.615462,14.249936,14.126471,14.356253,14.757515,13.862392,13.639469,13.282792,13.38568,14.153908,15.419425,16.462019,16.63007,16.37285,15.981877,15.597764,15.498305,15.206791,14.7026415,14.476289,15.553179,15.4914465,14.997586,14.874121,15.371411,16.194511,16.571766,16.444872,16.386568,16.729528,17.576635,18.152807,18.70154,19.408035,20.3546,21.510372,22.02481,23.211449,25.238335,27.697348,29.631636,32.59137,35.42078,38.25705,41.31624,44.931026,48.415485,55.346684,63.145565,69.3394,71.55492,77.100555,74.473495,64.58599,52.239475,46.114235,43.960453,40.7435,35.691715,29.991743,26.805656,27.85511,25.93111,21.819035,17.223389,14.79867,13.265644,11.279913,10.028113,9.654288,9.239308,10.189304,11.238758,11.286773,11.043272,13.035862,13.790371,14.87755,14.671775,13.166186,11.958971,10.463672,9.15014,7.630832,5.9914894,4.7945633,3.998899,3.0626216,2.452155,2.287535,2.3389788,1.5913286,1.0666018,0.91569984,1.0734608,1.2860953,0.6756287,0.75450927,1.0768905,1.4095604,1.7456601,1.5364552,1.3992717,1.2620882,1.1043272,0.97400284,0.89512235,0.75450927,0.58302987,0.48700142,0.6276145,0.7613684,0.7407909,0.71678376,0.7373613,0.7613684,0.5212973,0.45956472,0.45956472,0.4424168,0.36353627,0.5624523,0.6859175,0.8711152,1.2106444,1.7593783,2.8054025,5.6176643,9.458802,12.099585,9.849775,10.055551,10.940384,12.490558,13.749216,12.8197975,10.261326,8.488229,7.5416627,6.783724,4.897451,7.174697,6.5230756,6.1286726,7.0135064,8.045813,8.639131,9.568549,8.738589,6.169828,3.9886103,2.6133456,1.3306799,0.5761707,0.3806842,0.36353627,0.89169276,1.9239986,3.806842,4.698535,0.5761707,0.116605975,0.0,0.0,0.0,0.0,0.0,0.0,0.07545093,0.15433143,0.0,0.044584636,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08916927,0.24007112,0.39097297,0.607037,1.08032,0.6001778,0.6344737,0.53501564,0.24350071,0.28465575,0.37382504,0.33952916,0.4081209,0.5761707,0.59674823,0.7990939,0.7133542,0.6859175,0.83681935,1.0768905,1.5398848,2.061182,2.4658735,2.6956558,2.784825,2.7093742,2.942586,3.234101,3.525616,3.9440255,3.426158,3.9303071,4.863155,5.7136927,6.042933,6.433906,7.6033955,8.803751,9.729739,10.511685,10.264755,11.80121,13.46799,14.061309,12.8197975,14.191633,14.284232,14.819247,16.115631,17.093063,19.071936,20.563807,21.002794,20.495214,19.829874,19.630959,20.69413,21.644127,21.993944,22.134558,21.798458,20.776442,19.901896,19.03764,17.082775,17.586924,18.20425,19.164536,19.836735,18.728977,17.861292,18.639809,20.79016,23.132568,23.554407,23.280039,21.884197,21.897917,24.02083,27.114319,26.35295,25.368658,25.968836,28.228935,30.482174,34.74858,38.034126,43.03789,48.827038,50.840206,50.60699,46.203403,41.32653,37.16301,32.392452,28.84626,25.817934,27.062874,33.441906,42.948723,44.190235,36.267887,24.960537,14.7026415,8.567109,14.246507,8.872343,5.4084597,7.514226,9.534253,7.140401,6.601956,6.478491,7.2124224,11.118723,8.344186,7.1095347,7.0443726,7.4181976,7.130112,6.866034,6.728851,7.010077,7.6033955,7.98408,8.433355,8.851766,9.201583,9.427936,9.458802,9.095266,8.97866,8.635701,7.9875093,7.349606,6.807731,5.90575,5.453044,5.4599032,5.130663,4.8768735,4.791134,4.588788,4.273266,4.1429415,3.8960114,3.6970954,3.5564823,3.4776018,3.4638834,3.4638834,3.2683969,3.175798,3.275256,3.4364467,3.5153272,3.666229,3.9200184,4.3349986,4.996909,5.5902276,6.4407654,7.2192817,7.805741,8.282454,8.752307,9.006097,9.379922,9.692014,9.249598,9.102125,8.9100685,7.9909387,6.4407654,5.096367,4.383013,4.2698364,4.5819287,5.288424,6.5024977,8.23444,9.314759,10.14129,10.583707,9.97667,8.570539,7.6033955,7.4044795,7.949784,8.865483,9.153569,8.81404,8.450503,8.669997,10.076128,12.103014,12.809509,12.377381,11.249047,10.1481495,9.750318,9.592556,9.084977,8.213862,7.5450926,7.3358874,8.944365,10.364213,10.789482,10.6145735,10.9369545,10.947243,11.029553,10.803201,9.146709,8.299602,7.5245147,7.3290286,7.5107965,7.1369715,8.001227,7.864044,7.140401,6.427047,6.5024977,6.3207297,6.1904054,5.8337283,5.693115,6.9380555,7.8331776,8.855195,9.537683,10.048691,11.173596,13.443983,14.973578,16.105343,16.88729,17.086205,15.676644,14.54831,14.2533655,14.507155,14.195063,13.7526455,14.143619,14.205351,13.728639,13.419975,13.615462,14.315098,14.730078,14.445422,13.409687,13.653188,13.512574,13.145609,12.809509,12.833516,13.347955,13.121602,12.041282,10.72089,10.508256,9.829198,9.458802,9.283894,9.5033865,10.621432,11.05356,10.419086,9.6988735,9.386781,9.523964,9.342196,9.616563,9.777754,10.000677,11.180455,12.466551,13.293081,13.039291,11.856084,10.700313,9.914937,9.568549,10.39165,11.89038,12.322508,0.7579388,0.86082643,0.83338976,0.8848336,1.0940384,1.3855534,1.5570327,1.605047,1.6873571,1.8313997,1.9480057,2.0165975,1.9137098,1.786815,1.7388009,1.7936742,1.8931323,1.9994495,1.9445761,1.7490896,1.605047,1.6839274,1.845118,1.8382589,1.6427724,1.4575747,1.5433143,1.5673214,1.5227368,1.4267083,1.3306799,1.4095604,1.3306799,1.430138,1.6907866,1.7353712,2.4898806,2.6990852,2.9322972,3.74168,5.6793966,7.582818,11.602294,13.7697935,12.8197975,10.182446,8.501947,7.6514096,6.40304,4.6779575,3.5564823,2.8396983,1.879414,1.196926,0.97400284,1.0597426,1.0666018,1.1180456,1.2277923,1.3478279,1.3889829,1.3924125,1.5090185,1.8931323,2.2669573,1.9171394,1.2243627,1.1043272,1.0151579,0.89512235,1.1489118,1.0460242,0.84367853,0.6790583,0.5796003,0.5007198,0.5727411,0.47671264,0.33609957,0.22292319,0.14404267,0.20920484,0.21263443,0.17490897,0.14061308,0.17147937,0.3841138,0.42869842,0.33266997,0.16462019,0.048014224,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.058302987,0.274367,0.764798,0.85396725,0.8128122,0.5418748,0.16804978,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0034295875,0.017147938,0.037725464,0.030866288,0.030866288,0.030866288,0.0274367,0.0274367,0.01371835,0.0034295875,0.006859175,0.01371835,0.01371835,0.072021335,0.2503599,0.32581082,0.29837412,0.41498008,0.4424168,0.4115505,0.36696586,0.39097297,0.59674823,0.61046654,0.4972902,0.5555932,0.8093826,1.0117283,1.0082988,1.0048691,1.1866373,1.371835,0.9842916,0.97400284,0.96371406,0.9602845,0.91227025,0.70649505,0.66533995,0.77851635,0.7133542,0.5212973,0.61389613,0.6344737,0.70306545,0.67219913,0.52472687,0.3841138,0.6173257,0.45613512,0.29494452,0.28808534,0.34295875,0.36696586,0.42869842,0.4424168,0.4115505,0.4424168,0.38754338,0.36696586,0.38754338,0.37725464,0.216064,0.38754338,0.4081209,0.32924038,0.22978236,0.20577525,0.14061308,0.17147937,0.2469303,0.34295875,0.4698535,0.28122616,0.33266997,0.36696586,0.38754338,0.64476246,0.58988905,0.6276145,0.7133542,0.7613684,0.64476246,1.08032,1.0288762,1.0940384,1.4438564,1.8073926,1.937717,1.920569,2.0508933,2.5241764,3.457024,3.683377,3.6319332,3.8171308,4.3933015,5.1512403,6.118384,7.1026754,8.484799,9.928656,10.357354,11.523414,11.677745,12.22305,12.878101,11.701753,11.276484,11.677745,12.415107,13.107883,13.46799,14.589465,14.812388,15.0456,15.313108,14.743796,14.71636,14.850114,15.405707,16.221949,16.702091,16.691803,16.640358,16.520323,16.228807,15.594335,15.234227,14.808959,14.311668,14.05102,14.637479,15.889278,15.450292,15.337115,16.194511,17.288551,18.11165,18.139088,18.574646,19.342873,19.102802,19.685833,20.141968,20.999365,22.323185,23.753323,24.082563,25.413242,27.278938,29.388136,31.596788,35.537384,37.56427,39.471123,42.273094,46.210262,49.982807,57.26039,63.375347,67.40168,72.15509,74.74443,70.978745,62.054955,51.54327,45.38716,45.215683,44.155937,39.3991,32.478195,29.271528,29.93344,27.289227,23.135998,18.95533,15.885849,14.020154,11.441104,9.6817255,9.078118,8.769455,8.707723,9.081548,9.81205,10.899229,12.415107,12.343085,13.63604,12.243628,8.501947,7.1095347,6.591667,5.861165,4.8185706,3.6182148,2.6545007,2.1400626,1.6393428,1.7662375,2.3492675,2.4212887,1.6496316,1.1077567,0.9568549,1.1077567,1.2106444,0.64819205,0.66533995,0.89855194,1.2380811,1.8142518,1.2483698,1.0220171,0.9294182,0.8265306,0.65162164,0.50757897,0.39783216,0.34638834,0.34638834,0.32581082,0.44927597,0.4081209,0.4355576,0.52472687,0.45613512,0.48014224,0.5007198,0.4972902,0.4629943,0.41840968,0.66191036,0.8676856,1.08032,1.3512574,1.7216529,2.6545007,6.142391,11.22161,14.63062,10.816919,8.546532,10.875222,14.037301,14.997586,11.458252,9.156999,9.602845,11.218181,11.187314,5.4633327,9.019815,8.237869,8.100685,9.448513,8.971801,9.184435,10.422516,9.239308,5.5250654,2.510458,1.1934965,0.6241849,0.65162164,0.8711152,0.6379033,1.9068506,4.4721823,7.006647,6.8763227,0.14747226,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.05144381,0.23664154,0.5624523,0.84024894,1.0254467,1.214074,0.5007198,0.5761707,0.6379033,0.4629943,0.4081209,0.33952916,0.26064864,0.29494452,0.4355576,0.5212973,0.5590228,0.66876954,0.823101,1.0117283,1.2723769,1.6873571,2.0508933,2.5241764,2.8911421,2.551613,2.9871707,3.532475,3.707384,3.6319332,4.029765,4.461893,4.822,5.2472687,5.7651367,6.2727156,6.392751,7.764586,8.968371,9.692014,10.72089,10.38479,11.2593355,13.251926,14.788382,12.823228,15.049029,15.227368,15.415996,16.283682,17.096493,19.36688,21.599543,22.179142,21.232576,20.635828,19.949911,20.550089,21.582394,22.467228,22.913074,22.062536,22.096832,21.819035,20.683842,18.79414,17.466888,17.1205,17.62122,18.163095,17.267973,16.979887,18.399736,20.426622,21.908205,21.633839,21.86705,20.440342,20.526081,22.889067,25.886526,26.02371,26.10602,26.953129,28.287237,28.719366,28.623337,29.220085,33.188118,38.781776,39.848377,39.611736,37.701454,36.535397,35.564823,31.291555,29.978024,27.248072,27.539587,33.08866,43.926155,49.38263,40.79151,27.073164,15.069608,9.551401,14.644339,9.3079,5.662249,7.4456344,10.014396,7.140401,6.6876955,6.5162163,6.210983,7.099246,6.941485,6.667118,6.728851,6.8557453,6.0669403,7.0923867,7.56567,7.9943686,8.378482,8.220721,7.963502,8.327039,8.81404,9.136421,9.22902,9.194724,8.875772,8.303031,7.5725293,6.8626046,6.0052075,5.209543,5.0106273,5.2781353,5.212973,4.8082814,4.695105,4.523626,4.2286816,4.040054,3.6593697,3.450165,3.275256,3.1380725,3.1860867,3.316411,3.1483612,3.0420442,3.1415021,3.3815732,3.3884325,3.2855449,3.4227283,3.9097297,4.605936,5.2438393,5.895461,6.5985265,7.3050213,7.891481,8.299602,8.591117,8.824328,8.834618,8.220721,7.6959944,7.449064,6.831738,5.7719955,4.7945633,4.4927597,4.633373,4.9694724,5.552502,6.7391396,8.604835,9.026674,9.633711,10.504827,10.161868,9.328478,8.412778,8.025234,8.258447,8.683716,8.954653,8.117833,7.5210853,7.699424,8.371623,10.611144,11.979549,11.8869505,10.957532,11.036412,10.834066,10.065839,9.105555,8.182996,7.3873315,6.9380555,8.014946,9.270175,9.908078,9.692014,9.887501,10.316199,10.600855,10.357354,9.194724,8.30646,7.2707253,6.5950966,6.3893213,6.3824625,7.1198235,7.1232533,6.550512,5.8474464,5.73427,5.8200097,6.029215,5.7377,5.5490727,7.2878733,7.610255,8.498518,8.97523,9.287323,10.926665,14.027013,15.604623,16.6335,17.233677,16.657507,15.285671,14.778092,14.832966,14.918706,14.263655,13.653188,14.55174,15.354263,15.391989,14.928994,15.302819,16.187653,16.506605,15.848124,14.490007,13.814379,13.797231,13.834956,13.858963,14.318527,14.586036,14.291091,13.317088,12.096155,11.598865,10.412228,9.72631,9.671436,10.233889,11.231899,12.0138445,11.667457,11.105004,10.772334,10.655728,10.782623,10.950673,10.741467,10.714031,12.3911,12.932974,13.179905,12.994707,12.298501,11.039842,10.923236,10.14129,10.326488,11.712041,13.111313,0.61046654,0.64819205,0.78537554,1.1454822,1.5570327,1.5570327,1.3375391,1.2826657,1.2929544,1.313532,1.313532,1.862266,2.1194851,2.0577524,1.8554068,1.8931323,1.8073926,1.8862731,1.8382589,1.6667795,1.6770682,1.8245405,1.7250825,1.6256244,1.605047,1.5570327,1.728512,1.862266,1.762808,1.5261664,1.5261664,1.6359133,1.5364552,1.5398848,1.7010754,1.786815,2.3218307,2.603057,3.3061223,4.8254294,7.2775846,10.401938,13.584596,14.901558,12.987847,7.0203657,5.5559316,4.98662,4.479041,3.8102717,3.3712845,3.40901,2.5927682,1.6907866,1.1077567,0.90198153,0.6927767,0.88826317,1.0666018,1.0597426,0.9602845,0.7305021,0.9294182,1.4095604,1.9274281,2.136633,1.4644338,0.89512235,0.6756287,0.78537554,0.9294182,0.9911508,0.90541106,0.77851635,0.6824879,0.67219913,0.548734,0.30866286,0.17490897,0.18176813,0.16804978,0.15433143,0.116605975,0.14747226,0.24350071,0.30523327,0.6962063,0.78537554,0.58302987,0.24350071,0.061732575,0.037725464,0.01371835,0.0,0.0,0.0,0.0,0.0,0.006859175,0.106317215,0.47328308,0.5212973,0.4698535,0.29837412,0.08916927,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.030866288,0.0,0.0,0.0,0.01371835,0.024007112,0.024007112,0.01371835,0.01371835,0.0034295875,0.0,0.030866288,0.061732575,0.0,0.0,0.17490897,0.34638834,0.4629943,0.61046654,0.59674823,0.5590228,0.48357183,0.45270553,0.61046654,0.47671264,0.48700142,0.61046654,0.7579388,0.7922347,0.8162418,0.9534253,0.94656616,0.77508676,0.64133286,0.50757897,0.7476501,0.77851635,0.52472687,0.42869842,0.805953,0.84367853,0.65162164,0.45613512,0.6241849,0.72364295,0.41840968,0.26407823,0.37382504,0.39783216,0.3841138,0.34638834,0.2777966,0.24350071,0.36696586,0.5007198,0.4424168,0.40126175,0.41840968,0.3806842,0.4424168,0.40126175,0.34638834,0.31552204,0.29151493,0.12003556,0.17833854,0.20920484,0.1920569,0.34981793,0.18176813,0.2194936,0.22635277,0.18862732,0.33609957,0.32238123,0.40126175,0.432128,0.4355576,0.59674823,0.6207553,0.66191036,0.7956643,0.91227025,0.71678376,1.0940384,0.89855194,0.7339317,0.85396725,1.1592005,1.3169615,1.7422304,2.2429502,2.6887965,3.0043187,3.3472774,3.625074,4.338428,5.4084597,6.1629686,7.0923867,7.7371492,8.090397,8.330468,8.820899,10.700313,12.202472,13.430264,13.80066,12.055,11.701753,11.979549,12.617453,13.529722,14.784951,15.419425,15.2033615,14.860402,14.987297,16.03675,16.438013,17.051908,17.61436,17.995045,18.20425,17.274832,16.979887,17.158226,17.412016,17.1205,16.53404,15.223939,14.291091,14.332246,15.443433,16.13621,15.367981,14.928994,15.80011,18.142517,19.678972,20.45063,21.369759,22.669573,23.86307,23.400076,23.129137,23.959099,25.53328,26.229485,26.277498,27.68363,29.76882,32.11123,34.51537,37.224743,38.020405,39.474552,42.838978,48.06567,51.982258,61.78745,70.05276,73.61952,73.60924,69.99445,65.09014,58.903164,52.506985,48.04852,50.356632,48.71729,42.681217,34.728004,30.272968,30.650223,28.047167,23.962528,19.438902,15.0456,14.496866,12.325937,10.39165,9.170717,7.7680154,9.23245,9.184435,9.541112,10.693454,11.537132,9.654288,7.3564653,5.778855,5.0586414,4.3041325,3.865145,3.2683969,2.5310357,1.7525192,1.1283343,0.7990939,0.6790583,1.0768905,1.6770682,1.5398848,1.9308578,1.3512574,0.91912943,0.84367853,0.4424168,0.3566771,0.28122616,0.26407823,0.31552204,0.4115505,0.40126175,0.64476246,0.980862,1.1420527,0.7613684,0.53158605,0.3806842,0.33266997,0.33952916,0.29151493,0.216064,0.18176813,0.22978236,0.31209245,0.274367,0.432128,0.44584638,0.42869842,0.41840968,0.3806842,0.42869842,0.45956472,0.5521636,0.82996017,1.4644338,2.1743584,5.4084597,11.029553,15.189643,10.329918,8.779744,8.117833,7.6925645,7.0032177,5.7239814,4.7088237,5.453044,8.573969,10.834066,5.1580997,11.907528,9.887501,8.323608,9.1810055,7.140401,8.495089,10.216741,8.375052,3.7931237,2.061182,0.88826317,0.65162164,1.9754424,3.3472774,1.1146159,1.8965619,6.3001523,6.7665763,2.5996273,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05144381,0.26064864,0.490431,1.1180456,1.1180456,0.44584638,0.030866288,0.45613512,0.9568549,1.0494537,0.6790583,0.21263443,0.36010668,0.33266997,0.29494452,0.32581082,0.4115505,0.40126175,0.50757897,0.70306545,0.9431366,1.1763484,1.6873571,1.9445761,2.2600982,2.6373527,2.7470996,3.1140654,3.2683969,3.82399,4.32128,3.234101,4.431027,4.914599,5.504488,6.4098988,7.2021337,7.689135,7.822889,8.011517,8.889491,11.30735,13.673765,13.615462,14.006435,15.031882,14.191633,17.021042,18.070496,17.768692,17.20624,18.097933,18.903887,20.697561,20.814167,19.562366,20.234566,20.464348,20.649546,20.412905,20.018501,20.385468,21.1194,21.465788,21.174273,20.491785,20.186552,18.917604,18.04992,17.940172,18.255693,17.974468,17.37772,18.416885,19.737276,20.646116,21.133118,20.340883,19.792149,20.666695,22.823904,24.826784,25.056566,26.387245,27.285797,27.549875,28.304386,28.01287,25.035988,23.389786,24.404943,26.750782,30.557625,31.847149,32.282707,31.696247,28.105469,24.61415,27.697348,31.0069,33.57566,39.82437,44.097637,39.41625,30.687948,20.673553,9.9801,11.664027,9.026674,8.258447,9.1810055,5.2644167,7.7920227,8.110974,6.910619,5.363875,5.1580997,6.036074,6.8043017,7.349606,7.4936485,7.0203657,7.6033955,7.8434668,7.9600725,7.9909387,7.781734,7.2707253,7.5245147,7.8537555,8.069819,8.484799,9.825768,9.640571,9.06097,8.364764,6.9723516,5.9126086,5.6176643,5.6965446,5.7994323,5.6142344,5.113515,4.523626,4.1429415,4.029765,3.9680326,3.4776018,3.117495,2.976882,3.07634,3.357566,3.2718265,3.1689389,3.223812,3.4295874,3.6010668,3.5873485,3.391862,3.5221863,4.057202,4.65395,5.055212,5.3227196,5.6828265,6.169828,6.6225333,6.608815,7.0375133,7.548522,7.8434668,7.658269,7.8194594,7.5382333,6.615674,5.4153185,4.866585,5.3673043,5.7582774,6.142391,6.7871537,8.117833,7.98408,6.7974424,6.8283086,8.258447,9.184435,9.599416,9.870353,9.716022,9.194724,8.683716,9.06097,7.9292064,6.708273,6.210983,6.636252,7.689135,8.838047,9.441654,9.644,10.374502,10.97468,9.73317,8.766026,8.498518,7.6445503,7.0958166,7.4627824,8.512236,9.753747,10.436234,10.240748,10.477389,10.580277,10.158438,8.988949,8.107545,7.267296,6.1732574,5.6245236,7.4936485,6.941485,6.183546,5.470192,5.0003386,4.928317,4.770556,5.453044,6.001778,6.4579134,7.874333,7.2878733,6.8283086,7.4936485,9.301042,11.290202,13.478279,13.227919,13.591455,15.031882,15.412566,14.750656,15.193072,15.861842,16.300829,16.448301,15.302819,15.947581,16.938732,17.38115,16.96617,17.12736,16.808409,17.051908,17.418875,15.9921665,14.867262,15.3302555,15.323397,14.942713,16.417435,15.758954,15.127911,14.195063,13.004995,11.979549,11.074138,10.792912,10.696883,10.978109,12.466551,13.248496,13.9481325,13.965281,13.255356,12.329367,12.415107,12.096155,11.814929,12.048141,13.306799,13.293081,13.097594,12.548861,11.626302,10.467101,11.201033,11.05356,10.912948,11.461681,13.183334,0.70649505,0.6859175,0.764798,0.89169276,0.99801,1.0082988,1.2072148,1.2346514,1.4232788,1.7525192,1.8485477,2.153781,2.2120838,2.0680413,1.8348293,1.6976458,1.8073926,2.177788,2.2635276,2.0131679,1.8485477,1.9754424,1.99602,2.0406046,2.0577524,1.8142518,1.8382589,1.8554068,1.8005334,1.6599203,1.4644338,1.4369972,1.471293,1.5741806,1.704505,1.7593783,2.4041407,2.6545007,3.4433057,5.171818,7.6925645,10.515115,14.63062,15.532601,11.777204,4.9694724,3.542764,3.415869,3.7108135,3.82399,3.433017,3.1586502,2.6887965,2.07833,1.4610043,1.0597426,0.89855194,0.9602845,0.90541106,0.70306545,0.64476246,0.6173257,0.764798,1.0700313,1.3684053,1.3306799,0.83338976,0.59331864,0.5212973,0.53844523,0.5761707,0.65848076,0.64133286,0.5693115,0.4698535,0.39097297,0.37725464,0.32238123,0.29151493,0.2777966,0.216064,0.1371835,0.09259886,0.12003556,0.24350071,0.5007198,1.1043272,1.4472859,1.1660597,0.4698535,0.12346515,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.072021335,0.34981793,0.3806842,0.41840968,0.30523327,0.08573969,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.044584636,0.024007112,0.0274367,0.017147938,0.01371835,0.01371835,0.01371835,0.0034295875,0.01371835,0.01371835,0.006859175,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.0,0.0,0.034295876,0.1097468,0.22292319,0.37725464,0.42526886,0.3841138,0.42869842,0.5418748,0.52472687,0.48700142,0.47328308,0.45270553,0.4389872,0.47671264,0.607037,0.6379033,0.5761707,0.4664239,0.37382504,0.41498008,0.4355576,0.4424168,0.4389872,0.4389872,0.6893471,0.59674823,0.6893471,0.922559,0.6756287,0.6344737,0.42183927,0.39097297,0.53158605,0.45613512,0.37725464,0.31895164,0.32581082,0.37382504,0.37725464,0.4355576,0.3806842,0.3841138,0.48357183,0.5658819,0.4115505,0.33952916,0.30866286,0.33266997,0.48357183,0.28465575,0.20234565,0.19891608,0.21263443,0.16804978,0.16462019,0.24350071,0.2469303,0.17490897,0.21263443,0.28122616,0.37725464,0.45613512,0.4972902,0.51100856,0.4938606,0.5212973,0.6344737,0.78194594,0.7888051,0.8848336,0.9328478,1.0117283,1.1180456,1.1592005,1.4850113,1.8828435,2.0714707,2.1880767,2.7985435,2.9460156,3.333559,3.923448,4.7774153,6.090947,6.7940125,7.082098,7.699424,8.803751,9.966381,11.7086115,12.243628,12.840376,13.684054,13.862392,12.627741,12.751206,13.241637,13.88297,15.237658,16.37971,16.904436,16.763824,16.516893,17.343424,16.88729,17.034761,17.446312,17.655516,17.079346,16.777542,16.609491,17.021042,17.61779,17.168514,16.259674,14.688923,13.906977,14.068168,14.037301,14.421415,14.949572,15.638919,16.479168,17.436022,19.521212,20.498644,21.572105,22.985096,24.02426,23.852781,24.267761,24.998262,25.896814,26.973705,27.951138,29.614489,31.84372,34.103817,35.441357,37.224743,37.71517,39.8278,44.262257,49.506096,55.970867,67.43941,77.076546,81.36353,80.10145,74.370605,68.47514,64.321915,63.025528,64.904945,67.82009,61.8629,50.55555,38.857227,33.191547,31.50762,28.746801,24.76505,19.936192,15.141628,14.291091,12.668896,10.933525,9.554831,8.803751,9.527394,8.841476,8.501947,8.951223,9.314759,6.495639,4.664239,3.642222,3.1620796,2.8637056,2.5310357,2.1229146,1.7010754,1.3066728,0.9568549,0.6790583,0.5796003,0.5212973,0.5658819,0.96714365,1.4472859,0.881404,0.36353627,0.25378948,0.17490897,0.12689474,0.12003556,0.18862732,0.2777966,0.22978236,0.36353627,0.5418748,0.7956643,0.980862,0.7888051,0.59331864,0.58645946,0.58302987,0.53844523,0.5590228,0.5453044,0.4115505,0.32238123,0.31895164,0.31209245,0.45956472,0.4046913,0.36010668,0.37039545,0.28465575,0.53844523,0.58988905,0.86082643,1.5398848,2.5756202,4.7191124,6.392751,8.203573,9.47938,8.292743,8.7145815,7.9737906,6.042933,3.899441,3.5359046,3.4604537,8.23444,10.521975,8.114404,3.9131594,13.526293,15.522313,11.46854,5.4736214,4.187526,6.012067,7.3290286,5.7582774,2.1846473,0.75450927,3.8205605,3.974892,3.6970954,3.2512488,0.6859175,6.368744,6.8763227,4.249259,0.9774324,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.20577525,0.1920569,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22292319,0.20920484,0.2709374,0.4046913,0.2709374,0.31895164,0.66191036,0.64819205,0.39097297,0.77508676,0.6344737,0.5555932,0.490431,0.37725464,0.12689474,0.1371835,0.12689474,0.15090185,0.2469303,0.45956472,0.4081209,0.50757897,0.7305021,1.0117283,1.2243627,1.7182233,2.0714707,2.1400626,2.0303159,2.0989075,3.0214665,3.192946,4.012617,4.996909,3.782835,3.9165888,5.192395,6.0875177,6.368744,7.0923867,7.0032177,7.8777623,9.366203,11.122152,12.795791,13.22106,12.572867,13.145609,14.939283,15.680074,16.383139,16.640358,17.089634,17.809847,18.341434,19.157675,20.303158,20.505503,19.658396,18.804428,19.504065,19.726988,19.325726,18.54378,18.04306,19.281141,19.53836,19.263992,18.866161,18.69811,17.847572,17.768692,17.754974,17.676094,17.96418,17.490896,17.597214,17.933313,18.554068,19.912186,19.596663,20.35803,22.100262,23.815056,23.581844,23.996824,25.20061,25.876238,26.370098,28.657633,28.561604,27.203487,27.618467,29.981453,31.593359,33.448765,34.378185,32.536495,29.113768,28.338682,28.997162,28.084892,30.320982,33.49335,28.486153,32.16267,36.216442,37.35164,32.00834,16.362562,10.422516,7.517656,6.677407,6.5059276,5.2164025,5.857735,5.7891436,5.926327,6.2212715,5.6348124,5.535354,5.7239814,6.0326443,6.23499,6.042933,6.169828,6.550512,6.927767,7.085528,6.8283086,6.776865,7.082098,7.366754,7.4627824,7.4113383,7.9017696,7.7611566,7.4456344,6.8591747,5.3501563,4.7945633,4.928317,5.1512403,5.1992545,5.1512403,4.856296,4.712253,4.3521466,3.7931237,3.4192986,3.1552205,3.069481,3.0626216,3.0386145,2.9288676,2.9220085,2.976882,3.1723683,3.426158,3.4913201,3.4776018,3.4295874,3.6319332,4.125794,4.7019644,4.7945633,4.9008803,5.161529,5.435896,5.2918534,5.3878818,6.046363,6.958633,7.7097125,7.7714453,7.6274023,7.1232533,6.3481665,5.6073756,5.429037,5.892031,6.584808,7.058091,7.301592,7.764586,7.7268605,7.157549,7.085528,7.932636,9.513676,10.408798,9.956093,9.139851,8.4093485,7.682276,7.8366075,7.438775,6.5642304,5.6210938,5.3570156,6.3378778,7.5279446,8.141841,8.207003,8.556821,9.156999,9.105555,8.862054,8.519095,7.840037,7.349606,7.0272245,7.301592,8.2310095,9.510246,9.764035,10.161868,10.323058,9.956093,8.851766,7.936065,7.2295704,6.3618846,5.7377,6.540223,6.0497923,5.6999745,5.346727,4.976331,4.7088237,4.149801,4.7259717,5.4907694,6.012067,6.3721733,5.7754254,6.385892,7.675417,9.22216,10.707172,11.571428,11.204462,11.372512,12.284782,12.603734,13.145609,14.544881,15.748666,16.023033,14.946142,15.333686,16.921585,18.001905,18.104792,17.991615,17.682953,17.051908,17.027903,17.288551,16.273392,16.095055,17.079346,17.257685,16.39,15.954441,15.110763,14.520873,13.629181,12.466551,11.63659,11.533703,12.507706,12.854094,12.511135,13.063298,14.099034,15.0078745,15.354263,15.162207,14.915276,13.54687,12.778643,12.569438,12.908967,13.807519,13.725209,13.433694,12.775213,11.914387,11.31078,12.157887,12.408247,12.178465,11.955542,12.572867,0.6036074,0.65505123,0.70306545,0.71678376,0.7133542,0.77851635,0.90198153,0.9842916,1.2586586,1.6667795,1.8828435,1.9720128,1.9137098,1.7936742,1.6942163,1.704505,1.6770682,1.8999915,1.9651536,1.8245405,1.762808,1.8279701,1.8554068,1.9239986,1.9857311,1.8691251,1.9720128,1.8313997,1.6564908,1.5570327,1.5330256,1.4472859,1.6427724,1.8931323,2.0268862,1.9274281,2.7162333,2.7951138,3.474172,5.1100855,7.0923867,10.528833,16.084764,18.176813,14.321958,5.1512403,3.069481,2.8225505,3.2581081,3.6079261,3.4844608,2.976882,2.393852,1.879414,1.5055889,1.2346514,1.0082988,0.84024894,0.6756287,0.5521636,0.58302987,0.5178677,0.59331864,0.7682276,0.90884066,0.7888051,0.45613512,0.41840968,0.47328308,0.5041494,0.48014224,0.4972902,0.47328308,0.39440256,0.3018037,0.28465575,0.35324752,0.3806842,0.36696586,0.33266997,0.31209245,0.1920569,0.18862732,0.28808534,0.4698535,0.6859175,1.2792361,1.5673214,1.214074,0.45613512,0.1097468,0.034295876,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.17490897,0.2777966,0.4424168,0.37725464,0.116605975,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.030866288,0.01371835,0.006859175,0.006859175,0.006859175,0.006859175,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0,0.006859175,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.020577524,0.06516216,0.1371835,0.2503599,0.31552204,0.41840968,0.5555932,0.65162164,0.5555932,0.5144381,0.45270553,0.39097297,0.432128,0.4081209,0.39783216,0.3566771,0.31209245,0.38754338,0.34981793,0.31552204,0.28122616,0.2709374,0.36010668,0.5007198,0.5041494,0.61046654,0.7442205,0.5212973,0.78537554,0.764798,0.64476246,0.59674823,0.7922347,0.548734,0.5521636,0.65162164,0.67219913,0.39097297,0.44927597,0.37382504,0.35324752,0.4355576,0.5007198,0.47671264,0.39440256,0.34638834,0.36353627,0.39783216,0.28465575,0.22635277,0.18862732,0.16804978,0.18519773,0.1920569,0.26750782,0.26064864,0.20234565,0.3018037,0.32238123,0.38754338,0.4424168,0.4629943,0.45270553,0.58988905,0.53844523,0.6173257,0.8162418,0.8265306,0.7922347,1.0288762,1.1146159,1.0563129,1.2895249,1.4198492,1.611906,1.6599203,1.7010754,2.2155135,1.9754424,2.8225505,3.6627994,4.2389703,5.120374,6.200694,6.944915,7.8126,9.0644,10.7757635,11.979549,12.339656,13.275933,14.815818,15.611482,13.71492,14.071597,14.610043,14.956431,16.438013,17.525192,18.235117,18.324286,17.840714,17.137648,17.141079,17.350283,17.95389,18.564358,18.183672,17.669235,17.226818,17.319416,17.514904,16.486027,15.151917,13.817808,13.210771,13.327377,13.419975,14.116182,14.977009,15.7795315,16.414005,16.901007,18.938183,19.771572,20.797018,22.299177,23.44123,23.753323,24.346642,25.26577,26.60331,28.469006,29.144634,30.08777,32.100937,34.817173,36.68287,38.672028,39.947834,42.544033,46.745277,51.100853,58.76255,71.77784,82.99944,88.517654,87.667114,83.338974,77.30976,74.05165,75.51266,81.12346,82.364975,71.10221,56.018883,43.188793,36.0724,33.18469,30.537046,26.767931,21.69214,16.283682,14.023583,12.555719,11.087856,9.678296,9.239308,9.23245,8.169277,7.332458,7.006647,6.4887795,4.5339146,3.292404,2.5927682,2.2155135,1.879414,1.6256244,1.4507155,1.3238207,1.2106444,1.0631721,0.66876954,0.5041494,0.3841138,0.4081209,0.9602845,1.0151579,0.65505123,0.26064864,0.041155048,0.041155048,0.041155048,0.06516216,0.29494452,0.59674823,0.548734,0.4938606,0.47328308,0.52472687,0.58988905,0.5007198,0.5212973,0.45270553,0.36696586,0.32924038,0.39783216,0.50757897,0.51100856,0.4972902,0.5624523,0.805953,1.0185875,0.90198153,0.7613684,0.6859175,0.5418748,0.607037,0.6824879,0.864256,1.371835,2.5413244,5.4976287,7.281014,7.795452,7.2364297,6.0875177,7.6033955,6.8728933,4.5853586,2.1434922,1.6633499,8.831187,11.2421875,9.156999,4.9591837,3.1620796,9.139851,12.761495,11.087856,5.802862,3.199805,3.199805,3.3026927,2.4418662,0.89169276,0.26407823,4.0503426,4.3692946,4.5510626,5.171818,4.040054,8.539673,7.3564653,4.173808,1.371835,0.037725464,0.10288762,0.16462019,0.12346515,0.058302987,0.20920484,0.52472687,0.6241849,0.5007198,0.24007112,0.0,0.0,0.0,0.35324752,0.70649505,0.017147938,0.2777966,0.37725464,0.42183927,0.5007198,0.66876954,0.66876954,0.4424168,0.3018037,0.4389872,0.9534253,0.4355576,0.22978236,0.20577525,0.20920484,0.041155048,0.20920484,0.15090185,0.15776102,0.29151493,0.3806842,0.42183927,0.5761707,0.6859175,0.75450927,0.9259886,1.2380811,2.4624438,2.4727325,1.5536032,2.4041407,3.3952916,3.3781435,3.6525106,4.0674906,3.0351849,3.4192986,4.9831905,5.8234396,5.90575,7.0375133,6.9517736,8.327039,10.48082,12.5145645,13.313659,12.902108,12.212761,12.250486,13.275933,14.808959,15.909856,16.101913,16.400288,16.901007,16.79126,17.665806,18.564358,18.564358,17.892159,17.926455,19.05136,19.569225,19.270851,18.327715,17.29884,18.190533,17.943602,17.322845,16.770683,16.403717,16.04018,16.815268,17.247395,16.938732,16.606062,16.78783,17.12393,17.470318,18.019053,19.277712,19.95334,21.328604,23.163433,24.542128,23.86307,23.149715,23.959099,24.998262,26.058006,28.0163,28.77081,27.206917,27.60475,29.960876,29.967735,31.291555,30.814844,27.368109,22.319756,19.579515,23.11542,22.137987,24.202599,28.136335,24.048267,22.978235,29.68994,38.438816,40.5583,24.470106,14.195063,9.47595,6.8797526,5.223262,5.56965,5.90232,4.938606,5.06893,6.1492505,5.5319247,5.1821065,5.130663,5.0655007,4.962613,5.0655007,4.8082814,5.0106273,5.360445,5.761707,6.334448,6.478491,6.5882373,6.691125,6.7322803,6.5813785,6.842027,6.6568294,6.327589,5.892031,5.099797,4.9660425,5.103226,5.147811,5.0449233,5.055212,4.6916757,4.4859004,4.1635194,3.7108135,3.391862,3.2032347,3.0969174,3.0043187,2.942586,3.0043187,3.0626216,3.117495,3.2203827,3.3369887,3.3438478,3.5153272,3.789694,4.064061,4.2869844,4.4584637,4.3007026,4.372724,4.647091,4.9660425,5.0243454,5.761707,6.3961806,7.0375133,7.5725293,7.6514096,7.205563,7.0546613,6.948344,6.8557453,6.989499,7.0443726,7.394191,7.706283,7.73029,7.3084507,7.582818,7.6342616,7.7851634,8.580828,10.789482,11.646879,10.467101,9.129561,8.299602,7.421627,6.9620624,6.279575,5.521636,4.9831905,5.1100855,5.48734,6.327589,7.239859,7.840037,7.7714453,7.082098,6.7528577,6.9552035,7.390761,7.284444,7.116394,7.0546613,7.274155,7.939495,9.22216,9.602845,10.096705,10.268185,9.815479,8.553391,7.64798,6.9346256,6.1972647,5.5559316,5.442755,5.295283,5.188966,4.976331,4.6745276,4.479041,3.7759757,3.8274195,4.4721823,5.2781353,5.521636,5.0243454,5.6793966,7.010077,8.515666,9.6817255,9.866923,10.007536,10.4705305,11.204462,11.736049,13.193623,14.640909,15.611482,15.920145,15.662926,16.386568,17.820137,18.557497,18.45461,18.6158,18.20425,17.700102,17.665806,17.7927,16.901007,16.770683,17.271402,17.36057,16.70895,15.683503,15.127911,14.568888,13.893259,13.128461,12.411677,12.566009,13.924125,15.028452,15.227368,14.688923,15.244516,15.772673,16.314548,16.715809,16.643787,14.997586,13.9309845,13.509145,13.845244,15.076467,14.699212,14.846684,14.582606,13.732068,12.857523,12.922686,13.018714,12.891819,12.607163,12.538571,0.50757897,0.607037,0.6036074,0.6001778,0.65162164,0.78537554,0.86082643,0.97400284,1.1934965,1.5055889,1.7902447,1.8862731,1.920569,1.845118,1.7388009,1.7936742,1.5810398,1.6084765,1.670209,1.6564908,1.5741806,1.6187652,1.6667795,1.8039631,1.9445761,1.8691251,2.037175,1.8656956,1.6016173,1.4438564,1.5570327,1.5501735,1.8279701,2.0749004,2.1297739,1.9651536,2.935727,2.867135,3.457024,5.164959,7.226141,10.443094,17.305698,20.659836,17.04162,6.6876955,3.5187566,2.867135,3.292404,3.7142432,3.4124396,2.627064,1.9239986,1.471293,1.2758065,1.1934965,0.9568549,0.6824879,0.4938606,0.4424168,0.52815646,0.48357183,0.5212973,0.6001778,0.65162164,0.58988905,0.32924038,0.4081209,0.5418748,0.59674823,0.607037,0.51100856,0.41840968,0.32924038,0.26750782,0.30866286,0.37039545,0.3841138,0.37039545,0.36353627,0.41498008,0.26750782,0.2469303,0.36010668,0.5693115,0.7956643,1.2689474,1.371835,0.9842916,0.35324752,0.072021335,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.058302987,0.2503599,0.4355576,0.4046913,0.18862732,0.044584636,0.020577524,0.006859175,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.01371835,0.006859175,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.010288762,0.017147938,0.010288762,0.006859175,0.006859175,0.0034295875,0.006859175,0.01371835,0.0,0.01371835,0.010288762,0.006859175,0.01371835,0.020577524,0.1097468,0.21263443,0.30523327,0.39440256,0.5144381,0.45613512,0.4046913,0.36696586,0.3566771,0.39783216,0.31895164,0.29151493,0.26407823,0.26407823,0.38754338,0.35324752,0.32581082,0.31552204,0.32238123,0.32238123,0.5521636,0.50757897,0.5418748,0.65505123,0.51100856,0.823101,0.90884066,0.805953,0.7133542,1.0082988,0.7682276,0.7682276,0.7990939,0.7407909,0.53844523,0.51100856,0.39783216,0.37725464,0.44927597,0.42183927,0.42526886,0.37725464,0.37039545,0.4046913,0.36010668,0.32924038,0.2469303,0.16804978,0.13375391,0.19891608,0.18519773,0.22978236,0.2709374,0.29494452,0.32581082,0.29151493,0.33952916,0.37725464,0.37382504,0.36010668,0.5418748,0.5212973,0.5727411,0.7133542,0.69963586,0.7682276,0.94999576,1.0837497,1.1694894,1.371835,1.2792361,1.4027013,1.3958421,1.3443983,1.7525192,1.5947582,2.5756202,3.2581081,3.4638834,4.266407,5.5319247,6.684266,7.8537555,9.156999,10.72089,11.0981455,11.928105,13.375391,15.0078745,15.803539,14.640909,15.306249,16.019604,16.352274,17.240536,17.905876,18.752985,19.239986,19.054789,18.101362,18.62609,19.349733,20.11453,20.491785,19.775002,18.588364,17.86815,17.532051,17.069057,15.539461,14.102464,13.029003,12.562579,12.740917,13.38568,14.088745,14.754086,15.532601,16.383139,17.065628,18.639809,19.582945,20.683842,22.086544,23.27661,23.852781,24.233465,25.293207,27.467566,30.746252,31.058344,31.277838,33.16754,36.470234,38.89152,40.81895,43.07905,46.419468,50.596703,54.396687,61.969215,75.40977,87.36531,93.74435,93.679184,91.22017,85.605934,82.687355,84.37471,88.62054,85.56478,72.583786,58.67681,48.28516,41.30252,36.49767,33.363026,29.233803,23.5304,17.761833,14.778092,13.872682,12.898679,11.348505,10.347065,9.273604,7.6274023,6.3173003,5.439326,4.297273,3.1552205,2.3767042,1.879414,1.5330256,1.1729189,1.0254467,1.1180456,1.4164196,1.6667795,1.3855534,0.8128122,0.50757897,0.4355576,0.58645946,0.9602845,0.5624523,0.36696586,0.18176813,0.0,0.0,0.037725464,0.05144381,0.28122616,0.59674823,0.4938606,0.39440256,0.31552204,0.2777966,0.26750782,0.23321195,0.31895164,0.22978236,0.14061308,0.12346515,0.16462019,0.30523327,0.39097297,0.44927597,0.5590228,0.8471081,1.0700313,1.430138,1.471293,1.2037852,1.1111864,0.9774324,0.9911508,1.1077567,1.6770682,3.415869,5.4839106,6.4990683,6.358455,5.2438393,3.6216443,4.722542,4.297273,2.7882545,1.1900668,1.0357354,9.318189,8.748878,5.830299,3.8685746,2.9665933,4.715683,7.3255987,7.9292064,5.871454,2.719663,1.4198492,0.77851635,0.42526886,0.19891608,0.15776102,2.3286898,3.059192,4.537344,6.992929,8.690575,11.30049,8.076678,3.974892,1.4267083,0.32924038,0.17147937,0.17147937,0.12689474,0.10288762,0.44927597,0.97400284,0.9945804,0.72707254,0.34981793,0.0,0.08916927,0.044584636,0.47671264,0.9842916,0.15776102,0.34981793,0.34981793,0.28808534,0.30866286,0.59674823,0.8093826,0.490431,0.33266997,0.5212973,0.7579388,0.20234565,0.20577525,0.31209245,0.274367,0.048014224,0.30866286,0.29151493,0.28122616,0.34981793,0.36353627,0.4629943,0.5761707,0.6001778,0.6276145,0.9362774,1.2929544,2.6956558,2.750529,1.6736387,2.301253,3.1106358,3.2581081,3.5393343,3.8479972,3.192946,3.5290456,4.57164,5.1992545,5.6176643,7.3598948,7.936065,9.122703,10.967821,12.912396,13.821238,12.812939,12.185325,12.202472,12.902108,14.085316,14.96329,15.097044,15.46401,15.96816,15.453721,16.506605,17.782412,17.820137,17.117071,18.132229,19.171394,19.569225,19.1954,18.255693,17.28169,17.466888,16.822126,16.156786,15.827546,15.762384,15.340545,16.173935,17.099922,17.370861,16.695232,16.80498,17.597214,18.279701,18.677534,19.222837,20.656404,22.158566,23.540688,24.473536,24.480396,24.048267,24.326063,25.070284,26.037428,27.001143,28.729654,26.802225,25.838512,26.689049,26.414682,28.475864,25.93454,20.570665,15.391989,14.63062,19.329155,21.28059,22.751883,24.09971,23.753323,20.423193,24.332924,33.880894,41.446564,33.42133,19.994495,13.347955,8.838047,5.284994,4.976331,5.9434752,4.57164,4.331569,5.377593,4.57507,4.547633,4.5442033,4.1772375,3.7348208,4.1635194,3.8857226,3.9680326,4.2423997,4.7842746,5.909179,6.279575,6.358455,6.451054,6.5059276,6.118384,6.3035817,6.118384,5.8234396,5.593657,5.5250654,5.425607,5.284994,4.9660425,4.5922174,4.530485,4.15666,3.882293,3.6079261,3.340418,3.199805,3.0797696,2.959734,2.8739944,2.877424,3.0420442,3.0351849,3.0523329,3.1346428,3.2203827,3.1449318,3.3678548,3.799983,4.1017866,4.1463714,3.9886103,3.806842,3.9097297,4.2355404,4.6848164,5.1100855,6.4064693,7.0718093,7.5245147,7.936065,8.2310095,7.5245147,7.514226,7.623973,7.56224,7.301592,7.346176,7.5759587,7.8194594,7.764586,6.9654922,7.414768,7.8091707,8.320179,9.304471,11.283342,11.979549,10.820349,9.290752,8.1041155,7.1781263,6.7219915,5.892031,5.3501563,5.3330083,5.6656785,5.744559,6.7219915,7.8503256,8.539673,8.327039,7.3255987,6.56766,6.5710897,6.9826403,6.5813785,6.6053853,6.8145905,7.1712675,7.8263187,9.14328,9.630281,10.106995,10.360784,10.124143,9.067829,8.30646,7.579388,6.7802944,5.9228973,5.147811,4.9934793,4.955754,4.729401,4.297273,3.9200184,3.1895163,2.9803114,3.5153272,4.465323,4.9523244,4.681387,5.0655007,6.3310184,7.966932,8.738589,9.287323,9.884071,10.628291,11.375941,11.742908,13.917266,15.217079,15.951012,16.499744,17.322845,17.576635,18.646667,19.29143,19.428614,20.111101,19.61038,19.013634,18.584934,18.265984,17.676094,17.391438,17.480608,17.593784,17.388008,16.55119,16.523752,15.728088,14.747226,13.992717,13.687484,13.989287,15.062748,16.489456,17.29884,15.96816,15.597764,15.944152,17.051908,18.077356,17.267973,15.470869,14.280802,14.2190695,15.141628,16.242527,16.462019,16.938732,16.770683,15.806969,14.675205,13.824667,13.227919,12.902108,12.682614,12.22305,0.490431,0.5796003,0.53158605,0.5453044,0.67219913,0.8025235,0.9945804,1.1043272,1.2346514,1.4507155,1.7833855,1.9925903,2.1915064,2.1400626,1.8965619,1.8108221,1.5398848,1.529596,1.611906,1.6187652,1.3855534,1.4404267,1.4781522,1.6599203,1.8691251,1.7353712,1.9308578,1.9137098,1.7113642,1.4987297,1.5913286,1.6804979,1.8931323,1.99602,1.9445761,1.8999915,2.9185789,2.8225505,3.5221863,5.4599032,7.6033955,10.14129,17.95732,21.963078,18.324286,8.467651,4.3487167,3.357566,3.7622573,4.1017866,3.2066643,2.1194851,1.4850113,1.1489118,1.0048691,0.9877212,0.8093826,0.58645946,0.41840968,0.35324752,0.39440256,0.44927597,0.48014224,0.4972902,0.5178677,0.5658819,0.38754338,0.5212973,0.64476246,0.65848076,0.70649505,0.5453044,0.4115505,0.32924038,0.30866286,0.33952916,0.33266997,0.32581082,0.33609957,0.3806842,0.48357183,0.30523327,0.216064,0.274367,0.48700142,0.8162418,1.1489118,1.0666018,0.6962063,0.25378948,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.030866288,0.2194936,0.34295875,0.36353627,0.274367,0.09602845,0.037725464,0.010288762,0.0,0.0,0.0,0.017147938,0.006859175,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0,0.020577524,0.030866288,0.024007112,0.020577524,0.017147938,0.006859175,0.0,0.0,0.0,0.030866288,0.030866288,0.030866288,0.034295876,0.024007112,0.024007112,0.072021335,0.11317638,0.12689474,0.14061308,0.216064,0.18862732,0.19891608,0.26064864,0.2709374,0.31209245,0.29494452,0.28122616,0.31552204,0.4046913,0.47328308,0.39440256,0.41840968,0.5212973,0.3841138,0.7476501,0.5212973,0.48700142,0.7305021,0.6310441,0.64476246,0.6859175,0.71678376,0.764798,0.939707,0.8711152,0.84024894,0.72707254,0.59674823,0.72021335,0.5590228,0.42869842,0.432128,0.50757897,0.4115505,0.3018037,0.28122616,0.33609957,0.41498008,0.4046913,0.37725464,0.23664154,0.14404267,0.14061308,0.15776102,0.16462019,0.16119061,0.2709374,0.41498008,0.31209245,0.23664154,0.2777966,0.30866286,0.29837412,0.29151493,0.32581082,0.4424168,0.5178677,0.5144381,0.4938606,0.77851635,0.7579388,0.9568549,1.3443983,1.313532,1.1111864,1.3272504,1.371835,1.2586586,1.587899,1.9274281,2.5138876,2.7333813,2.8739944,4.1326528,4.8425775,5.9914894,7.4181976,8.745448,9.369633,9.692014,11.101575,12.644889,13.776653,14.369971,15.049029,16.060759,17.072487,17.78927,17.923023,18.38259,19.46291,20.364891,20.810738,21.064526,21.290878,22.065966,22.580404,22.271742,20.838173,19.023922,17.854433,16.88729,15.810398,14.455711,13.406258,12.672326,12.3533745,12.535142,13.3033695,13.738928,14.040731,14.901558,16.348843,17.734396,18.646667,19.802439,21.016512,22.20315,23.396646,24.048267,24.288338,25.540138,28.530739,33.25671,33.880894,33.798584,35.4928,38.946396,41.672916,43.199085,45.98391,50.04797,54.69506,58.53277,65.65602,78.767334,89.824326,95.07503,95.03387,94.341095,89.89977,87.64996,88.55195,88.56224,81.31209,71.60293,63.128418,56.409855,48.768734,40.839527,36.09984,30.904013,24.494114,19.027351,16.71238,16.842705,16.21852,14.123041,12.319078,9.537683,7.1781263,5.48734,4.3041325,3.0351849,2.1023371,1.5844694,1.2380811,0.939707,0.6927767,0.6756287,0.96371406,1.7079345,2.3732746,1.704505,1.0082988,0.5727411,0.4972902,0.65162164,0.6893471,0.16119061,0.037725464,0.024007112,0.0034295875,0.0034295875,0.05144381,0.034295876,0.1097468,0.21263443,0.037725464,0.08573969,0.09945804,0.106317215,0.11317638,0.10288762,0.08573969,0.072021335,0.06516216,0.061732575,0.05144381,0.116605975,0.15090185,0.19548649,0.2709374,0.39783216,0.5418748,1.4953002,1.903421,1.605047,1.6427724,1.4267083,1.3581166,1.529596,2.3767042,4.6608095,5.003768,4.5510626,3.8891523,3.0729103,1.6153357,1.3958421,1.3203912,1.0357354,0.84024894,1.7010754,4.2423997,2.6236343,3.2272418,5.861165,3.789694,3.2066643,3.2203827,3.7519686,3.882293,1.8519772,0.77165717,0.24350071,0.048014224,0.037725464,0.13375391,0.19891608,1.2449403,3.3781435,6.591667,10.762046,12.665466,7.548522,2.534465,0.6207553,0.6756287,0.16462019,0.024007112,0.010288762,0.1097468,0.5453044,0.939707,1.1317638,0.8265306,0.26064864,0.17833854,0.21263443,0.08916927,0.3566771,0.77165717,0.28808534,0.37039545,0.15776102,0.0,0.06859175,0.34638834,0.6756287,0.7099246,0.65848076,0.6036074,0.48357183,0.12003556,0.34638834,0.53844523,0.4355576,0.15776102,0.34981793,0.4046913,0.39097297,0.37382504,0.432128,0.5761707,0.607037,0.607037,0.7407909,1.2826657,1.8245405,2.4761622,2.503599,1.99602,1.8554068,2.3458378,2.7162333,3.4810312,4.3933015,4.437886,4.2115335,4.355576,4.8494368,5.9743414,8.275595,9.6645775,10.216741,11.249047,12.88496,14.071597,12.891819,12.329367,12.734058,13.618892,13.663476,13.227919,13.375391,14.184773,15.158776,15.22051,16.280252,17.87501,18.166525,17.532051,18.581505,19.28457,19.432043,18.9519,18.152807,17.734396,17.408587,16.815268,16.45516,16.503176,16.828985,15.752095,15.858413,16.925014,18.115082,17.96418,17.556059,18.941612,19.991066,20.066517,20.02193,21.314886,22.36091,23.11542,23.705309,24.45296,26.455837,26.579304,26.116308,25.673891,25.156025,27.474424,26.058006,23.842491,22.679861,23.341772,26.133457,22.227156,17.586924,15.560039,16.877,21.699,27.282368,27.409264,23.811626,26.1849,23.821915,24.658733,32.99949,44.498898,46.172535,26.781649,17.192522,11.379372,6.800872,4.389872,5.9640527,4.6848164,4.170378,4.8117113,3.7794054,4.064061,4.091498,3.5804894,3.0214665,3.6627994,3.415869,3.5290456,3.8685746,4.4927597,5.669108,6.166398,6.2864337,6.540223,6.728851,5.967482,6.077229,5.9297566,5.809721,5.8371577,6.0052075,5.56965,5.0826488,4.4275975,3.758828,3.5290456,3.2821152,3.083199,2.8877127,2.7402403,2.7711067,2.7985435,2.7333813,2.7368107,2.8122618,2.819121,2.651071,2.6716487,2.8637056,3.0523329,2.9254382,2.9734523,3.2889743,3.5599117,3.6147852,3.4535947,3.4021509,3.4947495,3.8171308,4.383013,5.127233,6.5367937,7.3255987,7.891481,8.491658,9.211872,8.549961,8.354475,8.134981,7.5931067,6.6122446,6.866034,7.14726,7.4696417,7.623973,7.160979,7.3839016,7.671987,8.364764,9.448513,10.566559,11.067279,10.443094,9.325048,8.282454,7.7885933,7.658269,6.8454566,6.4990683,6.7322803,6.619104,6.790583,8.025234,9.006097,9.301042,9.366203,9.218731,8.436785,8.014946,7.781734,6.3961806,6.0052075,6.118384,6.5539417,7.39762,8.988949,9.602845,10.014396,10.429376,10.662587,10.120712,9.493098,8.611694,7.5279446,6.3893213,5.435896,4.887162,4.8768735,4.6608095,4.0366244,3.340418,2.6716487,2.4967396,3.000889,3.9028704,4.4584637,4.57507,4.972902,6.0052075,7.3393173,7.9875093,9.47595,10.182446,11.067279,12.140739,12.452832,14.819247,16.009314,16.510035,17.031332,18.499195,18.183672,18.897026,19.79901,20.7833,22.467228,21.832754,20.841602,19.682402,18.687822,18.348293,18.145947,18.197392,18.502625,18.756414,18.362011,18.831865,17.833855,16.280252,15.13134,15.361122,15.6252,16.029892,16.95931,17.63494,16.108772,14.843254,15.45715,17.29541,18.722118,17.144508,15.409137,14.123041,14.55174,16.256245,17.069057,18.145947,18.516342,18.20082,17.367432,16.328266,15.079896,13.745787,12.833516,12.428825,12.175035,0.5041494,0.6001778,0.607037,0.58302987,0.5453044,0.47328308,0.64476246,0.7510797,0.9877212,1.4027013,1.8931323,1.9171394,1.9685832,1.9068506,1.7250825,1.5398848,1.4678634,1.5501735,1.5364552,1.3855534,1.2517995,1.2380811,1.0254467,0.94656616,1.0666018,1.1763484,1.5638919,1.8108221,1.8691251,1.8382589,1.9239986,1.8245405,1.8005334,1.7936742,1.8519772,2.1194851,2.719663,2.7230926,3.882293,5.7136927,5.4941993,9.386781,18.04306,22.247734,18.526632,9.139851,5.099797,4.245829,4.3795834,4.1360826,2.976882,1.7319417,1.255229,1.1454822,1.1111864,0.9774324,0.7579388,0.59331864,0.48700142,0.4046913,0.26064864,0.2469303,0.20920484,0.2194936,0.28465575,0.31895164,0.5144381,0.64819205,0.6173257,0.45270553,0.30523327,0.32924038,0.29837412,0.25721905,0.216064,0.16804978,0.1920569,0.2709374,0.34638834,0.39783216,0.45613512,0.2503599,0.12346515,0.19891608,0.4629943,0.7922347,1.039165,0.8505377,0.5144381,0.21263443,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.030866288,0.006859175,0.14747226,0.29837412,0.32924038,0.12346515,0.072021335,0.024007112,0.0,0.0,0.0,0.037725464,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.010288762,0.044584636,0.020577524,0.006859175,0.0,0.0,0.0,0.01371835,0.041155048,0.061732575,0.048014224,0.0,0.0,0.017147938,0.024007112,0.017147938,0.030866288,0.116605975,0.16462019,0.18176813,0.17490897,0.1371835,0.2469303,0.31209245,0.37382504,0.5041494,0.8093826,0.7476501,0.4389872,0.30523327,0.42183927,0.5178677,0.5796003,0.4389872,0.34295875,0.38754338,0.53501564,0.40126175,0.31209245,0.28808534,0.37725464,0.67219913,0.67219913,0.7888051,0.8025235,0.6824879,0.61046654,0.48700142,0.4389872,0.41498008,0.40126175,0.4115505,0.40126175,0.2777966,0.2469303,0.30866286,0.26064864,0.11317638,0.11317638,0.1371835,0.14747226,0.18176813,0.25721905,0.18176813,0.24350071,0.45613512,0.5796003,0.4081209,0.3566771,0.31895164,0.3018037,0.4115505,0.25378948,0.45956472,0.6310441,0.6173257,0.5178677,0.8128122,0.7922347,0.7510797,0.83681935,1.0666018,0.8471081,1.0597426,1.3821237,1.5981878,1.587899,2.0646117,1.9891608,2.452155,3.6559403,4.914599,4.0229063,4.880303,6.2830043,7.1232533,6.3790326,9.403929,10.628291,11.458252,12.332796,12.710052,14.5414505,16.163645,17.693241,19.106232,20.217419,21.647556,22.837624,23.69502,24.322634,24.994833,23.588703,22.175713,21.671564,21.78817,21.057667,19.312008,16.80498,14.376831,12.843805,13.015285,12.747777,13.035862,13.025573,12.545431,12.130451,12.9981365,13.066729,13.71492,15.46401,17.991615,18.307138,18.852442,19.713268,20.906765,22.384918,23.396646,24.35693,26.42497,30.036327,34.882336,36.772038,36.689728,37.334488,39.80379,43.56262,45.62723,48.06567,51.824497,56.481876,60.240704,68.32081,82.1249,90.12613,89.90664,88.13697,91.02811,89.26187,89.18299,91.515114,91.37107,85.82886,82.57418,78.9834,71.54805,55.861122,44.179947,36.535397,29.981453,23.835632,19.69955,19.065077,20.02193,18.684393,15.29939,14.2362175,8.879202,6.276145,4.6127954,3.117495,2.0440342,1.4815818,1.1043272,0.90884066,0.7888051,0.53501564,0.59674823,0.78537554,1.6393428,2.5207467,1.6187652,1.0323058,0.6276145,0.4389872,0.36010668,0.15433143,0.0548734,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.030866288,0.030866288,0.030866288,0.030866288,0.024007112,0.0274367,0.07545093,0.09945804,0.061732575,0.061732575,0.14061308,0.274367,0.31209245,0.59674823,1.0220171,1.4095604,1.4953002,1.1523414,1.2037852,1.4369972,1.9514352,3.1586502,3.7553983,4.0263357,3.841138,3.0797696,1.6016173,0.9911508,0.6379033,0.6241849,1.2106444,2.8225505,3.7622573,2.369845,5.353586,10.467101,6.4990683,4.557922,2.7470996,1.3478279,0.5212973,0.29151493,0.106317215,0.024007112,0.0,0.0,0.0,0.024007112,0.09602845,0.51100856,1.8485477,4.976331,5.754848,2.4830213,0.1920569,0.2709374,0.4424168,0.1371835,0.041155048,0.017147938,0.06859175,0.34981793,0.06859175,0.90541106,0.9294182,0.22978236,0.89855194,0.1920569,0.006859175,0.5418748,1.0940384,0.030866288,0.006859175,0.0,0.0,0.2709374,1.3581166,0.8711152,0.85739684,0.84367853,0.6790583,0.53501564,0.216064,0.16462019,0.24350071,0.32924038,0.30523327,0.42869842,0.31895164,0.26407823,0.34638834,0.45613512,0.823101,1.0082988,0.9259886,0.84367853,1.3443983,1.6736387,1.6084765,1.2792361,1.2586586,2.5619018,2.5756202,2.0920484,2.3081124,3.474172,4.914599,4.8151407,4.8288593,5.579939,7.3118806,9.887501,11.156448,11.55771,12.562579,13.718349,12.617453,12.922686,12.679185,12.428825,12.161317,11.30735,10.696883,11.780633,12.603734,13.255356,15.868701,16.12592,16.400288,16.558048,16.678083,17.04505,18.166525,19.181683,19.29143,18.78385,19.027351,19.017063,19.058218,18.78385,18.11165,17.257685,15.426285,14.904987,15.265094,16.108772,17.075916,17.514904,20.378609,21.918493,21.62012,22.230585,21.901346,21.527521,21.966507,22.94051,23.02625,28.34897,29.587051,27.76937,24.288338,20.920483,22.981665,23.341772,22.151705,20.62211,21.013083,22.12427,19.891607,25.498983,33.194977,20.29287,26.006561,32.2587,30.92802,25.536709,31.2504,27.94085,35.197857,54.53387,74.25743,69.48687,35.475655,18.684393,12.202472,10.031544,7.06495,7.8949103,6.262427,5.4941993,6.036074,5.4633327,5.0346346,4.5270553,3.981751,3.6868064,4.149801,3.0626216,3.1963756,3.8617156,4.8151407,6.2555676,6.193835,5.8680243,6.1321025,6.64997,5.90575,6.0635104,5.8645945,5.9331865,6.2144127,5.9812007,5.164959,4.5853586,3.882293,3.1140654,2.7470996,2.5893385,2.4212887,2.369845,2.4658735,2.6236343,2.952875,2.7882545,2.6304936,2.5996273,2.4418662,2.1846473,2.294394,2.534465,2.7299516,2.7916842,2.534465,2.609916,2.7813954,2.942586,3.1140654,3.0386145,2.8945718,3.0454736,3.7108135,4.945465,5.895461,6.6568294,7.346176,8.100685,9.0644,9.22216,9.115844,8.786603,8.285883,7.675417,7.2364297,6.742569,7.06495,8.052671,8.529384,7.932636,7.6274023,7.864044,8.601405,9.489669,9.56512,8.786603,9.043822,10.511685,11.657167,10.569988,8.844906,8.110974,8.255017,7.4010496,7.377043,7.407909,7.6205435,8.097256,8.865483,8.865483,8.213862,8.375052,8.899779,7.4456344,5.4941993,5.3158607,5.8165803,6.728851,8.621983,9.156999,9.623423,10.189304,10.607714,10.192734,9.314759,7.6925645,6.1801167,5.2266912,4.897451,4.15323,4.4241676,4.4996185,4.0606318,3.707384,3.2443898,2.760818,3.1277838,4.029765,3.981751,4.7019644,5.8988905,5.9228973,5.3741636,7.0958166,8.779744,9.328478,10.487679,12.600305,14.603184,15.885849,16.736387,16.259674,15.532601,17.607502,17.645227,17.53548,18.554068,21.03709,24.384367,23.797907,22.607841,21.129688,19.689262,18.6158,18.921034,18.821575,19.219408,19.949911,19.792149,20.436913,20.093952,18.903887,17.669235,17.851004,17.302269,17.03819,16.609491,15.851553,14.863832,13.419975,14.500296,16.280252,17.463459,17.243965,17.010754,15.323397,14.644339,15.80011,17.960749,17.775553,17.583494,17.816708,18.12194,17.364002,16.80155,15.635489,14.085316,13.104454,14.373401,0.4424168,0.5007198,0.5178677,0.5590228,0.66533995,0.8745448,0.78194594,0.7133542,0.7682276,0.9294182,1.0871792,1.2655178,1.4747226,1.6667795,1.7250825,1.4438564,1.2826657,1.4953002,1.646202,1.5604624,1.3375391,1.2277923,1.0837497,0.9568549,0.89855194,0.980862,1.1934965,1.2277923,1.1934965,1.2449403,1.5570327,1.5090185,1.605047,1.7765263,1.8759843,1.704505,1.9925903,2.8911421,4.245829,5.8337283,7.3598948,14.555169,20.776442,20.70785,14.102464,5.7582774,4.2081037,3.426158,2.8328393,2.153781,1.4267083,0.97057325,0.85396725,0.823101,0.7682276,0.7339317,0.70649505,0.7373613,0.6824879,0.5418748,0.45613512,0.5007198,0.47671264,0.41840968,0.39783216,0.5041494,0.5624523,0.42526886,0.33609957,0.32238123,0.19548649,0.26750782,0.29494452,0.2709374,0.22292319,0.20577525,0.2194936,0.17833854,0.15776102,0.18176813,0.21263443,0.18176813,0.16804978,0.216064,0.34295875,0.52472687,0.9945804,1.1043272,0.8025235,0.29494452,0.0548734,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.0034295875,0.07888051,0.18862732,0.2469303,0.14747226,0.08916927,0.05144381,0.0274367,0.010288762,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.09945804,0.0548734,0.01371835,0.01371835,0.020577524,0.017147938,0.01371835,0.01371835,0.020577524,0.048014224,0.020577524,0.0274367,0.0274367,0.01371835,0.01371835,0.01371835,0.017147938,0.01371835,0.0034295875,0.006859175,0.12003556,0.20577525,0.33266997,0.4389872,0.34638834,0.26064864,0.25378948,0.29494452,0.35324752,0.4046913,0.4046913,0.51100856,0.53844523,0.45613512,0.4081209,0.40126175,0.36696586,0.28122616,0.21263443,0.33952916,0.4389872,0.45270553,0.45270553,0.48014224,0.548734,0.5693115,0.6036074,0.53501564,0.39783216,0.40126175,0.28122616,0.29837412,0.32581082,0.31895164,0.3018037,0.26064864,0.23321195,0.26064864,0.31209245,0.2709374,0.22292319,0.14404267,0.106317215,0.106317215,0.072021335,0.1371835,0.16462019,0.23321195,0.33609957,0.36010668,0.30523327,0.26064864,0.26750782,0.32581082,0.38754338,0.37382504,0.70649505,0.8745448,0.83338976,1.0185875,0.8711152,0.8265306,1.0357354,1.2963841,1.0185875,1.0528834,1.3409687,1.6427724,1.7490896,1.5124481,2.0886188,2.411,2.7882545,3.3026927,3.8274195,4.040054,5.06893,6.451054,7.5931067,7.795452,9.921797,10.31277,10.768905,11.8869505,13.077017,15.367981,17.175373,18.310568,19.03421,20.045938,21.486366,22.210009,22.323185,22.10712,22.02824,21.12283,20.742146,20.567236,20.423193,20.27572,18.149376,16.149927,14.4145565,13.155897,12.672326,13.029003,13.440554,13.629181,13.55373,13.413116,12.950122,13.186764,14.123041,15.402277,16.317978,18.265984,19.322296,20.011642,20.95135,22.847912,24.134007,26.157463,28.520449,31.26412,34.868614,37.941525,39.670036,40.520576,41.38826,43.57634,46.49835,49.818188,54.074306,58.481327,60.912903,69.97044,81.15433,85.235535,82.025444,80.37238,81.27436,79.775635,77.73503,75.20742,70.47116,64.16758,61.19413,59.314716,55.778812,47.31802,35.84948,29.871706,25.61216,22.144846,21.397196,19.970488,19.003344,17.017612,14.582606,14.321958,9.266746,6.108095,4.0229063,2.527606,1.4815818,1.1660597,0.864256,0.7373613,0.764798,0.7407909,0.5693115,0.8745448,1.5638919,2.0508933,1.2758065,0.7888051,0.65162164,0.48014224,0.274367,0.4081209,0.08573969,0.010288762,0.010288762,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.017147938,0.006859175,0.01371835,0.017147938,0.020577524,0.041155048,0.044584636,0.044584636,0.058302987,0.1097468,0.22635277,0.7407909,1.1214751,1.5398848,1.9651536,2.1674993,1.670209,1.5638919,1.646202,2.0234566,3.1346428,4.8940215,6.800872,8.014946,7.8023114,5.545643,3.7519686,1.9823016,1.4095604,2.0920484,2.9700227,3.2649672,2.8499873,3.1346428,4.1635194,4.6093655,4.0434837,2.201795,0.71678376,0.18862732,0.18176813,0.044584636,0.18862732,0.2709374,0.17833854,0.01371835,0.0274367,0.116605975,0.2194936,0.8779744,3.2409601,1.6599203,0.548734,0.06859175,0.15090185,0.48014224,0.23321195,0.25378948,0.4115505,0.58302987,0.66876954,0.13375391,0.18176813,0.18519773,0.044584636,0.18176813,0.037725464,0.4115505,0.5624523,0.30523327,0.006859175,0.14747226,0.24007112,0.70649505,1.2895249,1.0768905,1.3786942,1.5055889,1.2792361,0.8505377,0.6927767,0.97057325,0.7682276,0.52472687,0.6001778,1.2689474,0.5041494,0.37039545,0.3841138,0.39097297,0.5693115,0.5727411,0.9362774,1.1454822,1.1797781,1.5124481,1.3169615,2.270387,2.5173173,1.99602,2.4418662,2.6887965,2.527606,2.877424,3.7691166,4.338428,4.2526884,4.846007,5.9812007,7.6514096,9.97324,9.640571,10.755186,12.048141,12.662037,12.120162,11.612583,10.960961,10.847785,10.844356,9.403929,9.47595,10.511685,11.465111,12.181894,13.368532,14.287662,15.2033615,15.728088,16.029892,16.825556,17.851004,19.167965,20.104242,20.430052,20.382038,19.949911,19.740705,19.442331,18.914175,18.183672,16.578627,16.355703,16.554619,16.674654,16.671225,17.099922,19.071936,19.672113,18.962189,19.9602,21.623549,24.03798,26.476416,28.17749,28.359259,27.460707,25.629307,24.43924,23.537258,20.62554,19.085653,17.929884,16.314548,15.189643,17.288551,16.369421,12.048141,12.699762,15.731518,7.56224,20.395756,28.18435,28.451859,24.298628,24.415234,24.182022,34.463924,60.26471,90.56512,98.33313,43.47002,21.260014,14.870691,12.583157,7.7714453,8.484799,6.8385973,5.888602,5.960623,4.6436615,4.4413157,3.9680326,3.4673128,3.1415021,3.1380725,2.9700227,3.6285036,4.383013,5.0346346,5.926327,5.9914894,5.9469047,5.9983487,6.046363,5.672538,6.036074,5.9469047,5.970912,5.9434752,4.979761,4.2423997,3.899441,3.4673128,2.9048605,2.6373527,2.4487255,2.3321195,2.4247184,2.6304936,2.6133456,2.435007,2.4418662,2.4795918,2.4452958,2.294394,2.0303159,1.99602,2.1263442,2.318401,2.4384367,2.5138876,2.7711067,2.8739944,2.784825,2.7711067,2.9906003,2.983741,3.3644254,4.266407,5.3330083,5.857735,6.81802,7.840037,8.546532,8.56368,8.440215,8.296172,7.915488,7.4113383,7.2604365,6.4098988,6.3481665,6.711703,7.0375133,6.773435,7.1026754,7.425057,7.915488,8.549961,9.088407,9.091836,9.081548,9.033533,9.132992,9.753747,9.156999,8.378482,8.176137,8.539673,8.683716,8.951223,8.608265,8.690575,9.290752,9.561689,9.424506,9.14328,8.759167,8.289313,7.7131424,6.9620624,6.917478,7.0958166,7.64798,9.366203,10.381361,10.803201,10.611144,9.997248,9.386781,7.932636,6.927767,6.0395036,5.1992545,4.616225,4.1463714,4.046913,4.1635194,4.2355404,3.8925817,3.8857226,3.6936657,3.7485392,4.2766957,5.312431,5.48734,6.2830043,6.420188,6.1732574,7.3873315,9.170717,10.690024,12.291641,14.126471,16.12935,17.185663,18.78042,18.067066,15.824117,16.424294,17.984756,18.45461,18.78042,19.44576,20.464348,20.553518,20.467777,19.408035,17.799559,17.322845,18.54378,19.174824,19.288,19.586374,21.400625,22.196291,21.712719,20.488356,18.9519,17.425734,17.130789,17.322845,17.254255,16.798119,16.47231,15.354263,15.635489,16.321407,17.192522,18.766703,17.87158,16.266533,15.422854,15.71437,16.420864,15.848124,15.45715,15.13134,14.908417,14.973578,16.060759,16.180794,15.916716,15.789821,16.228807,0.5453044,0.5658819,0.5693115,0.58645946,0.65162164,0.7922347,0.7888051,0.764798,0.77165717,0.8093826,0.8025235,0.9259886,1.1351935,1.2963841,1.3478279,1.2895249,1.2998136,1.5330256,1.646202,1.5536032,1.4404267,1.255229,1.0837497,0.9534253,0.88826317,0.90198153,0.9877212,0.96371406,0.94656616,1.0734608,1.5193073,1.6221949,1.5090185,1.5673214,1.7353712,1.529596,2.1229146,3.57363,4.773986,6.368744,10.765475,17.833855,20.639257,17.329706,9.832627,3.8342788,3.3747141,2.767677,2.0989075,1.4918705,1.1214751,0.8196714,0.67219913,0.5796003,0.5178677,0.5418748,0.5178677,0.5658819,0.5727411,0.52815646,0.5590228,0.4664239,0.42869842,0.34981793,0.2709374,0.3566771,0.52815646,0.42183927,0.30866286,0.28465575,0.2503599,0.32924038,0.33266997,0.30523327,0.2777966,0.29494452,0.2503599,0.20920484,0.17833854,0.16462019,0.18862732,0.18519773,0.20577525,0.23321195,0.29151493,0.4389872,1.3443983,1.4987297,1.0631721,0.4081209,0.106317215,0.0274367,0.0034295875,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.006859175,0.006859175,0.05144381,0.116605975,0.16462019,0.13375391,0.12346515,0.18176813,0.21263443,0.17833854,0.09259886,0.061732575,0.0274367,0.006859175,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.024007112,0.082310095,0.0548734,0.020577524,0.01371835,0.006859175,0.006859175,0.006859175,0.006859175,0.010288762,0.024007112,0.024007112,0.017147938,0.006859175,0.0,0.006859175,0.006859175,0.006859175,0.0034295875,0.006859175,0.0274367,0.15090185,0.26750782,0.40126175,0.50757897,0.48014224,0.35324752,0.3806842,0.4115505,0.4081209,0.42526886,0.3841138,0.48700142,0.52472687,0.44927597,0.36353627,0.28122616,0.20920484,0.16119061,0.14747226,0.18862732,0.37725464,0.31552204,0.33952916,0.47328308,0.42869842,0.36353627,0.31209245,0.29151493,0.2777966,0.21263443,0.15090185,0.17147937,0.20920484,0.22292319,0.18176813,0.17833854,0.17490897,0.18862732,0.20920484,0.20234565,0.15433143,0.08916927,0.058302987,0.058302987,0.044584636,0.08573969,0.16462019,0.22292319,0.26064864,0.33266997,0.31552204,0.26750782,0.29151493,0.37039545,0.3806842,0.53158605,0.89855194,1.0631721,0.980862,0.980862,0.86082643,0.864256,0.9945804,1.1111864,0.89855194,1.2723769,1.2895249,1.3546871,1.5261664,1.5055889,1.9274281,2.2463799,2.5481834,2.9460156,3.5633414,4.1463714,5.06893,6.276145,7.4696417,8.131552,9.266746,9.493098,9.832627,10.662587,11.694893,14.009865,15.316538,16.067617,16.691803,17.607502,17.7927,18.362011,18.6158,18.434032,18.272842,18.262554,18.564358,18.999914,19.20569,18.643238,17.960749,16.756964,15.275383,13.937843,13.347955,13.488567,13.982429,14.164196,13.903547,13.594885,12.912396,13.183334,14.016724,14.623761,13.838386,15.940722,17.302269,18.437462,19.644676,20.995934,22.679861,25.18346,27.800236,30.399864,33.438477,35.780888,37.99983,40.259926,42.458294,44.22796,48.319458,51.70789,55.075745,58.717968,62.555676,70.971886,79.43268,82.11462,79.161736,76.67186,77.92366,79.95055,78.48268,73.36916,68.571175,65.12787,60.69684,55.490726,49.64328,43.202515,33.81916,27.676771,23.972816,22.000803,21.12283,18.9519,17.12736,15.337115,13.708061,12.795791,8.2481575,5.219832,3.216953,1.9548649,1.3443983,0.9328478,0.8745448,0.9431366,1.0014396,0.9945804,0.91569984,1.1249046,1.5741806,1.8005334,0.91569984,0.5555932,0.45956472,0.33266997,0.15776102,0.216064,0.044584636,0.0034295875,0.0034295875,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.010288762,0.0034295875,0.0034295875,0.006859175,0.006859175,0.017147938,0.017147938,0.01371835,0.017147938,0.020577524,0.037725464,0.037725464,0.058302987,0.14061308,0.32238123,1.4987297,2.0406046,2.6647894,3.3781435,3.4776018,2.3767042,2.2292318,2.270387,2.5447538,3.9165888,5.826869,8.683716,10.535692,10.494537,8.7283,7.284444,5.06893,3.4535947,3.3438478,5.1752477,4.0709205,4.9420357,4.5201964,3.100347,4.5099077,3.6456516,1.762808,0.41498008,0.07888051,0.14404267,0.29837412,0.38754338,0.31895164,0.14061308,0.01371835,0.048014224,0.16119061,0.22292319,0.4046913,1.1866373,0.28808534,0.07888051,0.06516216,0.14747226,0.65162164,0.34638834,0.32238123,0.48014224,0.65848076,0.6379033,0.4355576,0.31209245,0.4972902,0.77851635,0.5212973,0.6310441,0.4698535,0.22978236,0.05144381,0.0,0.072021335,0.4389872,0.7579388,0.94656616,1.1729189,1.3341095,1.3238207,1.1626302,0.9431366,0.84367853,0.764798,0.5727411,0.39097297,0.45613512,1.1180456,0.50757897,0.42183927,0.4081209,0.36353627,0.5212973,0.5761707,0.8505377,1.1592005,1.3684053,1.3821237,1.5570327,2.1674993,2.2841053,1.9857311,2.3561265,2.170929,2.3081124,2.8534167,3.5050385,3.5633414,3.9714622,4.835718,5.9434752,7.3050213,9.153569,9.637141,11.324498,12.229909,11.900668,11.417097,10.878652,9.993818,9.321619,8.882631,8.165848,8.944365,10.39165,11.550851,12.22305,12.977559,13.831526,14.71636,15.560039,16.239098,16.578627,17.007324,18.235117,19.274282,19.819586,20.255144,20.224277,20.001354,19.558937,19.013634,18.608942,17.916164,18.605513,18.907316,18.269413,17.367432,17.398296,18.108221,18.45461,18.45461,19.164536,20.821026,25.032558,29.01774,30.969175,30.043186,26.905113,23.571554,22.751883,23.266321,20.03222,17.346853,16.098484,14.102464,12.123591,13.865822,13.413116,12.099585,13.2690735,15.199932,11.087856,19.52807,23.825344,23.60242,20.913624,20.268862,19.267422,23.972816,39.24477,59.50677,68.74265,33.218983,18.04649,12.826657,10.628291,7.966932,9.55826,7.9875093,7.301592,7.658269,5.329579,4.465323,4.15666,3.6353626,2.9871707,3.1586502,3.2478194,3.7142432,4.40702,5.113515,5.56965,5.8062916,6.0806584,6.0806584,5.7925735,5.4976287,5.8165803,5.3913116,5.0277753,4.787704,3.9714622,3.3815732,3.199805,2.9494452,2.6064866,2.5893385,2.2566686,2.3389788,2.503599,2.585909,2.5824795,2.510458,2.4007113,2.2258022,2.0303159,1.9274281,1.9239986,1.9342873,2.0337453,2.1983654,2.3046827,2.486451,2.784825,2.884283,2.750529,2.6407824,2.9460156,3.117495,3.6216443,4.5442033,5.579939,6.111525,6.742569,7.3393173,7.781734,7.970361,8.529384,8.361334,7.630832,6.6568294,5.90232,5.5490727,6.1972647,6.931196,7.233,6.9723516,7.630832,8.045813,8.299602,8.467651,8.601405,8.275595,8.152129,8.131552,8.30646,8.947794,9.187865,8.707723,8.340756,8.40249,8.683716,8.868914,8.81747,9.184435,9.743458,9.369633,9.571979,9.455373,9.102125,8.762596,8.824328,8.529384,8.323608,8.423067,9.095266,10.6488695,11.427385,11.574858,10.8958,9.695444,8.766026,7.8846216,7.373613,6.4236174,5.0757895,4.2081037,3.8274195,3.7622573,3.8960114,4.016047,3.799983,4.400161,4.5030484,4.331569,4.4687524,5.8474464,5.9571934,6.4887795,6.636252,6.56766,7.4353456,9.342196,11.183885,12.80608,14.2190695,15.611482,17.134218,19.294859,19.634388,17.837284,15.724659,18.063637,18.934752,19.11995,19.003344,18.578075,19.229696,19.548649,18.969048,17.751545,16.997036,17.936743,18.523201,19.05136,19.847023,21.246294,22.5221,22.480946,21.225718,19.315437,17.748116,16.756964,16.252815,16.194511,16.444872,16.774113,16.911295,17.072487,17.62465,18.646667,19.95677,17.71382,16.37971,15.947581,15.909856,15.251375,15.083325,15.3817,15.577187,15.46401,15.206791,16.173935,16.335125,16.331696,16.317978,15.971589,0.6379033,0.65848076,0.69963586,0.72707254,0.72364295,0.6962063,0.6962063,0.7373613,0.7922347,0.823101,0.7888051,0.8745448,1.039165,1.1214751,1.1146159,1.1866373,1.3066728,1.4850113,1.5227368,1.4369972,1.4472859,1.2277923,1.0768905,0.980862,0.9328478,0.922559,0.980862,0.9774324,0.9911508,1.1454822,1.6187652,1.821111,1.5707511,1.5193073,1.704505,1.5604624,2.7230926,4.3658648,5.9434752,8.639131,15.343974,19.414894,17.895588,12.607163,6.3618846,2.952875,2.469303,1.9685832,1.5124481,1.1729189,0.99801,0.7579388,0.5796003,0.45613512,0.40126175,0.4389872,0.39440256,0.432128,0.45956472,0.4664239,0.5144381,0.33952916,0.28808534,0.24350071,0.1920569,0.23664154,0.4629943,0.48014224,0.41840968,0.35324752,0.32238123,0.37725464,0.37382504,0.34638834,0.33609957,0.36353627,0.28808534,0.25721905,0.22635277,0.18519773,0.17833854,0.19548649,0.20234565,0.20577525,0.25378948,0.45613512,1.4507155,1.6084765,1.1351935,0.4355576,0.13032432,0.030866288,0.0034295875,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0,0.006859175,0.034295876,0.0548734,0.08916927,0.14061308,0.21263443,0.3566771,0.5521636,0.66533995,0.6207553,0.4081209,0.23321195,0.09602845,0.024007112,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.017147938,0.034295876,0.024007112,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.030866288,0.09945804,0.20234565,0.30866286,0.39783216,0.47328308,0.5521636,0.4698535,0.4938606,0.48357183,0.44584638,0.5144381,0.4389872,0.41840968,0.3806842,0.30866286,0.26407823,0.216064,0.14404267,0.13375391,0.17147937,0.13375391,0.28465575,0.21263443,0.24350071,0.37382504,0.29151493,0.2503599,0.15090185,0.15090185,0.20577525,0.10288762,0.06859175,0.08916927,0.11317638,0.116605975,0.116605975,0.12003556,0.106317215,0.11317638,0.13032432,0.09602845,0.07545093,0.041155048,0.030866288,0.041155048,0.058302987,0.09602845,0.17147937,0.22292319,0.26064864,0.3806842,0.37039545,0.29494452,0.32581082,0.42526886,0.34638834,0.607037,1.039165,1.2689474,1.2037852,1.0288762,0.85396725,0.823101,0.90884066,0.9945804,0.86082643,1.2895249,1.0837497,1.0357354,1.3169615,1.4850113,1.7216529,2.0646117,2.3835633,2.7745364,3.5770597,4.307562,5.1752477,6.138962,7.0958166,7.874333,8.158989,8.635701,9.139851,9.688584,10.491108,12.082437,13.022143,13.694343,14.287662,14.822677,14.850114,15.5085945,15.827546,15.63206,15.577187,16.441442,16.938732,17.432592,17.689812,16.86671,17.278261,16.80155,15.758954,14.668345,14.239647,14.2190695,14.452282,13.88983,12.668896,12.106443,11.945253,12.315649,12.627741,12.356804,11.032983,12.898679,14.448852,16.431154,18.523201,19.360022,21.064526,23.650434,26.496992,29.237232,31.76141,33.160683,34.961216,37.711742,41.000717,43.442585,48.731007,52.071426,55.1169,58.7797,63.25188,72.309425,80.33123,83.12634,80.55758,76.56211,79.7722,84.20666,83.63049,78.94567,78.15687,75.392624,66.66432,56.69451,48.54581,43.62435,34.738293,28.414133,24.418663,21.939072,19.593233,17.36057,15.340545,13.368532,11.379372,9.407358,6.029215,3.782835,2.3149714,1.4369972,1.1214751,0.7956643,0.8676856,1.0631721,1.2037852,1.214074,1.2929544,1.4987297,1.7422304,1.7113642,0.86082643,0.5007198,0.33952916,0.23664154,0.14061308,0.08916927,0.030866288,0.010288762,0.006859175,0.01371835,0.024007112,0.030866288,0.034295876,0.0274367,0.020577524,0.010288762,0.01371835,0.006859175,0.0034295875,0.006859175,0.006859175,0.020577524,0.01371835,0.01371835,0.020577524,0.01371835,0.024007112,0.030866288,0.061732575,0.16119061,0.37725464,1.3889829,2.085189,3.0283258,3.998899,4.0091877,2.7711067,3.0214665,3.2135234,3.2992632,4.7328305,7.1129646,9.256456,10.686595,11.067279,10.233889,8.659708,6.475061,5.3707337,5.9571934,7.73372,5.2335505,6.6225333,6.307011,3.9611735,4.554492,3.0729103,1.4541451,0.4081209,0.09602845,0.106317215,0.42526886,0.61046654,0.52815646,0.28465575,0.23664154,0.10288762,0.15776102,0.37725464,0.51100856,0.07545093,0.037725464,0.3841138,0.40126175,0.18176813,0.6241849,0.42869842,0.35324752,0.3806842,0.45270553,0.48357183,0.9431366,0.83338976,0.823101,1.0048691,0.9259886,1.0254467,0.64819205,0.22978236,0.037725464,0.15776102,0.274367,0.607037,0.75450927,0.7510797,1.0425946,1.08032,1.0494537,0.9568549,0.88826317,1.0117283,0.58988905,0.36010668,0.24007112,0.26407823,0.6173257,0.47671264,0.51100856,0.53158605,0.51100856,0.5761707,0.64133286,0.84367853,1.1832076,1.4987297,1.4747226,1.8588364,1.862266,1.8005334,1.8416885,2.0097382,1.7250825,1.9925903,2.6716487,3.3815732,3.508468,3.9783216,5.4187484,6.756287,7.6925645,8.669997,10.021255,11.080997,11.355364,10.912948,10.39165,9.914937,9.1981535,8.495089,8.035523,8.038953,9.338767,10.254466,11.002116,11.742908,12.590015,13.680624,14.493437,15.227368,15.933864,16.523752,16.63007,17.63494,18.560926,19.075365,19.504065,20.063087,20.004784,19.661825,19.45262,19.8676,19.555508,20.145397,19.836735,18.386019,17.134218,16.770683,16.722668,17.069057,17.744686,18.512913,19.644676,23.653864,27.18634,28.486153,27.381826,24.826784,21.685282,21.064526,21.891056,18.883308,17.000465,17.103354,14.387119,10.055551,11.303921,11.80121,12.576297,14.994157,17.12736,13.745787,17.04505,17.53891,16.523752,15.275383,15.0456,13.039291,13.361672,18.879879,28.324963,36.288464,19.86074,12.511135,9.379922,8.117833,8.903209,10.563129,9.362774,9.054111,9.379922,6.0497923,4.770556,4.479041,3.9131594,3.0454736,3.1106358,3.3850029,3.7691166,4.3658648,5.0106273,5.271276,5.3158607,5.6656785,5.751418,5.4496145,5.0757895,5.003768,4.2835546,3.782835,3.5976372,3.0557625,2.7402403,2.6613598,2.49331,2.2806756,2.4384367,2.1091962,2.287535,2.4418662,2.4075704,2.386993,2.5207467,2.411,2.1332035,1.8485477,1.786815,1.8965619,1.937717,2.0714707,2.2635276,2.2806756,2.4418662,2.6476414,2.74367,2.6990852,2.5893385,2.9082901,3.2409601,3.8479972,4.763697,5.7925735,6.355026,6.461343,6.334448,6.327589,6.9346256,8.001227,7.829748,6.9723516,5.936616,5.1752477,5.7274113,6.636252,7.3255987,7.4936485,7.1266828,7.5107965,7.7542973,7.8366075,7.822889,7.857185,7.414768,7.2535777,7.5553813,8.282454,9.174147,9.853205,9.31133,8.868914,8.851766,8.567109,8.47451,8.951223,9.489669,9.633711,8.97866,9.39707,9.448513,9.119273,8.80718,9.314759,9.016385,8.597976,8.721441,9.613133,11.067279,11.979549,12.003556,10.971251,9.39021,8.405919,8.049242,7.966932,7.208993,5.874883,5.0826488,4.8185706,4.6745276,4.5647807,4.4413157,4.2869844,4.839148,5.1066556,4.9934793,4.931747,5.8645945,6.101236,6.800872,7.14726,7.1884155,7.829748,9.427936,11.365653,12.939834,13.999576,14.959861,16.095055,18.02934,19.167965,18.392878,15.055889,17.504614,18.694681,19.428614,19.78186,19.11652,19.329155,19.325726,19.157675,18.656956,17.425734,18.331144,18.907316,19.510923,20.241425,20.941061,22.834194,22.789608,21.623549,20.059656,18.71183,16.664366,15.391989,15.608052,16.901007,17.744686,18.265984,18.338005,18.656956,19.329155,19.871029,17.511473,16.6335,16.657507,16.726099,15.707511,15.638919,16.55119,17.610931,18.176813,17.799559,18.190533,17.943602,17.339994,16.736387,16.554619,0.72707254,0.7579388,0.85396725,0.90541106,0.8745448,0.7990939,0.6893471,0.70649505,0.78194594,0.864256,0.9259886,1.0494537,1.1934965,1.2655178,1.2449403,1.196926,1.2826657,1.3752645,1.371835,1.3032433,1.3203912,1.1283343,1.0871792,1.0563129,1.0082988,1.0494537,1.1797781,1.1934965,1.2277923,1.3855534,1.762808,1.9548649,1.7490896,1.7182233,1.978872,2.170929,3.8308492,5.130663,7.5279446,12.168177,19.87789,19.260563,13.577737,7.671987,3.9851806,2.5550427,1.5810398,1.097468,0.864256,0.7339317,0.65162164,0.5555932,0.490431,0.42526886,0.36353627,0.36353627,0.3566771,0.39783216,0.4081209,0.37725464,0.35324752,0.22978236,0.18176813,0.19891608,0.24007112,0.23321195,0.37382504,0.45956472,0.48357183,0.4389872,0.33609957,0.33952916,0.36353627,0.37382504,0.36353627,0.36353627,0.30523327,0.26750782,0.22635277,0.17833854,0.1371835,0.18519773,0.17147937,0.15776102,0.25721905,0.64133286,1.1866373,1.3032433,0.9362774,0.34638834,0.1097468,0.030866288,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.024007112,0.09602845,0.13375391,0.15776102,0.216064,0.3566771,0.65162164,1.0185875,1.2792361,1.2792361,0.8745448,0.48014224,0.19548649,0.0548734,0.024007112,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.048014224,0.14747226,0.20577525,0.26750782,0.31209245,0.36353627,0.47328308,0.4698535,0.4698535,0.432128,0.39440256,0.48357183,0.4046913,0.31552204,0.19891608,0.106317215,0.14061308,0.19548649,0.18519773,0.18862732,0.20577525,0.16119061,0.23664154,0.25721905,0.274367,0.2709374,0.18176813,0.25378948,0.16804978,0.116605975,0.13032432,0.072021335,0.037725464,0.06859175,0.06859175,0.041155048,0.09602845,0.06859175,0.037725464,0.058302987,0.09259886,0.01371835,0.044584636,0.030866288,0.034295876,0.06516216,0.08916927,0.15090185,0.20234565,0.24350071,0.29494452,0.40126175,0.39097297,0.29494452,0.34638834,0.4698535,0.31552204,0.5693115,1.039165,1.3375391,1.3238207,1.1214751,0.85396725,0.7407909,0.8779744,1.1008976,0.980862,1.1660597,0.939707,0.9328478,1.2517995,1.471293,1.6907866,2.153781,2.551613,2.9734523,3.8925817,4.664239,5.501058,6.2487082,6.831738,7.2364297,7.2021337,7.881192,8.628842,9.242738,9.966381,10.566559,11.393089,12.168177,12.6757555,12.761495,13.642899,14.356253,14.544881,14.318527,14.2362175,15.752095,16.04361,16.03675,16.029892,15.6869335,16.407146,16.540901,16.064188,15.309678,14.973578,14.706071,14.116182,12.46998,10.408798,9.945804,10.179015,10.847785,10.751757,9.897789,9.510246,10.837497,12.603734,15.37827,18.313997,19.150816,20.567236,23.053686,25.913963,28.571894,30.571342,31.524769,32.707977,34.937206,38.215893,41.73122,47.657547,50.79562,54.314377,58.92031,62.840332,73.34173,83.20865,86.80629,84.007744,80.19747,85.307556,89.66313,89.88263,88.10267,91.95067,86.188965,71.46917,57.69252,49.63642,46.940765,35.93522,29.837412,25.468117,21.349182,17.71382,15.566897,13.670336,11.039842,7.8846216,5.6210938,3.5770597,2.3218307,1.5604624,1.0837497,0.77851635,0.70649505,0.7442205,0.9259886,1.1729189,1.2895249,1.5433143,1.9651536,2.1469216,1.8759843,1.1351935,0.6344737,0.39097297,0.32924038,0.32238123,0.20577525,0.08916927,0.06516216,0.061732575,0.048014224,0.05144381,0.048014224,0.048014224,0.037725464,0.020577524,0.0,0.010288762,0.0034295875,0.0034295875,0.01371835,0.01371835,0.01371835,0.0034295875,0.010288762,0.024007112,0.017147938,0.0034295875,0.020577524,0.072021335,0.17833854,0.36010668,0.64476246,1.371835,2.3286898,3.0900583,3.0420442,2.4967396,3.3301294,3.7794054,3.806842,5.1238036,7.8194594,8.399059,8.961512,9.904649,9.938945,7.73029,5.936616,6.7322803,9.177576,9.211872,6.036074,6.8797526,6.790583,4.8288593,4.0366244,2.510458,1.3443983,0.5590228,0.15433143,0.08916927,0.29837412,0.90198153,1.2929544,1.2106444,0.7579388,0.32238123,0.17490897,0.44584638,0.71678376,0.024007112,0.0034295875,0.66533995,0.72364295,0.19548649,0.37725464,0.45956472,0.4664239,0.40126175,0.36010668,0.5144381,1.2277923,1.1317638,0.7888051,0.6173257,0.8711152,0.8471081,0.90884066,0.64819205,0.25721905,0.51100856,0.78194594,0.72364295,0.84367853,1.0837497,0.7990939,0.8711152,1.0460242,1.039165,0.90541106,1.0494537,0.64133286,0.3566771,0.25378948,0.3018037,0.35324752,0.53844523,0.6962063,0.7510797,0.72364295,0.7339317,0.72707254,0.97057325,1.2998136,1.5741806,1.6770682,1.8725548,1.6770682,1.6804979,1.8416885,1.4815818,1.4918705,1.7799559,2.534465,3.4810312,3.865145,3.9268777,5.785714,7.4799304,8.351046,9.043822,10.264755,10.155008,9.9869585,10.086417,9.822338,9.270175,8.841476,8.488229,8.323608,8.628842,10.124143,9.918367,9.918367,10.734609,11.688034,13.461131,14.352823,14.572317,14.843254,16.424294,16.492886,17.353712,18.255693,18.756414,18.725548,19.281141,19.229696,19.233126,19.908754,21.836184,21.081675,20.344313,18.831865,16.877,15.940722,15.29939,15.069608,15.402277,16.331696,17.768692,18.571217,20.759293,22.336903,22.673002,22.498095,21.356041,19.44919,18.9519,19.36688,17.545769,17.367432,18.694681,15.086755,8.694004,10.261326,9.993818,10.484249,13.176475,15.46401,10.714031,12.075578,11.015835,9.777754,9.239308,8.934075,7.291303,7.0272245,10.357354,17.418875,26.274069,13.71492,8.505377,6.941485,7.442205,10.583707,11.718901,11.369082,10.813489,9.709162,6.108095,5.127233,4.5030484,3.8788633,3.2546785,2.983741,3.415869,3.9028704,4.3007026,4.5990767,4.9180284,4.605936,4.804852,4.931747,4.73969,4.314421,3.7931237,3.07634,2.7711067,2.8156912,2.4761622,2.417859,2.3664153,2.2052248,2.0440342,2.2223728,2.0165975,2.1023371,2.177788,2.136633,2.037175,2.2463799,2.270387,2.1194851,1.9239986,1.8965619,1.862266,1.8554068,2.037175,2.2978237,2.277246,2.3972816,2.4967396,2.5619018,2.5756202,2.534465,2.8019729,3.2889743,4.0606318,4.996909,5.796003,6.1801167,5.885172,5.2747054,4.955754,5.778855,6.601956,6.540223,6.036074,5.5490727,5.5730796,6.7391396,7.349606,7.5862474,7.4765005,6.90033,6.615674,6.478491,6.451054,6.526505,6.759717,6.5333643,6.7494283,7.500508,8.611694,9.661148,10.240748,9.637141,9.352485,9.441654,8.543102,8.275595,9.084977,9.719451,9.6645775,9.126132,9.352485,9.386781,8.8929205,8.303031,8.803751,8.628842,8.189855,8.241299,9.057541,10.429376,11.921246,12.089295,11.005547,9.386781,8.587687,8.169277,8.320179,8.165848,7.5931067,7.267296,6.7391396,6.1801167,5.73427,5.4667625,5.3741636,5.3261495,5.518206,5.610805,5.5559316,5.6005163,5.970912,7.1061053,7.9189177,8.2310095,8.796892,9.678296,11.410237,12.833516,13.697772,14.640909,14.71636,15.906426,16.842705,16.486027,14.150477,16.228807,17.741257,19.507494,21.095392,20.807306,19.733847,19.03421,19.164536,19.493774,18.28999,19.665255,20.649546,20.96164,20.882757,21.273731,23.52354,22.926792,21.904776,21.174273,19.730417,16.63007,15.155347,15.999025,18.296848,19.600092,19.6241,19.459478,19.20912,19.047928,19.229696,17.899017,17.350283,17.46003,17.686382,17.089634,17.113642,18.221397,19.836735,21.20171,21.37319,21.211998,20.4472,19.20569,18.245405,18.95876,1.0082988,0.97057325,0.9602845,0.89855194,0.86082643,1.0666018,1.1043272,0.9774324,0.8848336,0.94999576,1.2037852,1.3409687,1.5021594,1.6359133,1.6359133,1.3443983,1.3924125,1.4232788,1.3786942,1.2620882,1.1146159,1.0288762,1.1180456,1.1729189,1.1832076,1.3443983,1.5501735,1.5193073,1.5810398,1.8005334,1.9823016,2.0577524,1.8999915,2.0063086,2.6956558,4.1360826,5.953764,6.025785,8.580828,14.7026415,22.309467,17.106783,9.493098,4.3109913,2.6647894,1.9068506,1.0048691,0.59674823,0.37382504,0.2469303,0.31895164,0.29494452,0.37382504,0.37382504,0.26407823,0.16804978,0.22978236,0.24350071,0.22635277,0.19548649,0.18176813,0.14747226,0.12689474,0.19548649,0.28122616,0.18176813,0.20920484,0.21263443,0.274367,0.34638834,0.274367,0.18862732,0.26064864,0.33266997,0.33952916,0.29151493,0.24007112,0.22978236,0.19891608,0.16119061,0.19891608,0.18519773,0.17490897,0.20577525,0.44584638,1.1900668,0.94656616,0.7476501,0.47328308,0.17147937,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.061732575,0.23321195,0.3566771,0.4115505,0.4046913,0.3806842,0.5761707,1.1489118,1.728512,1.8999915,1.2037852,0.6927767,0.29837412,0.07888051,0.01371835,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.116605975,0.13032432,0.044584636,0.12003556,0.26407823,0.34638834,0.32238123,0.274367,0.22635277,0.12346515,0.061732575,0.07888051,0.15090185,0.17833854,0.17490897,0.14404267,0.12346515,0.19891608,0.31895164,0.33266997,0.33952916,0.32924038,0.18176813,0.24350071,0.21263443,0.13375391,0.061732575,0.061732575,0.072021335,0.09602845,0.09602845,0.072021335,0.061732575,0.01371835,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.061732575,0.11317638,0.1371835,0.19891608,0.28808534,0.29837412,0.25721905,0.30523327,0.29151493,0.2709374,0.34638834,0.45956472,0.4115505,0.45956472,0.7099246,0.881404,0.8265306,0.53501564,0.8162418,0.8025235,0.8265306,1.0048691,1.2346514,1.2346514,1.0906088,1.0357354,1.1900668,1.5570327,2.1194851,2.5070283,2.9391565,3.6970954,5.127233,5.5662203,5.9983487,6.636252,7.051232,6.1492505,6.8557453,7.034084,7.716572,8.831187,9.184435,9.832627,10.196163,10.707172,11.345076,11.626302,11.869802,12.096155,12.706621,13.368532,13.015285,14.932424,14.925565,14.675205,15.001016,15.868701,17.418875,18.310568,17.785841,16.314548,15.594335,13.824667,11.7257595,9.9869585,9.163857,9.688584,8.81061,10.065839,10.72432,10.593996,12.024134,11.585147,13.780083,16.643787,18.95533,20.248285,21.712719,24.185452,26.42497,28.18092,30.18037,30.890295,32.27585,34.875473,38.49712,42.221653,47.28715,49.286602,52.60644,58.066345,62.912354,71.77441,83.38356,87.86946,85.83572,88.36332,92.73261,96.13134,98.43259,100.23998,102.88763,93.31908,74.291725,58.84829,51.81421,49.7736,35.407063,28.976585,24.826784,20.471207,16.602633,12.953552,11.252477,8.519095,5.086078,4.6093655,2.644212,1.7216529,1.3238207,1.0700313,0.71678376,0.5453044,0.5761707,0.6790583,0.8265306,1.0837497,1.7182233,2.5173173,2.8911421,2.5378947,1.4644338,0.8162418,0.5453044,0.6241849,0.764798,0.4115505,0.17833854,0.22292319,0.22292319,0.09945804,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.017147938,0.030866288,0.006859175,0.0274367,0.12003556,0.26407823,0.39783216,0.9328478,1.3992717,1.3375391,0.8471081,0.5658819,1.3443983,2.1194851,2.6750782,3.3301294,4.928317,5.5147767,6.293293,7.0923867,7.8263187,8.498518,7.1198235,6.355026,8.06296,10.532263,8.467651,6.0154963,5.6656785,5.7719955,5.171818,3.2203827,2.620205,1.5364552,0.6241849,0.18519773,0.19891608,0.12346515,1.3615463,3.0386145,3.7485392,1.5261664,0.96371406,0.4115505,0.082310095,0.0,0.0,0.0,0.0274367,0.082310095,0.15776102,0.24350071,0.45270553,0.7682276,0.96371406,1.0151579,1.1146159,0.48014224,0.44927597,0.6927767,0.8093826,0.31895164,0.30866286,0.70649505,0.97057325,0.9602845,0.9602845,1.1454822,0.7407909,0.7407909,1.2037852,1.2517995,0.8848336,1.3169615,1.6873571,1.5021594,0.61046654,0.32924038,0.21263443,0.42183927,0.7682276,0.7339317,0.91569984,1.0425946,0.85396725,0.5418748,0.7476501,0.9568549,1.2346514,1.4678634,1.5158776,1.2346514,1.4438564,1.6976458,1.9342873,1.920569,1.2346514,1.0528834,1.5090185,2.4315774,3.2683969,3.0969174,3.0969174,3.7211025,4.945465,6.941485,10.055551,10.398509,10.978109,11.002116,10.714031,11.396519,10.837497,10.045261,8.9100685,8.032094,8.7283,9.997248,10.196163,10.343636,10.820349,11.382801,13.505715,14.387119,14.105893,13.786942,15.594335,15.155347,16.108772,17.19938,17.87158,18.248835,17.261114,16.46545,16.702091,18.674105,22.933651,21.554956,19.45262,17.384579,15.978448,15.748666,14.771234,14.225929,14.4317045,15.597764,17.806417,18.392878,18.924463,19.613811,20.27572,20.323736,18.6158,17.556059,17.189093,17.21653,16.983316,17.861292,17.137648,13.183334,8.858624,11.519984,6.358455,7.3187394,10.63858,12.593445,9.506817,9.225591,9.266746,8.320179,6.6533995,6.1046658,5.7994323,4.1463714,8.632272,20.29287,33.719704,20.27915,10.285333,7.0443726,9.410788,11.780633,14.037301,15.169065,12.55915,7.5759587,5.5833683,5.4153185,3.9783216,3.2786856,3.6696587,3.875434,3.9371665,4.0057583,3.8479972,3.6868064,4.2115335,4.149801,4.280125,4.0674906,3.5461934,3.3266997,2.959734,2.5756202,2.3972816,2.4624438,2.609916,2.4761622,2.2841053,2.1332035,2.0886188,2.1983654,1.903421,1.7765263,1.7525192,1.7593783,1.7079345,1.9171394,1.821111,1.7662375,1.8382589,1.862266,1.6290541,1.5536032,1.6942163,1.9823016,2.2292318,2.386993,2.5893385,2.5961976,2.435007,2.411,2.4830213,3.1723683,4.245829,5.171818,5.1100855,5.0757895,4.8014226,4.557922,4.6676683,5.5250654,5.3398676,5.641671,5.967482,6.183546,6.4990683,7.1095347,7.3530354,7.507367,7.6445503,7.6445503,6.7048435,5.8200097,5.161529,4.9180284,5.295283,5.381023,6.1149545,7.130112,8.134981,8.940934,9.345626,9.115844,8.683716,8.261876,7.857185,7.9429245,8.460793,9.736599,11.043272,10.604284,10.261326,9.482809,8.879202,8.536243,8.011517,8.937505,8.913498,8.567109,8.601405,9.794902,11.345076,11.760056,11.399949,10.624862,9.794902,8.820899,8.7317295,8.958082,9.194724,9.414218,7.2158523,5.9640527,5.658819,5.970912,6.2418494,6.0566516,5.857735,5.826869,5.796003,5.2335505,5.672538,6.90033,8.292743,9.445084,10.179015,10.484249,11.118723,11.842365,12.641459,13.701202,13.920695,15.049029,14.808959,13.296511,12.953552,14.455711,16.352274,19.109661,21.527521,20.721567,18.732407,17.686382,18.019053,19.095943,19.181683,20.594673,22.36091,23.005672,22.494663,22.20315,23.983105,23.091412,22.011093,21.328604,19.730417,15.71437,14.781522,16.204802,18.770132,20.797018,21.211998,20.968498,20.37175,19.936192,20.402617,19.167965,18.190533,17.734396,17.518333,16.722668,18.554068,19.726988,21.013083,22.474087,23.437801,22.374628,20.920483,20.45063,21.181131,22.172283,0.8471081,0.8505377,0.823101,0.7510797,0.7099246,0.8471081,0.9534253,1.0117283,1.0666018,1.1934965,1.4987297,1.6633499,1.5227368,1.4198492,1.4369972,1.4267083,1.7216529,1.8142518,1.6736387,1.4027013,1.2483698,1.2998136,1.605047,1.6016173,1.3272504,1.4164196,1.8588364,2.0989075,2.2909644,2.4384367,2.386993,2.6853669,2.386993,2.417859,3.216953,4.746549,6.574519,7.2775846,10.347065,15.690363,19.6241,13.906977,7.6171136,3.3850029,1.7113642,0.9431366,0.70306545,0.4972902,0.34638834,0.2777966,0.33266997,0.33609957,0.37039545,0.36353627,0.33952916,0.38754338,0.41840968,0.28122616,0.17490897,0.15090185,0.1097468,0.12346515,0.10288762,0.16804978,0.28122616,0.23321195,0.274367,0.25721905,0.28122616,0.34638834,0.36010668,0.42183927,0.39440256,0.41498008,0.45270553,0.31552204,0.28465575,0.2709374,0.26407823,0.28465575,0.3806842,0.4664239,0.5144381,0.5658819,0.7922347,1.5090185,1.6359133,1.0837497,0.51100856,0.20577525,0.08573969,0.0274367,0.0034295875,0.0034295875,0.017147938,0.037725464,0.07545093,0.08573969,0.08573969,0.08573969,0.072021335,0.1371835,0.26407823,0.38754338,0.45956472,0.45613512,0.53158605,0.89169276,1.1832076,1.2037852,0.90198153,0.5624523,0.33952916,0.216064,0.16462019,0.12346515,0.106317215,0.07545093,0.048014224,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.06859175,0.08573969,0.044584636,0.010288762,0.034295876,0.058302987,0.082310095,0.106317215,0.116605975,0.16462019,0.09259886,0.030866288,0.034295876,0.06859175,0.072021335,0.1097468,0.12003556,0.11317638,0.1371835,0.26064864,0.28465575,0.3566771,0.44927597,0.39097297,0.31552204,0.16804978,0.14061308,0.19548649,0.09602845,0.05144381,0.044584636,0.072021335,0.09945804,0.048014224,0.020577524,0.01371835,0.006859175,0.0034295875,0.01371835,0.01371835,0.030866288,0.06859175,0.11317638,0.1371835,0.22635277,0.22978236,0.26064864,0.32581082,0.31895164,0.33609957,0.3806842,0.45270553,0.5212973,0.5212973,0.51100856,0.7339317,0.939707,1.0563129,1.1934965,1.0254467,0.8505377,0.8848336,1.0288762,0.8711152,1.0151579,1.0220171,1.0700313,1.2586586,1.605047,2.644212,3.234101,3.5359046,3.8788633,4.7602673,5.24041,5.5387836,6.0737996,6.694555,6.697984,6.694555,6.81802,7.682276,8.680285,7.9909387,9.074688,9.578837,9.983529,10.635151,11.7257595,11.694893,11.934964,12.205902,12.370522,12.356804,13.598314,13.886399,14.733508,16.026463,16.002455,18.54035,20.62897,19.661825,16.513464,15.556609,13.320518,12.133881,10.933525,9.55826,8.772884,9.760606,9.949233,10.117283,10.88551,12.744347,14.150477,15.697222,17.014183,18.262554,20.100813,22.463799,24.332924,26.174612,28.18435,30.303835,30.612497,31.905453,34.817173,38.716614,41.707214,45.38716,47.71242,50.78533,55.36726,60.885468,72.15852,83.740234,88.64455,88.14383,91.79291,95.47971,98.09306,101.41633,105.53184,108.834526,85.83914,68.87984,57.397575,49.81476,43.535183,31.60022,26.466127,22.669573,18.670673,16.87014,12.185325,9.465661,7.8091707,6.1801167,3.3987212,2.5001693,1.7765263,1.3203912,1.1420527,1.1694894,0.90884066,0.881404,0.9945804,1.2483698,1.7182233,2.2841053,3.083199,3.5118976,3.1860867,1.9171394,1.6804979,1.8691251,1.5673214,0.7579388,0.32581082,0.17147937,0.13375391,0.09259886,0.030866288,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0274367,0.048014224,0.06859175,0.07888051,0.15090185,0.3018037,0.5178677,0.939707,1.8245405,2.5001693,1.8965619,1.2998136,1.2449403,1.529596,0.91227025,1.1832076,1.704505,2.294394,3.2203827,3.765687,4.9831905,6.121814,6.5470824,5.717122,7.8023114,9.132992,9.832627,9.517105,7.3084507,5.5079174,5.501058,4.7602673,2.819121,1.2655178,0.9602845,0.53844523,0.20920484,0.058302987,0.05144381,0.06516216,0.38754338,1.2826657,2.1915064,1.6976458,0.9774324,0.40126175,0.082310095,0.0,0.0,0.0,0.006859175,0.32924038,0.84367853,0.9877212,0.61046654,0.8779744,1.0082988,0.8676856,0.9568549,1.0151579,0.83338976,0.6927767,0.6859175,0.7339317,1.1523414,1.0220171,0.89855194,0.939707,0.90198153,1.0048691,0.9259886,0.72364295,0.64819205,1.1660597,1.1008976,1.1454822,1.2072148,1.1489118,0.805953,1.0117283,0.58645946,0.65162164,1.2449403,1.3066728,1.4027013,1.3306799,1.0700313,0.8093826,0.96714365,0.922559,1.1180456,1.2689474,1.3958421,1.7971039,1.5364552,1.3786942,1.371835,1.4438564,1.3958421,1.4541451,1.4027013,1.8999915,2.760818,2.9494452,4.40702,5.5593615,6.615674,7.7028537,8.872343,10.230459,11.266195,11.619442,11.585147,12.144169,11.201033,10.22703,9.633711,9.290752,8.532814,10.299051,10.439664,10.864933,11.718901,11.382801,12.199042,13.327377,14.013294,14.46257,15.837835,15.584045,15.8138275,16.39,16.80498,16.187653,16.828985,16.153357,16.568336,18.30028,19.408035,18.056778,16.084764,14.500296,13.958421,14.781522,13.718349,13.88297,13.7526455,13.574307,15.354263,16.554619,16.228807,15.981877,16.540901,17.761833,16.441442,15.666355,15.206791,15.141628,15.834405,16.520323,14.239647,15.937293,18.37916,8.1384115,8.865483,9.253027,8.536243,7.548522,8.738589,6.7665763,6.2967224,5.9400454,6.2384195,9.644,12.404818,12.3533745,14.390549,19.150816,23.01596,19.8676,15.316538,10.604284,7.932636,10.436234,12.315649,14.788382,12.048141,6.0532217,6.5230756,6.6568294,4.479041,3.3541365,3.8720043,3.8137012,3.99204,4.2595477,4.2835546,4.098357,4.1120753,4.0229063,3.8685746,3.4810312,2.9940298,2.8637056,2.3389788,2.2258022,2.253239,2.2738166,2.2566686,2.1400626,2.1263442,2.07833,1.9823016,1.9171394,1.7422304,1.8039631,1.8725548,1.8416885,1.7456601,1.7662375,1.903421,1.9514352,1.8519772,1.6907866,1.7696671,1.920569,2.054323,2.1503513,2.2292318,2.3286898,2.5756202,2.6304936,2.534465,2.702515,2.942586,3.2032347,3.6559403,4.149801,4.197815,3.8171308,3.9714622,4.1360826,4.2286816,4.5853586,4.791134,5.394741,5.967482,6.4236174,7.023795,7.0306544,6.667118,6.5230756,6.701414,6.8283086,7.3221693,7.2878733,6.632822,5.8200097,5.857735,5.874883,6.4373355,7.332458,8.14527,8.258447,8.083538,8.14527,7.9463544,7.490219,7.2707253,7.016936,7.0718093,7.864044,9.191295,10.22703,10.882081,11.372512,11.413667,10.786053,9.352485,10.377932,10.100135,9.445084,9.383351,10.930096,11.417097,11.859513,12.061859,11.794352,10.796341,10.405369,10.868362,10.912948,10.240748,9.513676,7.284444,5.7822843,4.99005,5.007198,6.0566516,5.3261495,5.305572,5.4016004,5.295283,4.928317,5.504488,5.9880595,7.421627,9.421077,10.203023,10.576848,10.100135,9.918367,10.669447,12.4802685,12.926115,13.917266,14.63062,14.682064,14.112752,14.277372,14.5585985,16.506605,19.312008,19.792149,18.145947,17.69667,18.639809,20.27572,21.03709,21.582394,22.44665,22.470657,21.77445,21.77445,22.882208,23.067406,22.299177,20.899906,19.53493,16.434584,16.084764,17.528622,19.761284,21.750444,23.502962,23.893936,23.612709,23.201159,23.050257,20.382038,19.294859,18.886738,18.650097,18.482046,19.11995,18.427174,17.761833,17.851004,18.787281,19.277712,20.018501,21.078245,22.213438,22.892496,0.69963586,0.8128122,0.77165717,0.77851635,0.8676856,0.90198153,0.8196714,0.9602845,1.1454822,1.371835,1.8279701,2.1880767,2.0886188,1.8725548,1.7250825,1.6599203,2.0508933,1.8965619,1.6290541,1.4747226,1.4541451,1.3958421,1.6976458,1.6530612,1.3203912,1.5261664,1.8142518,2.0920484,2.3835633,2.5207467,2.1469216,2.311542,2.194936,2.3389788,3.3061223,5.686256,6.615674,7.9600725,12.428825,18.176813,18.79414,11.177026,5.967482,2.952875,1.5536032,0.82996017,0.6893471,0.48014224,0.3806842,0.38754338,0.32581082,0.32581082,0.32924038,0.31895164,0.29494452,0.31552204,0.35324752,0.26750782,0.2194936,0.22292319,0.14747226,0.17833854,0.16462019,0.16804978,0.1920569,0.17147937,0.2709374,0.32581082,0.33609957,0.32581082,0.31895164,0.37039545,0.42183927,0.4424168,0.41498008,0.32924038,0.36353627,0.33609957,0.33266997,0.3806842,0.45613512,0.5212973,0.58302987,0.66533995,0.8745448,1.4232788,1.7662375,1.1660597,0.5007198,0.16462019,0.06516216,0.024007112,0.006859175,0.010288762,0.030866288,0.0548734,0.09602845,0.13032432,0.15090185,0.15090185,0.10288762,0.10288762,0.20577525,0.32924038,0.42526886,0.48357183,0.53158605,0.6276145,0.66876954,0.6036074,0.44927597,0.35324752,0.28465575,0.23321195,0.18862732,0.16119061,0.16804978,0.16119061,0.14747226,0.12346515,0.09259886,0.061732575,0.037725464,0.020577524,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0274367,0.030866288,0.010288762,0.0,0.01371835,0.006859175,0.006859175,0.020577524,0.030866288,0.058302987,0.034295876,0.010288762,0.006859175,0.017147938,0.017147938,0.048014224,0.061732575,0.058302987,0.07545093,0.15433143,0.18519773,0.24007112,0.29837412,0.23321195,0.22292319,0.1097468,0.07888051,0.13375391,0.06859175,0.024007112,0.01371835,0.0274367,0.041155048,0.017147938,0.006859175,0.006859175,0.006859175,0.010288762,0.01371835,0.044584636,0.06516216,0.09259886,0.15433143,0.26407823,0.28122616,0.274367,0.2709374,0.274367,0.26407823,0.36353627,0.42526886,0.432128,0.4629943,0.6962063,0.64133286,0.66876954,0.7579388,0.8779744,0.9842916,0.8471081,0.8128122,0.9431366,1.1043272,0.9534253,1.039165,1.1763484,1.3821237,1.7456601,2.4315774,3.2855449,3.6216443,3.8617156,4.2081037,4.623084,5.2644167,5.5833683,5.8165803,6.025785,6.111525,6.169828,6.5059276,7.1129646,7.6274023,7.3427467,8.412778,9.304471,9.712592,9.97324,11.05356,11.914387,12.21619,12.535142,13.111313,13.831526,14.994157,15.752095,16.702091,17.494326,16.87014,18.900457,20.546658,19.390888,16.12935,14.55174,13.203912,12.367092,11.218181,9.9869585,9.935514,10.333347,10.278474,10.851214,12.147599,13.310229,14.5243025,16.12249,17.765263,19.270851,20.642687,23.009102,24.343212,25.8488,27.642475,28.76052,30.029469,31.67567,34.028366,36.68287,38.49369,43.23338,45.514053,48.87162,54.85968,63.059826,75.464645,86.10665,92.14616,94.27936,96.75209,97.7501,99.41345,102.263435,104.468666,101.87247,77.94766,64.983826,56.36527,48.518375,40.89783,28.945719,24.655304,21.356041,17.168514,15.0250225,11.399949,9.218731,8.128122,6.944915,3.683377,3.4295874,2.5721905,2.020027,1.961724,1.8965619,1.5055889,1.3958421,1.4507155,1.6633499,2.1503513,2.4144297,3.0146074,3.450165,3.4192986,2.836269,3.3438478,2.6647894,1.5090185,0.50757897,0.18519773,0.09602845,0.058302987,0.034295876,0.017147938,0.0274367,0.0274367,0.017147938,0.010288762,0.006859175,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.0274367,0.08573969,0.17147937,0.28808534,0.4389872,0.5007198,0.97400284,1.4507155,1.762808,1.9823016,2.386993,2.061182,1.8416885,2.0028791,2.2566686,1.3341095,1.2243627,1.5673214,2.1812177,3.0866287,3.899441,4.3761535,5.312431,6.2247014,5.360445,7.274155,9.544542,9.081548,6.4098988,5.672538,5.2609873,4.4516044,3.0146074,1.3581166,0.51100856,0.34638834,0.16804978,0.05144381,0.037725464,0.13375391,0.06859175,0.8265306,1.2346514,1.3443983,2.417859,1.4918705,0.53844523,0.034295876,0.0,0.0,0.0,0.037725464,0.31552204,0.7579388,1.0117283,1.0288762,1.1694894,1.0700313,0.864256,1.1900668,0.7476501,0.864256,0.89169276,0.69963586,0.65505123,0.9842916,1.138623,1.1763484,1.1420527,1.0871792,1.1660597,1.3478279,1.1866373,0.8676856,1.2072148,1.1317638,1.1146159,0.96714365,0.7407909,0.71678376,0.9431366,0.9362774,1.0597426,1.3512574,1.5330256,1.546744,1.4850113,1.3684053,1.1866373,0.89512235,0.90198153,1.0768905,1.3101025,1.6530612,2.3218307,1.7456601,1.5844694,1.4438564,1.2860953,1.4267083,1.6221949,1.8005334,2.095478,2.3561265,2.1469216,3.532475,4.8151407,6.0703697,7.160979,7.73372,8.1212635,9.541112,10.820349,11.159878,10.14129,9.410788,9.112414,8.879202,8.680285,8.793462,10.569988,10.6317215,10.47396,10.6488695,10.768905,11.616013,12.329367,12.744347,13.351384,15.285671,15.254805,15.930434,16.434584,16.12249,14.589465,15.275383,15.940722,17.237106,18.516342,17.837284,16.187653,14.46257,13.265644,12.960411,13.680624,12.812939,12.679185,12.38424,12.202472,13.567448,14.359683,14.30481,14.318527,14.579176,14.503725,14.153908,13.88297,13.886399,14.538021,16.383139,15.9921665,14.1299,15.721229,18.104792,11.046701,10.930096,10.000677,8.553391,7.455923,8.131552,8.669997,8.958082,8.453933,7.514226,7.39762,9.637141,15.169065,24.343212,31.061773,22.77589,16.115631,13.029003,14.7369375,20.320305,26.689049,13.258785,10.333347,8.862054,6.0395036,5.295283,5.137522,3.99204,3.216953,3.2272418,3.5153272,4.0023284,4.046913,4.098357,4.190956,3.9783216,3.6559403,3.3438478,2.935727,2.510458,2.335549,2.2360911,2.0989075,1.9342873,1.8176813,1.8725548,1.762808,1.7971039,1.8142518,1.7971039,1.8656956,1.7902447,1.786815,1.762808,1.6907866,1.6187652,1.6942163,1.845118,1.862266,1.7388009,1.6496316,1.7113642,1.8485477,1.9994495,2.1434922,2.2841053,2.2498093,2.3149714,2.435007,2.620205,2.942586,3.1723683,3.1586502,3.069481,3.000889,2.9803114,2.7333813,3.0283258,3.3026927,3.415869,3.6353626,4.064061,4.6436615,5.2575574,5.8817425,6.5985265,6.4373355,6.3378778,6.5127864,6.9037595,7.1712675,7.630832,7.5450926,7.14726,6.835168,7.160979,6.8728933,7.2535777,7.8091707,8.1212635,7.8503256,7.3255987,7.407909,7.56224,7.6205435,7.747438,7.3050213,7.380472,8.035523,9.002667,9.674867,9.983529,10.525404,10.714031,10.268185,9.23245,9.73317,9.839486,9.904649,10.22703,11.087856,11.204462,11.698323,12.247057,12.205902,10.624862,10.103564,10.076128,9.6645775,8.748878,7.9909387,6.186976,4.928317,4.434457,4.698535,5.4907694,4.9180284,5.2918534,5.5833683,5.4736214,5.346727,5.267846,5.8062916,6.927767,8.371623,9.640571,9.613133,8.776315,8.745448,9.904649,11.406808,11.4754,12.891819,14.345964,14.928994,14.1299,14.325387,15.385129,17.29198,19.45262,20.697561,18.578075,18.11165,19.37374,21.558388,22.981665,22.44665,23.043398,23.492674,23.338343,22.957659,23.180582,23.087982,22.309467,20.94792,19.569225,18.310568,18.224829,19.095943,20.766151,23.122278,23.986534,23.719027,23.386356,23.11542,22.100262,20.251715,19.154245,18.386019,17.998474,18.499195,19.157675,18.46147,17.943602,18.04992,18.135658,18.173384,19.308577,20.851892,22.306036,23.372639,0.6756287,0.75450927,0.6893471,0.7305021,0.88826317,0.94656616,0.805953,0.9911508,1.2106444,1.4610043,2.037175,2.2052248,2.1091962,1.903421,1.6873571,1.4953002,1.8965619,1.7388009,1.587899,1.6084765,1.5638919,1.3615463,1.5261664,1.4541451,1.2243627,1.587899,1.8519772,2.2086544,2.4487255,2.3801336,1.8554068,2.0714707,2.1057668,2.3732746,3.4878905,6.252138,6.807731,8.735159,13.653188,18.838724,17.233677,8.433355,4.1772375,2.3252604,1.488441,1.039165,0.8162418,0.61389613,0.5658819,0.6036074,0.44927597,0.44584638,0.45270553,0.5007198,0.5418748,0.45613512,0.42183927,0.33609957,0.29837412,0.31895164,0.29837412,0.29151493,0.23664154,0.1920569,0.1920569,0.20920484,0.28465575,0.34295875,0.34295875,0.29494452,0.274367,0.26064864,0.3566771,0.40126175,0.3566771,0.30523327,0.34295875,0.36010668,0.39097297,0.4424168,0.5144381,0.53158605,0.5727411,0.64133286,0.78537554,1.0940384,1.3684053,0.94999576,0.4355576,0.13032432,0.034295876,0.01371835,0.0034295875,0.010288762,0.030866288,0.048014224,0.07888051,0.11317638,0.13032432,0.12003556,0.07888051,0.06516216,0.1371835,0.2469303,0.36696586,0.5007198,0.5041494,0.4629943,0.3841138,0.28808534,0.20577525,0.19548649,0.18862732,0.17833854,0.19548649,0.3018037,0.41498008,0.48700142,0.53158605,0.53844523,0.48357183,0.37039545,0.2469303,0.15433143,0.09945804,0.06859175,0.0274367,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.017147938,0.01371835,0.034295876,0.082310095,0.12689474,0.16804978,0.17490897,0.1097468,0.18519773,0.13375391,0.07545093,0.058302987,0.05144381,0.024007112,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.05144381,0.09602845,0.14061308,0.20577525,0.30866286,0.29151493,0.29494452,0.26750782,0.216064,0.216064,0.3841138,0.44927597,0.45956472,0.5041494,0.70306545,0.67219913,0.70306545,0.77851635,0.8471081,0.82996017,0.75450927,0.88826317,1.039165,1.0700313,0.91569984,0.97400284,1.2792361,1.5776103,1.9445761,2.7916842,3.3129816,3.765687,4.2595477,4.6676683,4.647091,5.086078,5.5079174,5.693115,5.6210938,5.470192,5.9160385,6.3035817,6.6396813,6.944915,7.2707253,8.213862,9.273604,9.794902,9.949233,10.748327,12.38767,13.169616,13.982429,15.196502,16.688372,17.991615,18.821575,19.414894,19.418324,17.902447,18.749556,20.124819,19.147387,16.04018,14.13676,13.22106,12.641459,11.701753,10.717461,11.012405,10.933525,10.9541025,11.72233,13.077017,14.016724,14.778092,16.084764,17.638369,19.099373,20.097382,22.014523,22.837624,24.000254,25.739054,27.11089,28.777668,30.605639,32.454185,34.179268,35.636845,40.338806,43.034462,47.307728,54.256073,62.493942,74.68955,84.05233,90.53082,94.70463,97.77411,96.20679,97.873566,100.62067,99.82157,88.40105,69.84012,59.880596,52.729908,45.013336,35.794605,25.841942,22.391777,19.325726,15.001016,12.253916,10.110424,8.779744,8.018375,7.1026754,4.8322887,4.5922174,3.4398763,3.0386145,3.474172,3.2443898,2.609916,2.7779658,3.1895163,3.4707425,3.433017,2.8225505,2.7573884,3.1277838,3.5393343,3.309552,3.5221863,2.2909644,0.97400284,0.23664154,0.06516216,0.030866288,0.020577524,0.017147938,0.030866288,0.06859175,0.06859175,0.041155048,0.020577524,0.01371835,0.0,0.024007112,0.05144381,0.058302987,0.048014224,0.058302987,0.07888051,0.11317638,0.23664154,0.4424168,0.64819205,0.84367853,1.5021594,2.061182,2.218943,1.9308578,2.1640697,2.2223728,2.3424082,2.585909,2.8156912,2.136633,1.9308578,2.1126258,2.620205,3.426158,4.0434837,4.4447455,5.5593615,6.9654922,6.8797526,7.332458,8.340756,7.082098,4.1463714,3.525616,4.4859004,3.357566,1.7525192,0.6276145,0.28808534,0.18519773,0.09945804,0.07888051,0.13375391,0.23321195,0.16119061,1.646202,1.728512,0.6241849,1.7216529,1.097468,0.37725464,0.024007112,0.08573969,0.18176813,0.12346515,0.22292319,0.432128,0.7579388,1.2346514,1.5261664,1.5707511,1.3752645,1.138623,1.2689474,0.823101,0.8196714,0.8471081,0.77165717,0.7476501,1.0220171,1.2209331,1.2620882,1.2209331,1.3478279,1.8759843,2.386993,2.1674993,1.4335675,1.3306799,1.3272504,1.2586586,0.9945804,0.6756287,0.7099246,0.939707,1.2380811,1.3752645,1.4129901,1.7216529,1.6153357,1.5330256,1.5158776,1.4507155,1.0666018,1.2517995,1.3341095,1.488441,1.7971039,2.2600982,1.7250825,1.7010754,1.6976458,1.6221949,1.786815,1.6256244,1.8313997,2.1126258,2.2669573,2.1743584,2.6922262,3.9063,5.295283,6.416758,6.9037595,6.759717,7.915488,9.362774,9.9801,8.56025,8.436785,8.303031,7.8537555,7.5382333,8.556821,9.966381,10.106995,9.709162,9.47938,10.086417,11.201033,11.753197,11.684605,11.869802,14.102464,14.860402,16.143068,16.798119,16.146498,13.992717,14.1299,15.1862135,16.46545,17.04162,15.755525,14.328816,13.519434,12.867812,12.329367,12.253916,11.797781,11.598865,11.578287,11.753197,12.212761,12.202472,12.6757555,13.399398,13.862392,13.2690735,13.344524,12.867812,12.737488,13.704632,16.386568,15.1862135,13.845244,14.287662,15.80011,15.0078745,12.6757555,10.655728,9.609704,9.537683,9.80519,12.343085,13.38911,14.860402,16.2974,14.860402,9.146709,14.140189,25.471546,33.963203,25.656744,16.729528,12.181894,16.695232,28.911423,41.449993,19.157675,8.597976,5.394741,5.446185,4.911169,3.7931237,3.3850029,3.0489032,2.7985435,3.3026927,4.0263357,3.9440255,3.9543142,4.1429415,3.7519686,3.2443898,2.760818,2.3904223,2.1400626,1.9754424,2.1469216,1.9754424,1.7593783,1.6496316,1.6599203,1.5604624,1.6221949,1.6427724,1.6290541,1.7799559,1.8142518,1.6976458,1.5433143,1.4369972,1.4404267,1.5673214,1.7388009,1.7765263,1.6907866,1.6839274,1.6907866,1.7833855,1.9480057,2.1469216,2.318401,2.1846473,2.0989075,2.1572106,2.3595562,2.6236343,2.8328393,2.7299516,2.4247184,2.1057668,2.0440342,2.0886188,2.335549,2.603057,2.8122618,3.0043187,3.5393343,4.0709205,4.523626,4.979761,5.693115,5.796003,6.23156,6.914048,7.56224,7.7028537,7.7851634,7.723431,7.699424,7.8434668,8.22758,7.8983397,8.06296,8.340756,8.464222,8.31332,7.6959944,7.6274023,7.891481,8.279024,8.591117,8.165848,8.460793,9.108984,9.6817255,9.705732,9.746887,9.551401,9.246168,9.0369625,9.218731,9.2153015,9.239308,9.626852,10.264755,10.593996,10.220171,10.367643,10.834066,10.960961,9.619993,9.544542,9.126132,8.193284,7.1712675,7.0786686,5.8680243,4.880303,4.588788,4.911169,5.2164025,4.887162,5.267846,5.686256,5.8645945,5.9126086,5.4496145,5.909179,6.4716315,7.1884155,8.958082,9.057541,8.443645,8.608265,9.633711,10.199594,10.556271,12.199042,14.061309,15.285671,15.21022,15.484588,17.55263,19.408035,20.433481,21.37319,19.414894,18.53692,19.288,21.36633,23.616138,22.9508,23.883648,24.888515,25.173172,24.679312,24.202599,23.760181,23.019392,21.973368,20.94792,19.987637,19.682402,20.176264,21.52066,23.647005,23.746464,22.933651,22.26831,21.880768,20.982216,20.189981,18.989626,17.88873,17.412016,18.097933,19.603521,19.421753,18.831865,18.45804,18.269413,17.923023,18.643238,19.973917,21.4555,22.628418,0.6859175,0.65162164,0.61389613,0.65162164,0.764798,0.90198153,0.91569984,1.08032,1.2072148,1.3786942,1.9823016,1.7353712,1.5501735,1.4507155,1.3649758,1.1351935,1.4438564,1.4781522,1.5741806,1.7079345,1.5193073,1.3203912,1.3855534,1.3306799,1.255229,1.728512,2.16064,2.5413244,2.5481834,2.177788,1.7388009,2.218943,2.2806756,2.7402403,4.0949273,6.543653,7.4696417,9.671436,13.828096,17.391438,14.592895,6.0154963,2.6167753,1.5810398,1.2483698,1.1214751,0.8779744,0.7442205,0.7442205,0.7888051,0.6927767,0.6962063,0.70649505,0.8265306,0.9602845,0.7922347,0.6790583,0.5796003,0.53501564,0.5453044,0.5658819,0.432128,0.32238123,0.26407823,0.2709374,0.32238123,0.31209245,0.29837412,0.28122616,0.26064864,0.24007112,0.19548649,0.26064864,0.31209245,0.30866286,0.28122616,0.25721905,0.33609957,0.41840968,0.48357183,0.61389613,0.5727411,0.5658819,0.59331864,0.65848076,0.7476501,0.7339317,0.548734,0.30523327,0.106317215,0.01371835,0.0034295875,0.01371835,0.0274367,0.030866288,0.030866288,0.05144381,0.06516216,0.058302987,0.037725464,0.0274367,0.024007112,0.07888051,0.18519773,0.32924038,0.48357183,0.42526886,0.39783216,0.32924038,0.22635277,0.19891608,0.1371835,0.106317215,0.12346515,0.23321195,0.51100856,0.7990939,1.0220171,1.1763484,1.2449403,1.2037852,0.9328478,0.66876954,0.45613512,0.3018037,0.18176813,0.07888051,0.024007112,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.01371835,0.05144381,0.106317215,0.14747226,0.15090185,0.12346515,0.19548649,0.18176813,0.106317215,0.037725464,0.072021335,0.06516216,0.024007112,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.09602845,0.16804978,0.22635277,0.23664154,0.25378948,0.26064864,0.23321195,0.19548649,0.22978236,0.40126175,0.4629943,0.5453044,0.6241849,0.5658819,0.65162164,0.8471081,0.9945804,1.0425946,1.0357354,0.90541106,1.0460242,1.0940384,0.9362774,0.7133542,0.8471081,1.2620882,1.5810398,1.8382589,2.486451,2.7711067,3.673088,4.547633,4.955754,4.7019644,4.870014,5.267846,5.6039457,5.693115,5.4633327,6.077229,6.3824625,6.574519,6.8797526,7.548522,8.519095,9.55826,10.347065,10.858074,11.365653,12.908967,14.483148,16.071047,17.754974,19.713268,21.081675,21.575535,21.77102,21.386908,19.281141,19.054789,20.299728,19.675543,16.921585,14.832966,13.756075,13.498857,12.953552,12.0138445,11.55428,11.63659,11.7257595,12.332796,13.478279,14.688923,15.367981,15.951012,16.698662,17.700102,18.8593,20.19684,20.917053,22.103691,23.931662,25.69104,26.812515,28.451859,30.163221,31.850578,33.74028,36.974384,40.58574,45.774704,52.335506,58.666523,68.86612,76.6307,82.60504,87.57452,92.46511,90.26674,91.734604,93.39452,89.59797,72.53235,60.737995,52.438393,45.942753,38.884663,28.19464,22.686722,19.744135,16.434584,12.487128,10.257896,9.174147,8.467651,7.8331776,7.0375133,5.909179,5.504488,4.2355404,4.32128,5.586798,5.435896,4.2252517,4.7534084,5.6656785,5.9297566,4.839148,3.3644254,2.551613,2.7470996,3.3815732,2.9391565,2.0920484,1.1420527,0.4389872,0.09945804,0.01371835,0.024007112,0.020577524,0.0274367,0.05144381,0.09602845,0.09259886,0.05144381,0.024007112,0.01371835,0.010288762,0.09602845,0.16119061,0.16119061,0.12346515,0.15433143,0.18519773,0.14747226,0.2503599,0.4972902,0.66533995,1.0768905,1.6907866,2.0680413,2.0749004,1.8965619,2.253239,2.301253,2.386993,2.6647894,3.069481,2.7711067,2.8225505,3.018037,3.2649672,3.5839188,4.1600895,5.06893,6.4304767,7.936065,8.841476,7.98408,6.6122446,5.3398676,4.0023284,1.6599203,3.1277838,2.4144297,1.1763484,0.36010668,0.18176813,0.12689474,0.15433143,0.2469303,0.32924038,0.2709374,0.6001778,2.0268862,1.7525192,0.0,0.0,0.0,0.21263443,0.30523327,0.29494452,0.53844523,0.61046654,0.66191036,0.805953,1.1351935,1.7113642,1.9823016,2.0131679,1.9514352,1.7525192,1.1489118,1.2929544,0.8711152,0.6310441,0.77508676,0.94999576,1.3203912,1.2620882,1.1489118,1.2072148,1.5364552,2.5653315,3.1723683,2.8328393,1.8999915,1.6084765,1.6633499,1.5741806,1.2895249,0.9945804,1.0940384,1.1900668,1.4987297,1.6256244,1.611906,1.9171394,1.7319417,1.5844694,1.546744,1.5741806,1.4953002,1.7593783,1.6633499,1.587899,1.6736387,1.821111,1.5741806,1.6667795,1.8931323,2.1160555,2.3081124,1.7696671,1.704505,1.978872,2.4658735,3.0214665,2.9151495,4.149801,5.435896,6.1904054,6.5299344,6.917478,7.514226,8.419638,9.132992,8.546532,8.762596,8.06296,7.1678376,6.842027,7.9017696,8.735159,9.129561,9.170717,9.177576,9.736599,10.5597,11.303921,11.252477,11.129011,13.097594,14.503725,16.098484,16.986746,16.486027,14.13676,13.96871,14.2533655,14.757515,14.839825,13.454271,12.579727,12.792361,12.723769,11.97269,11.084427,11.05699,11.283342,11.616013,11.7257595,11.111863,10.796341,11.523414,12.572867,13.457702,13.917266,13.756075,12.593445,11.924676,12.648318,15.073037,13.975569,12.764925,12.908967,14.55174,16.503176,13.231348,11.005547,10.593996,11.626302,12.617453,15.059319,15.371411,19.497204,27.296087,32.539925,14.164196,11.598865,16.87357,24.223177,30.084341,27.35096,18.567787,17.007324,26.555296,41.700356,26.058006,10.882081,3.3061223,3.649081,5.4153185,3.5530527,3.1655092,3.0969174,2.9974594,3.333559,4.081209,4.040054,4.0091877,4.033195,3.4227283,2.884283,2.2463799,1.8897027,1.8519772,1.8108221,1.8931323,1.7971039,1.7593783,1.7765263,1.6359133,1.5398848,1.605047,1.587899,1.4953002,1.5776103,1.7250825,1.5604624,1.3375391,1.2277923,1.3272504,1.4335675,1.6496316,1.7456601,1.7182233,1.7662375,1.786815,1.8656956,2.0303159,2.218943,2.2806756,2.1297739,1.9891608,1.8931323,1.8828435,2.0028791,2.1640697,2.0920484,1.9068506,1.728512,1.6907866,1.862266,2.0165975,2.287535,2.5961976,2.6819375,3.2066643,3.758828,4.0229063,4.139512,4.715683,5.3158607,6.1492505,7.1541195,7.970361,7.939495,7.8091707,7.9737906,8.258447,8.539673,8.735159,8.724871,8.621983,8.659708,8.889491,9.1810055,8.831187,8.656279,8.831187,9.242738,9.462232,9.054111,9.530824,10.206452,10.607714,10.491108,10.542552,9.671436,8.769455,8.539673,9.510246,9.239308,8.868914,9.129561,9.925226,10.31277,9.431366,9.047252,9.14328,9.3936405,9.139851,9.668007,9.5205345,8.508806,7.3084507,7.449064,6.4716315,5.6176643,5.2164025,5.2781353,5.4839106,5.377593,5.4324665,5.8234396,6.3824625,6.5813785,6.2658563,6.262427,6.1972647,6.560801,8.718011,9.318189,9.033533,9.129561,9.616563,9.23245,10.607714,12.048141,13.937843,16.04361,17.518333,17.665806,19.576086,20.917053,21.11597,21.325174,20.467777,19.45262,19.294859,20.522652,23.170294,23.44809,24.727325,25.756203,26.03057,25.804216,25.063425,24.730755,24.134007,23.314335,23.022821,21.074816,20.296299,20.762722,21.997374,22.974806,23.578413,23.142857,22.271742,21.469217,21.157125,20.827885,19.469769,18.217968,17.751545,18.30028,20.512363,20.474638,19.020493,17.53548,17.95732,17.765263,18.21111,19.178253,20.35803,21.263443,0.4424168,0.5521636,0.7442205,0.89855194,0.9534253,0.91569984,1.0734608,1.0117283,0.90198153,0.980862,1.5398848,1.529596,1.4335675,1.4953002,1.6496316,1.5261664,1.5501735,1.3546871,1.313532,1.4335675,1.371835,1.4575747,1.7079345,1.7833855,1.786815,2.287535,2.6922262,2.5447538,2.2155135,1.9102802,1.6770682,2.1194851,2.2738166,3.2683969,5.2609873,7.4456344,8.508806,10.247607,13.745787,16.571766,12.785502,5.1100855,2.411,1.5673214,1.0117283,0.7339317,0.6241849,0.5041494,0.5041494,0.65505123,0.89855194,0.8745448,0.83338976,0.8505377,0.89169276,0.7922347,0.85396725,1.0700313,1.2415106,1.2243627,0.9294182,0.5658819,0.5178677,0.432128,0.26407823,0.274367,0.26407823,0.2503599,0.23664154,0.20577525,0.106317215,0.18176813,0.23664154,0.22978236,0.2194936,0.36696586,0.30523327,0.30866286,0.38754338,0.5418748,0.7476501,0.6001778,0.52815646,0.5761707,0.6859175,0.6859175,0.42869842,0.2469303,0.11317638,0.024007112,0.0,0.0,0.072021335,0.1097468,0.07888051,0.030866288,0.030866288,0.041155048,0.058302987,0.07545093,0.07545093,0.06516216,0.116605975,0.21263443,0.31209245,0.33609957,0.28808534,0.32924038,0.29837412,0.18519773,0.1371835,0.12346515,0.12346515,0.15776102,0.28122616,0.548734,1.0014396,1.4815818,1.8108221,1.9720128,2.1057668,1.5810398,1.2380811,0.9328478,0.61046654,0.30523327,0.13375391,0.044584636,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.010288762,0.034295876,0.061732575,0.061732575,0.037725464,0.01371835,0.01371835,0.048014224,0.12346515,0.12346515,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.034295876,0.08916927,0.16119061,0.19891608,0.2469303,0.23321195,0.18862732,0.1920569,0.34981793,0.42526886,0.48014224,0.53501564,0.5761707,0.5658819,0.85739684,0.91227025,0.94999576,1.0700313,1.2655178,1.155771,1.0014396,0.922559,0.90884066,0.823101,1.0563129,1.2586586,1.6256244,2.095478,2.3664153,2.4624438,3.2478194,4.040054,4.496189,4.5922174,5.521636,5.377593,5.4941993,6.108095,6.3790326,6.3310184,6.893471,6.924337,6.6568294,7.706283,9.047252,10.401938,11.701753,12.682614,12.878101,13.231348,15.29939,17.569777,19.44576,21.239435,22.36434,22.717587,22.741594,22.552967,21.942501,21.503513,20.851892,20.303158,19.239986,16.12935,15.87213,15.7795315,15.230798,14.116182,12.847235,12.188754,12.21619,13.077017,14.273943,14.664916,15.127911,15.443433,16.335125,17.87158,19.469769,20.347742,22.172283,24.576424,25.982555,23.588703,24.418663,25.697899,27.357819,29.213226,30.945168,34.16898,38.442245,43.199085,48.988228,57.493603,63.073544,68.38597,73.8253,78.75705,81.52815,82.10089,79.7482,74.76157,67.03815,56.077183,48.912777,43.099625,37.955246,32.224403,24.092852,21.897917,18.015623,13.978998,11.2593355,11.245617,10.7586155,10.652299,9.73317,7.798882,5.675967,6.0532217,5.353586,6.135532,8.193284,8.56025,6.0703697,6.135532,6.6396813,6.1458206,3.875434,3.0454736,2.435007,2.277246,2.3149714,1.8142518,1.0940384,0.6310441,0.33952916,0.16119061,0.07545093,0.06516216,0.041155048,0.048014224,0.06859175,0.044584636,0.034295876,0.020577524,0.01371835,0.020577524,0.044584636,0.22978236,0.34638834,0.32238123,0.22978236,0.29151493,0.38754338,0.32924038,0.39097297,0.6276145,0.8848336,1.1900668,1.6976458,1.7696671,1.4061309,1.2346514,1.9548649,1.8073926,1.7593783,2.1434922,2.6545007,2.6304936,3.2478194,3.758828,3.789694,3.3266997,6.0737996,6.0635104,6.135532,7.3393173,8.927217,7.425057,5.7582774,5.576509,5.6142344,1.7079345,1.8691251,1.155771,0.4664239,0.15776102,0.061732575,0.072021335,0.31552204,0.53501564,0.5658819,0.31895164,1.8691251,1.3512574,0.44927597,0.0,0.0,0.0,1.0631721,1.2826657,0.61389613,0.8711152,1.8108221,1.4781522,1.2998136,1.6016173,1.6016173,2.3218307,2.4212887,2.633923,2.6887965,1.2963841,1.1249046,1.0666018,0.8505377,0.53501564,0.47328308,0.764798,1.0768905,1.3581166,1.5364552,1.5261664,1.8313997,1.5673214,1.4781522,1.7902447,2.2429502,1.7319417,2.0063086,1.8348293,1.3649758,2.1194851,1.2792361,1.7559488,2.1263442,1.978872,1.8931323,1.903421,1.8245405,1.7593783,1.728512,1.6770682,1.6290541,1.3889829,1.2792361,1.4678634,1.9685832,1.845118,1.978872,1.9994495,1.9274281,2.1983654,2.5893385,2.6956558,2.6407824,2.668219,3.1449318,4.0229063,5.761707,6.800872,6.800872,6.6533995,7.4696417,8.443645,9.571979,10.244178,9.23245,8.40249,7.3255987,6.848886,7.191845,7.949784,8.207003,8.920357,9.530824,9.832627,9.9801,9.465661,10.014396,10.882081,11.952112,13.732068,13.670336,15.37827,16.55119,16.064188,13.975569,14.417986,14.507155,15.361122,16.12935,13.992717,12.747777,12.418536,12.47341,12.367092,11.537132,11.646879,12.037852,11.787492,10.868362,10.1481495,11.159878,11.670886,11.766914,12.010415,13.426835,13.255356,12.325937,12.277924,13.094165,13.107883,13.193623,12.627741,12.346515,12.758065,13.732068,10.755186,9.523964,10.38479,12.168177,12.1921835,13.9481325,10.323058,12.027563,24.106571,45.942753,19.500635,10.652299,9.798331,16.657507,40.253067,51.55356,34.99208,19.493774,16.61292,20.508932,23.743034,12.9809885,3.5187566,1.4987297,3.8925817,3.3061223,3.4878905,3.6593697,3.5873485,3.6010668,4.1155047,3.9474552,3.8891523,3.875434,3.0214665,2.568761,1.9891608,1.605047,1.529596,1.6633499,1.5913286,1.6530612,1.6976458,1.6736387,1.6496316,1.5124481,1.4438564,1.3821237,1.3341095,1.3581166,1.6016173,1.471293,1.2826657,1.2312219,1.3889829,1.5364552,1.5913286,1.5913286,1.6324836,1.8759843,1.9239986,1.937717,2.1023371,2.3046827,2.1194851,2.0474637,1.8176813,1.6839274,1.7696671,2.0749004,1.9651536,1.8828435,1.9239986,2.020027,1.9239986,1.7525192,1.9480057,2.311542,2.5619018,2.3046827,2.6716487,3.199805,3.590778,3.7862647,3.981751,4.9351764,5.813151,6.6636887,7.414768,7.905199,7.5862474,7.4696417,7.7748747,8.416207,9.002667,9.3936405,8.913498,8.443645,8.433355,8.9100685,9.362774,9.47595,9.846346,10.401938,10.39165,9.513676,9.925226,10.710602,11.334786,11.626302,10.9541025,10.72432,10.333347,9.630281,8.9100685,8.385342,8.759167,9.753747,10.923236,11.64345,11.252477,11.015835,10.943813,11.091286,11.581717,10.703742,11.509696,11.653738,10.316199,8.193284,6.327589,5.6039457,5.23698,5.178677,6.118384,6.6053853,6.7391396,6.9209075,7.31531,7.8263187,7.658269,7.267296,6.742569,6.9620624,9.599416,9.767465,9.132992,9.297611,10.086417,9.537683,11.537132,12.644889,14.181344,16.540901,19.164536,19.812727,19.771572,19.997925,20.752434,21.606401,21.959648,22.213438,22.158566,22.230585,23.513252,24.891945,25.35837,25.471546,25.447538,25.132017,24.655304,24.672453,24.082563,23.118849,23.376068,22.144846,21.249723,21.548098,22.398636,21.668133,24.010542,25.073713,24.830214,23.612709,22.11055,22.02481,20.721567,19.390888,18.910746,19.850452,21.047379,20.330595,18.406595,16.822126,17.943602,17.322845,18.547209,19.744135,20.423193,21.482935,0.6756287,0.6276145,0.72364295,0.8265306,0.85739684,0.78194594,0.90198153,0.78537554,0.7682276,0.9568549,1.2346514,1.3306799,1.4472859,1.4781522,1.4472859,1.5021594,1.5536032,1.3958421,1.4335675,1.6530612,1.6290541,1.4610043,1.5673214,1.7182233,2.0303159,2.959734,2.4075704,1.9823016,1.762808,1.6770682,1.5433143,1.6804979,2.1503513,3.9200184,6.608815,8.471081,8.7317295,11.430815,16.204802,19.161106,12.847235,5.960623,3.2032347,2.0646117,1.3855534,1.3684053,1.4027013,1.1832076,0.91912943,0.7305021,0.6310441,0.5693115,0.5453044,0.5693115,0.59674823,0.548734,0.805953,0.7133542,0.6790583,0.7922347,0.8196714,0.42526886,0.34981793,0.34295875,0.33609957,0.44584638,0.4424168,0.3806842,0.32238123,0.2777966,0.22978236,0.3018037,0.2777966,0.28122616,0.33952916,0.37725464,0.36696586,0.3806842,0.40126175,0.45613512,0.6241849,0.5658819,0.4938606,0.4938606,0.5521636,0.5521636,0.33609957,0.18519773,0.08916927,0.034295876,0.0,0.0,0.01371835,0.020577524,0.017147938,0.006859175,0.024007112,0.0548734,0.06859175,0.06516216,0.07545093,0.13375391,0.18519773,0.20577525,0.19891608,0.21263443,0.23321195,0.20577525,0.14404267,0.07888051,0.041155048,0.106317215,0.17490897,0.28465575,0.40126175,0.41498008,0.65162164,1.1008976,1.6084765,2.0165975,2.1434922,1.7936742,1.546744,1.1694894,0.66876954,0.30523327,0.12346515,0.034295876,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0034295875,0.01371835,0.0034295875,0.0034295875,0.006859175,0.01371835,0.01371835,0.006859175,0.0034295875,0.006859175,0.020577524,0.024007112,0.072021335,0.15090185,0.15776102,0.07888051,0.01371835,0.0034295875,0.006859175,0.017147938,0.020577524,0.01371835,0.044584636,0.13032432,0.18519773,0.17833854,0.1371835,0.18519773,0.28122616,0.32581082,0.31895164,0.34981793,0.3841138,0.39440256,0.4938606,0.58988905,0.39440256,0.75450927,0.96714365,1.1111864,1.2312219,1.3409687,1.1626302,1.1420527,1.3032433,1.4232788,1.0563129,1.0425946,1.0631721,1.471293,2.0714707,2.095478,2.136633,2.253239,2.7093742,3.4878905,4.2869844,4.863155,5.7102633,6.3618846,6.4579134,5.7308407,6.0052075,6.6876955,7.2878733,8.018375,9.781183,10.967821,12.185325,12.977559,13.450842,14.270514,15.786391,18.025911,19.764713,20.968498,22.803328,23.163433,23.10856,23.245745,23.35549,22.395206,22.18943,22.847912,24.082563,24.219748,20.231136,20.45063,19.380598,17.717249,15.834405,13.776653,13.954991,14.054449,14.270514,14.678635,15.223939,15.981877,17.103354,18.30028,19.167965,19.21255,19.497204,22.131128,24.332924,25.368658,26.521,24.216316,22.5221,22.847912,25.35837,28.956007,35.293884,41.30595,48.97108,56.6122,58.910023,62.41849,65.604576,69.781815,73.44462,72.25112,73.653824,71.18452,64.73347,56.132057,49.14256,41.792953,37.23846,33.373314,28.678211,22.237446,19.980776,16.846134,14.908417,13.663476,10.038403,8.680285,9.369633,9.31133,7.9086285,6.7631464,7.239859,6.8385973,7.0306544,7.716572,7.2535777,6.677407,6.200694,5.411889,4.0880685,2.2292318,2.1400626,1.9582944,1.8485477,1.6976458,1.1214751,0.7613684,0.6276145,0.6036074,0.5727411,0.42869842,0.41840968,0.39783216,0.3841138,0.36010668,0.2777966,0.16804978,0.12346515,0.15776102,0.19891608,0.106317215,0.2503599,0.490431,1.0494537,1.546744,1.0220171,0.89512235,0.7579388,0.6927767,0.7682276,1.0425946,1.2792361,1.5433143,1.4953002,1.255229,1.4061309,1.5501735,1.6221949,1.5398848,1.4918705,1.9480057,1.8554068,2.5996273,3.316411,3.7039545,4.0091877,6.6876955,5.8337283,5.994919,8.06296,9.266746,9.290752,7.4113383,5.192395,3.5942078,2.976882,2.4041407,1.2175035,0.36696586,0.11317638,0.024007112,0.0274367,0.06859175,0.19548649,0.28808534,0.06516216,0.39440256,0.30866286,0.2469303,0.25378948,0.0,0.020577524,0.5144381,0.8093826,0.86082643,1.2723769,1.430138,1.5844694,1.5776103,1.6633499,2.49331,2.2258022,2.4007113,2.7745364,2.6990852,1.1146159,1.9480057,1.670209,1.4267083,1.5090185,1.3512574,1.2723769,1.5364552,1.670209,1.587899,1.587899,1.9411465,1.529596,1.6564908,2.253239,1.8656956,1.5261664,2.2258022,2.1434922,1.3272504,1.6942163,1.9171394,2.3081124,2.3972816,2.1503513,1.978872,1.6667795,1.670209,1.5193073,1.1866373,1.0666018,2.1915064,2.644212,2.2978237,1.6324836,1.7730967,2.0406046,2.74367,3.525616,3.7931237,2.6853669,2.527606,2.4041407,2.5138876,3.117495,4.523626,4.3452873,4.8185706,5.4084597,6.0052075,6.9346256,7.6445503,8.423067,8.858624,8.769455,8.207003,7.795452,7.006647,6.848886,7.1884155,6.7528577,8.378482,8.694004,8.381912,8.48137,10.405369,11.115293,11.293632,11.619442,12.360233,13.392539,13.7697935,14.88098,15.254805,14.898128,15.319967,16.023033,16.266533,16.588915,16.815268,16.0539,14.027013,12.843805,12.133881,11.770344,11.876661,11.489118,11.640019,11.63659,11.129011,10.134431,10.573419,10.9369545,11.074138,11.30049,12.401388,12.212761,11.921246,12.531713,13.478279,12.63117,14.153908,13.13189,11.670886,11.201033,12.500846,11.406808,10.875222,13.272504,17.014183,16.54776,12.291641,10.738038,24.720467,51.093994,70.735245,25.876238,17.233677,17.700102,22.62156,49.7736,55.13062,42.273094,27.008001,16.750105,10.497967,10.278474,12.723769,9.825768,2.9254382,2.719663,3.4707425,3.5702004,3.415869,3.5187566,4.5167665,4.180667,3.7725463,3.707384,3.683377,2.6922262,2.4727325,2.0714707,1.7216529,1.6016173,1.8348293,1.6427724,1.6187652,1.5501735,1.4472859,1.5501735,1.6221949,1.529596,1.3649758,1.2929544,1.5536032,1.4541451,1.2037852,1.1729189,1.371835,1.4129901,1.704505,1.7902447,1.6599203,1.4815818,1.6084765,1.7662375,2.0303159,2.0920484,1.920569,1.7662375,1.7422304,1.6359133,1.5810398,1.6564908,1.903421,2.352697,2.2841053,2.1297739,2.0508933,1.9342873,1.6084765,1.7490896,2.1023371,2.3732746,2.2566686,2.6304936,3.4124396,4.190956,4.6265135,4.4721823,4.602506,5.336438,6.042933,6.667118,7.720001,7.2878733,6.9346256,7.3290286,8.344186,9.074688,8.635701,8.05953,8.141841,8.899779,9.571979,10.772334,10.556271,10.151579,10.31277,11.30735,11.773774,11.952112,12.247057,12.507706,12.017275,10.9369545,10.947243,10.477389,9.256456,8.31332,7.3873315,7.579388,8.56025,9.870353,10.923236,11.653738,12.185325,12.706621,13.368532,14.267084,12.929544,12.5145645,11.907528,10.6145735,8.755736,7.7851634,7.6376915,7.4627824,7.058091,6.8763227,6.1629686,6.3824625,6.866034,7.56224,9.012956,8.656279,8.035523,7.613684,7.8331776,9.122703,10.151579,9.798331,9.938945,10.792912,10.926665,12.05157,13.368532,15.409137,17.528622,17.909306,18.907316,18.677534,18.163095,18.12194,19.102802,20.395756,21.836184,22.679861,23.060547,23.989964,25.399525,25.752771,25.159454,24.404943,24.936531,26.167753,26.586163,25.979126,24.703318,23.681301,22.69358,21.897917,21.647556,21.795029,21.668133,23.297188,23.904224,23.44123,22.309467,21.352612,20.838173,20.385468,19.802439,19.802439,22.011093,21.558388,21.733295,21.421204,20.148827,18.077356,17.161655,18.03277,19.277712,20.244854,21.033659,0.6310441,0.6927767,0.7613684,0.8093826,0.8471081,0.9294182,1.0185875,0.97400284,0.91569984,0.89855194,0.89512235,1.0528834,1.2895249,1.3684053,1.3306799,1.4850113,1.3409687,1.2620882,1.4198492,1.6770682,1.5844694,1.5570327,1.7765263,2.194936,2.6373527,2.8259802,2.2360911,1.9411465,1.7456601,1.6256244,1.7216529,1.6873571,2.417859,4.3795834,6.914048,8.23444,8.697433,12.46998,16.969599,18.293419,11.2250395,5.4667625,2.9974594,1.8897027,1.214074,1.0494537,1.0494537,0.94999576,0.7888051,0.6893471,0.8676856,0.86082643,0.82996017,0.8128122,0.7682276,0.5693115,0.64819205,0.45270553,0.39097297,0.51100856,0.51100856,0.31895164,0.3018037,0.30866286,0.31209245,0.38754338,0.490431,0.4081209,0.31895164,0.28122616,0.26064864,0.35324752,0.3806842,0.42869842,0.52472687,0.61046654,0.5727411,0.48014224,0.4046913,0.4081209,0.53158605,0.53844523,0.4664239,0.42869842,0.42869842,0.36353627,0.23664154,0.13375391,0.072021335,0.037725464,0.010288762,0.017147938,0.006859175,0.0,0.0,0.0,0.010288762,0.034295876,0.05144381,0.061732575,0.10288762,0.1097468,0.17147937,0.19548649,0.18519773,0.20920484,0.23321195,0.18176813,0.11317638,0.0548734,0.024007112,0.116605975,0.17147937,0.26064864,0.37382504,0.42869842,0.61046654,0.939707,1.4267083,1.9102802,2.0680413,1.6907866,1.3409687,0.9431366,0.52815646,0.22292319,0.09945804,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06859175,0.08916927,0.044584636,0.037725464,0.030866288,0.044584636,0.061732575,0.072021335,0.06516216,0.041155048,0.024007112,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.044584636,0.044584636,0.048014224,0.106317215,0.13032432,0.116605975,0.13375391,0.09945804,0.07888051,0.058302987,0.044584636,0.061732575,0.11317638,0.15776102,0.16462019,0.15090185,0.18519773,0.21263443,0.28122616,0.30866286,0.3018037,0.36010668,0.39783216,0.44927597,0.53501564,0.58302987,0.4424168,0.7682276,0.8471081,0.89169276,0.97057325,1.0185875,1.0151579,1.1592005,1.2312219,1.1797781,1.1146159,1.3478279,1.3375391,1.5261664,1.845118,1.7010754,1.7696671,1.845118,2.2909644,3.0660512,3.7348208,4.15666,5.1409516,6.1286726,6.5813785,5.970912,6.2384195,6.7185616,7.486789,8.663138,10.429376,12.140739,13.437123,14.407697,15.199932,16.047039,17.339994,19.219408,20.889618,22.004232,22.652426,23.022821,23.26975,23.61957,23.921373,23.643576,22.806757,23.482386,25.255482,26.068295,22.216867,21.20514,20.111101,18.725548,17.175373,15.913286,15.700651,15.29253,15.117621,15.426285,16.300829,16.763824,17.38115,18.567787,19.768143,19.469769,20.814167,22.237446,23.60242,25.625877,29.871706,28.414133,25.982555,24.751333,26.572443,32.9892,43.291683,49.95537,55.13062,59.170673,60.621387,59.890884,62.93979,67.08616,69.55889,67.50457,70.1625,70.207085,63.625706,52.016552,42.56804,38.06156,35.012657,31.521338,26.665043,20.491785,17.730967,14.517444,12.106443,10.460241,8.251588,7.31531,7.932636,8.570539,8.790032,9.239308,9.287323,8.8929205,8.567109,8.244728,7.2947326,7.4010496,6.090947,4.3761535,2.8911421,1.879414,2.16064,2.1572106,1.9514352,1.6359133,1.3409687,1.0048691,0.8505377,0.7682276,0.6859175,0.6001778,0.6036074,0.58988905,0.5727411,0.52472687,0.39097297,0.30866286,0.274367,0.34981793,0.42526886,0.22292319,0.3566771,0.5144381,0.8162418,1.1146159,0.9774324,0.66876954,0.7133542,0.864256,0.99801,1.1111864,1.3443983,1.4747226,1.4747226,1.4335675,1.5330256,1.430138,1.5810398,1.6221949,1.5776103,1.8691251,1.8485477,2.510458,3.1552205,3.8137012,5.2506986,8.200144,8.419638,9.115844,10.55284,10.05898,9.23245,7.06838,5.079219,4.2698364,5.137522,3.1620796,1.3992717,0.37382504,0.08916927,0.024007112,0.048014224,0.2469303,0.31552204,0.18519773,0.010288762,0.010288762,0.020577524,0.09259886,0.18862732,0.16462019,0.36353627,0.7476501,1.039165,1.2620882,1.7216529,1.9274281,1.6839274,1.7388009,2.1400626,2.2498093,2.469303,2.4555845,2.620205,2.719663,1.845118,2.603057,2.5893385,2.393852,2.2223728,1.8931323,1.4781522,1.3958421,1.4747226,1.6016173,1.704505,1.6530612,1.5707511,1.8245405,2.2223728,2.0268862,1.6530612,1.8073926,2.0577524,2.3458378,2.9871707,2.2086544,2.469303,2.3595562,1.7833855,1.961724,1.5124481,1.4164196,1.4918705,1.5913286,1.5638919,2.335549,2.3767042,2.4555845,2.603057,2.1194851,2.3801336,3.018037,3.590778,3.6970954,2.952875,2.7985435,2.2292318,2.428148,3.7142432,5.5250654,5.6519604,6.495639,7.373613,7.7440085,7.233,8.083538,9.709162,9.932085,8.724871,8.179566,8.436785,7.720001,7.1129646,6.6739774,5.4187484,6.6396813,7.4696417,7.582818,7.750868,9.853205,10.604284,10.971251,11.105004,11.30735,12.024134,13.011855,13.526293,13.670336,13.680624,13.951562,14.538021,14.874121,14.856973,14.613472,14.520873,12.699762,11.499407,10.8958,10.854645,11.321068,11.218181,11.31078,11.588576,11.609154,10.487679,10.422516,10.4705305,10.731179,11.338216,12.466551,12.672326,13.121602,13.7526455,14.003006,12.785502,14.308239,13.032433,11.664027,11.327928,11.540562,10.669447,10.744898,13.1421795,16.78783,18.180243,12.22648,14.339106,31.363577,55.72051,65.409096,23.03311,14.205351,18.279701,26.19176,40.42798,37.780334,27.155474,17.473747,11.80121,7.363324,6.108095,12.710052,14.033872,7.8023114,2.5824795,3.74168,4.1120753,3.99204,4.0194764,5.1752477,4.479041,4.1017866,3.8925817,3.525616,2.5070283,2.253239,1.8382589,1.6599203,1.7182233,1.5947582,1.6016173,1.6221949,1.488441,1.2758065,1.3169615,1.4095604,1.3101025,1.1592005,1.1180456,1.3443983,1.6016173,1.4815818,1.4369972,1.5776103,1.6942163,2.1400626,2.3149714,2.0886188,1.670209,1.605047,1.5981878,1.7593783,1.728512,1.5090185,1.4507155,1.5021594,1.4095604,1.3409687,1.3752645,1.5055889,1.8931323,2.0577524,2.1332035,2.1126258,1.8725548,1.529596,1.6359133,1.879414,2.0680413,2.1160555,2.4212887,3.2306714,4.197815,4.7979927,4.3281393,4.091498,4.588788,5.137522,5.6176643,6.475061,6.9552035,7.2192817,7.548522,8.100685,8.882631,8.999237,8.882631,9.009526,9.431366,9.80862,12.020704,12.648318,12.603734,12.586586,13.101024,13.210771,13.001566,12.864383,12.812939,12.4802685,11.026124,10.854645,10.398509,9.3079,8.447074,8.608265,8.793462,8.985519,9.427936,10.6145735,11.626302,12.205902,11.941824,11.31078,11.650309,11.372512,11.026124,10.244178,9.301042,9.132992,9.253027,9.856634,9.918367,9.325048,8.868914,7.613684,6.9963584,7.051232,7.9875093,10.213311,10.508256,10.096705,9.455373,9.067829,9.431366,11.430815,11.396519,11.118723,11.701753,13.584596,13.008426,13.783512,15.436573,16.911295,16.558048,17.19938,17.648657,18.025911,18.550638,19.548649,20.70785,21.825895,22.714157,23.420652,24.226606,24.888515,25.159454,24.816494,24.60386,26.250063,27.52244,27.374968,26.315224,25.059996,24.545557,23.485815,22.796469,22.117409,21.61669,21.969936,23.259462,24.10314,23.310905,21.465788,20.899906,20.604961,20.488356,20.934202,21.78817,22.36091,22.151705,22.429502,21.956219,20.337454,18.012194,17.768692,18.334574,19.102802,20.066517,21.798458,0.607037,0.6927767,0.83681935,0.939707,0.9842916,1.0220171,1.1283343,1.08032,0.9774324,0.89169276,0.85739684,1.0151579,1.2380811,1.3341095,1.3272504,1.4541451,1.2723769,1.2415106,1.3341095,1.4472859,1.3821237,1.605047,1.8897027,2.352697,2.7059445,2.270387,2.0097382,1.8965619,1.7662375,1.6907866,2.0028791,1.9582944,2.8465576,4.629943,6.728851,8.018375,8.416207,12.562579,16.37628,16.084764,8.241299,4.3692946,2.5241764,1.6427724,1.1351935,0.90884066,1.0151579,0.9534253,0.75450927,0.65162164,1.0871792,1.3821237,1.2209331,1.0220171,0.9259886,0.77165717,0.59674823,0.36010668,0.33609957,0.45956472,0.32581082,0.25378948,0.26750782,0.28808534,0.29837412,0.34638834,0.51100856,0.39440256,0.26407823,0.22978236,0.24007112,0.3806842,0.51100856,0.6344737,0.7339317,0.7682276,0.65505123,0.5693115,0.5761707,0.64476246,0.64133286,0.5521636,0.45956472,0.44927597,0.4664239,0.33952916,0.2469303,0.16804978,0.11317638,0.07545093,0.041155048,0.0274367,0.010288762,0.0,0.0,0.0,0.01371835,0.037725464,0.06516216,0.106317215,0.17147937,0.12003556,0.14061308,0.16462019,0.18519773,0.24007112,0.274367,0.23321195,0.15776102,0.08573969,0.0548734,0.12003556,0.13375391,0.17490897,0.26750782,0.36010668,0.4698535,0.65505123,1.0014396,1.4232788,1.6839274,1.3341095,0.9568549,0.59674823,0.3018037,0.12003556,0.058302987,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.08573969,0.044584636,0.037725464,0.048014224,0.061732575,0.07545093,0.08573969,0.082310095,0.05144381,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.037725464,0.044584636,0.0274367,0.037725464,0.06516216,0.106317215,0.15776102,0.12003556,0.08916927,0.06516216,0.0548734,0.072021335,0.12346515,0.14404267,0.14747226,0.17147937,0.26064864,0.2503599,0.274367,0.31552204,0.3566771,0.37382504,0.38754338,0.48014224,0.53844523,0.5555932,0.6241849,0.7510797,0.7339317,0.7579388,0.8196714,0.72707254,0.88826317,1.155771,1.1694894,1.0014396,1.155771,1.4438564,1.4164196,1.4472859,1.5536032,1.4061309,1.5055889,1.8142518,2.335549,2.9254382,3.2786856,3.8479972,4.681387,5.501058,5.9983487,5.8508763,6.355026,6.807731,7.5519514,8.800322,10.628291,12.63803,13.71492,14.706071,15.87213,16.852993,17.604073,18.807858,20.313446,21.657845,22.041958,22.28546,23.314335,23.986534,23.972816,23.739605,22.85477,22.933651,24.758192,26.496992,23.712168,21.013083,19.802439,19.023922,18.20082,17.436022,17.04848,16.571766,16.365992,16.657507,17.562918,17.919594,18.670673,19.658396,20.35803,19.87446,20.855322,21.229147,22.258022,24.53184,27.947708,28.153484,27.141756,25.965406,27.275509,35.33504,47.270004,52.87395,57.20895,61.293587,62.10297,62.751163,68.2728,72.031624,72.17567,71.63036,77.15886,75.13197,64.60314,49.8079,40.167328,37.279617,35.42078,31.689388,25.392666,18.063637,14.407697,11.153018,8.577398,6.948344,6.4887795,6.444195,7.2021337,8.210432,9.506817,11.705182,12.010415,11.55428,10.960961,10.13786,8.2653055,7.5210853,5.785714,4.0023284,3.0420442,3.6936657,3.6010668,4.482471,4.0537724,2.510458,2.5241764,1.7456601,1.2895249,0.980862,0.75450927,0.66876954,0.66191036,0.61389613,0.5624523,0.4972902,0.37725464,0.34295875,0.34981793,0.4081209,0.44584638,0.28465575,0.64133286,0.72021335,0.66533995,0.64476246,0.83681935,0.59674823,0.96714365,1.3615463,1.6256244,2.0337453,1.862266,1.8897027,1.7216529,1.4267083,1.5330256,1.6256244,1.762808,1.9411465,2.1057668,2.1469216,2.352697,3.357566,4.2835546,5.5250654,8.748878,10.88551,11.739478,11.934964,11.502836,9.877212,9.736599,8.186425,6.6293926,5.8234396,5.8817425,2.9563043,1.1592005,0.29837412,0.06516216,0.030866288,0.048014224,0.2503599,0.2777966,0.09602845,0.010288762,0.0034295875,0.22635277,0.25721905,0.16804978,0.53158605,0.922559,1.2758065,1.6427724,1.8999915,1.786815,2.2086544,1.8313997,1.762808,2.136633,2.095478,3.0111778,3.100347,3.3952916,3.923448,3.7142432,3.8685746,3.8445675,3.5804894,3.1586502,2.8259802,2.2120838,1.6667795,1.4918705,1.6016173,1.5364552,1.7490896,2.2360911,2.534465,2.551613,2.568761,2.627064,2.417859,2.5310357,2.942586,3.0111778,2.3561265,2.4555845,2.3252604,1.8245405,1.6770682,1.529596,1.2517995,1.3272504,1.704505,1.8039631,2.1194851,2.16064,2.393852,2.8088322,2.8980014,3.3198407,3.5873485,3.6319332,3.3678548,2.702515,2.4624438,2.1229146,2.510458,3.8685746,5.857735,6.48535,6.9860697,7.7440085,8.340756,7.5553813,7.846896,9.674867,10.271614,9.31133,8.916927,8.755736,7.4765005,6.5230756,6.012067,4.7602673,5.267846,6.310441,7.0443726,7.5862474,9.043822,10.024684,10.652299,10.738038,10.655728,11.31078,12.30536,12.408247,12.517994,12.744347,12.397959,12.566009,12.569438,12.277924,11.842365,11.677745,10.477389,10.072699,10.230459,10.666017,11.039842,11.362224,11.444533,11.8115,12.168177,11.396519,10.906088,10.679735,10.861504,11.567999,12.912396,13.437123,14.435134,15.093615,14.822677,13.245067,13.989287,12.644889,11.88352,12.168177,11.773774,10.48082,10.748327,11.290202,12.761495,17.772121,11.945253,13.327377,24.699888,39.868954,43.66208,22.340332,13.663476,14.7095,21.290878,27.927132,23.420652,14.428274,8.625413,7.466212,6.1732574,6.2658563,13.437123,17.36057,13.6086035,3.6696587,4.48933,4.5819287,4.341858,4.3761535,5.4804807,4.6916757,4.355576,3.974892,3.2958336,2.277246,1.9754424,1.5604624,1.5638919,1.8245405,1.5021594,1.5330256,1.5193073,1.3581166,1.138623,1.1626302,1.2449403,1.2175035,1.1111864,1.0597426,1.2792361,1.7902447,1.7593783,1.6736387,1.7730967,2.061182,2.5756202,2.6407824,2.2669573,1.7388009,1.587899,1.3615463,1.2963841,1.2072148,1.1146159,1.2620882,1.4198492,1.2895249,1.1729189,1.1866373,1.2483698,1.5741806,1.8142518,2.0063086,2.07833,1.8691251,1.6153357,1.7422304,1.9342873,2.0680413,2.2120838,2.4041407,3.1072063,3.9714622,4.482471,3.974892,3.7931237,4.0674906,4.5201964,5.0106273,5.5422134,6.5813785,7.5279446,8.107545,8.467651,9.177576,9.818909,9.97324,10.168727,10.532263,10.762046,13.354814,14.424845,14.688923,14.640909,14.54831,13.71492,13.361672,13.227919,13.186764,13.245067,12.175035,11.770344,11.05356,9.97667,9.400499,10.000677,9.897789,9.534253,9.451943,10.319629,11.523414,12.377381,12.020704,10.686595,9.685155,10.209882,10.028113,9.441654,9.002667,9.513676,9.73317,10.323058,10.652299,10.460241,9.849775,7.864044,6.948344,6.9792104,8.128122,10.868362,12.130451,11.880091,11.173596,10.611144,10.323058,12.147599,12.439114,12.006986,12.178465,14.784951,14.123041,14.555169,15.422854,16.005884,15.553179,16.400288,17.638369,19.03421,20.244854,20.79016,21.44178,21.860191,22.52896,23.509823,24.4461,24.44953,24.504402,24.326063,24.384367,25.910534,26.795366,25.728765,24.254042,23.396646,23.677872,23.454948,23.434372,23.101702,22.70044,23.252604,23.725885,24.243753,23.35549,21.558388,21.314886,21.356041,20.652975,20.893047,21.69557,20.62554,21.53781,22.5221,22.10712,20.124819,17.700102,17.926455,18.238546,18.903887,20.19341,22.384918,0.66533995,0.6379033,0.85739684,1.0494537,1.0837497,0.9568549,1.1111864,0.96714365,0.8779744,0.94656616,1.0357354,1.138623,1.2380811,1.3032433,1.3409687,1.4027013,1.4095604,1.4267083,1.3443983,1.2175035,1.2723769,1.5398848,1.6976458,1.9720128,2.1640697,1.6839274,1.762808,1.7319417,1.7353712,1.8965619,2.3149714,2.318401,3.4398763,5.0106273,6.6739774,8.364764,8.385342,12.466551,15.63206,14.164196,5.593657,3.5187566,2.2155135,1.5261664,1.2620882,1.1900668,1.5913286,1.4644338,1.0117283,0.66876954,1.1111864,1.7216529,1.3649758,0.9328478,0.823101,0.9568549,0.64476246,0.36353627,0.33952916,0.4698535,0.3018037,0.23664154,0.2777966,0.32924038,0.36010668,0.38754338,0.51100856,0.37382504,0.22635277,0.18862732,0.26407823,0.4389872,0.6276145,0.7990939,0.8848336,0.7922347,0.5796003,0.6344737,0.8745448,1.0734608,0.8711152,0.5727411,0.4629943,0.5658819,0.7305021,0.64133286,0.4938606,0.35324752,0.22635277,0.13032432,0.06859175,0.030866288,0.020577524,0.017147938,0.01371835,0.010288762,0.044584636,0.09602845,0.15433143,0.20234565,0.2469303,0.17833854,0.1371835,0.14061308,0.18862732,0.2709374,0.31552204,0.28808534,0.20920484,0.12003556,0.09259886,0.11317638,0.1371835,0.16804978,0.19891608,0.20920484,0.19891608,0.274367,0.45613512,0.72707254,1.039165,0.82996017,0.5693115,0.30523327,0.10288762,0.044584636,0.020577524,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.034295876,0.024007112,0.0274367,0.037725464,0.017147938,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0274367,0.06516216,0.061732575,0.05144381,0.034295876,0.034295876,0.048014224,0.041155048,0.06859175,0.106317215,0.15433143,0.216064,0.26750782,0.2709374,0.3018037,0.39440256,0.47671264,0.3806842,0.35324752,0.45613512,0.4972902,0.52815646,0.8265306,0.70649505,0.6927767,0.78537554,0.85739684,0.66876954,0.8676856,1.1180456,1.1900668,1.1283343,1.2517995,1.1866373,1.1283343,1.1489118,1.2312219,1.2449403,1.3752645,1.8759843,2.4418662,2.8705647,3.0557625,3.9028704,4.479041,4.839148,5.113515,5.4941993,6.3035817,6.941485,7.6857057,8.851766,10.799771,12.744347,13.375391,14.009865,15.103903,16.280252,16.828985,17.339994,18.272842,19.70298,21.328604,21.225718,22.810186,23.650434,23.129137,22.44322,22.487804,22.065966,23.69502,26.34609,25.450968,21.904776,20.296299,19.744135,19.377169,18.317427,18.145947,18.022482,18.02934,18.221397,18.636377,19.157675,20.502073,21.20514,20.848463,20.04251,19.432043,19.428614,20.467777,21.901346,22.004232,23.705309,25.035988,25.327503,26.798796,34.525658,44.88987,49.430645,55.933144,63.903503,64.589424,70.95131,79.37094,82.21064,80.46498,83.77796,93.34308,83.46244,65.55313,49.48552,43.55576,40.455414,38.17817,32.65996,23.705309,14.997586,10.686595,7.73372,5.9434752,5.099797,4.9351764,5.892031,7.425057,8.759167,10.216741,13.22106,14.812388,14.30481,13.598314,12.747777,9.949233,7.7577267,6.111525,4.6848164,4.2081037,6.4819202,5.4770513,8.848335,8.553391,4.4550343,4.3281393,2.719663,1.7765263,1.2003556,0.83338976,0.66876954,0.6276145,0.5212973,0.42526886,0.36696586,0.31552204,0.33266997,0.36010668,0.3566771,0.33266997,0.33952916,0.9259886,1.0288762,0.89512235,0.7682276,0.91569984,0.89855194,1.6496316,2.3286898,2.836269,3.7965534,3.1895163,2.9220085,2.2498093,1.4061309,1.5844694,2.1229146,2.318401,2.6956558,3.192946,3.1517909,3.4021509,5.1066556,6.914048,9.023245,13.183334,13.186764,13.906977,13.495427,11.694893,9.846346,11.595435,10.792912,8.738589,6.40304,4.420738,1.7422304,0.5453044,0.13375391,0.05144381,0.106317215,0.10288762,0.048014224,0.006859175,0.0034295875,0.01371835,0.0034295875,0.4698535,0.5521636,0.36010668,0.97400284,1.3649758,1.7113642,2.2738166,2.6167753,1.6084765,1.9171394,1.8759843,1.6633499,1.670209,2.5001693,3.5564823,3.899441,4.7191124,5.936616,6.2212715,5.662249,5.3227196,4.8734436,4.341858,4.1120753,3.6696587,2.7333813,1.9857311,1.6359133,1.3752645,2.287535,3.2272418,3.4913201,3.1895163,3.2581081,3.7691166,3.8171308,3.4433057,2.760818,1.961724,2.4761622,2.3767042,2.3081124,2.218943,1.3409687,1.6084765,1.2620882,1.1317638,1.3855534,1.5638919,1.7593783,2.3595562,2.4212887,2.2463799,3.3850029,3.9543142,3.9851806,3.8479972,3.4707425,2.3149714,1.7662375,2.1091962,2.8019729,3.789694,5.5113473,6.2212715,5.878313,6.2144127,7.390761,7.9909387,7.2295704,8.419638,9.47938,9.647429,9.5033865,8.196714,6.3035817,5.411889,5.470192,4.7945633,5.113515,5.9160385,6.842027,7.654839,8.220721,9.72288,10.525404,10.700313,10.700313,11.345076,11.756626,11.694893,11.828648,12.089295,11.667457,11.533703,10.991828,10.494537,10.172156,9.818909,8.916927,9.431366,10.415657,11.180455,11.303921,11.794352,11.753197,11.993267,12.46998,12.284782,11.667457,11.465111,11.444533,11.825217,13.282792,13.728639,14.692352,15.4914465,15.357693,13.440554,13.529722,12.267634,11.893809,12.63117,12.672326,11.358793,11.55771,9.619993,8.165848,16.084764,12.13731,8.800322,10.443094,16.695232,22.480946,28.599329,21.129688,12.768354,11.214751,19.164536,19.315437,12.939834,7.7748747,6.166398,5.051782,7.9257765,16.945591,22.875349,19.802439,5.137522,5.0174866,4.4859004,4.139512,4.386442,5.4187484,4.6848164,4.2423997,3.7108135,2.9322972,1.9651536,1.7388009,1.4027013,1.4747226,1.8142518,1.6221949,1.4678634,1.3203912,1.1592005,1.0494537,1.1249046,1.2586586,1.371835,1.2895249,1.1489118,1.4027013,1.8176813,1.7422304,1.6736387,1.8313997,2.1743584,2.6236343,2.469303,2.0097382,1.546744,1.3821237,1.0151579,0.8025235,0.7373613,0.85739684,1.2655178,1.4610043,1.2963841,1.1694894,1.214074,1.3032433,1.6393428,1.7319417,1.8005334,1.8897027,1.862266,1.7422304,1.8965619,2.1057668,2.2841053,2.4761622,2.6750782,3.2786856,3.8479972,4.057202,3.7039545,3.7931237,3.9303071,4.372724,5.0140567,5.3878818,6.2247014,7.473071,8.385342,8.9100685,9.688584,10.463672,10.655728,11.105004,11.921246,12.47341,14.623761,15.29596,15.29939,15.114192,14.904987,13.450842,13.279363,13.560589,13.896688,14.335675,14.150477,13.560589,12.394529,11.163307,11.077567,10.950673,10.336777,9.966381,10.089847,10.487679,11.924676,13.114742,13.402828,12.476839,10.374502,10.755186,10.216741,9.849775,9.938945,9.959522,9.496528,9.383351,9.839486,10.39165,9.873782,7.301592,6.550512,6.9552035,8.399059,11.303921,13.056439,12.706621,12.151029,11.958971,11.362224,11.921246,12.583157,12.545431,12.356804,13.951562,14.620332,15.13134,15.45715,15.529172,15.244516,16.770683,18.471758,20.320305,21.736725,21.572105,22.052248,22.323185,22.889067,23.797907,24.627867,24.072275,23.917942,23.574984,23.218307,23.77733,24.497543,22.906214,21.410915,21.04052,21.431492,22.631847,23.660725,24.27462,24.569565,25.008553,24.175161,23.70188,22.916504,22.076254,22.336903,22.559826,20.807306,19.79901,19.740705,18.362011,20.409475,22.36091,22.53925,20.659836,17.806417,17.511473,17.590355,18.639809,20.52951,22.415783,0.64133286,0.6036074,0.65848076,0.70306545,0.7339317,0.8711152,1.0151579,0.83338976,0.8196714,0.99801,0.90198153,0.9362774,0.90884066,0.9568549,1.1214751,1.3443983,1.5261664,1.7079345,1.7079345,1.5776103,1.6016173,1.371835,1.2312219,1.4438564,1.7696671,1.4644338,1.7593783,1.7216529,1.8862731,2.3389788,2.7299516,2.5961976,4.431027,6.2144127,7.425057,9.047252,9.585697,14.507155,16.815268,13.663476,6.3618846,3.8479972,2.1846473,1.3615463,1.1763484,1.2517995,1.8965619,1.8691251,1.3066728,0.7442205,1.097468,1.4164196,1.0460242,0.58988905,0.44584638,0.823101,0.5693115,0.26407823,0.106317215,0.12003556,0.16804978,0.2777966,0.48014224,0.5761707,0.5212973,0.4115505,0.38754338,0.35324752,0.29837412,0.28808534,0.45613512,0.6036074,0.66876954,0.764798,0.8779744,0.85396725,0.5624523,0.67219913,1.0117283,1.2517995,0.8848336,0.50757897,0.42183927,0.7133542,1.1900668,1.371835,1.1283343,0.7579388,0.39783216,0.14404267,0.044584636,0.044584636,0.072021335,0.08573969,0.06859175,0.044584636,0.06859175,0.23321195,0.34295875,0.33266997,0.26064864,0.20920484,0.18862732,0.20234565,0.2469303,0.31895164,0.29494452,0.24350071,0.16462019,0.09259886,0.09259886,0.15090185,0.33266997,0.4115505,0.32924038,0.18176813,0.13375391,0.19548649,0.29837412,0.39097297,0.42869842,0.31895164,0.19891608,0.09945804,0.044584636,0.044584636,0.020577524,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.0,0.048014224,0.024007112,0.0,0.0034295875,0.01371835,0.01371835,0.05144381,0.106317215,0.14747226,0.12346515,0.28122616,0.40126175,0.44584638,0.41840968,0.3806842,0.3806842,0.490431,0.5144381,0.53501564,0.89855194,0.77851635,0.6927767,0.66876954,0.71678376,0.84024894,0.9602845,0.9294182,0.9945804,1.2037852,1.371835,0.7990939,0.77508676,0.8162418,0.8162418,1.039165,1.3066728,1.6839274,2.2463799,2.8225505,3.0043187,3.8377085,3.7965534,4.15666,5.23698,6.4098988,6.6533995,7.281014,8.241299,9.445084,10.789482,12.950122,13.588025,13.838386,14.267084,14.87755,15.817257,16.016174,15.889278,16.582056,19.973917,20.045938,20.79016,21.10568,20.930773,21.208569,22.504953,22.388348,23.334913,25.60873,27.282368,25.0257,23.417223,22.371199,21.53781,20.29287,19.682402,19.274282,19.404606,19.69955,19.089085,19.442331,19.521212,19.949911,20.395756,19.576086,19.613811,18.752985,18.691252,19.6241,20.234566,24.494114,26.713057,27.645905,29.384705,35.355618,42.362263,49.873062,57.21924,64.19845,71.06105,77.12799,83.90829,86.50791,87.69798,97.91472,110.573326,91.85807,69.0959,55.898846,52.14002,50.0514,43.716953,32.725124,20.073376,12.175035,8.64942,6.111525,4.4447455,3.5564823,3.3712845,5.521636,8.244728,10.569988,12.157887,13.306799,16.674654,16.071047,15.031882,14.404267,12.329367,10.254466,8.7283,6.7391396,5.212973,7.0203657,5.3227196,13.63261,14.760944,7.380472,6.012067,3.4844608,1.9925903,1.1797781,0.77851635,0.59674823,0.5453044,0.45270553,0.3841138,0.36353627,0.34981793,0.4972902,0.45956472,0.41840968,0.45956472,0.59674823,0.7407909,0.97057325,1.0494537,1.0117283,1.1592005,1.1214751,2.2498093,3.6044965,4.6882463,5.4324665,5.5662203,4.437886,3.0866287,2.2052248,2.1194851,2.867135,3.4638834,4.331569,5.360445,5.936616,5.3261495,7.31531,10.4705305,13.293081,14.222499,11.694893,13.231348,15.446862,16.009314,13.639469,13.896688,11.489118,7.81603,4.1155047,1.4815818,0.6379033,0.20920484,0.041155048,0.09602845,0.4115505,0.44927597,0.18176813,0.0,0.01371835,0.061732575,0.01371835,0.082310095,0.32581082,0.7305021,1.2037852,1.155771,1.7319417,2.5893385,3.0111778,1.8759843,1.4267083,1.4850113,1.4918705,1.6942163,3.1586502,3.5599117,3.4707425,4.605936,6.831738,8.162418,7.0272245,6.7631464,6.2247014,5.305572,4.928317,5.4153185,4.32128,2.7711067,1.7559488,2.1194851,2.5721905,3.3987212,3.5393343,3.1860867,3.782835,3.210094,3.8377085,3.57363,2.5721905,3.2203827,2.620205,2.2326615,2.0440342,1.9137098,1.5707511,1.4507155,1.4472859,1.488441,1.5741806,1.7696671,1.6221949,2.1194851,2.503599,2.4795918,2.2120838,2.0303159,2.486451,3.2066643,3.5976372,2.8534167,2.1572106,2.294394,3.2649672,4.4859004,4.791134,5.07236,6.159539,7.1095347,7.7577267,8.697433,7.781734,8.779744,9.304471,8.759167,8.330468,7.2192817,6.210983,5.5559316,5.195825,4.746549,5.610805,6.615674,7.226141,7.3187394,7.1712675,8.282454,9.3764925,9.959522,10.1481495,10.635151,10.6488695,10.6317215,10.9369545,11.38623,11.276484,11.691463,11.180455,10.652299,10.621432,11.245617,9.427936,9.602845,10.511685,11.290202,11.4754,11.732618,11.235329,11.334786,11.993267,11.8115,11.797781,12.21619,12.325937,12.332796,13.38225,13.210771,13.039291,13.663476,14.29452,12.572867,13.2690735,12.144169,11.283342,11.489118,12.284782,12.394529,12.895248,10.6317215,8.200144,13.96185,15.999025,10.768905,7.274155,10.64201,22.141417,40.037003,35.547672,20.834743,8.632272,12.205902,16.029892,15.608052,11.818358,7.040943,5.171818,10.422516,26.802225,35.50652,27.817385,5.1100855,3.549623,3.3781435,3.782835,4.3452873,5.0655007,4.5167665,3.782835,3.083199,2.4418662,1.7079345,1.6976458,1.4267083,1.3478279,1.4987297,1.5090185,1.3752645,1.1694894,1.0528834,1.0528834,1.0528834,1.3203912,1.5707511,1.4747226,1.1729189,1.2826657,1.5364552,1.4095604,1.4027013,1.5776103,1.5398848,1.786815,1.7559488,1.5536032,1.2620882,0.9294182,0.5521636,0.4115505,0.5453044,0.9362774,1.5090185,1.4507155,1.3238207,1.2998136,1.4267083,1.6324836,1.6084765,1.5638919,1.546744,1.5673214,1.6187652,1.5570327,1.6221949,1.8176813,2.1091962,2.4247184,3.0351849,3.765687,4.1635194,4.0846386,3.6936657,3.8891523,4.0023284,4.4756117,5.2164025,5.56965,6.0566516,7.040943,7.449064,7.589677,9.139851,10.323058,11.012405,11.653738,12.55915,13.900118,15.278812,15.422854,14.726648,13.893259,13.917266,12.840376,12.956982,13.653188,14.568888,15.594335,15.532601,14.640909,13.344524,12.46998,13.214201,12.284782,11.485688,11.314209,11.784062,12.404818,13.625751,13.9481325,13.63261,12.867812,11.780633,11.4376745,10.007536,9.39021,9.935514,10.436234,10.069269,9.657719,9.788043,10.494537,11.276484,9.798331,8.083538,8.083538,10.093276,12.754636,13.416546,12.782072,12.229909,12.130451,11.8869505,11.458252,12.651748,13.426835,13.1593275,12.634601,13.245067,13.718349,14.5585985,15.584045,15.913286,17.099922,18.86959,20.70099,21.891056,21.561817,22.926792,24.322634,25.084003,25.042849,24.504402,22.662714,22.731306,22.43979,21.726437,22.751883,23.581844,22.762173,21.877338,21.421204,20.797018,22.151705,23.69159,24.843931,25.413242,25.557285,23.739605,22.645567,21.801888,21.517231,22.87192,23.11542,21.174273,19.775002,19.53493,18.934752,21.45207,22.53582,22.487804,21.506943,19.69955,17.490896,17.29541,18.557497,20.584383,22.53582,0.8471081,0.7442205,1.039165,1.1249046,0.9328478,0.9294182,0.8711152,0.7613684,0.84367853,1.0357354,0.9362774,1.2860953,1.2415106,1.1934965,1.3443983,1.7079345,1.7662375,2.0714707,2.2360911,2.1126258,1.786815,1.6496316,1.6016173,1.6667795,1.728512,1.5021594,1.7079345,1.5673214,1.6153357,1.9823016,2.4007113,2.4247184,4.149801,6.1972647,7.7371492,8.512236,11.763485,17.62808,18.886738,13.807519,6.166398,3.4192986,1.8931323,1.2758065,1.1729189,1.1283343,1.5433143,1.4027013,0.980862,0.607037,0.64819205,0.8471081,0.6241849,0.37039545,0.32238123,0.5555932,0.5727411,0.4355576,0.29151493,0.26064864,0.4355576,0.78194594,0.96714365,0.96714365,0.8196714,0.6310441,0.51100856,0.3841138,0.28808534,0.2709374,0.432128,0.64819205,0.8025235,0.8711152,0.86082643,0.805953,0.6893471,0.9294182,1.2655178,1.3615463,0.7990939,0.50757897,0.607037,1.0254467,1.546744,1.786815,1.5330256,0.91912943,0.37725464,0.09945804,0.020577524,0.08916927,0.14061308,0.18176813,0.2194936,0.25378948,0.22978236,0.20234565,0.19891608,0.24007112,0.33266997,0.34295875,0.31209245,0.26750782,0.22292319,0.19891608,0.1920569,0.13032432,0.082310095,0.1097468,0.274367,0.3566771,0.45270553,0.4389872,0.31895164,0.23321195,0.24007112,0.25721905,0.28465575,0.32581082,0.40126175,0.33266997,0.29494452,0.22635277,0.1371835,0.106317215,0.05144381,0.024007112,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.010288762,0.01371835,0.006859175,0.0,0.0034295875,0.024007112,0.048014224,0.07545093,0.116605975,0.2194936,0.31895164,0.39783216,0.36696586,0.31895164,0.5144381,0.5555932,0.5555932,0.5041494,0.47671264,0.65505123,0.52472687,0.5624523,0.66876954,0.7476501,0.70649505,0.9842916,1.2963841,1.3375391,1.1592005,1.1660597,1.0425946,0.85739684,0.7888051,0.91912943,1.2449403,1.2106444,1.7319417,2.3767042,2.8294096,2.884283,3.069481,3.8788633,4.7534084,5.329579,5.456474,6.228131,7.1712675,8.035523,8.81061,9.712592,11.571428,12.898679,14.345964,15.402277,14.400838,14.5585985,14.1299,13.642899,13.978998,16.396858,17.065628,18.79071,19.884748,20.255144,21.404055,22.738165,23.043398,24.521551,27.52244,30.540476,29.456726,28.932,27.42984,25.080574,23.69845,20.978786,18.969048,17.724108,17.367432,18.073925,18.118511,18.691252,19.54179,20.21056,20.028791,20.584383,21.287449,22.480946,24.500973,27.6802,29.165213,29.806545,30.571342,33.311584,40.726353,44.48861,53.216908,63.41307,72.19968,77.32348,79.9917,81.3361,81.3018,82.41642,89.81061,87.684265,75.46121,62.68943,53.882248,48.501225,42.90071,35.215004,25.567575,15.906426,10.028113,7.9737906,6.447624,5.137522,4.173808,4.1155047,4.9180284,7.9737906,11.0981455,13.087306,13.697772,15.443433,14.531162,13.536582,13.55373,14.171056,11.413667,10.851214,10.052121,8.570539,7.9463544,6.1149545,12.812939,15.806969,12.607163,10.48082,5.0414934,2.2669573,1.0837497,0.72707254,0.7305021,0.67219913,0.6893471,0.71678376,0.7579388,0.91227025,0.8162418,0.6893471,0.64133286,0.72364295,0.9362774,1.0734608,1.2620882,1.4987297,1.7147937,1.7936742,2.1572106,3.3712845,4.911169,6.0737996,5.970912,6.3173003,5.593657,5.305572,5.4907694,4.7328305,4.372724,4.338428,5.038064,6.3378778,7.548522,6.427047,9.712592,12.603734,13.433694,13.646329,13.13189,15.752095,17.854433,17.95389,16.715809,14.699212,11.026124,6.5059276,2.4555845,0.6859175,0.26407823,0.09259886,0.034295876,0.072021335,0.3018037,0.13375391,0.037725464,0.0,0.0034295875,0.01371835,0.0034295875,0.017147938,0.36696586,0.94999576,1.2415106,1.0871792,0.922559,1.2517995,1.6290541,0.66876954,2.218943,2.1057668,2.2258022,3.450165,5.6485305,5.504488,7.0718093,7.9600725,8.080108,9.616563,9.613133,8.320179,7.0752387,6.4819202,6.4064693,7.051232,6.697984,5.830299,4.804852,3.841138,2.8980014,3.175798,3.5770597,3.6799474,3.758828,4.1429415,3.9371665,3.5839188,3.2512488,2.8534167,3.2203827,2.4761622,2.1400626,2.4212887,2.2052248,2.3081124,2.1640697,1.8656956,1.7182233,2.2463799,2.1880767,2.5001693,2.767677,2.7813954,2.5413244,2.767677,3.1620796,3.2821152,3.093488,2.9631636,2.8225505,2.1983654,2.6613598,3.9543142,3.9851806,3.758828,4.770556,6.2864337,8.131552,10.662587,11.379372,9.523964,9.839486,11.1393,6.3173003,6.0086374,5.909179,5.4976287,4.791134,4.331569,5.501058,6.3310184,6.701414,6.6225333,6.23156,6.5127864,7.5382333,8.4264965,8.707723,8.327039,8.879202,9.595985,9.952662,9.846346,9.626852,10.072699,10.792912,11.478829,11.924676,12.037852,11.080997,10.923236,11.156448,11.382801,11.204462,10.816919,10.237319,10.871792,12.260776,12.065289,12.308789,12.490558,12.202472,11.742908,12.099585,12.22305,12.9809885,13.862392,14.140189,12.878101,13.924125,13.474849,12.555719,12.044711,12.662037,12.21619,13.1593275,11.982979,9.3936405,10.31277,18.36544,14.249936,10.065839,12.5145645,22.909645,32.67025,28.119188,18.392878,10.755186,10.583707,16.894148,15.913286,10.960961,5.8474464,4.880303,16.96617,25.811075,26.812515,18.746124,3.806842,3.2992632,3.7142432,4.0229063,4.0023284,4.2355404,3.6182148,2.976882,2.428148,2.037175,1.8313997,1.4781522,1.3341095,1.3786942,1.471293,1.3752645,1.2895249,1.1832076,1.1008976,1.1351935,1.4198492,1.5227368,1.670209,1.5090185,1.2037852,1.4404267,1.529596,1.704505,1.8416885,1.7319417,1.0906088,1.4027013,1.2209331,0.85739684,0.5521636,0.4664239,0.35324752,0.39440256,0.5624523,0.8505377,1.2792361,1.3924125,1.3272504,1.3203912,1.3992717,1.3512574,1.4850113,1.4815818,1.4164196,1.4198492,1.6530612,1.6221949,1.7936742,1.8862731,1.9342873,2.2806756,2.7642474,3.2992632,3.6182148,3.6044965,3.3026927,3.4878905,4.2423997,5.1100855,5.7102633,5.7411294,6.8626046,7.7131424,7.857185,7.7028537,8.491658,9.784613,10.521975,11.105004,12.05157,14.009865,15.059319,15.227368,14.946142,14.596324,14.500296,14.256795,14.184773,14.064738,14.054449,14.678635,15.234227,14.7197895,14.21564,14.174485,14.421415,13.505715,12.3911,11.832077,12.123591,13.125031,13.293081,13.320518,12.46312,11.461681,12.572867,13.080446,12.8197975,12.380811,11.876661,10.960961,11.231899,10.799771,10.679735,11.369082,12.864383,13.516005,12.38424,11.753197,11.849225,10.827208,10.401938,10.707172,11.046701,11.393089,12.397959,12.812939,13.125031,12.442543,11.365653,11.976119,11.862943,12.250486,13.152468,14.441993,15.865272,17.04162,18.4649,19.524641,20.124819,20.69413,22.28546,24.651875,25.488693,24.569565,23.749893,23.485815,23.022821,22.350622,21.7916,22.007662,23.177153,23.550978,22.837624,21.77788,22.151705,23.633287,24.744474,25.450968,25.622448,24.998262,23.050257,22.134558,22.261452,23.03311,23.667583,23.20802,21.644127,20.728426,20.985645,21.69557,23.417223,23.297188,23.070835,22.895926,21.335464,20.100813,19.87789,19.94305,20.169403,21.047379,0.70649505,0.65848076,0.82996017,0.8745448,0.78194594,0.85396725,0.7373613,0.6756287,0.764798,0.91569984,0.85396725,1.2243627,1.4232788,1.4369972,1.4404267,1.7902447,1.961724,2.2978237,2.2978237,1.9651536,1.786815,1.7113642,1.7113642,1.7490896,1.8656956,2.170929,2.1332035,1.8142518,1.7182233,1.9582944,2.2566686,2.534465,4.0709205,5.861165,7.284444,8.093826,13.649758,17.267973,15.721229,9.719451,3.9028704,2.3424082,2.0131679,1.7593783,1.2895249,1.2072148,2.2669573,1.5638919,0.69963586,0.36353627,0.34295875,0.44584638,0.4046913,0.31209245,0.31552204,0.607037,0.6036074,0.52472687,0.48357183,0.5624523,0.805953,1.0185875,1.0563129,0.9911508,0.8471081,0.59674823,0.50757897,0.53501564,0.53158605,0.48357183,0.51100856,0.6962063,0.8676856,0.85396725,0.70306545,0.6927767,0.7373613,0.97057325,1.2620882,1.3272504,0.7339317,0.53844523,0.6207553,0.9568549,1.3375391,1.3992717,1.1043272,0.6001778,0.20920484,0.05144381,0.041155048,0.12003556,0.17833854,0.26407823,0.39097297,0.53501564,0.37382504,0.2503599,0.22978236,0.3018037,0.4046913,0.42183927,0.39440256,0.3566771,0.34295875,0.39783216,0.29494452,0.22635277,0.2503599,0.34981793,0.44927597,0.42526886,0.490431,0.5144381,0.44584638,0.30866286,0.274367,0.28122616,0.30523327,0.31552204,0.2777966,0.32581082,0.32924038,0.274367,0.18176813,0.08573969,0.048014224,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.006859175,0.006859175,0.010288762,0.010288762,0.020577524,0.044584636,0.0548734,0.06516216,0.12346515,0.25378948,0.31552204,0.30523327,0.274367,0.34638834,0.4389872,0.44927597,0.47328308,0.5658819,0.72364295,0.6344737,0.6824879,0.70649505,0.6962063,0.7990939,1.2483698,1.5330256,1.3375391,0.89512235,0.9774324,0.8779744,0.83338976,0.89512235,1.1043272,1.5158776,1.371835,1.8931323,2.4898806,2.8945718,3.1449318,3.3609958,4.1772375,4.955754,5.4976287,6.060081,6.8111606,7.531374,8.285883,9.270175,10.81006,12.202472,13.413116,14.579176,15.189643,14.061309,13.807519,13.111313,12.127021,11.640019,13.049581,14.520873,16.160215,17.388008,18.416885,20.244854,22.487804,23.904224,26.147175,30.228384,36.49081,35.7363,35.16356,32.11123,27.17262,24.175161,20.913624,18.21111,16.925014,17.20967,18.516342,18.584934,19.44919,20.910194,22.456938,23.245745,25.838512,26.798796,25.255482,22.44665,21.705858,22.923363,24.960537,27.278938,31.106358,39.423107,46.46405,56.149204,66.91811,76.603264,82.450714,84.31298,83.38699,81.09946,79.27492,80.159744,69.356544,60.237274,52.13659,44.65666,37.66716,30.866287,23.983105,17.346853,11.667457,8.06296,7.06838,6.2075534,5.5490727,5.192395,5.302142,5.6828265,7.740579,10.302481,12.020704,11.369082,12.71691,12.751206,12.260776,12.394529,14.634049,13.512574,14.040731,15.71437,16.657507,13.6086035,10.405369,12.075578,13.347955,12.116733,9.455373,5.669108,3.1072063,1.7250825,1.2415106,1.1283343,1.1283343,1.1626302,1.4369972,1.920569,2.3424082,2.2292318,1.8931323,1.670209,1.6770682,1.7902447,1.8656956,1.9891608,2.1263442,2.2223728,2.1743584,2.352697,3.3198407,4.8905916,6.4133286,6.800872,6.416758,6.842027,7.490219,7.658269,6.5127864,5.950334,6.252138,7.0306544,8.320179,10.5597,14.483148,15.79325,17.37429,19.675543,20.70785,18.79071,18.173384,18.142517,17.658945,15.343974,13.306799,9.650859,5.4667625,1.961724,0.4698535,0.15090185,0.06859175,0.06859175,0.09259886,0.14747226,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.32581082,0.823101,0.8471081,0.5761707,0.7339317,1.1694894,1.5604624,1.4369972,1.7662375,2.3561265,3.5976372,5.717122,8.769455,9.39021,9.057541,8.673427,9.3936405,12.644889,11.540562,9.441654,8.501947,8.927217,8.961512,8.718011,8.436785,7.840037,6.8111606,5.3981705,4.170378,3.974892,3.724532,3.2958336,3.532475,3.2615378,3.2272418,3.2443898,3.059192,2.3424082,3.4055803,2.843128,2.5378947,2.750529,2.0989075,2.318401,2.5756202,2.8156912,2.983741,3.0248961,2.760818,2.7128036,2.4967396,2.386993,3.3198407,3.0489032,3.3232703,3.433017,3.2581081,3.2821152,2.9322972,2.8534167,3.0729103,3.5118976,3.9954693,4.173808,4.945465,6.5024977,9.033533,12.699762,11.979549,8.988949,7.7783046,8.200144,5.90575,5.305572,5.254128,5.0003386,4.479041,4.3452873,4.57164,5.0826488,5.5387836,5.751418,5.703404,6.4887795,7.431916,7.675417,7.3187394,7.394191,8.107545,8.988949,9.609704,9.801761,9.674867,9.547972,10.583707,11.948683,12.6757555,11.688034,11.4205265,10.995257,10.899229,11.238758,11.760056,11.177026,10.782623,10.950673,11.506266,11.729189,12.253916,12.507706,12.233338,11.574858,11.084427,11.739478,12.655178,13.512574,13.992717,13.759505,13.402828,12.9638405,12.487128,12.243628,12.737488,11.955542,12.528283,11.986408,10.295622,9.884071,16.002455,12.46312,9.369633,12.566009,23.650434,32.99606,26.167753,18.12194,14.147048,9.866923,16.410576,14.603184,9.235879,6.8969,15.964729,20.179693,19.829874,15.553179,9.112414,3.3781435,3.57363,3.7725463,3.9474552,4.016047,3.8548563,2.976882,2.4727325,2.2052248,2.0406046,1.8416885,1.4198492,1.2860953,1.3546871,1.4678634,1.3889829,1.2483698,1.08032,1.0666018,1.2415106,1.4644338,1.5638919,1.6804979,1.6290541,1.4987297,1.6633499,1.6256244,1.5055889,1.4164196,1.255229,0.7099246,0.8128122,0.6859175,0.45956472,0.26064864,0.22292319,0.18862732,0.40126175,0.65505123,0.8848336,1.1660597,1.5947582,1.4027013,1.2106444,1.2346514,1.2723769,1.546744,1.6427724,1.5707511,1.4815818,1.6907866,1.5330256,1.7182233,1.845118,1.8759843,2.1434922,2.2566686,2.5070283,2.9151495,3.2683969,3.1037767,3.6319332,4.341858,5.0826488,5.720552,6.1492505,6.601956,6.941485,7.010077,7.0375133,7.6342616,8.587687,9.482809,10.374502,11.516555,13.37882,15.155347,16.11906,16.269962,15.71437,14.640909,14.38369,14.932424,14.452282,13.125031,13.1593275,13.96185,13.958421,14.376831,15.199932,15.145059,14.099034,12.205902,10.967821,10.909517,11.574858,12.898679,13.210771,12.706621,12.096155,12.607163,12.823228,12.960411,13.505715,14.044161,13.272504,12.271064,11.646879,11.4376745,11.736049,12.682614,13.639469,12.857523,11.406808,9.97324,8.844906,8.999237,9.541112,10.079557,10.827208,12.600305,13.070158,12.6929035,11.777204,11.187314,12.349944,11.742908,12.034423,12.8197975,13.855534,15.083325,16.403717,18.11165,19.315437,19.925903,20.670124,21.232576,23.11199,24.130577,23.972816,24.171732,22.666143,22.398636,23.153145,24.079134,23.68816,23.502962,23.472097,23.334913,23.067406,22.875349,23.643576,24.727325,25.34122,25.300066,24.994833,23.623,23.808197,24.696459,25.44068,25.173172,25.059996,24.02426,22.648996,21.963078,23.44809,24.284908,24.336353,24.147726,23.743034,22.6147,21.740154,21.318316,21.04395,20.7833,20.567236,0.6276145,0.65162164,0.6893471,0.6893471,0.6824879,0.77508676,0.6824879,0.66876954,0.7339317,0.8128122,0.7510797,1.1008976,1.3203912,1.3855534,1.4232788,1.704505,1.8485477,2.1434922,2.0920484,1.7490896,1.7250825,1.845118,1.8176813,1.8519772,2.07833,2.5241764,2.2429502,1.9171394,1.9102802,2.1846473,2.3046827,3.0626216,4.2389703,5.521636,6.619104,7.239859,13.663476,15.758954,12.55915,6.3001523,2.4075704,1.5638919,1.9274281,1.8313997,1.1249046,1.196926,2.411,1.4404267,0.4424168,0.23321195,0.30523327,0.34638834,0.4046913,0.3806842,0.34981793,0.58302987,0.6790583,0.61046654,0.59674823,0.71678376,0.90198153,1.0871792,1.0871792,1.0254467,0.90198153,0.607037,0.5590228,0.5796003,0.5693115,0.52815646,0.58302987,0.75450927,0.823101,0.7579388,0.6927767,0.90541106,0.922559,0.9945804,1.1351935,1.155771,0.6790583,0.53501564,0.64476246,0.922559,1.1832076,1.1523414,0.72021335,0.32238123,0.106317215,0.09602845,0.19548649,0.274367,0.36353627,0.4664239,0.5693115,0.65505123,0.48357183,0.36696586,0.3566771,0.432128,0.47328308,0.41840968,0.5144381,0.58302987,0.5761707,0.5796003,0.4046913,0.3566771,0.45956472,0.61046654,0.59674823,0.47328308,0.53158605,0.6790583,0.77165717,0.607037,0.47671264,0.36696586,0.29151493,0.22978236,0.1371835,0.22635277,0.24350071,0.216064,0.15776102,0.072021335,0.037725464,0.024007112,0.020577524,0.024007112,0.030866288,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.020577524,0.017147938,0.010288762,0.010288762,0.01371835,0.01371835,0.020577524,0.041155048,0.05144381,0.044584636,0.05144381,0.17147937,0.2194936,0.216064,0.1920569,0.19548649,0.31895164,0.4115505,0.52815646,0.66191036,0.7407909,0.6207553,0.6756287,0.66191036,0.6859175,1.1900668,1.2586586,1.255229,1.0220171,0.69963586,0.72021335,0.71678376,0.82996017,0.97057325,1.1489118,1.4507155,1.4267083,2.020027,2.5824795,2.9254382,3.3472774,3.9337368,4.2423997,4.6608095,5.425607,6.6225333,7.2535777,7.7577267,8.580828,10.086417,12.555719,13.920695,14.760944,15.134769,15.055889,14.527733,13.924125,12.758065,11.303921,10.401938,11.451392,13.461131,14.493437,15.810398,17.689812,19.438902,22.20658,24.696459,27.741934,32.289566,39.375095,40.82924,39.80379,35.31446,28.67478,23.506393,20.985645,18.015623,16.45516,16.743246,17.919594,18.938183,20.604961,22.275171,23.739605,25.217756,27.254932,27.309805,24.19231,19.260563,16.400288,20.69413,22.669573,24.92624,29.662502,38.65488,47.24257,55.1169,63.114697,70.98217,77.37835,80.41697,80.17347,77.6973,74.08252,70.44716,59.42446,52.397236,45.72669,37.533405,27.690489,21.211998,15.71437,11.447963,8.381912,6.183546,5.7582774,5.638242,5.8474464,6.252138,6.557371,7.191845,8.285883,9.743458,10.813489,10.096705,11.327928,12.006986,12.103014,12.555719,15.285671,16.664366,18.598652,20.60839,20.958208,16.6335,12.730629,11.197603,10.6488695,9.750318,7.2021337,5.360445,3.724532,2.6647894,2.1332035,1.6530612,1.5398848,1.529596,1.9514352,2.7882545,3.673088,3.707384,3.6285036,3.5976372,3.707384,3.9954693,4.15323,4.1017866,3.9954693,3.8925817,3.758828,3.6799474,4.554492,6.142391,7.8503256,8.738589,8.635701,9.513676,10.113853,9.89436,9.026674,10.580277,10.710602,11.163307,12.895248,16.074476,19.085653,19.298288,20.179693,22.271742,23.18744,20.337454,18.324286,17.583494,17.12393,14.531162,11.375941,7.6274023,4.170378,1.6427724,0.432128,0.16804978,0.16119061,0.24007112,0.2777966,0.18862732,0.072021335,0.017147938,0.0,0.0,0.0,0.0,0.0,0.1920569,0.47671264,0.48357183,0.5624523,0.97057325,1.2415106,1.3889829,1.8828435,1.529596,2.9734523,4.846007,6.807731,9.541112,10.823778,9.928656,9.342196,10.542552,14.016724,12.024134,10.302481,10.31277,11.492548,11.276484,10.813489,10.302481,9.386781,8.045813,6.601956,4.7431192,4.170378,3.6044965,2.8396983,2.702515,2.5173173,2.603057,2.8465576,2.942586,2.4007113,3.1037767,2.983741,2.8911421,2.860276,2.0817597,2.3458378,2.5207467,2.9700227,3.5016088,3.3781435,3.2306714,3.0900583,2.620205,2.2258022,3.0454736,3.093488,4.0846386,4.3452873,3.8548563,4.2355404,3.789694,3.9543142,3.7553983,3.3815732,4.1772375,5.535354,6.111525,7.250148,9.14328,10.847785,9.304471,7.7851634,6.90033,6.464772,5.5079174,4.8837323,4.8185706,4.7362604,4.523626,4.5099077,4.033195,4.496189,5.288424,5.8371577,5.610805,6.869464,7.431916,7.1198235,6.5642304,7.2158523,7.8023114,8.656279,9.386781,9.781183,9.794902,9.626852,10.412228,11.766914,12.6929035,11.616013,11.125582,10.666017,10.696883,11.327928,12.312219,11.674315,11.413667,11.012405,10.710602,11.482259,11.506266,11.543991,11.55428,11.444533,11.039842,12.092726,12.6757555,13.166186,13.642899,13.900118,12.737488,12.408247,12.459691,12.610593,12.761495,12.247057,12.291641,11.262765,10.065839,12.161317,15.0456,11.245617,8.584257,11.159878,19.342873,29.724234,25.574434,19.109661,14.764374,9.211872,13.176475,11.029553,7.407909,8.23444,20.721567,19.95334,14.534592,8.1212635,3.8205605,4.1600895,4.1463714,3.6799474,3.5839188,3.7862647,3.3232703,2.4418662,2.1194851,2.0577524,2.0097382,1.8005334,1.4404267,1.2723769,1.313532,1.4198492,1.3032433,1.1797781,1.0631721,1.0425946,1.1420527,1.3306799,1.4781522,1.670209,1.7525192,1.7319417,1.7799559,1.5844694,1.196926,0.94999576,0.83681935,0.490431,0.48014224,0.39097297,0.26750782,0.15776102,0.12003556,0.11317638,0.35324752,0.6344737,0.8471081,0.9842916,1.4335675,1.2963841,1.08032,1.0425946,1.1797781,1.4541451,1.5330256,1.5158776,1.5158776,1.6667795,1.5158776,1.6530612,1.7799559,1.821111,1.9411465,1.8862731,2.037175,2.5378947,3.1106358,3.0489032,3.765687,4.396731,5.1340923,5.8543057,6.125243,5.919468,6.0395036,6.3035817,6.6293926,7.006647,7.9875093,9.016385,9.873782,10.803201,12.507706,14.747226,15.741806,15.803539,15.038741,13.344524,13.55373,14.699212,14.671775,13.519434,13.4474125,13.38911,13.437123,14.102464,14.96672,14.682064,13.9481325,11.996697,10.779194,10.799771,11.129011,12.360233,13.039291,13.152468,12.785502,12.099585,11.842365,12.487128,13.858963,15.066177,14.500296,12.63803,11.694893,11.30735,11.238758,11.399949,12.065289,11.4754,10.072699,8.697433,8.601405,8.779744,9.129561,9.784613,10.902658,12.672326,12.71691,11.965831,11.166737,10.967821,11.9040985,11.619442,12.397959,13.248496,13.982429,15.223939,16.163645,17.676094,18.680964,19.178253,20.272291,19.977346,21.006224,21.925352,22.326614,22.830763,21.78131,22.419212,23.931662,25.01884,23.866499,23.1943,23.334913,23.68473,23.911083,23.948809,24.789059,25.461258,25.643026,25.509272,25.708187,25.320644,26.082012,27.121178,27.625326,26.822803,26.668472,25.800787,24.456388,23.458378,24.233465,25.008553,25.663603,25.365229,24.319204,23.773901,23.643576,22.913074,22.065966,21.28402,20.460918,0.7099246,0.77851635,0.7922347,0.764798,0.72707254,0.7373613,0.67219913,0.6962063,0.7579388,0.7990939,0.7579388,1.1317638,1.1214751,1.1797781,1.3992717,1.5364552,1.5364552,1.7525192,1.8348293,1.7422304,1.7456601,2.054323,1.9514352,1.961724,2.177788,2.277246,1.9171394,1.8039631,2.054323,2.4452958,2.3972816,4.280125,4.90431,5.4187484,6.0840883,6.2692857,12.600305,15.107333,12.288212,6.210983,2.510458,1.4335675,1.587899,1.3889829,0.7305021,1.0014396,1.6324836,0.8779744,0.24350071,0.2469303,0.42183927,0.44584638,0.52472687,0.5007198,0.39783216,0.4389872,0.71678376,0.65505123,0.6344737,0.764798,0.864256,1.1008976,1.1660597,1.1420527,1.0323058,0.7613684,0.66876954,0.51100856,0.40126175,0.432128,0.6927767,0.84367853,0.7442205,0.6859175,0.86082643,1.3306799,1.1934965,1.0460242,0.97400284,0.91569984,0.65162164,0.5796003,0.7888051,1.0768905,1.2620882,1.196926,0.6276145,0.25378948,0.1371835,0.24007112,0.4355576,0.52815646,0.64133286,0.7099246,0.6962063,0.59331864,0.53501564,0.4972902,0.4938606,0.5144381,0.5041494,0.37039545,0.6207553,0.7990939,0.7407909,0.58302987,0.4389872,0.4389872,0.5693115,0.72707254,0.69963586,0.5144381,0.53844523,0.8128122,1.138623,1.0940384,0.85739684,0.5624523,0.30523327,0.1371835,0.06859175,0.09602845,0.12689474,0.12689474,0.10288762,0.082310095,0.037725464,0.037725464,0.072021335,0.12003556,0.16119061,0.13032432,0.072021335,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.037725464,0.0274367,0.017147938,0.01371835,0.01371835,0.017147938,0.017147938,0.034295876,0.041155048,0.05144381,0.061732575,0.06516216,0.1097468,0.1371835,0.11317638,0.07888051,0.15433143,0.26064864,0.42526886,0.58302987,0.6859175,0.6859175,0.5418748,0.6173257,0.64819205,0.78537554,1.6153357,1.0494537,0.7442205,0.65848076,0.64819205,0.42869842,0.6379033,0.77851635,0.90541106,1.0323058,1.1420527,1.371835,2.0646117,2.627064,2.9391565,3.340418,4.2595477,4.166949,4.383013,5.411889,6.924337,7.706283,8.31332,9.283894,10.998687,13.680624,15.323397,16.0539,15.96816,15.549749,15.676644,14.860402,13.210771,11.5645685,10.748327,11.595435,13.594885,14.277372,15.820687,18.245405,19.432043,22.161995,25.149164,28.619907,32.86231,38.22618,43.668938,42.739517,37.262466,29.638494,22.841053,21.047379,17.88873,15.570327,14.96672,15.638919,17.86815,20.172834,21.489796,22.179142,24.0174,23.160004,22.134558,19.857311,17.20281,16.997036,24.555847,24.830214,25.745913,30.979464,39.98556,46.244556,49.97252,53.566727,58.35443,64.56884,69.877846,72.22025,70.84156,66.43111,61.128967,56.553898,52.02684,44.591496,33.77458,21.568676,16.540901,12.315649,9.108984,6.835168,5.137522,5.1066556,5.6793966,6.5779486,7.5553813,8.388771,9.791472,10.611144,11.129011,11.605724,12.253916,12.905538,13.529722,13.992717,14.822677,17.195951,19.812727,22.12084,22.069395,19.270851,15.014734,11.814929,10.05898,8.80718,7.4113383,5.4804807,4.372724,3.875434,3.5187566,3.059192,2.4898806,1.9823016,1.8416885,2.1915064,3.069481,4.4516044,4.8837323,5.528495,6.135532,6.7219915,7.589677,8.018375,7.8366075,7.5107965,7.281014,7.157549,7.1061053,7.9600725,9.469091,11.146159,12.253916,13.615462,14.088745,14.003006,13.776653,13.896688,17.233677,17.089634,17.820137,20.272291,21.767591,18.560926,19.102802,20.015072,20.145397,20.553518,18.732407,18.53692,18.770132,18.180243,15.46744,9.709162,5.4907694,2.7093742,1.1317638,0.35324752,0.19891608,0.29151493,0.45613512,0.5453044,0.41840968,0.20234565,0.058302987,0.0,0.0,0.0,0.0,0.0,0.030866288,0.13032432,0.35324752,1.1420527,1.4610043,1.3203912,1.1420527,1.7730967,2.2429502,4.4516044,6.341307,7.366754,8.498518,9.736599,10.449953,10.858074,11.509696,13.262215,11.849225,11.646879,12.46312,13.419975,12.946692,13.018714,12.319078,11.05356,9.496528,7.9875093,5.0003386,3.8685746,3.3266997,2.702515,1.9068506,2.4452958,2.4007113,2.5961976,3.0557625,2.9871707,2.6167753,2.8088322,2.9185789,2.6990852,2.2978237,2.5001693,2.1674993,2.3492675,3.0454736,3.2306714,3.3472774,3.3850029,3.0729103,2.527606,2.2806756,3.2478194,4.9934793,5.3501563,4.6265135,5.6245236,5.5387836,5.3227196,4.57164,3.8205605,4.523626,6.914048,7.473071,7.956643,8.22758,6.2555676,5.4633327,6.5196457,7.4765005,7.1026754,4.8597255,4.4756117,4.605936,4.7362604,4.6745276,4.5270553,4.2183924,4.7534084,5.7754254,6.5779486,6.101236,7.239859,7.373613,7.0546613,6.917478,7.7028537,7.949784,8.7317295,9.290752,9.441654,9.544542,9.945804,10.323058,11.156448,12.085866,11.924676,10.868362,10.525404,10.792912,11.523414,12.517994,11.838936,11.598865,10.991828,10.374502,11.276484,10.360784,9.9801,10.38479,11.255906,11.742908,12.710052,12.850664,12.812939,12.850664,12.809509,12.082437,12.199042,12.72034,13.080446,12.600305,12.586586,12.370522,10.429376,9.040393,14.308239,15.9750185,12.147599,9.153569,9.445084,11.588576,19.696121,24.504402,21.304598,12.614022,8.189855,8.320179,6.701414,5.857735,8.272165,16.403717,18.259123,11.862943,5.597087,3.5804894,5.638242,4.57507,3.4810312,3.0729103,3.1792276,2.7093742,2.0165975,1.8554068,1.8656956,1.845118,1.7559488,1.5364552,1.3546871,1.3203912,1.3409687,1.1146159,1.097468,1.1592005,1.0768905,0.9568549,1.2243627,1.4027013,1.7010754,1.8108221,1.7010754,1.6359133,1.3443983,0.96714365,0.7682276,0.70649505,0.42869842,0.4629943,0.34981793,0.216064,0.1371835,0.10288762,0.12689474,0.274367,0.4938606,0.6893471,0.7099246,0.89855194,0.97400284,0.939707,0.89512235,1.0357354,1.214074,1.1694894,1.2415106,1.4610043,1.5741806,1.5364552,1.6324836,1.704505,1.704505,1.670209,1.6873571,1.9548649,2.5138876,3.1209247,3.2581081,3.7965534,4.386442,5.2438393,5.994919,5.693115,5.3878818,5.5833683,6.121814,6.697984,6.8557453,8.093826,9.139851,9.774324,10.401938,12.061859,14.160767,14.044161,13.536582,12.97413,11.211322,12.332796,13.687484,14.514014,14.733508,14.946142,13.87954,13.7697935,13.958421,14.023583,13.756075,14.003006,12.826657,11.955542,11.845795,11.688034,11.753197,12.778643,13.46799,13.128461,11.670886,11.0981455,12.401388,13.975569,14.733508,14.088745,12.336226,11.105004,10.525404,10.377932,10.103564,10.511685,10.127572,9.496528,9.132992,9.523964,8.961512,9.043822,9.8429165,11.115293,12.312219,11.965831,11.105004,10.316199,9.983529,10.268185,11.008976,12.6757555,13.972139,14.836395,16.46545,16.619781,17.412016,17.826996,18.03963,19.380598,19.147387,19.754423,20.382038,20.62554,20.512363,21.664703,23.334913,24.463247,24.295198,22.36434,22.336903,23.406935,24.09971,24.408375,25.780209,27.549875,27.495003,26.946268,26.661613,26.822803,27.18291,27.563595,28.153484,28.541027,27.711067,26.977135,26.171183,25.670462,25.382378,24.720467,25.859089,26.586163,26.033998,24.789059,24.878227,25.780209,24.77534,22.889067,21.102251,20.361462,0.7476501,0.84367853,0.8162418,0.7407909,0.6893471,0.70306545,0.5693115,0.58988905,0.70649505,0.8676856,1.039165,1.3924125,1.3443983,1.4027013,1.5707511,1.3272504,1.5364552,1.6427724,1.7525192,1.8931323,2.0131679,2.037175,1.9239986,1.8691251,1.8862731,1.8005334,1.7147937,1.8588364,2.1640697,2.4075704,2.2120838,6.6053853,6.5230756,5.7068334,5.802862,6.3790326,13.615462,16.973028,15.436573,9.870353,3.0351849,1.6942163,1.5124481,1.196926,0.59674823,0.7339317,0.91569984,0.5041494,0.20577525,0.23664154,0.33609957,0.4081209,0.53844523,0.5555932,0.47671264,0.48700142,0.5624523,0.4972902,0.6756287,1.0837497,1.3272504,1.1934965,1.1592005,1.1111864,1.0151579,0.9294182,0.66191036,0.5212973,0.5041494,0.64476246,1.0220171,0.99801,0.84367853,0.8093826,0.9877212,1.3443983,1.2449403,0.9842916,0.7990939,0.7510797,0.70306545,0.8711152,1.097468,1.313532,1.3306799,0.85396725,0.45270553,0.21263443,0.21263443,0.40126175,0.59674823,0.70649505,0.7133542,0.6962063,0.65162164,0.5178677,0.48357183,0.5658819,0.53501564,0.4046913,0.4424168,0.4046913,0.5418748,0.6036074,0.5212973,0.4115505,0.42526886,0.45613512,0.5041494,0.58988905,0.7476501,0.4664239,0.34295875,0.6276145,1.1900668,1.4953002,1.1900668,0.85739684,0.5521636,0.31209245,0.15090185,0.15090185,0.18862732,0.17833854,0.106317215,0.044584636,0.020577524,0.034295876,0.15090185,0.34638834,0.5041494,0.34638834,0.23321195,0.1097468,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.006859175,0.017147938,0.030866288,0.0548734,0.05144381,0.05144381,0.06516216,0.07545093,0.06516216,0.06859175,0.06859175,0.06859175,0.106317215,0.14404267,0.216064,0.37382504,0.61389613,0.8711152,0.980862,1.0528834,1.0048691,1.0048691,1.4815818,1.2003556,0.9568549,0.78537554,0.61389613,0.26064864,0.37039545,0.4424168,0.6310441,0.9328478,1.1900668,1.5570327,2.0406046,2.5893385,3.0729103,3.2821152,4.0606318,4.5853586,5.2575574,6.375603,8.131552,9.595985,10.703742,11.509696,12.21619,13.169616,14.54831,15.861842,16.407146,16.324837,16.616352,16.139639,14.949572,13.749216,12.80608,11.962401,13.2690735,14.867262,16.571766,18.159666,19.394318,22.456938,24.998262,27.875687,31.706535,36.8955,45.16081,46.03535,39.529427,29.312685,22.721018,19.315437,15.827546,13.330807,12.356804,12.895248,14.651197,15.374841,16.05733,17.401728,19.805868,18.355152,17.88873,16.194511,14.973578,19.8676,23.712168,24.737614,27.01486,32.16267,39.351086,43.34313,43.98446,46.049072,51.20374,58.0149,65.52227,70.49174,68.22821,59.712547,51.605003,54.228638,53.083157,42.694935,26.586163,17.274832,14.781522,11.928105,9.403929,7.589677,6.5162163,7.394191,7.953213,8.635701,9.89093,12.161317,14.832966,16.005884,16.335125,16.818697,18.78385,17.905876,18.471758,18.886738,19.161106,20.920483,20.711279,19.497204,17.86815,15.6869335,12.085866,10.597425,8.64942,6.7459984,5.079219,3.5393343,3.223812,3.875434,3.9680326,3.5290456,4.149801,2.976882,2.5481834,2.627064,3.2546785,4.746549,6.0635104,7.291303,8.615124,10.127572,11.825217,12.607163,12.699762,12.439114,12.13731,12.099585,12.586586,12.857523,13.862392,15.6697855,17.439453,19.857311,20.169403,20.340883,21.270302,22.796469,20.86904,22.638706,26.93941,29.285248,21.86705,19.984205,19.20569,19.456049,20.906765,23.972816,24.240324,25.653315,25.622448,22.484375,15.501736,8.251588,4.0674906,1.821111,0.6962063,0.18176813,0.14747226,0.26407823,0.45956472,0.61389613,0.5658819,0.3566771,0.12346515,0.0,0.0,0.0,0.0,0.0,0.0,0.08573969,0.42869842,1.587899,2.0886188,2.2086544,2.335549,2.9460156,3.9200184,7.0478024,9.589127,10.353925,9.719451,10.39165,11.657167,12.415107,12.493987,12.665466,13.361672,14.760944,15.059319,14.325387,14.496866,14.277372,13.780083,13.433694,12.843805,10.816919,7.363324,4.897451,3.4638834,2.8945718,2.8225505,2.1880767,2.3767042,2.609916,2.74367,3.2821152,2.5961976,2.5001693,2.4144297,2.2120838,2.2120838,2.1023371,1.9925903,2.3767042,3.0626216,3.1586502,2.7059445,2.7573884,2.7779658,2.8396983,3.6456516,3.9886103,4.064061,4.4241676,5.305572,6.636252,7.1369715,6.9071894,5.994919,5.120374,5.645101,7.257007,8.008087,7.9772205,7.1095347,5.219832,4.962613,5.785714,6.2864337,5.9228973,5.020916,3.7759757,4.0777793,4.3761535,4.184097,4.07435,4.5853586,4.5956473,5.0895076,6.245279,7.431916,8.090397,8.539673,8.673427,8.7283,9.277034,9.043822,9.654288,9.873782,9.55826,9.644,10.278474,10.545981,10.851214,11.238758,11.399949,11.30049,10.909517,10.683165,11.077567,12.542002,11.835506,11.749766,11.314209,10.518545,10.299051,9.530824,9.321619,9.9869585,11.204462,12.024134,12.120162,12.1921835,11.910957,11.317638,10.816919,10.696883,11.324498,12.38767,13.004995,11.732618,11.317638,11.334786,10.089847,8.718011,11.183885,13.601744,12.428825,10.549411,9.328478,8.621983,7.888051,23.424082,25.543568,11.756626,6.773435,5.518206,5.305572,4.588788,5.7822843,15.244516,19.150816,9.990388,3.7485392,4.9077396,6.468202,4.2218223,3.1415021,2.651071,2.503599,2.7470996,1.8691251,1.6667795,1.7388009,1.8142518,1.7559488,1.7902447,1.6359133,1.4644338,1.3101025,1.0528834,1.1146159,1.2037852,1.1900668,1.1626302,1.4198492,1.5913286,1.8348293,1.7353712,1.3306799,1.097468,1.0117283,0.8162418,0.70306545,0.65162164,0.4424168,0.41840968,0.33952916,0.26407823,0.21263443,0.15090185,0.16462019,0.29494452,0.42526886,0.490431,0.5041494,0.61389613,0.64133286,0.7133542,0.8505377,0.9602845,1.1694894,1.1111864,1.196926,1.4404267,1.4644338,1.3306799,1.4815818,1.5844694,1.5227368,1.3889829,1.3752645,1.7490896,2.4144297,3.234101,4.029765,4.0777793,4.170378,4.6402316,5.3261495,5.56965,5.521636,5.425607,5.8234396,6.6465406,7.233,7.8537555,8.779744,9.993818,11.417097,12.895248,14.88441,13.275933,12.343085,12.517994,10.405369,11.516555,12.80265,13.687484,14.016724,14.054449,14.493437,15.086755,14.819247,14.05102,14.527733,16.2974,15.741806,13.824667,11.492548,9.674867,11.321068,12.9707,14.191633,14.29452,12.329367,11.327928,12.624311,13.814379,14.003006,13.807519,11.917816,10.676306,10.316199,10.494537,10.299051,10.532263,10.618003,10.1481495,9.266746,8.683716,8.40249,8.577398,9.184435,10.014396,10.710602,10.748327,9.8429165,8.906639,8.450503,8.56025,10.209882,12.212761,14.363112,16.29397,17.501184,17.405157,17.947031,18.571217,18.941612,18.965618,19.795578,20.882757,21.596113,21.78474,21.757303,22.381487,24.10314,25.238335,24.85422,22.765602,22.436361,23.417223,24.717037,26.123167,28.198069,30.24896,30.111778,29.305824,28.506731,27.543016,27.44356,27.035439,27.004572,27.196629,26.610168,25.879667,26.016851,26.407824,26.579304,26.198618,26.407824,25.708187,25.135447,25.18346,25.817934,26.8571,25.804216,23.063976,20.237995,20.141968,0.7339317,0.823101,0.7407909,0.67219913,0.70306545,0.8128122,0.7373613,0.77851635,0.8505377,0.91227025,0.96371406,1.3478279,1.5193073,1.6427724,1.8313997,2.1332035,1.978872,1.8656956,1.8554068,1.978872,2.2086544,2.2738166,2.0234566,1.99602,2.2360911,2.277246,2.3458378,2.428148,2.301253,2.1126258,2.3458378,6.310441,5.9812007,4.955754,5.0929375,6.5367937,16.62664,20.234566,17.597214,10.72432,3.391862,1.9514352,1.7388009,1.4061309,0.66876954,0.30523327,0.32238123,0.20577525,0.15433143,0.2194936,0.29837412,0.36353627,0.36353627,0.38754338,0.432128,0.41498008,0.5453044,0.44584638,0.44584638,0.6824879,1.0837497,1.0563129,1.1523414,1.1626302,0.9877212,0.65162164,0.53844523,0.5761707,0.7476501,0.97400284,1.1077567,0.89855194,0.6927767,0.65162164,0.7922347,1.0014396,0.97057325,0.8505377,0.7305021,0.6790583,0.7373613,0.823101,1.0117283,1.1763484,1.155771,0.7579388,0.432128,0.2194936,0.1371835,0.17147937,0.29151493,0.40126175,0.48357183,0.4698535,0.3806842,0.33609957,0.45613512,0.490431,0.48357183,0.44927597,0.37039545,0.6173257,0.47328308,0.29494452,0.2469303,0.31552204,0.4424168,0.65848076,0.7888051,0.7510797,0.5418748,0.38754338,0.33609957,0.58988905,1.2209331,2.177788,2.6647894,2.2669573,1.6256244,1.0597426,0.5796003,0.39440256,0.28808534,0.19548649,0.09259886,0.020577524,0.006859175,0.01371835,0.041155048,0.1097468,0.2469303,0.3806842,0.37725464,0.2469303,0.07888051,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.006859175,0.017147938,0.017147938,0.034295876,0.041155048,0.048014224,0.048014224,0.05144381,0.06859175,0.07545093,0.11317638,0.16462019,0.14404267,0.15090185,0.20920484,0.40126175,0.6241849,0.58988905,0.9328478,0.7956643,0.72707254,1.0082988,1.6496316,1.0871792,0.881404,0.83338976,0.7442205,0.42869842,0.4046913,0.53844523,0.7373613,0.9431366,1.1420527,1.7799559,2.369845,2.750529,3.1209247,4.0606318,5.096367,6.358455,7.4010496,8.303031,9.671436,10.909517,11.814929,12.662037,13.601744,14.668345,15.258235,15.738377,16.12935,16.2974,15.944152,15.391989,15.059319,14.863832,14.733508,14.623761,16.009314,17.61779,18.938183,20.141968,22.127699,24.998262,28.18435,31.373867,34.882336,39.690617,47.71928,48.20285,40.63032,28.523878,19.411465,16.640358,13.3033695,10.799771,9.740028,9.962952,12.171606,13.519434,15.223939,17.902447,21.575535,20.522652,20.364891,20.36832,20.148827,19.682402,20.724997,23.681301,27.296087,31.617367,37.98611,43.675797,47.115673,50.38407,54.653904,60.18583,65.24447,77.36463,74.89876,58.141796,49.334614,52.338936,45.66496,33.116096,20.642687,16.307688,15.234227,13.186764,10.943813,9.102125,8.076678,8.255017,8.440215,8.477941,8.783174,10.329918,13.834956,15.234227,15.525743,16.194511,19.222837,20.306587,21.27716,23.557837,25.732195,23.557837,17.782412,17.549198,17.765263,15.618341,10.569988,8.868914,7.1026754,5.439326,4.0263357,2.9665933,2.7368107,3.2512488,3.7382503,3.940596,4.1120753,3.275256,2.8534167,2.8054025,3.1037767,3.7451096,5.2575574,7.390761,9.736599,12.085866,14.424845,16.280252,16.973028,16.935303,16.777542,17.288551,18.849012,20.522652,21.921923,23.520111,26.668472,26.887966,28.136335,29.18579,30.067194,32.059784,34.371326,35.85291,31.572783,23.297188,19.497204,22.11055,24.85422,24.874798,23.149715,24.497543,25.927681,25.420103,22.350622,17.069057,10.88894,6.2658563,3.3609958,1.611906,0.64819205,0.29151493,0.14061308,0.20577525,0.34981793,0.45613512,0.45613512,0.35324752,0.2503599,0.116605975,0.0,0.0,0.0,0.0,0.0,0.0274367,0.13375391,0.84367853,1.7147937,2.1743584,2.3458378,3.0557625,2.7813954,4.695105,7.596536,9.829198,9.294182,10.422516,11.173596,11.47197,11.7257595,12.836946,12.710052,13.972139,14.925565,15.055889,15.031882,13.865822,13.347955,13.512574,14.201921,15.066177,11.688034,8.14527,5.552502,4.0366244,2.7128036,2.2052248,2.7059445,2.668219,2.452155,4.307562,2.9185789,2.5721905,2.4384367,2.201795,2.054323,2.0303159,2.843128,3.2718265,3.1243541,3.2306714,2.819121,3.0420442,3.1483612,2.942586,2.7813954,4.0023284,4.091498,4.506478,5.586798,6.5642304,7.455923,7.7885933,7.5725293,7.1987042,7.438775,10.192734,9.523964,7.864044,6.4236174,5.206114,5.5833683,6.0635104,6.138962,5.7719955,5.3878818,3.758828,3.7313912,4.057202,3.99204,3.316411,4.4550343,4.540774,5.020916,6.2041235,7.2707253,8.069819,8.690575,9.023245,9.352485,10.350495,9.6817255,9.654288,9.589127,9.445084,9.801761,10.593996,10.233889,10.30934,11.008976,11.118723,11.146159,11.146159,11.105004,11.159878,11.592006,11.372512,11.091286,10.449953,9.637141,9.349055,8.375052,9.033533,10.48082,11.842365,12.21962,11.790922,11.362224,10.871792,10.31277,9.743458,9.836057,10.374502,11.0981455,11.454823,10.573419,9.613133,9.616563,11.101575,13.22106,13.773223,12.977559,12.363663,11.660598,10.398509,7.9120584,9.386781,22.957659,26.119738,15.371411,6.200694,6.341307,6.3207297,5.4667625,5.0929375,8.519095,17.754974,9.578837,3.2615378,4.420738,5.0174866,3.1312134,2.5927682,2.352697,2.201795,2.7573884,1.7147937,1.5433143,1.6427724,1.7490896,1.961724,1.7147937,1.5124481,1.2929544,1.0631721,0.89512235,0.89512235,1.0940384,1.1763484,1.1420527,1.3101025,1.4198492,1.4232788,1.2586586,1.0082988,0.90198153,0.8162418,0.66533995,0.5693115,0.5453044,0.5041494,0.42869842,0.39783216,0.32924038,0.28465575,0.45613512,0.29494452,0.31552204,0.40126175,0.45270553,0.4046913,0.5727411,0.72707254,0.8093826,0.864256,1.0220171,1.3169615,1.1866373,1.1832076,1.371835,1.3169615,1.1660597,1.1934965,1.1900668,1.1729189,1.3992717,1.4164196,1.8416885,2.534465,3.316411,3.9440255,4.0503426,4.1155047,4.633373,5.3981705,5.4976287,5.1821065,5.192395,5.504488,6.217842,7.5382333,8.618553,9.997248,11.64345,13.152468,13.711491,15.29939,14.126471,12.655178,11.760056,10.710602,11.218181,12.072148,12.987847,13.629181,13.625751,12.706621,13.138749,13.162757,12.507706,12.377381,13.581166,14.774663,15.107333,14.325387,12.751206,11.72233,12.641459,13.985858,14.579176,13.598314,12.744347,14.393978,15.12448,14.126471,13.200482,12.000127,10.251037,9.373062,9.527394,9.616563,10.14129,10.652299,10.624862,10.124143,9.791472,8.742019,8.64599,8.652849,8.625413,9.136421,10.268185,10.607714,10.381361,9.56512,7.8777623,8.862054,10.81006,13.344524,15.71094,16.780972,16.400288,16.732958,18.248835,20.152256,20.382038,20.217419,21.246294,22.408924,23.434372,24.84736,24.463247,24.4461,24.936531,25.334362,24.291767,24.312346,24.326063,25.632736,28.25637,30.955456,31.387585,31.58993,31.291555,30.475315,29.374416,29.247522,27.951138,27.045727,26.949697,26.93941,25.865948,26.812515,27.560165,27.254932,26.407824,26.428402,25.76992,24.933102,24.415234,24.706749,24.76848,24.346642,23.177153,21.510372,20.104242,0.6790583,0.7613684,0.7956643,0.7476501,0.66191036,0.66533995,0.69963586,0.8779744,0.8779744,0.764798,0.96371406,1.4953002,1.6770682,1.7936742,2.0063086,2.369845,2.352697,2.1469216,2.0577524,2.177788,2.369845,2.5790498,2.3424082,2.1674993,2.2155135,2.3046827,2.2669573,2.2669573,2.1503513,2.1126258,2.719663,5.206114,5.2164025,5.0140567,6.0326443,8.855195,18.598652,20.491785,15.786391,8.05953,3.2306714,2.527606,2.435007,1.8828435,0.82996017,0.26407823,0.17147937,0.106317215,0.11317638,0.16804978,0.19891608,0.3018037,0.2777966,0.30523327,0.4115505,0.45956472,0.45270553,0.432128,0.5178677,0.7099246,0.8848336,0.83338976,0.9328478,0.9362774,0.7442205,0.4046913,0.4355576,0.65162164,0.89512235,1.0151579,0.89169276,0.70649505,0.6173257,0.66533995,0.8162418,0.9431366,0.7990939,0.66876954,0.67219913,0.805953,0.94999576,1.0700313,1.1763484,1.2106444,1.1146159,0.83338976,0.45613512,0.23321195,0.12346515,0.10288762,0.14061308,0.25721905,0.31209245,0.34295875,0.37382504,0.40126175,0.39097297,0.36353627,0.4664239,0.59674823,0.4046913,0.5418748,0.37382504,0.1920569,0.116605975,0.12346515,0.26064864,0.6790583,1.0460242,1.1283343,0.8093826,0.5693115,0.4972902,0.5521636,0.939707,2.1297739,3.450165,3.673088,3.0351849,1.9891608,1.2072148,0.823101,0.52472687,0.29494452,0.13032432,0.034295876,0.01371835,0.006859175,0.006859175,0.020577524,0.072021335,0.16462019,0.33609957,0.4046913,0.33266997,0.21263443,0.12346515,0.061732575,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.006859175,0.010288762,0.01371835,0.01371835,0.020577524,0.024007112,0.030866288,0.041155048,0.0548734,0.06516216,0.06859175,0.09259886,0.14061308,0.17147937,0.14747226,0.16119061,0.23321195,0.33952916,0.40126175,0.69963586,0.6790583,0.7339317,1.0357354,1.529596,0.980862,0.7442205,0.6379033,0.5555932,0.4629943,0.4115505,0.5555932,0.8093826,1.0837497,1.313532,2.136633,2.8328393,3.426158,4.105216,5.2266912,6.310441,7.610255,8.721441,9.510246,10.127572,11.101575,11.934964,13.272504,14.942713,15.96816,16.681513,17.237106,17.288551,16.859852,16.362562,15.944152,16.05733,16.588915,17.350283,18.080786,19.586374,21.568676,23.35206,24.843931,26.510712,29.206367,31.898594,34.66284,38.31535,44.416588,48.353752,48.017654,39.683758,26.051146,16.259674,13.224489,10.460241,8.803751,8.200144,7.6925645,9.184435,11.050131,13.375391,16.63007,21.661274,20.409475,20.652975,21.53781,22.686722,24.19574,21.44864,24.17859,28.654203,34.052376,42.458294,51.131718,52.088573,52.56186,55.55589,59.84973,60.405323,63.059826,57.726818,45.80214,40.181046,40.805233,32.845158,23.091412,16.191082,14.640909,13.838386,12.63117,11.008976,9.108984,7.233,7.15069,6.9552035,6.495639,6.125243,6.6876955,8.594546,9.709162,10.4705305,11.948683,15.844694,22.158566,25.76649,25.721907,23.163433,21.304598,18.62266,18.145947,17.63151,15.419425,10.429376,8.107545,6.591667,5.2815647,3.9783216,2.867135,2.9322972,3.6216443,5.0620713,6.355026,5.586798,4.5682106,4.0606318,4.057202,4.4413157,4.976331,5.6245236,7.8263187,10.323058,12.71691,15.46058,17.388008,18.766703,19.689262,20.62897,22.43979,22.813616,23.753323,26.051146,29.59048,33.352737,32.965195,35.684856,38.46625,39.378525,37.601997,36.66229,34.00779,28.980015,23.928232,24.216316,25.752771,24.874798,24.230036,25.111439,27.44699,26.318655,21.410915,15.690363,10.950673,7.8023114,5.3158607,3.4844608,1.9685832,0.7922347,0.36696586,0.2777966,0.32238123,0.36010668,0.34638834,0.34638834,0.28465575,0.22292319,0.13032432,0.037725464,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.4115505,1.1832076,1.9857311,2.4795918,2.3321195,2.0303159,2.8294096,5.5559316,9.081548,10.31277,11.602294,11.667457,11.780633,12.9707,16.019604,15.697222,15.271953,14.123041,12.929544,13.684054,12.682614,12.6757555,12.991278,13.474849,14.490007,12.240198,8.738589,6.121814,4.8185706,3.5564823,3.216953,3.1037767,2.7470996,2.5001693,3.5290456,3.9200184,3.3644254,2.8122618,2.568761,2.287535,2.2463799,3.0317552,3.210094,2.7642474,3.0866287,2.6304936,3.1140654,3.666229,3.8891523,3.8445675,4.3692946,4.0537724,4.434457,5.826869,7.332458,8.879202,9.918367,10.007536,9.369633,8.89635,10.213311,8.886061,7.051232,5.6005163,4.170378,4.5442033,5.377593,5.5319247,4.976331,4.8014226,3.4981792,3.782835,4.187526,4.0949273,3.7313912,4.695105,5.051782,5.98463,7.257007,7.233,7.133542,8.049242,8.577398,8.697433,9.788043,9.575408,9.517105,9.379922,9.383351,10.189304,10.5597,9.832627,9.626852,10.192734,10.443094,10.731179,10.81006,10.967821,11.365653,12.010415,11.780633,11.122152,10.096705,9.1810055,9.256456,8.742019,9.547972,10.672876,11.434244,11.461681,10.950673,10.412228,9.928656,9.445084,8.769455,9.349055,9.990388,10.419086,10.497967,10.220171,9.369633,8.196714,8.652849,11.736049,17.487467,17.652086,15.841265,12.956982,10.065839,8.39563,9.301042,17.017612,19.167965,13.070158,5.7479887,7.1952744,8.025234,7.682276,7.2192817,9.297611,11.410237,7.2467184,3.8925817,3.4364467,2.9803114,2.5824795,2.5790498,2.2566686,1.7696671,2.1469216,1.670209,1.670209,1.7113642,1.670209,1.7388009,1.6427724,1.529596,1.4267083,1.2929544,1.0288762,1.039165,1.1146159,1.1832076,1.2346514,1.3375391,1.2003556,1.155771,1.1077567,1.0151579,0.881404,0.7613684,0.58302987,0.48357183,0.4698535,0.42869842,0.53844523,0.64476246,0.5693115,0.4355576,0.64476246,0.37725464,0.37382504,0.5041494,0.607037,0.4629943,0.5144381,0.6173257,0.71678376,0.86082643,1.1832076,1.3684053,1.1832076,1.0837497,1.2106444,1.371835,1.1626302,1.214074,1.1934965,1.138623,1.4404267,1.7593783,2.3218307,2.9117198,3.4810312,4.1772375,4.48933,4.530485,4.914599,5.5113473,5.442755,4.9523244,5.1580997,5.7822843,6.7871537,8.347616,9.764035,11.197603,12.517994,13.392539,13.282792,14.335675,13.855534,12.682614,11.629731,11.492548,11.605724,11.989838,12.812939,13.72178,13.838386,12.627741,13.149038,12.723769,11.026124,10.093276,10.751757,12.109874,12.9809885,12.956982,12.411677,11.087856,11.849225,12.926115,13.516005,13.780083,12.507706,12.991278,14.044161,14.5585985,13.522863,11.718901,10.611144,10.549411,11.204462,11.567999,11.653738,11.71547,11.777204,11.941824,12.377381,11.958971,11.619442,11.05356,10.336777,9.904649,11.0981455,11.598865,11.63659,10.950673,8.786603,9.06097,10.515115,12.579727,14.38369,14.760944,15.409137,15.512024,17.309128,20.11453,20.344313,20.910194,22.11398,24.226606,26.500422,27.148615,26.133457,25.4544,24.6896,23.849352,23.393215,24.000254,25.306927,26.651323,28.300955,31.463036,32.08036,31.2504,30.790836,31.109787,31.202387,30.461596,28.414133,27.080023,26.747353,25.989414,25.114868,25.444109,25.728765,25.43382,24.747904,25.330933,25.478405,24.696459,23.314335,22.487804,22.408924,22.470657,22.659285,22.491234,21.03023,0.6173257,0.7133542,0.78194594,0.7510797,0.6344737,0.5418748,0.6276145,0.84367853,0.8779744,0.7922347,1.0323058,1.4232788,1.5398848,1.6667795,1.903421,2.1743584,2.335549,2.294394,2.2635276,2.2978237,2.311542,2.6373527,2.4967396,2.2258022,2.1229146,2.4452958,2.3595562,2.2223728,2.1674993,2.5138876,3.7622573,5.7239814,5.892031,5.809721,7.040943,11.177026,18.217968,17.38115,11.530273,4.839148,2.7985435,2.4075704,2.1091962,1.4781522,0.6379033,0.2503599,0.17833854,0.13032432,0.1371835,0.17490897,0.18519773,0.32924038,0.33609957,0.32238123,0.34638834,0.4046913,0.39440256,0.44584638,0.58988905,0.7442205,0.7442205,0.6824879,0.6962063,0.6344737,0.45956472,0.22978236,0.3806842,0.6241849,0.823101,0.8676856,0.6824879,0.548734,0.5521636,0.64819205,0.78537554,0.881404,0.65505123,0.53158605,0.6173257,0.85739684,1.039165,1.2517995,1.3032433,1.2277923,1.0425946,0.7339317,0.39783216,0.2194936,0.1371835,0.10288762,0.09259886,0.23321195,0.26064864,0.31552204,0.4424168,0.5693115,0.4664239,0.41498008,0.5144381,0.65505123,0.51100856,0.47671264,0.31209245,0.15090185,0.061732575,0.041155048,0.274367,0.67219913,1.0117283,1.138623,0.97400284,0.7579388,0.66191036,0.64133286,0.91569984,1.9582944,3.923448,5.302142,5.079219,3.4981792,2.0920484,1.5261664,1.0185875,0.6310441,0.38754338,0.2469303,0.24350071,0.75450927,0.72707254,0.15776102,0.09602845,0.061732575,0.22978236,0.59674823,0.84024894,0.31209245,0.20577525,0.12003556,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.006859175,0.010288762,0.01371835,0.01371835,0.010288762,0.010288762,0.01371835,0.024007112,0.048014224,0.048014224,0.048014224,0.0548734,0.07888051,0.12689474,0.12003556,0.106317215,0.10288762,0.13375391,0.2469303,0.42183927,0.5007198,0.64133286,0.9362774,1.4267083,1.0288762,0.72364295,0.61046654,0.64133286,0.59674823,0.48700142,0.6859175,1.0288762,1.3924125,1.7216529,2.6304936,3.4947495,4.3658648,5.3227196,6.492209,7.2775846,8.128122,9.030104,9.856634,10.367643,11.036412,11.773774,13.334236,15.422854,16.684942,17.38115,17.905876,17.730967,17.051908,16.760393,16.815268,17.415445,18.650097,20.337454,22.03167,23.341772,26.198618,29.127487,31.161232,31.857437,34.138115,35.90435,37.48539,40.613174,48.415485,51.81078,50.2023,39.868954,24.315775,14.287662,10.371073,7.939495,7.051232,7.0546613,6.5813785,7.64798,9.72288,12.456262,15.923574,20.598103,20.186552,19.994495,20.687271,22.419212,24.833643,22.453508,25.77335,31.054914,37.385933,46.690403,56.478447,53.47756,50.46295,52.12973,55.072315,52.843082,47.866753,41.09675,34.43649,30.732533,28.311245,21.86362,16.341984,13.845244,13.6086035,13.279363,12.449403,10.871792,8.639131,6.138962,5.7239814,5.161529,4.506478,3.981751,4.0023284,4.8151407,5.4324665,5.994919,7.2947326,10.772334,19.274282,22.8582,22.913074,21.469217,21.187992,21.62012,21.61326,18.763273,13.701202,10.100135,7.473071,6.3001523,5.8680243,5.336438,3.7519686,3.3644254,4.033195,5.9812007,8.128122,8.107545,7.7611566,7.531374,7.2467184,7.116394,7.716572,7.8606143,9.023245,10.710602,12.771784,15.391989,17.37772,19.342873,21.500084,23.835632,26.119738,26.34266,26.236343,27.42984,30.272968,33.83974,35.053814,37.50597,40.987,43.428867,40.914978,40.513718,36.305614,31.58307,28.575323,28.458717,27.069735,24.216316,23.574984,25.632736,27.6802,23.475527,16.894148,11.159878,7.805741,6.64997,5.206114,3.923448,2.5584722,1.2586586,0.5693115,0.40126175,0.3566771,0.33266997,0.28808534,0.26407823,0.21263443,0.15776102,0.09602845,0.037725464,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.17490897,0.6824879,1.5501735,2.335549,2.1469216,1.7902447,1.8725548,3.7313912,7.421627,11.729189,12.895248,12.826657,12.950122,14.695783,19.473198,19.047928,17.247395,15.155347,13.762935,13.951562,11.516555,11.657167,11.825217,11.46854,12.006986,11.194174,8.790032,6.8728933,5.874883,4.5853586,3.9954693,3.3129816,2.935727,3.018037,3.4776018,4.8014226,3.9440255,3.000889,2.7162333,2.4658735,2.352697,2.884283,3.0317552,2.8122618,3.275256,2.8122618,2.9665933,3.666229,4.6127954,5.2918534,5.171818,4.547633,4.8151407,6.0566516,7.06495,9.527394,11.019264,10.926665,9.836057,9.523964,9.259886,8.200144,6.660259,5.055212,3.858286,4.32128,5.0174866,4.996909,4.3281393,4.0674906,3.6147852,4.0606318,4.396731,4.4241676,4.770556,5.686256,6.042933,6.9654922,8.032094,7.3050213,6.2247014,7.0786686,7.675417,7.6342616,8.371623,8.611694,8.7283,8.899779,9.342196,10.329918,10.360784,9.73317,9.613133,10.134431,10.401938,10.741467,10.868362,10.926665,11.173596,11.986408,11.825217,10.868362,9.654288,8.793462,8.934075,8.796892,9.637141,10.401938,10.573419,10.185875,9.736599,9.054111,8.752307,8.735159,8.196714,8.635701,9.167287,9.424506,9.373062,9.349055,9.355915,8.014946,6.5539417,8.2653055,18.492336,21.726437,18.903887,14.599753,12.0138445,12.984418,11.567999,12.871242,13.55373,11.835506,7.4970784,8.275595,9.225591,8.882631,8.193284,10.511685,8.508806,5.73427,3.5153272,2.3629858,1.9480057,2.0989075,2.294394,2.0508933,1.5673214,1.7216529,1.6873571,1.7216529,1.6976458,1.6427724,1.7456601,1.6427724,1.4953002,1.4472859,1.4232788,1.1249046,1.1351935,1.0871792,1.1180456,1.2209331,1.2380811,0.97400284,1.0597426,1.1077567,0.97400284,0.7476501,0.65505123,0.5144381,0.47328308,0.53501564,0.548734,0.6824879,0.77165717,0.6893471,0.52472687,0.5761707,0.4389872,0.4629943,0.5212973,0.5624523,0.59331864,0.7510797,0.66191036,0.64476246,0.85739684,1.2929544,1.3443983,1.1832076,1.1077567,1.2072148,1.371835,1.1934965,1.2415106,1.2415106,1.214074,1.5021594,2.2052248,2.8294096,3.3815732,3.9097297,4.506478,4.846007,5.144381,5.6142344,6.060081,5.892031,5.4633327,5.926327,6.992929,8.299602,9.421077,10.515115,11.592006,12.445972,12.723769,11.934964,12.586586,12.55915,11.945253,11.207891,11.194174,10.940384,11.177026,12.024134,13.05301,13.313659,12.991278,13.409687,12.734058,11.026124,10.251037,9.822338,10.446524,11.211322,11.581717,11.417097,10.635151,11.101575,11.537132,11.893809,13.368532,12.284782,11.55428,12.205902,13.54687,13.200482,11.2593355,11.101575,11.461681,11.8869505,12.723769,12.79922,12.466551,12.3533745,12.737488,13.567448,13.780083,13.365103,12.662037,11.873232,11.070708,11.842365,12.319078,12.686044,12.586586,11.129011,10.672876,11.396519,12.778643,14.033872,14.109323,15.004445,15.001016,16.647217,19.500635,20.111101,21.78131,24.027689,27.11089,29.460155,27.656193,26.496992,26.860529,25.85223,23.461807,22.573545,23.122278,25.258911,26.908543,28.01973,30.554195,31.133795,30.139215,29.484163,29.731094,30.098059,29.329832,27.618467,26.469557,25.9414,24.645016,24.27119,24.134007,23.797907,23.413794,23.739605,24.504402,24.981115,24.710178,23.626429,22.072824,21.78817,21.674994,22.052248,22.470657,21.705858,0.6379033,0.6859175,0.66876954,0.6379033,0.6001778,0.53501564,0.6173257,0.75450927,0.89512235,1.0082988,1.0940384,1.1523414,1.2758065,1.4507155,1.6599203,1.8588364,2.0920484,2.311542,2.3561265,2.2258022,2.0920484,2.4384367,2.4144297,2.194936,2.16064,2.8945718,2.7162333,2.4555845,2.4590142,3.1277838,4.914599,7.1849856,7.205563,6.461343,7.1266828,12.055,16.139639,13.107883,7.373613,2.6853669,2.1194851,1.4953002,0.85396725,0.4081209,0.20920484,0.17490897,0.20234565,0.22635277,0.25378948,0.28122616,0.30523327,0.42183927,0.47671264,0.4081209,0.28122616,0.31552204,0.45270553,0.5521636,0.6241849,0.66876954,0.6790583,0.64476246,0.53844523,0.4046913,0.2777966,0.17833854,0.39783216,0.51100856,0.5796003,0.607037,0.5521636,0.45956472,0.490431,0.5796003,0.67219913,0.72707254,0.5178677,0.45613512,0.5693115,0.805953,1.0254467,1.3032433,1.3238207,1.1866373,0.922559,0.490431,0.29837412,0.216064,0.17147937,0.13375391,0.09945804,0.26064864,0.31552204,0.36696586,0.48357183,0.7099246,0.70306545,0.67219913,0.64819205,0.6276145,0.5727411,0.5212973,0.32924038,0.15090185,0.07545093,0.14061308,0.53501564,0.6927767,0.7339317,0.75450927,0.8196714,0.7956643,0.7956643,0.91569984,1.2758065,2.0337453,3.940596,6.0395036,6.420188,4.9180284,3.1209247,2.5550427,2.0028791,1.546744,1.2209331,1.0082988,0.805953,1.9548649,1.9925903,0.78194594,0.5178677,0.41498008,0.40126175,0.8505377,1.3306799,0.5658819,0.32924038,0.1920569,0.08916927,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.006859175,0.01371835,0.017147938,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.0274367,0.024007112,0.0274367,0.030866288,0.034295876,0.041155048,0.08916927,0.07545093,0.08916927,0.13032432,0.13375391,0.20234565,0.26407823,0.38754338,0.67219913,1.2449403,1.0631721,0.78537554,0.764798,0.94656616,0.86082643,0.72707254,1.0220171,1.4095604,1.7833855,2.2566686,3.0454736,3.9714622,4.9488945,5.9640527,7.099246,7.517656,7.970361,8.604835,9.465661,10.508256,10.847785,11.543991,12.950122,14.853543,16.462019,16.825556,17.12736,17.175373,17.04162,17.072487,17.79613,18.972477,20.910194,23.465237,26.037428,27.35439,31.219534,35.10183,37.358498,37.25218,38.672028,39.31679,39.344227,41.56317,51.46096,59.156956,56.056606,42.29024,24.02426,13.46799,9.054111,6.677407,6.108095,6.684266,7.301592,8.971801,10.950673,14.081886,17.851004,20.388897,21.819035,20.172834,19.771572,21.45207,22.559826,24.624437,29.480734,35.444786,41.947285,49.523243,58.656235,52.945972,47.307728,46.98192,47.53408,44.666946,39.553432,33.65797,28.19121,24.096281,20.11453,16.359133,14.095605,13.526293,13.7697935,14.04759,12.898679,10.796341,8.237869,5.7479887,4.787704,3.9371665,3.3266997,3.0111778,2.9803114,3.9783216,4.3109913,4.15323,4.2938433,6.1321025,12.068718,13.29994,15.930434,20.4472,21.705858,22.727877,24.837072,20.807306,12.277924,9.72631,7.1987042,6.121814,6.3961806,7.010077,6.025785,4.98662,4.8014226,6.0806584,8.601405,11.324498,12.411677,12.926115,12.312219,11.293632,11.866373,12.13731,12.607163,13.790371,15.6526375,17.600643,18.468328,19.970488,22.2786,24.933102,26.829662,29.213226,29.487593,28.506731,28.208357,31.624226,34.055805,35.564823,38.877804,43.06876,43.524895,46.89618,44.852146,39.96841,34.443348,30.080912,27.18634,26.075153,26.119738,26.078583,24.11,18.11165,13.186764,9.716022,7.689135,6.7185616,5.3707337,4.197815,3.0557625,1.9308578,0.939707,0.5212973,0.30523327,0.23664154,0.23321195,0.20234565,0.14747226,0.09602845,0.044584636,0.0,0.0,0.0,0.010288762,0.010288762,0.0034295875,0.01371835,0.09945804,0.37039545,0.9877212,1.8073926,2.3767042,1.8897027,1.8348293,2.8122618,5.8405876,12.370522,13.649758,14.040731,14.349394,15.858413,20.337454,20.364891,18.718689,17.765263,17.54234,15.769243,10.278474,9.952662,9.956093,9.050681,9.585697,9.8429165,8.844906,7.720001,6.742569,5.3261495,4.4927597,3.6765177,3.4981792,4.029765,4.7979927,5.2815647,4.2526884,3.1586502,2.644212,2.5138876,2.3561265,2.6853669,3.0043187,3.1792276,3.4467354,3.3747141,2.9494452,3.2958336,4.5819287,6.0223556,6.0497923,5.754848,6.138962,6.9037595,6.4373355,9.22902,10.587136,10.199594,9.122703,9.788043,8.882631,8.100685,6.5950966,4.8768735,4.839148,5.1683884,5.127233,4.6882463,4.081209,3.7794054,4.201245,4.355576,4.6265135,5.120374,5.686256,6.8557453,6.989499,7.4113383,7.9943686,7.157549,5.785714,6.228131,6.7974424,6.924337,7.15069,7.39762,7.706283,8.399059,9.383351,10.168727,10.206452,10.096705,10.323058,10.840926,11.094715,11.2250395,11.30735,11.05356,10.738038,11.190743,11.201033,10.161868,9.040393,8.385342,8.309891,8.186425,8.999237,9.592556,9.458802,8.759167,8.330468,7.490219,7.377043,7.8983397,7.723431,7.689135,7.953213,8.213862,8.272165,8.008087,8.872343,8.491658,6.0840883,5.6176643,15.789821,21.44521,19.03078,15.6869335,15.371411,18.852442,15.1862135,11.814929,11.701753,13.145609,9.770895,9.084977,9.609704,8.659708,7.1884155,9.764035,9.623423,5.8817425,2.6064866,1.529596,2.0474637,1.6221949,1.7422304,1.7559488,1.5707511,1.6564908,1.7319417,1.6256244,1.5536032,1.6633499,2.0406046,1.6839274,1.3855534,1.2929544,1.3032433,1.0871792,1.097468,1.0254467,1.0460242,1.1454822,1.1077567,0.8711152,1.1008976,1.1146159,0.77851635,0.5212973,0.548734,0.53501564,0.59331864,0.71678376,0.7956643,0.7682276,0.7476501,0.69963586,0.6001778,0.44927597,0.4938606,0.5693115,0.48357183,0.37382504,0.70306545,1.1763484,0.864256,0.6379033,0.83681935,1.2860953,1.3066728,1.2277923,1.2380811,1.3238207,1.255229,1.138623,1.1489118,1.1934965,1.2998136,1.611906,2.6853669,3.2443898,3.806842,4.4447455,4.8117113,4.99005,5.717122,6.4579134,6.8557453,6.742569,6.615674,7.1987042,8.443645,9.863494,10.532263,10.7757635,11.149589,11.382801,11.180455,10.203023,10.683165,10.703742,10.477389,10.113853,9.623423,9.156999,9.609704,10.487679,11.355364,11.825217,12.836946,13.049581,12.63117,12.085866,12.260776,10.906088,10.429376,10.7586155,11.338216,11.125582,10.81006,10.700313,10.432805,10.607714,12.79922,12.504276,11.396519,11.067279,11.701753,12.085866,10.899229,11.4033785,11.369082,10.796341,11.907528,12.46312,12.3533745,12.157887,12.271064,12.895248,13.399398,13.1593275,12.655178,12.157887,11.712041,12.267634,12.860953,13.454271,13.869251,13.786942,13.001566,12.88839,13.601744,14.682064,15.031882,15.193072,15.313108,16.770683,19.154245,20.251715,22.721018,26.18147,29.67279,30.976034,26.630747,25.951689,28.084892,27.851679,24.734184,22.844482,23.142857,25.005123,26.925692,28.27352,29.295536,29.305824,29.072613,28.328392,27.357819,26.980564,26.634176,25.979126,25.378946,24.77534,23.69845,23.643576,23.653864,23.242313,22.981665,24.511261,24.789059,25.049707,25.26577,25.063425,23.743034,22.899355,22.271742,21.908205,21.819035,21.956219,0.8711152,0.6756287,0.6241849,0.5590228,0.47328308,0.53501564,0.70649505,0.78537554,0.91912943,1.0666018,1.0082988,1.1180456,1.4918705,1.7113642,1.7353712,1.9068506,2.2841053,2.3904223,2.194936,1.9068506,1.9685832,2.2978237,2.3252604,2.253239,2.452155,3.4776018,2.6373527,2.4452958,2.760818,3.4981792,4.6093655,5.8165803,5.861165,5.2644167,5.8543057,10.772334,14.983868,12.428825,6.8557453,1.8897027,1.0220171,0.6207553,0.34638834,0.23664154,0.23664154,0.19891608,0.23664154,0.37382504,0.45613512,0.4629943,0.48700142,0.4389872,0.5178677,0.48357183,0.37382504,0.53501564,0.6790583,0.8711152,0.84367853,0.65505123,0.71678376,0.6310441,0.45613512,0.32581082,0.3018037,0.34981793,0.51100856,0.48357183,0.3806842,0.29494452,0.31895164,0.39440256,0.4938606,0.6241849,0.70306545,0.5796003,0.42183927,0.40126175,0.5521636,0.85396725,1.2209331,1.4404267,1.3958421,1.1934965,0.89512235,0.5041494,0.37039545,0.30866286,0.26064864,0.19891608,0.1371835,0.26064864,0.40126175,0.45613512,0.48014224,0.6859175,0.9431366,0.97057325,0.8711152,0.6962063,0.42869842,0.548734,0.4698535,0.30523327,0.21263443,0.39783216,0.7510797,0.70306545,0.5727411,0.5144381,0.5041494,0.61389613,1.0151579,1.371835,1.7147937,2.4727325,2.8396983,3.415869,4.091498,4.5030484,4.012617,3.9165888,3.806842,3.5530527,3.1689389,2.8396983,1.7388009,2.2600982,2.6887965,2.3492675,1.6187652,1.5433143,1.3889829,1.2037852,1.1660597,1.5570327,0.7510797,0.3841138,0.19548649,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.010288762,0.006859175,0.030866288,0.006859175,0.010288762,0.010288762,0.0034295875,0.01371835,0.0034295875,0.017147938,0.037725464,0.041155048,0.030866288,0.116605975,0.09259886,0.12346515,0.19548649,0.12346515,0.12346515,0.19548649,0.2503599,0.30523327,0.48700142,0.59674823,0.67219913,0.6962063,0.7613684,1.0666018,1.2277923,1.5501735,1.8073926,2.0646117,2.6853669,2.9665933,3.4227283,4.170378,5.096367,5.830299,6.4990683,7.473071,8.176137,8.724871,9.932085,9.921797,10.960961,12.343085,13.690913,14.983868,15.388559,16.13621,17.182234,18.132229,18.279701,19.46291,20.923914,23.36578,26.59988,29.539038,32.471333,36.56283,39.65289,41.048733,41.549454,41.525444,40.623463,39.498558,42.122192,55.77195,67.782364,63.471375,45.97705,24.185452,12.710052,9.89093,7.8949103,7.4113383,8.522525,10.696883,14.016724,15.806969,19.524641,24.209457,24.490685,27.052586,23.492674,21.702429,24.161444,27.906553,33.14353,37.766617,43.768394,50.510963,54.746506,64.77119,59.27356,51.663307,47.105385,42.540604,38.25705,33.369884,28.314674,23.61957,19.898466,18.053349,16.386568,15.090185,14.466,14.891269,14.428274,12.315649,10.010965,7.9909387,5.7822843,4.355576,3.3678548,2.7745364,2.469303,2.2738166,3.3472774,4.1463714,4.2218223,3.8479972,4.0434837,5.5593615,7.6651278,8.838047,9.657719,12.816368,15.443433,21.225718,21.767591,16.194511,11.153018,8.628842,6.677407,5.6828265,6.4064693,9.993818,10.1652975,7.507367,6.475061,9.102125,14.997586,16.719238,18.221397,18.28313,17.432592,17.943602,18.091074,21.404055,25.029129,27.42984,28.379837,23.633287,21.904776,21.04395,20.838173,23.009102,29.113768,32.845158,32.99263,32.27242,37.337917,34.800022,39.097298,43.614063,45.757557,46.96477,44.97561,44.65323,42.90071,38.551994,32.365017,32.19354,31.902023,32.24498,30.34499,19.713268,13.612033,9.678296,7.7440085,7.034084,6.1801167,4.8734436,3.8685746,3.1380725,2.452155,1.4027013,0.82996017,0.42183927,0.18862732,0.10288762,0.09259886,0.06859175,0.024007112,0.0,0.0,0.0,0.0,0.0548734,0.0548734,0.0,0.0,0.24350071,0.37725464,0.65162164,1.0700313,1.3889829,1.8759843,2.311542,3.9200184,7.0135064,10.957532,13.581166,14.417986,15.103903,15.88242,15.6252,18.104792,18.732407,18.897026,18.406595,15.488017,8.004657,7.0135064,7.3050213,7.143831,8.255017,8.56025,7.8777623,6.7974424,5.861165,5.56965,5.8508763,5.1512403,4.8940215,5.470192,6.2247014,5.627953,5.0929375,4.105216,2.952875,2.7470996,2.6373527,2.6545007,2.8088322,2.860276,2.335549,3.690236,3.789694,3.5393343,3.799983,5.3878818,6.217842,7.438775,8.800322,9.599416,8.697433,9.517105,9.866923,9.904649,10.069269,11.094715,10.22703,7.7577267,5.518206,4.8288593,6.4990683,5.120374,4.729401,4.3692946,3.9646032,4.3178506,4.804852,4.40702,5.144381,6.526505,5.5387836,6.711703,6.931196,7.2295704,7.425057,6.118384,5.7651367,5.9331865,6.5367937,7.2364297,7.431916,7.298162,7.8126,8.7283,9.654288,10.069269,10.302481,10.871792,11.043272,10.97468,11.718901,11.585147,11.101575,10.840926,10.871792,10.789482,10.542552,9.630281,8.673427,8.1384115,8.347616,8.06639,8.23444,8.241299,7.905199,7.4765005,6.989499,6.427047,6.2075534,6.3447366,6.4544835,7.1129646,7.4627824,7.9429245,8.31332,7.630832,7.750868,7.5450926,6.012067,5.4016004,11.201033,15.2033615,15.114192,14.249936,14.71636,17.425734,14.225929,9.170717,9.585697,12.994707,7.1095347,8.405919,9.72631,8.577398,6.5539417,9.338767,7.4936485,6.6396813,4.2355404,1.2037852,1.937717,1.5227368,1.7388009,1.7079345,1.3752645,1.5090185,1.7902447,1.5673214,1.4472859,1.6633499,2.0920484,1.6153357,1.3409687,1.2346514,1.196926,1.039165,1.1489118,1.1214751,1.1797781,1.3409687,1.3889829,1.0837497,1.1729189,1.0117283,0.59674823,0.53501564,0.71678376,0.84367853,0.91227025,0.881404,0.6859175,0.6859175,0.8162418,0.91227025,0.89855194,0.77851635,0.5590228,0.6859175,0.6756287,0.5178677,0.70306545,1.2620882,0.8711152,0.5693115,0.7476501,1.1763484,1.3821237,1.3066728,1.2380811,1.2415106,1.1454822,0.91227025,0.96371406,1.1420527,1.4027013,1.8313997,3.2478194,3.7005248,4.0606318,4.616225,5.0826488,5.2266912,6.0532217,6.776865,7.1198235,7.2775846,7.582818,7.750868,8.4093485,9.736599,11.458252,11.118723,10.583707,9.410788,8.2481575,8.834618,9.287323,9.115844,8.81747,8.512236,7.949784,7.8777623,8.608265,9.091836,9.31133,10.299051,11.495977,12.041282,12.048141,11.921246,12.360233,12.22648,10.652299,9.781183,10.30934,11.506266,11.297061,10.72432,10.302481,10.63858,12.421966,12.360233,12.0138445,11.928105,12.000127,11.4754,11.012405,11.526843,11.159878,10.028113,10.2236,10.710602,11.592006,12.05843,12.055,12.298501,13.495427,13.684054,13.121602,12.298501,11.931535,13.29994,13.896688,13.780083,13.615462,14.678635,14.802099,13.780083,13.642899,14.654627,15.289101,15.412566,15.981877,17.775553,20.069946,20.62897,23.595562,26.44212,29.072613,29.85113,25.6053,26.178041,28.225504,28.187778,25.725336,23.712168,25.348082,27.296087,28.5959,29.000591,28.976585,29.329832,28.630196,27.556736,26.713057,26.627317,25.721907,25.149164,24.751333,24.37065,23.835632,23.211449,23.321196,24.120289,25.402954,26.795366,26.466127,27.059444,26.644464,25.303495,25.145735,23.705309,23.393215,22.78275,21.980227,22.628418,0.7099246,0.5144381,0.4972902,0.48357183,0.45956472,0.5590228,0.72021335,0.83338976,0.9328478,1.039165,1.1523414,1.3032433,1.5124481,1.5947582,1.6084765,1.8588364,1.9137098,2.020027,2.136633,2.2429502,2.335549,2.194936,1.9445761,2.0131679,2.3389788,2.369845,2.7573884,3.1415021,3.3541365,3.6593697,4.7774153,6.046363,5.2781353,4.7602673,7.449064,16.997036,22.467228,17.477179,9.15014,2.6545007,1.1934965,0.70306545,0.5007198,0.5041494,0.6276145,0.7956643,0.8025235,0.6927767,0.6001778,0.59331864,0.64819205,0.5007198,0.5555932,0.5693115,0.5418748,0.7305021,0.7579388,0.7373613,0.7476501,0.7888051,0.7888051,0.75450927,0.66876954,0.6207553,0.6276145,0.65505123,0.5521636,0.40126175,0.34295875,0.37382504,0.37039545,0.4115505,0.41840968,0.4355576,0.45613512,0.42183927,0.36010668,0.4081209,0.5727411,0.86082643,1.2449403,1.2003556,1.1832076,1.0117283,0.67219913,0.31895164,0.23664154,0.18519773,0.12689474,0.07545093,0.11317638,0.35324752,0.5212973,0.5761707,0.59674823,0.78537554,0.85396725,0.83681935,0.8848336,0.91227025,0.5727411,0.5007198,0.5418748,0.6207553,0.6859175,0.7133542,0.66876954,0.53501564,0.35324752,0.24007112,0.39440256,0.77851635,1.2037852,1.4267083,1.5193073,1.8862731,1.7936742,1.8142518,2.386993,3.3747141,4.0846386,4.5339146,6.2487082,7.6616983,7.671987,5.6348124,2.836269,2.0406046,2.2360911,2.9048605,4.0091877,3.974892,4.064061,3.7211025,2.901431,2.0817597,1.5981878,0.83681935,0.30866286,0.13032432,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0034295875,0.0,0.006859175,0.0,0.010288762,0.010288762,0.0,0.0034295875,0.010288762,0.017147938,0.024007112,0.030866288,0.017147938,0.044584636,0.041155048,0.14061308,0.2709374,0.15776102,0.13032432,0.22292319,0.2709374,0.25378948,0.32924038,0.5453044,0.72021335,0.8848336,1.0734608,1.2998136,1.3992717,1.6564908,1.9925903,2.3321195,2.6133456,2.7162333,3.1209247,3.724532,4.461893,5.2918534,6.608815,7.3530354,7.8263187,8.2653055,8.848335,9.637141,10.590566,11.434244,12.236768,13.423406,14.616901,15.769243,16.726099,17.514904,18.351723,20.28944,22.998814,26.215767,29.902573,34.241,38.438816,42.496017,45.301422,46.203403,45.016766,42.598907,39.72834,38.33593,42.969303,60.786007,77.01824,72.93361,53.563297,30.221525,20.484926,20.45063,19.332584,17.974468,16.767254,15.638919,16.654078,18.118511,21.69557,26.147175,27.333813,24.02083,21.963078,22.933651,27.416122,34.621685,39.742058,46.261703,56.718517,68.632904,74.4975,77.909935,67.55944,57.6205,51.766193,43.175076,37.211025,31.970613,27.038868,23.002243,21.44864,20.971928,17.902447,15.717799,15.117621,14.003006,14.102464,11.797781,9.513676,7.840037,5.501058,3.974892,3.1106358,2.6647894,2.486451,2.5070283,3.5804894,4.1155047,4.280125,4.3041325,4.4721823,4.7842746,7.164408,10.690024,18.993055,40.270218,21.19485,18.025911,16.098484,11.746337,12.30193,10.203023,7.922347,6.0635104,5.2747054,6.2487082,5.3844523,5.6828265,8.467651,12.507706,13.999576,15.63206,21.843042,25.9414,26.277498,26.243204,21.565247,27.02858,28.887415,25.430391,26.977135,24.182022,24.576424,26.27064,27.378397,26.02371,29.443008,32.255272,36.206154,39.766068,38.130154,41.840965,45.273983,48.031372,49.279743,47.736427,47.660976,47.623253,44.80413,39.779785,36.549114,38.438816,38.613724,35.83233,29.048605,17.418875,11.989838,8.3922,6.307011,5.1855364,4.262977,3.474172,2.9082901,2.4144297,1.9102802,1.3786942,0.9911508,0.61389613,0.32238123,0.1371835,0.017147938,0.01371835,0.0034295875,0.0,0.0,0.0,0.07888051,0.058302987,0.024007112,0.024007112,0.072021335,0.4938606,0.89169276,1.039165,1.1351935,1.8039631,2.7711067,3.5221863,5.874883,8.985519,9.345626,10.7586155,11.05356,11.598865,12.195613,11.06042,13.087306,13.612033,14.225929,14.788382,13.413116,8.742019,7.5382333,7.023795,6.5024977,7.3393173,7.157549,6.9723516,6.3961806,5.6142344,5.3981705,6.1766872,5.778855,4.619654,3.9165888,5.689686,5.6965446,5.2472687,4.6745276,4.016047,3.0283258,2.8980014,2.6922262,2.8534167,3.2512488,3.175798,3.5839188,3.6387923,3.6627994,3.923448,4.6402316,5.6965446,7.963502,10.281903,11.523414,10.600855,9.80862,9.9698105,9.410788,8.522525,9.764035,8.093826,5.6519604,3.9165888,3.5359046,4.338428,4.0846386,4.331569,4.3349986,4.0777793,4.307562,5.195825,5.1512403,5.768566,6.7631464,5.977771,6.094377,6.7700057,7.4044795,7.425057,6.2658563,5.675967,5.909179,6.759717,7.747438,8.128122,8.244728,8.577398,9.163857,9.80862,10.045261,9.908078,10.340206,10.624862,10.6488695,10.926665,11.338216,11.022695,10.861504,10.871792,10.203023,10.024684,9.482809,8.745448,8.162418,8.272165,8.1384115,7.9772205,7.723431,7.2775846,6.4887795,6.0875177,5.453044,5.188966,5.456474,5.967482,6.509357,6.869464,7.2878733,7.8331776,8.399059,7.671987,7.2432885,6.0052075,5.669108,10.786053,13.323947,12.699762,11.917816,11.55428,9.770895,14.599753,12.788932,11.790922,12.542002,9.441654,9.914937,10.930096,10.933525,9.904649,9.338767,6.5882373,4.232111,2.2738166,1.2517995,2.218943,1.5604624,1.7147937,1.9445761,1.8965619,1.6187652,1.5707511,1.4815818,1.5261664,1.6942163,1.7971039,1.6839274,1.4267083,1.3306799,1.3752645,1.2072148,1.0631721,1.0460242,1.1797781,1.3615463,1.3512574,1.2517995,1.1660597,0.9431366,0.70306545,0.8265306,0.922559,0.9328478,0.97057325,0.97400284,0.7099246,0.7510797,0.6962063,0.67219913,0.7305021,0.8505377,0.6310441,0.66533995,0.7442205,0.75450927,0.65162164,1.155771,1.1008976,0.9294182,0.8848336,1.0288762,1.2346514,1.1592005,1.0940384,1.1454822,1.2415106,0.89169276,0.9534253,1.1592005,1.4610043,2.0131679,3.2821152,3.9440255,4.3761535,4.787704,5.2026844,5.086078,5.501058,6.1492505,6.7631464,7.1061053,7.548522,7.936065,8.477941,9.242738,10.151579,10.093276,9.829198,8.906639,7.949784,8.652849,9.434795,8.958082,8.333898,7.956643,7.5210853,7.654839,8.06296,8.423067,8.796892,9.626852,10.161868,9.949233,9.685155,9.705732,9.9801,10.714031,10.106995,9.102125,8.755736,10.237319,10.134431,9.616563,9.860064,10.943813,11.845795,12.157887,12.123591,12.068718,11.934964,11.303921,11.317638,11.7257595,11.526843,11.032983,11.88352,13.193623,13.745787,13.416546,12.572867,12.055,13.125031,13.72178,13.443983,12.744347,12.932974,14.280802,14.668345,14.2362175,13.529722,13.505715,13.042721,12.511135,12.874671,14.267084,15.995596,16.208231,15.978448,16.37285,17.62122,19.140528,19.401176,22.336903,25.282919,26.332373,24.308916,26.445549,27.903124,27.697348,26.411253,26.215767,27.234354,27.337242,27.591032,28.390125,29.439579,29.480734,28.661062,27.577312,26.459267,25.173172,24.758192,24.936531,25.732195,26.404394,25.457829,24.055126,22.724447,23.180582,25.207468,26.647894,27.285797,27.549875,26.582733,24.84736,24.120289,25.111439,25.169743,24.624437,23.959099,23.825344,0.7339317,0.5693115,0.5521636,0.5624523,0.5590228,0.61046654,0.72364295,0.864256,1.0048691,1.1420527,1.2723769,1.4678634,1.5673214,1.5055889,1.4747226,1.9102802,1.7765263,2.0680413,2.2909644,2.2738166,2.16064,2.0646117,1.8725548,1.8999915,2.1126258,2.1263442,2.867135,3.4810312,3.82399,4.262977,5.672538,5.7479887,4.99005,6.186976,11.451392,22.254593,25.008553,19.250275,10.964391,4.417309,2.170929,1.0425946,0.6276145,0.5590228,0.6001778,0.64476246,0.7990939,0.7888051,0.72364295,0.67219913,0.66876954,0.5555932,0.65162164,0.65848076,0.58988905,0.77851635,0.9602845,1.371835,1.8828435,2.0886188,1.3203912,1.2106444,1.0323058,0.8471081,0.69963586,0.61389613,0.4355576,0.33609957,0.33609957,0.39783216,0.4355576,0.40126175,0.36696586,0.37039545,0.39783216,0.4081209,0.33609957,0.41840968,0.58302987,0.77851635,0.9945804,0.89855194,0.84024894,0.6927767,0.44927597,0.20234565,0.20234565,0.20234565,0.18862732,0.18176813,0.24350071,0.42526886,0.66191036,0.7613684,0.7339317,0.8093826,0.8471081,0.7613684,0.72021335,0.6893471,0.40126175,0.490431,0.548734,0.66876954,0.7956643,0.7099246,0.65162164,0.5727411,0.41498008,0.31552204,0.61389613,1.0734608,1.4644338,1.6324836,1.6530612,1.8416885,2.095478,2.16064,2.527606,3.3301294,4.341858,5.2506986,7.0786686,9.462232,10.515115,6.81802,3.7485392,2.4590142,1.9480057,2.0303159,3.3369887,7.0375133,7.099246,6.23156,5.254128,3.0900583,2.5790498,1.6736387,0.89512235,0.45613512,0.274367,0.16462019,0.09259886,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.01371835,0.01371835,0.017147938,0.020577524,0.01371835,0.020577524,0.08573969,0.19891608,0.274367,0.16804978,0.14747226,0.20234565,0.24007112,0.28808534,0.48357183,0.6824879,0.8265306,0.99801,1.2723769,1.7147937,1.7113642,2.037175,2.4247184,2.7711067,3.1449318,3.0866287,3.4638834,3.9954693,4.636802,5.586798,6.866034,7.442205,7.966932,8.663138,9.325048,9.801761,10.55284,11.578287,12.761495,13.862392,15.745236,16.46545,17.069057,18.022482,19.20569,22.580404,25.663603,29.552755,34.631973,40.55144,45.442036,49.286602,51.9754,52.736767,50.168007,44.985897,40.705772,41.100178,49.46837,68.643196,87.99979,83.99746,63.17643,38.462822,29.141205,33.966633,37.770046,39.038994,37.574562,34.470783,33.66483,33.325302,35.681427,39.00813,37.612286,29.17893,29.75167,32.450756,35.605976,42.74638,49.557537,61.0398,78.78105,96.60462,100.603516,84.78969,65.22047,52.932255,48.94707,44.258827,36.110126,30.029469,25.224615,22.011093,21.825895,20.930773,17.741257,16.167076,16.427725,15.05246,14.503725,12.212761,9.685155,7.7542973,6.5950966,4.7362604,3.8788633,3.542764,3.4776018,3.6525106,4.537344,4.513337,4.4859004,4.8494368,5.4941993,6.6396813,8.56025,12.830087,20.62554,32.707977,28.228935,20.800447,15.868701,14.54831,13.622321,10.659158,7.7542973,5.7102633,4.822,4.863155,5.0277753,5.751418,7.5553813,10.028113,11.814929,15.405707,20.766151,22.793037,21.963078,24.346642,20.015072,21.928782,23.098272,22.429502,24.703318,24.895376,24.295198,24.542128,25.502413,25.258911,29.521889,33.802013,41.014435,47.516933,43.109913,50.514393,50.267464,48.576675,47.523792,45.07164,50.006813,47.510075,42.763527,40.167328,43.30883,38.22961,34.230713,29.134346,22.487804,15.584045,11.513125,8.289313,5.970912,4.4241676,3.316411,2.5790498,2.0165975,1.587899,1.2620882,1.0357354,0.823101,0.5693115,0.33952916,0.15433143,0.0,0.0,0.061732575,0.061732575,0.0034295875,0.010288762,0.0548734,0.037725464,0.01371835,0.020577524,0.044584636,0.4355576,0.9259886,1.1420527,1.1454822,1.4507155,3.5770597,5.3570156,6.948344,8.354475,9.434795,10.635151,11.46854,11.962401,11.996697,11.31078,10.765475,10.39508,10.316199,10.449953,10.532263,8.261876,7.284444,6.8626046,6.711703,6.992929,6.159539,5.744559,5.888602,6.3207297,6.3447366,6.2658563,6.4990683,6.0737996,5.442755,6.4887795,6.0326443,5.5559316,5.096367,4.5510626,3.683377,3.4913201,3.2306714,3.2821152,3.649081,3.9543142,3.8617156,3.7279615,3.7382503,3.940596,4.273266,5.610805,8.069819,10.014396,10.645439,10.024684,9.23245,8.913498,8.371623,7.829748,8.405919,6.728851,4.712253,3.542764,3.5839188,4.40359,3.724532,4.0674906,4.307562,4.1463714,4.1292233,5.2575574,5.967482,6.210983,6.090947,5.885172,6.773435,7.274155,7.407909,7.1541195,6.447624,6.3207297,6.9037595,7.723431,8.275595,8.045813,8.272165,8.457363,8.80718,9.355915,9.97667,9.129561,9.39707,9.863494,10.038403,9.877212,10.851214,10.72432,10.549411,10.460241,9.671436,9.283894,8.793462,8.169277,7.6685576,7.8331776,7.6205435,7.438775,7.016936,6.3207297,5.5730796,5.377593,5.055212,5.0895076,5.4804807,5.751418,6.200694,6.8454566,7.130112,7.2158523,7.9772205,7.5862474,7.2535777,6.138962,5.7754254,10.05898,13.982429,16.064188,16.94902,15.6526375,9.561689,14.099034,16.146498,14.671775,11.334786,10.47396,11.729189,10.038403,7.846896,6.557371,6.509357,5.90232,3.292404,1.5055889,1.4335675,2.0406046,1.5193073,1.5810398,1.9411465,2.287535,2.287535,1.5981878,1.4404267,1.5810398,1.8485477,2.136633,2.0680413,1.704505,1.488441,1.4369972,1.1489118,1.0460242,1.0871792,1.2792361,1.4644338,1.3512574,1.3924125,1.2380811,0.9945804,0.8093826,0.864256,0.90198153,0.91227025,0.939707,0.9259886,0.72707254,0.78194594,0.66876954,0.5624523,0.548734,0.61389613,0.5761707,0.6276145,0.72021335,0.7339317,0.47671264,0.6859175,0.8676856,0.91227025,0.8779744,0.96371406,1.1489118,1.1454822,1.1317638,1.2312219,1.4953002,1.138623,1.0631721,1.1626302,1.4061309,1.821111,3.07634,3.9028704,4.5442033,5.086078,5.453044,5.4667625,5.638242,5.9812007,6.4236174,6.807731,7.407909,8.049242,8.577398,8.947794,9.22216,9.095266,8.899779,8.707723,8.4093485,7.7371492,7.723431,7.781734,7.905199,8.080108,8.275595,7.596536,7.455923,7.6033955,7.891481,8.289313,8.340756,8.364764,8.241299,8.117833,8.385342,9.39021,10.024684,9.465661,8.361334,8.827758,8.944365,8.934075,9.445084,10.545981,11.72233,12.843805,13.684054,14.369971,14.5585985,13.430264,12.356804,11.921246,11.516555,11.2421875,11.9040985,13.368532,13.780083,13.443983,12.696333,11.928105,12.329367,13.1593275,13.203912,12.836946,14.016724,14.376831,14.562028,14.273943,13.63604,13.197053,12.257345,11.808069,12.521424,14.407697,16.842705,15.71094,16.019604,17.058767,18.331144,19.54522,20.766151,23.022821,24.367218,24.43924,24.490685,26.747353,27.121178,26.332373,25.571005,26.493563,27.865398,27.340672,26.68562,26.740494,27.422981,28.235794,27.84482,27.244642,26.569014,25.084003,23.890507,24.226606,25.035988,25.663603,25.845371,25.564144,24.418663,23.660725,23.931662,25.238335,25.670462,26.575872,26.514141,25.43382,24.669024,25.324074,25.306927,24.981115,24.572994,24.168303,0.7407909,0.6276145,0.5761707,0.5796003,0.6310441,0.6962063,0.77508676,0.84367853,0.96714365,1.1489118,1.3341095,1.4815818,1.5570327,1.529596,1.5398848,1.8965619,1.7696671,2.0817597,2.2258022,2.0920484,2.0920484,2.1194851,1.9342873,1.8965619,2.1640697,2.6716487,3.4535947,3.82399,4.4550343,5.4187484,6.1904054,5.5662203,5.4016004,8.769455,15.638919,22.875349,20.436913,14.661487,8.790032,4.57164,2.2806756,1.0700313,0.59674823,0.48357183,0.4698535,0.40126175,0.5796003,0.64133286,0.6379033,0.61389613,0.6207553,0.6824879,0.8128122,1.0220171,1.2312219,1.255229,1.4232788,2.318401,3.0557625,2.976882,1.6633499,1.4781522,1.1832076,0.89512235,0.66533995,0.490431,0.38754338,0.34981793,0.3566771,0.3841138,0.38754338,0.3018037,0.274367,0.31209245,0.3841138,0.4081209,0.32581082,0.4081209,0.5453044,0.67219913,0.7922347,0.70306545,0.5658819,0.47671264,0.4115505,0.23321195,0.26750782,0.22635277,0.21263443,0.25378948,0.32924038,0.40126175,0.5590228,0.6241849,0.58988905,0.61389613,0.7305021,0.6173257,0.5007198,0.47671264,0.53844523,0.52472687,0.5418748,0.6756287,0.8128122,0.65162164,1.1626302,1.0871792,0.77851635,0.58302987,0.8505377,1.2620882,1.7422304,1.9754424,2.0063086,2.2360911,3.0626216,3.0489032,2.884283,3.0386145,3.7931237,5.288424,6.866034,9.112414,10.449953,7.160979,4.746549,3.5153272,2.4384367,1.5673214,2.0303159,6.166398,6.262427,5.593657,5.127233,3.532475,2.9117198,2.1229146,1.4061309,0.91569984,0.7133542,0.6036074,0.42869842,0.25721905,0.12346515,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.017147938,0.024007112,0.0274367,0.041155048,0.17490897,0.2777966,0.29151493,0.216064,0.274367,0.22978236,0.2194936,0.36010668,0.7510797,0.8676856,1.0906088,1.3203912,1.587899,2.037175,2.1434922,2.5310357,2.9322972,3.2786856,3.7039545,3.4913201,3.9337368,4.5201964,5.127233,6.001778,7.3701835,8.049242,8.779744,9.712592,10.412228,10.786053,11.297061,12.274493,13.63261,14.894698,16.660936,17.600643,18.399736,19.572655,21.486366,25.742483,29.062325,33.77115,40.201626,46.680115,50.174866,52.681892,54.163475,54.016003,51.076847,46.446903,44.53662,48.268013,58.75912,75.29659,89.41963,80.79765,58.44017,34.786304,25.68761,29.322973,33.719704,36.264458,36.274746,34.99208,36.233593,37.018967,39.08015,40.860104,37.5094,30.523329,33.91862,37.217884,38.682316,45.335716,54.54416,68.53345,89.224144,107.69933,104.232025,75.17656,54.406975,43.871284,41.278515,40.08502,33.32873,28.122618,24.68617,23.341772,24.518122,22.724447,19.95334,19.675543,21.112541,19.257133,18.938183,16.839275,13.618892,10.371073,8.628842,6.560801,6.1629686,6.358455,6.276145,5.2506986,6.228131,6.135532,6.138962,6.8145905,8.128122,14.939283,16.067617,17.583494,21.674994,26.630747,27.669912,22.28546,17.367432,15.251375,13.690913,15.031882,10.055551,5.8062916,4.65395,4.2938433,5.535354,7.2535777,8.656279,9.743458,11.321068,15.549749,18.176813,19.78186,21.383478,24.418663,20.255144,19.589804,21.002794,22.62156,22.103691,25.125158,25.402954,24.11686,23.156574,25.111439,31.123507,36.271317,43.284824,49.770172,48.23029,51.95482,49.173424,44.97561,42.784103,44.368572,49.80104,45.027054,39.15903,37.40994,41.113895,31.661951,25.52985,20.481497,15.899568,12.751206,10.079557,7.6651278,5.693115,4.190956,3.0248961,2.1434922,1.5227368,1.1008976,0.82996017,0.66191036,0.5144381,0.37382504,0.22978236,0.09602845,0.0,0.0,0.1371835,0.18519773,0.09602845,0.020577524,0.0274367,0.020577524,0.01371835,0.010288762,0.01371835,0.24350071,0.89855194,1.1351935,1.08032,1.821111,5.6245236,7.956643,8.309891,8.128122,10.816919,12.610593,13.728639,13.533153,13.035862,14.911846,12.590015,11.561139,10.326488,8.844906,8.522525,7.4284863,6.461343,6.1766872,6.5230756,6.852316,6.1561093,5.1340923,5.1821065,6.23156,6.759717,6.8728933,7.0478024,6.7974424,6.334448,6.543653,6.0806584,6.2967224,6.217842,5.4187484,4.0057583,4.1463714,3.9165888,3.8720043,4.046913,3.9783216,4.2526884,3.8479972,3.6113555,3.8445675,4.3041325,5.689686,7.582818,8.81061,9.156999,9.373062,8.7145815,7.73029,7.414768,7.6514096,7.233,5.888602,4.8254294,4.389872,4.5442033,4.856296,4.1463714,4.2526884,4.4447455,4.513337,4.7499785,5.9983487,6.783724,6.632822,5.98463,6.1732574,7.699424,7.936065,7.6445503,7.233,6.776865,7.1884155,7.73372,8.224151,8.467651,8.268735,8.258447,8.203573,8.351046,8.776315,9.403929,8.697433,8.718011,9.102125,9.3936405,9.043822,9.990388,9.8429165,9.72288,9.777754,9.187865,8.621983,8.1487,7.582818,7.1541195,7.517656,7.1884155,6.9346256,6.4990683,5.871454,5.267846,5.422178,5.0757895,5.103226,5.576509,5.751418,5.7582774,6.385892,6.6396813,6.5196457,7.006647,6.756287,6.557371,6.0566516,5.785714,7.164408,11.293632,15.46744,17.024471,15.055889,10.377932,13.368532,15.0456,13.87954,10.587136,8.134981,9.325048,6.8763227,4.537344,3.8514268,4.1600895,5.7068334,3.5804894,1.6564908,1.371835,1.704505,1.605047,1.6427724,1.8691251,2.2360911,2.5996273,1.7319417,1.5193073,1.6187652,1.8485477,2.1915064,2.2463799,1.9239986,1.5638919,1.2963841,1.0460242,0.9842916,1.08032,1.2346514,1.3341095,1.2415106,1.3306799,1.2106444,1.0288762,0.91227025,0.96714365,0.96371406,0.9328478,0.91912943,0.881404,0.70306545,0.7339317,0.67219913,0.5761707,0.490431,0.4424168,0.5418748,0.6276145,0.65848076,0.607037,0.44584638,0.39097297,0.58645946,0.71678376,0.7373613,0.8711152,0.9945804,1.0597426,1.1454822,1.2826657,1.4541451,1.2380811,1.1660597,1.2003556,1.3272504,1.5536032,2.7779658,3.6970954,4.437886,5.007198,5.271276,5.446185,5.627953,5.871454,6.186976,6.5779486,7.226141,7.997798,8.519095,8.772884,9.081548,8.690575,8.124693,8.004657,7.9875093,6.7528577,6.8385973,7.298162,7.7748747,8.189855,8.735159,7.9737906,7.675417,7.589677,7.473071,7.1061053,7.4181976,7.970361,8.165848,7.9772205,7.922347,8.7145815,9.743458,9.849775,9.15014,8.999237,9.472521,9.15014,8.882631,9.283894,10.703742,12.336226,13.910407,14.788382,14.843254,14.438563,13.2862215,12.778643,12.545431,12.185325,11.269625,12.994707,13.179905,12.6929035,12.061859,11.47197,11.273054,12.157887,12.281353,11.958971,13.649758,13.992717,13.924125,13.7697935,13.522863,12.878101,12.120162,12.373952,13.375391,14.822677,16.37285,14.79867,15.776102,17.566347,19.281141,20.875898,23.11199,23.996824,23.712168,23.321196,24.778769,27.083452,25.9414,24.295198,24.079134,26.219196,28.369547,28.400414,27.261791,26.071724,26.099161,26.462696,26.10945,26.02371,26.082012,25.042849,24.216316,24.11686,23.746464,23.307476,24.185452,24.813065,24.535269,23.640146,23.26975,25.420103,24.730755,25.701328,26.565584,26.620459,26.202047,26.44212,25.426962,24.713608,24.648445,24.36036,0.67219913,0.6241849,0.5418748,0.5521636,0.66876954,0.77851635,0.84024894,0.84024894,0.91569984,1.1077567,1.3581166,1.371835,1.4369972,1.5398848,1.6496316,1.704505,1.7593783,1.8725548,1.8485477,1.8245405,2.270387,2.1915064,1.9274281,1.9137098,2.3904223,3.3815732,4.249259,4.383013,5.305572,6.6705475,6.2864337,5.8165803,6.40304,11.362224,18.416885,19.682402,11.996697,6.557371,3.7759757,2.7642474,1.3169615,0.7407909,0.4972902,0.4389872,0.44927597,0.432128,0.45613512,0.4081209,0.39783216,0.4629943,0.5658819,0.9294182,1.2929544,1.8108221,2.2566686,2.0234566,1.9582944,2.8808534,3.3026927,2.7230926,1.6187652,1.4267083,1.1043272,0.8265306,0.6344737,0.44584638,0.4424168,0.4115505,0.37725464,0.33609957,0.25378948,0.18176813,0.1920569,0.2709374,0.37039545,0.3806842,0.32924038,0.40126175,0.50757897,0.6173257,0.7510797,0.64819205,0.4389872,0.4046913,0.50757897,0.39783216,0.33266997,0.19548649,0.14061308,0.1920569,0.2709374,0.2709374,0.26407823,0.2469303,0.23664154,0.2777966,0.45613512,0.38754338,0.32581082,0.45270553,0.8779744,0.5212973,0.52472687,0.6962063,0.86082643,0.82996017,2.1263442,1.9720128,1.3409687,0.90541106,1.0117283,1.4027013,2.0920484,2.4624438,2.534465,2.9494452,3.8342788,3.4364467,2.7230926,2.352697,2.6785078,4.5167665,6.0875177,7.599966,8.3922,6.9346256,5.3844523,4.417309,3.234101,1.8965619,1.2963841,2.2258022,2.3492675,2.6064866,3.1655092,3.433017,2.8877127,2.2360911,1.670209,1.2895249,1.097468,1.1111864,0.91912943,0.64133286,0.36696586,0.15090185,0.041155048,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.034295876,0.0548734,0.09259886,0.23321195,0.31895164,0.32238123,0.31895164,0.42183927,0.33266997,0.29151493,0.4629943,0.9294182,0.99801,1.3443983,1.6564908,1.8554068,2.0817597,2.4418662,2.901431,3.4021509,3.858286,4.149801,3.8171308,4.338428,5.0929375,5.8337283,6.697984,8.134981,9.091836,10.055551,11.015835,11.502836,12.123591,12.531713,13.183334,14.284232,15.803539,17.141079,19.017063,20.663265,22.28546,25.077143,29.278389,33.09895,38.291344,44.577778,49.660427,50.500675,51.073418,50.62757,49.070538,46.97849,46.364594,50.061687,57.53476,67.82695,79.56643,81.52473,64.74375,41.32996,21.397196,13.059869,10.371073,10.443094,11.653738,13.279363,15.498305,20.659836,24.61415,27.258362,27.875687,25.135447,23.976246,28.962866,32.1661,33.393894,40.187904,50.973957,65.77263,86.08951,101.24485,88.37361,58.501904,45.15738,39.762638,37.128716,35.461933,32.972054,30.197517,29.18236,30.410152,32.807434,31.288126,28.287237,28.091751,29.655643,26.589592,27.491573,26.421541,22.762173,17.576635,13.622321,11.211322,11.080997,11.794352,12.027563,10.5597,10.347065,9.873782,9.959522,11.005547,12.994707,26.143745,28.126047,25.35837,23.976246,29.8477,20.745575,21.43835,19.11995,13.070158,14.654627,20.430052,13.708061,7.140401,5.528495,5.8234396,5.8405876,8.951223,11.694893,13.365103,16.002455,16.62664,17.504614,22.556396,29.292107,28.84283,24.483826,23.845922,25.114868,25.797358,22.703869,26.59645,27.927132,25.968836,23.221737,25.416672,31.404732,36.06897,40.98014,46.021633,49.38263,45.78842,42.56461,39.268776,38.25362,44.687523,44.951603,39.4917,34.546234,32.15924,30.17351,22.186,17.384579,14.044161,11.255906,8.940934,7.3530354,6.0086374,4.9214582,3.9543142,2.8568463,1.937717,1.3649758,0.96714365,0.65162164,0.4046913,0.2503599,0.16804978,0.082310095,0.0,0.0,0.0,0.18519773,0.3018037,0.24350071,0.061732575,0.037725464,0.024007112,0.0274367,0.041155048,0.037725464,0.13375391,1.0357354,1.3101025,1.2792361,3.0317552,7.7783046,9.613133,9.369633,9.225591,12.710052,15.429714,16.352274,15.100473,13.852104,17.315987,15.066177,14.517444,13.334236,10.978109,8.721441,6.7459984,5.3844523,4.98662,5.456474,6.262427,6.368744,5.06893,4.4516044,5.15467,6.327589,7.4044795,6.989499,6.159539,5.6313825,5.778855,5.9914894,6.948344,7.3221693,6.40304,4.1155047,5.1580997,4.822,4.57507,4.5682106,3.6593697,4.619654,4.0229063,3.532475,3.789694,4.40359,5.802862,7.06495,7.8434668,8.40249,9.630281,9.06097,7.3839016,6.944915,7.5382333,6.385892,5.73427,5.6485305,5.7479887,5.672538,5.0895076,5.038064,4.928317,4.972902,5.329579,6.101236,7.051232,7.1678376,6.776865,6.3961806,6.7528577,8.011517,8.141841,7.922347,7.6651278,7.1884155,7.840037,7.9429245,7.9875093,8.255017,8.81404,8.292743,8.100685,8.196714,8.423067,8.464222,8.591117,8.337327,8.368194,8.628842,8.347616,8.769455,8.519095,8.584257,8.951223,8.594546,7.966932,7.6033955,7.1266828,6.756287,7.3358874,7.0306544,6.667118,6.3618846,6.046363,5.446185,5.8165803,5.164959,4.9694724,5.4976287,5.8165803,5.15467,5.377593,5.627953,5.6828265,5.953764,5.4324665,5.188966,5.518206,5.641671,3.7176728,5.857735,9.9698105,10.779194,8.687145,9.760606,11.626302,9.695444,9.098696,9.277034,3.9714622,3.8960114,3.1655092,3.1517909,3.7108135,3.2032347,5.103226,3.899441,2.1400626,1.2483698,1.5124481,1.7490896,1.8382589,1.8108221,1.8519772,2.311542,1.8382589,1.6770682,1.6633499,1.7388009,1.9239986,2.1160555,1.9102802,1.4747226,1.0597426,0.9842916,0.922559,1.0151579,1.0700313,1.0494537,1.0666018,1.08032,1.0460242,0.9945804,0.9842916,1.1283343,1.0940384,0.980862,0.91227025,0.864256,0.67219913,0.6207553,0.6276145,0.6001778,0.5212973,0.4389872,0.5453044,0.61389613,0.58988905,0.5212973,0.5693115,0.39440256,0.45613512,0.5624523,0.65162164,0.823101,0.8471081,0.922559,1.0768905,1.2106444,1.1180456,1.1043272,1.1797781,1.2415106,1.2929544,1.430138,2.4590142,3.3952916,4.105216,4.523626,4.6436615,4.9180284,5.212973,5.5593615,5.9640527,6.4133286,7.051232,7.8366075,8.320179,8.597976,9.328478,8.762596,7.7920227,7.267296,7.1678376,6.6293926,7.4696417,7.8846216,8.042382,8.207003,8.742019,8.748878,8.597976,8.309891,7.8194594,6.9654922,7.829748,8.7317295,9.1981535,8.985519,8.052671,8.381912,9.146709,9.863494,10.31277,10.535692,11.2421875,10.072699,8.64599,8.110974,9.129561,10.5597,12.370522,12.946692,12.528283,13.200482,13.495427,13.978998,14.2533655,13.567448,10.80663,12.22648,12.13731,11.451392,10.827208,10.693454,10.487679,11.262765,11.170166,10.535692,11.828648,13.2862215,13.207341,13.344524,13.903547,13.540011,13.543441,14.771234,15.659496,15.614912,15.028452,14.417986,15.361122,16.997036,19.061647,21.897917,23.78076,23.142857,22.059107,22.127699,24.466677,26.69591,24.250612,22.275171,23.125708,26.35981,28.554745,29.559614,28.571894,26.593021,26.414682,24.936531,23.821915,23.825344,24.566135,24.511261,25.44068,24.621008,22.683292,20.889618,21.150267,21.506943,22.035099,22.275171,22.998814,26.195189,24.85422,25.042849,25.958548,26.867388,27.121178,27.52244,25.725336,24.6896,25.053137,25.135447,0.61046654,0.6241849,0.6344737,0.7133542,0.8162418,0.77851635,0.7888051,1.0117283,1.2209331,1.3341095,1.4198492,1.3341095,1.2209331,1.2072148,1.2758065,1.2517995,1.5810398,1.4987297,1.430138,1.6599203,2.318401,1.7216529,1.6359133,1.8005334,2.2086544,3.1140654,4.2252517,5.195825,6.210983,7.0203657,6.958633,6.468202,7.373613,12.445972,18.814716,17.960749,8.354475,3.7279615,1.7422304,0.90198153,0.53501564,0.53501564,0.6344737,0.66533995,0.65162164,0.823101,0.6893471,0.42869842,0.31209245,0.4046913,0.5658819,1.3203912,2.609916,3.0420442,2.5241764,2.2429502,2.0714707,2.1297739,1.8999915,1.4472859,1.4335675,1.313532,1.1180456,0.89855194,0.6893471,0.5178677,0.45613512,0.39783216,0.32238123,0.25378948,0.22978236,0.216064,0.30523327,0.39097297,0.41840968,0.3806842,0.37039545,0.44927597,0.59674823,0.7373613,0.7613684,0.64133286,0.3806842,0.30866286,0.45613512,0.5796003,0.21263443,0.10288762,0.08573969,0.07545093,0.07545093,0.07545093,0.15090185,0.18176813,0.14404267,0.106317215,0.12003556,0.15090185,0.3018037,0.51100856,0.548734,0.32924038,0.42869842,0.61389613,0.90198153,1.587899,2.942586,2.750529,1.8999915,1.1694894,1.2037852,1.8519772,2.6545007,3.093488,3.2546785,3.8308492,3.3644254,2.609916,2.2120838,2.301253,2.4727325,3.450165,5.1100855,6.742569,7.39762,5.919468,4.530485,3.5770597,2.7470996,1.9068506,1.1146159,1.5055889,1.1729189,2.020027,3.7622573,3.9200184,3.8720043,2.8980014,1.879414,1.2689474,1.097468,1.1592005,1.2312219,1.039165,0.6173257,0.274367,0.10288762,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.041155048,0.09259886,0.14061308,0.17147937,0.2194936,0.30866286,0.4424168,0.30866286,0.4389872,0.5624523,0.6241849,0.8093826,1.0048691,1.1523414,1.3238207,1.5330256,1.7388009,2.1297739,2.8225505,3.7622573,4.6127954,4.7602673,4.417309,4.8288593,5.761707,7.0786686,8.711152,9.102125,10.079557,11.173596,12.0138445,12.343085,12.5145645,13.207341,14.147048,15.241087,16.571766,18.866161,21.006224,23.568125,26.493563,29.069183,32.790287,37.437378,41.57003,44.313698,45.36315,45.448895,45.500336,44.38915,42.609196,42.266235,45.733547,53.998856,63.800617,73.50978,83.12977,76.13684,54.53044,32.19011,16.856422,10.117283,5.953764,3.9783216,3.590778,4.108646,4.791134,8.3922,11.351934,13.368532,14.369971,14.527733,13.430264,16.825556,20.21399,23.26975,29.861418,39.443684,60.388176,86.19582,102.65441,87.85917,63.896645,55.398125,52.987125,50.64472,45.71297,44.89673,43.593487,44.423447,47.37289,49.787323,51.718178,46.193115,41.89584,40.32166,35.780888,37.015537,39.200184,36.91608,30.50275,26.061436,22.312897,20.406046,20.28601,22.168854,26.565584,20.265432,16.739817,16.101913,17.730967,20.29287,29.35041,37.40308,34.635403,24.048267,21.424633,18.787281,23.44466,21.86362,15.789821,22.247734,16.023033,12.590015,10.120712,9.349055,13.5503,7.39762,8.824328,11.602294,16.235666,29.967735,20.237995,22.456938,31.442457,38.25362,30.197517,30.283257,28.856548,27.10403,27.3441,33.02007,33.387035,27.580742,23.797907,23.499533,21.424633,22.902784,27.196629,34.155262,41.007576,42.372555,40.126175,36.480522,35.791176,38.020405,38.74405,33.517357,28.787956,27.669912,28.023159,22.44665,16.599203,12.792361,9.801761,7.257007,5.645101,4.7808447,4.012617,3.590778,3.223812,2.0749004,1.5364552,1.1111864,0.7579388,0.4664239,0.26064864,0.20920484,0.16119061,0.082310095,0.0,0.0,0.0,0.15433143,0.2709374,0.26750782,0.18176813,0.072021335,0.037725464,0.10288762,0.19548649,0.12346515,0.36696586,1.371835,2.054323,2.4727325,3.8137012,6.451054,6.800872,7.795452,10.477389,13.992717,17.189093,18.320856,16.928444,13.786942,10.8958,9.746887,11.595435,14.315098,15.436573,12.116733,6.3790326,4.4584637,3.957744,3.8102717,4.273266,4.664239,4.448175,4.1635194,4.448175,6.0566516,5.9228973,5.73427,5.336438,5.144381,6.135532,6.5985265,6.1904054,6.1321025,6.2418494,4.9591837,7.377043,6.4407654,5.5147767,5.429037,4.4996185,4.9660425,4.513337,4.139512,4.098357,3.8925817,5.953764,7.81603,8.628842,8.875772,10.374502,10.9369545,8.752307,7.1781263,6.90033,5.936616,6.8145905,6.632822,6.1972647,5.909179,5.7377,5.675967,5.871454,6.1629686,6.526505,7.06495,6.6876955,6.3618846,5.967482,5.7891436,6.5470824,7.023795,7.1678376,7.473071,7.8126,7.4456344,7.9086285,7.805741,7.6651278,7.8606143,8.604835,7.6651278,7.953213,8.447074,8.515666,7.905199,8.038953,7.630832,7.3530354,7.3221693,7.1266828,7.332458,7.394191,7.73029,8.093826,7.5690994,6.8728933,6.697984,6.4544835,6.2384195,6.835168,6.824879,6.728851,6.5779486,6.217842,5.3261495,5.164959,4.7774153,4.9488945,5.5833683,5.7068334,4.7431192,4.602506,4.557922,4.537344,5.1100855,4.856296,4.2252517,4.3933015,5.1340923,4.791134,4.7534084,7.4284863,7.7885933,6.355026,9.184435,6.6465406,4.722542,4.0674906,4.1292233,3.1277838,2.3595562,2.5070283,2.750529,2.6545007,2.1674993,2.0337453,2.1091962,2.037175,1.8073926,1.7696671,1.6221949,1.7525192,1.7593783,1.6496316,1.845118,1.786815,1.7250825,1.7353712,1.8759843,2.1812177,2.0097382,1.5741806,1.214074,1.0425946,0.94656616,1.0425946,1.0494537,1.0494537,1.0666018,1.0666018,0.83681935,0.8505377,0.9259886,0.97057325,1.0082988,0.9328478,0.8711152,0.8162418,0.7682276,0.7339317,0.52472687,0.42869842,0.42183927,0.45270553,0.42869842,0.4629943,0.4355576,0.51100856,0.64133286,0.5796003,0.39783216,0.4424168,0.6927767,0.9945804,1.0666018,0.9842916,0.9877212,1.0494537,1.08032,0.94656616,0.9842916,1.0563129,1.1729189,1.3443983,1.6016173,2.1023371,3.0248961,3.7691166,4.0949273,4.1189346,4.6093655,4.695105,4.938606,5.4976287,6.135532,6.927767,7.8023114,8.213862,8.268735,8.742019,8.498518,8.182996,8.2310095,8.556821,8.543102,8.31332,8.584257,8.663138,8.656279,9.47595,9.561689,9.06097,8.64599,8.601405,8.834618,9.054111,9.887501,10.374502,9.736599,7.3701835,7.3084507,8.683716,9.753747,10.230459,11.290202,11.561139,10.858074,9.856634,9.105555,9.033533,9.434795,10.984968,12.13731,12.113303,10.878652,12.614022,14.198492,14.500296,13.272504,11.183885,9.585697,9.578837,9.73317,9.668007,10.069269,10.899229,11.4205265,10.991828,10.045261,10.069269,12.181894,12.950122,14.369971,16.616352,18.019053,18.667244,19.442331,19.020493,17.250826,15.151917,15.604623,15.350834,15.837835,17.768692,21.102251,22.03167,20.742146,19.497204,20.02193,23.513252,24.061985,21.747015,21.44864,24.19917,27.18977,26.874247,27.800236,27.728214,26.709627,27.1006,24.339783,21.7916,21.013083,22.10712,23.743034,25.889956,24.662163,22.391777,20.378609,18.890167,17.988186,18.71526,19.829874,20.985645,22.703869,23.705309,23.2869,23.002243,23.557837,24.826784,24.593573,24.967398,25.76649,26.689049,27.299517,0.6824879,0.65505123,0.64476246,0.6790583,0.7305021,0.70649505,0.6790583,0.8162418,0.9534253,1.0323058,1.1249046,1.313532,1.3649758,1.5090185,1.7216529,1.7147937,1.6427724,1.6599203,1.6564908,1.7936742,2.4898806,1.9308578,1.8691251,1.9068506,1.920569,2.0646117,3.2135234,3.998899,5.4667625,7.1026754,6.835168,7.5862474,8.766026,12.504276,16.732958,15.165636,6.9723516,3.4707425,2.0131679,1.1763484,0.7407909,0.67219913,0.72707254,0.72707254,0.66876954,0.7133542,0.6790583,0.78537554,0.7990939,0.7682276,1.0151579,1.8691251,2.4727325,2.6750782,2.5310357,2.2806756,2.0303159,1.6873571,1.3581166,1.2346514,1.5913286,1.3649758,1.0906088,0.85739684,0.6859175,0.5555932,0.5041494,0.3806842,0.3018037,0.3018037,0.32581082,0.3841138,0.42869842,0.45613512,0.44927597,0.39440256,0.4115505,0.45270553,0.5212973,0.5693115,0.4938606,0.490431,0.42869842,0.4081209,0.45956472,0.5418748,0.34295875,0.22978236,0.14747226,0.09259886,0.11317638,0.09259886,0.08916927,0.07888051,0.061732575,0.044584636,0.09602845,0.1097468,0.14404267,0.216064,0.29151493,0.3566771,0.607037,0.8265306,1.1214751,1.9411465,2.1812177,2.1091962,2.0063086,2.2463799,3.2821152,3.5873485,3.6936657,3.6765177,3.5118976,3.1106358,2.2155135,2.170929,2.5241764,3.0248961,3.642222,4.2286816,4.7979927,5.7102633,6.3310184,5.0277753,3.7931237,2.9700227,2.8122618,2.9151495,2.201795,3.3438478,3.2135234,3.865145,5.5559316,6.728851,5.470192,3.8720043,2.767677,2.0714707,0.7682276,0.6241849,0.6276145,0.7476501,0.7510797,0.21263443,0.082310095,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.041155048,0.07888051,0.12689474,0.20920484,0.33266997,0.42526886,0.34638834,0.26064864,0.4629943,0.764798,0.9568549,0.7956643,0.65162164,0.6927767,0.980862,1.4164196,1.7525192,2.054323,2.8054025,3.532475,3.9508848,3.9783216,4.5956473,5.346727,6.560801,8.285883,10.261326,10.456812,11.297061,12.061859,12.4974165,12.809509,13.097594,13.738928,15.035312,16.835844,18.547209,20.666695,23.890507,27.371538,30.732533,34.059235,36.720592,39.868954,42.039883,42.602337,41.789524,42.90757,42.0879,41.31281,42.355404,46.758995,53.398678,65.12101,74.92963,80.25921,82.99602,73.441185,50.751034,29.172071,15.5085945,9.091836,7.116394,5.7925735,5.346727,5.754848,6.7322803,10.038403,13.313659,15.05246,15.2033615,15.1862135,15.364552,19.87446,23.972816,27.885975,36.782326,46.258274,77.20687,106.21775,117.631424,103.570114,79.14802,67.964134,61.235283,54.10517,45.616943,43.38428,41.72779,41.751797,42.88356,42.869843,43.216232,36.387924,31.50419,30.358707,27.409264,31.140654,29.885426,27.570454,26.781649,28.77081,24.60386,22.62156,24.295198,29.394995,35.97637,31.620796,26.18833,24.315775,26.202047,27.594461,32.94119,38.07185,36.60056,29.130917,23.252604,19.86417,22.089973,22.20658,19.78872,21.685282,16.513464,12.6929035,10.97468,11.910957,15.858413,13.728639,14.366542,15.114192,17.991615,29.724234,26.03057,31.596788,41.957573,50.56241,48.775593,37.766617,34.67656,33.558514,31.905453,30.626217,27.117748,23.074265,20.793589,21.321745,24.44953,30.019178,29.998602,30.643364,33.884323,37.32077,40.465702,38.620583,38.994408,41.3814,38.15759,29.278389,22.77246,19.394318,17.960749,15.3302555,13.018714,11.046701,8.790032,6.392751,4.791134,3.7691166,2.8739944,2.277246,1.8999915,1.4164196,1.0631721,0.77851635,0.5418748,0.33609957,0.15090185,0.061732575,0.030866288,0.09945804,0.16462019,0.0,0.0,0.030866288,0.058302987,0.19891608,0.72021335,0.5796003,0.4424168,0.45613512,0.5590228,0.47671264,0.72021335,0.823101,1.8828435,3.923448,5.888602,3.8308492,5.425607,10.031544,15.103903,16.239098,18.986197,17.974468,15.848124,13.673765,10.9541025,8.498518,11.345076,13.941273,14.280802,13.910407,8.954653,6.3447366,5.0140567,4.201245,3.4535947,2.527606,2.7299516,3.175798,3.8342788,5.5319247,5.6519604,6.711703,6.6431108,5.377593,4.852866,5.4907694,6.1046658,6.2487082,6.0737996,6.3138704,7.226141,6.8900414,6.2384195,5.610805,4.7808447,4.846007,4.4859004,4.48933,5.0174866,5.6005163,7.466212,9.403929,10.285333,10.155008,10.240748,8.937505,7.222711,6.3001523,6.018926,4.897451,5.8543057,6.1458206,6.5196457,6.8385973,6.090947,6.0978065,6.742569,6.9346256,6.584808,6.625963,6.0532217,6.0978065,6.1286726,6.200694,7.034084,6.7494283,6.8454566,7.5210853,8.39563,8.508806,8.279024,7.723431,7.191845,7.181556,8.337327,7.720001,7.6033955,7.764586,7.932636,7.7714453,7.455923,6.6293926,6.2658563,6.4098988,6.186976,5.6313825,5.4736214,5.6999745,6.1149545,6.310441,5.857735,5.967482,6.018926,6.001778,6.495639,6.492209,6.159539,5.9743414,5.8165803,4.9351764,5.0586414,4.9488945,4.972902,5.0929375,4.863155,3.841138,3.8171308,3.7313912,3.333559,3.1963756,3.2718265,3.292404,3.590778,3.8960114,3.340418,2.8739944,3.5633414,3.9200184,3.7382503,4.1189346,3.7485392,3.4192986,3.3541365,3.4535947,3.309552,3.7142432,3.6182148,3.1243541,2.4658735,2.0097382,2.527606,2.2909644,2.0028791,1.9102802,1.8073926,1.7182233,1.7353712,1.6976458,1.6084765,1.6256244,1.6736387,1.6016173,1.5810398,1.7490896,2.2292318,2.2841053,1.7216529,1.1934965,0.97057325,0.922559,0.9328478,0.90884066,0.88826317,0.8848336,0.8848336,0.88826317,0.9842916,1.0906088,1.1489118,1.1180456,1.1008976,0.9568549,0.8505377,0.7990939,0.6962063,0.5658819,0.44584638,0.41498008,0.4698535,0.52472687,0.36696586,0.36353627,0.48014224,0.6036074,0.5418748,0.4972902,0.52472687,0.5624523,0.61389613,0.77508676,1.0494537,1.214074,1.1900668,1.0528834,1.0082988,0.88826317,0.94999576,1.1249046,1.3546871,1.6016173,2.0063086,2.7128036,3.4673128,4.108646,4.57164,4.540774,4.5339146,4.7191124,5.254128,6.2692857,6.759717,7.2947326,7.7577267,8.189855,8.793462,8.683716,8.687145,9.0369625,9.5205345,9.458802,8.865483,9.019815,9.695444,10.30934,9.914937,9.3764925,8.916927,8.793462,9.067829,9.602845,10.048691,10.425946,10.600855,10.316199,9.187865,8.738589,9.619993,10.611144,11.30735,12.133881,11.993267,11.276484,9.945804,8.604835,8.484799,8.995808,10.443094,11.633161,12.21619,12.723769,13.155897,13.663476,13.642899,12.535142,9.8429165,9.678296,10.991828,11.993267,12.13731,12.109874,12.46998,12.322508,11.581717,10.748327,10.88894,12.854094,13.927555,14.675205,15.481158,16.54433,17.610931,17.79613,17.096493,15.985307,15.409137,15.223939,15.450292,15.806969,16.914726,20.28601,19.668684,19.123379,18.79071,19.486916,22.69701,23.27318,22.20315,22.055677,23.358921,24.60386,23.19087,23.406935,23.749893,23.214878,21.290878,20.718138,20.841602,21.386908,22.254593,23.509823,24.185452,23.986534,22.86163,21.407484,20.855322,19.102802,19.178253,19.884748,21.016512,23.35206,23.297188,23.166862,23.372639,23.61957,22.895926,21.70929,22.60441,23.69159,24.600431,26.479845,0.72021335,0.66876954,0.6790583,0.6859175,0.6893471,0.7682276,0.7476501,0.77508676,0.90198153,1.0734608,1.1351935,1.2963841,1.3752645,1.4061309,1.4678634,1.6942163,1.6839274,1.7490896,1.7388009,1.8039631,2.3972816,2.3149714,2.2669573,2.136633,1.978872,2.0028791,3.4535947,4.2938433,5.435896,6.478491,5.7068334,6.8283086,8.124693,11.581717,15.258235,13.282792,6.701414,3.8445675,2.633923,1.8725548,1.2586586,0.91912943,0.7373613,0.5796003,0.4629943,0.58645946,1.1146159,1.08032,0.89169276,0.8711152,1.2483698,2.2086544,2.3835633,2.2566686,2.0577524,1.7765263,1.3821237,1.0906088,0.9568549,0.9945804,1.1763484,0.83681935,0.64133286,0.5178677,0.4389872,0.3806842,0.4355576,0.36010668,0.29837412,0.31895164,0.4046913,0.48014224,0.5041494,0.4698535,0.40126175,0.37725464,0.39440256,0.36010668,0.3566771,0.37382504,0.32581082,0.31552204,0.32581082,0.30866286,0.28808534,0.37039545,0.32924038,0.22635277,0.14404267,0.1097468,0.10288762,0.13032432,0.12346515,0.08916927,0.041155048,0.030866288,0.07545093,0.06859175,0.07545093,0.116605975,0.17490897,0.34638834,0.72021335,1.0014396,1.1900668,1.5913286,1.5913286,1.937717,2.4487255,3.0626216,3.8548563,4.139512,4.636802,4.5819287,3.8377085,2.884283,2.8568463,3.2032347,3.350707,3.357566,3.899441,4.5339146,5.003768,5.1512403,5.051782,5.0174866,4.671098,3.6010668,3.2992632,3.6765177,3.07634,4.173808,3.765687,3.57363,4.1772375,5.003768,4.0503426,2.6853669,1.6736387,1.097468,0.33952916,0.25378948,0.23664154,0.29837412,0.33266997,0.09602845,0.041155048,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.024007112,0.041155048,0.0548734,0.08573969,0.07545093,0.14404267,0.2777966,0.40126175,0.37382504,0.29494452,0.59674823,0.8471081,0.9431366,1.0871792,0.71678376,0.59674823,0.7990939,1.2003556,1.471293,1.7353712,2.417859,3.1586502,3.7519686,4.1326528,5.096367,5.9880595,7.373613,9.280463,11.180455,11.327928,11.897239,12.394529,12.761495,13.371962,13.96871,14.781522,16.417435,18.656956,20.460918,23.290329,26.881107,30.660511,34.289017,37.653442,38.435387,39.687187,40.030144,39.32365,38.685745,39.378525,37.7186,37.766617,41.635193,49.475227,56.54361,66.31107,74.59353,79.23033,80.06029,66.90096,43.130493,22.78275,11.907528,8.56025,7.2192817,7.133542,7.6274023,8.344186,9.239308,12.452832,14.812388,15.7795315,15.937293,16.990177,17.511473,20.570665,24.257473,29.425861,39.711193,39.83123,69.600044,93.28821,96.2548,84.96803,58.95461,49.588406,43.528324,35.437927,27.988863,27.577312,26.956558,27.800236,29.473875,29.028028,29.271528,25.93111,24.401514,25.221186,24.068846,28.835972,26.929121,23.866499,23.266321,26.822803,24.284908,23.712168,25.512701,29.065754,32.707977,31.75455,27.611609,27.066305,30.327843,30.993181,31.048056,31.939749,30.554195,26.802225,23.629858,20.323736,20.776442,21.925352,22.738165,24.19231,18.735836,14.805529,11.89038,11.094715,15.162207,15.927004,17.593784,19.480057,23.85964,35.962654,43.40143,40.359386,39.111015,44.31713,53.055717,46.30286,40.75036,37.855785,36.357056,32.282707,28.26323,24.826784,21.825895,20.834743,25.135447,29.34012,28.774239,28.784527,31.830002,37.4751,37.653442,35.57511,35.921497,38.31535,37.33106,27.659622,21.808746,18.245405,15.885849,14.088745,12.178465,10.556271,8.766026,6.807731,5.171818,3.789694,2.6956558,1.8999915,1.3546871,0.94999576,0.6790583,0.48357183,0.33609957,0.2194936,0.13032432,0.08573969,0.116605975,0.13032432,0.082310095,0.0,0.0,0.0,0.1920569,0.4664239,0.4046913,0.5144381,0.7442205,1.0185875,1.1523414,0.8471081,1.1283343,0.85739684,1.9274281,4.65395,7.7714453,2.8088322,4.434457,8.282454,10.998687,10.254466,15.638919,16.901007,15.46401,12.836946,10.6317215,10.432805,10.329918,9.887501,9.575408,10.762046,8.519095,6.3653145,5.096367,4.2526884,2.1434922,1.8073926,2.2978237,2.8088322,3.549623,5.7411294,5.638242,6.8969,6.9552035,5.562791,4.7602673,5.7068334,6.4990683,6.3824625,5.977771,7.267296,8.090397,7.3873315,6.3824625,5.627953,5.0003386,4.6779575,4.6127954,5.2609873,6.4064693,7.1712675,9.253027,10.401938,10.39508,9.3593445,7.764586,6.7631464,6.2658563,5.4633327,4.6745276,5.360445,5.8474464,6.046363,6.5950966,7.116394,6.2247014,6.447624,7.473071,7.3701835,6.3824625,6.917478,6.228131,6.1458206,6.2967224,6.5367937,6.9826403,6.8866115,6.783724,7.208993,8.083538,8.718011,8.182996,7.7371492,7.143831,6.7871537,7.658269,7.281014,7.0889573,7.1026754,7.284444,7.534804,7.349606,6.012067,5.2609873,5.2987127,4.7979927,4.6676683,4.6127954,4.7602673,5.113515,5.5559316,5.3432975,5.5730796,5.645101,5.552502,5.9160385,5.6348124,5.2506986,5.2335505,5.4153185,4.9831905,5.164959,4.9214582,4.57507,4.2938433,4.0880685,3.2032347,3.1209247,3.093488,2.884283,2.7711067,2.6887965,2.627064,2.7573884,2.8945718,2.4795918,2.352697,2.3595562,2.4144297,2.4075704,2.2120838,2.8156912,3.175798,3.1483612,2.9494452,3.1449318,3.316411,3.3129816,3.3815732,3.316411,2.452155,2.294394,2.287535,2.435007,2.4967396,1.9720128,1.7456601,1.6736387,1.6907866,1.7147937,1.6530612,1.646202,1.5913286,1.5673214,1.6427724,1.8588364,1.9754424,1.5981878,1.255229,1.1043272,0.91569984,0.823101,0.89855194,0.939707,0.88826317,0.8196714,0.8745448,1.0151579,1.1694894,1.2415106,1.1249046,1.0666018,0.9911508,0.89855194,0.77851635,0.6036074,0.58302987,0.53501564,0.5178677,0.5178677,0.4664239,0.3841138,0.40126175,0.4424168,0.44584638,0.37725464,0.38754338,0.47328308,0.48357183,0.432128,0.490431,0.6962063,0.8676856,1.0117283,1.097468,1.0494537,0.91227025,1.0014396,1.1454822,1.2895249,1.4747226,1.9239986,2.5378947,3.3369887,4.1326528,4.5030484,4.554492,4.588788,4.6848164,5.0243454,5.871454,6.6465406,7.174697,7.73029,8.261876,8.419638,8.433355,8.752307,9.290752,9.753747,9.644,9.071259,9.489669,10.501397,11.417097,11.231899,10.192734,9.208443,8.958082,9.441654,9.9801,9.6817255,9.712592,9.637141,9.366203,9.15014,9.253027,9.911508,10.72432,11.4033785,11.777204,11.677745,11.458252,10.7757635,9.729739,8.841476,8.954653,10.30591,11.862943,12.9981365,13.474849,11.732618,11.026124,11.122152,11.303921,10.347065,10.851214,12.250486,12.682614,12.017275,11.869802,12.096155,12.003556,11.766914,11.499407,11.276484,13.512574,14.87755,14.894698,13.941273,13.262215,14.96329,15.388559,15.165636,14.802099,14.695783,14.932424,16.441442,17.54234,17.802988,18.056778,17.312557,17.737827,18.605513,19.740705,21.503513,21.77445,21.764162,21.657845,21.606401,21.723007,20.742146,21.44178,21.95279,21.061096,18.20768,18.708399,19.562366,21.146837,23.142857,24.52498,24.058556,23.328054,22.384918,21.61669,21.723007,20.680412,20.409475,20.992504,22.415783,24.576424,25.070284,23.811626,22.77246,22.501524,22.12084,21.009653,21.825895,23.02625,23.78419,24.003683,0.7888051,0.7133542,0.72707254,0.7339317,0.7407909,0.8711152,0.88826317,0.8162418,0.91569984,1.1420527,1.1351935,1.1900668,1.3066728,1.371835,1.4472859,1.7730967,1.6839274,1.6976458,1.6427724,1.6256244,2.0097382,2.287535,2.3081124,2.2566686,2.270387,2.4247184,3.6593697,4.523626,5.381023,5.826869,4.6676683,5.802862,7.257007,10.401938,13.786942,13.138749,7.7097125,4.712253,3.4638834,2.9665933,1.920569,1.0494537,0.6173257,0.50757897,0.6379033,0.96371406,1.3615463,1.1317638,0.84024894,0.823101,1.1866373,2.5138876,2.4075704,1.845118,1.3684053,1.0734608,0.78537554,0.64819205,0.66533995,0.7305021,0.64476246,0.37039545,0.29494452,0.26750782,0.22635277,0.20577525,0.33609957,0.29837412,0.2709374,0.31552204,0.37382504,0.4046913,0.39097297,0.33609957,0.28122616,0.30523327,0.34295875,0.30523327,0.25378948,0.22635277,0.23664154,0.20920484,0.22978236,0.23664154,0.23321195,0.30866286,0.2469303,0.1920569,0.15090185,0.11317638,0.08573969,0.15776102,0.15776102,0.10288762,0.030866288,0.017147938,0.05144381,0.037725464,0.037725464,0.08573969,0.20577525,0.31209245,0.5761707,0.805953,0.980862,1.255229,1.4164196,2.1434922,2.9803114,3.6216443,3.9028704,4.1600895,4.7808447,4.897451,4.2526884,3.1895163,3.5976372,3.9680326,3.9200184,3.5702004,3.5530527,4.496189,4.57507,4.3795834,4.434457,5.1992545,5.9331865,4.7019644,3.875434,3.9714622,3.642222,3.6182148,2.8877127,2.2498093,2.1434922,2.668219,1.9994495,1.1934965,0.59674823,0.30866286,0.17490897,0.14061308,0.1097468,0.10288762,0.09945804,0.037725464,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.010288762,0.006859175,0.010288762,0.010288762,0.010288762,0.034295876,0.037725464,0.034295876,0.041155048,0.061732575,0.09259886,0.13032432,0.12003556,0.19548649,0.3841138,0.61389613,0.5521636,0.6241849,0.70649505,0.7888051,0.9774324,0.72364295,0.6001778,0.69963586,0.94656616,1.1111864,1.488441,2.0714707,2.8911421,3.7862647,4.431027,5.470192,6.4373355,7.8537555,9.657719,11.218181,11.763485,12.295071,12.854094,13.54687,14.55174,15.522313,16.46888,18.063637,20.303158,22.52553,26.531288,29.875137,33.18469,36.41193,38.82979,38.596577,38.606865,37.81806,36.545685,36.470234,36.57998,35.355618,36.885212,42.24909,49.49238,55.312386,61.83546,69.59662,76.42493,77.46752,59.53764,35.2493,16.54433,7.9429245,6.557371,5.593657,6.667118,7.7131424,8.2653055,9.462232,12.620882,14.2190695,15.316538,16.520323,17.995045,19.178253,20.70099,23.297188,29.233803,42.31082,34.779446,55.267803,67.77208,63.745743,62.10983,36.874924,30.368998,26.28093,19.809298,17.672665,16.955881,17.158226,18.581505,20.436913,20.827885,21.94593,20.910194,21.805317,24.27462,23.502962,26.702768,25.577864,22.799898,21.225718,23.897366,22.069395,21.548098,22.477516,24.161444,25.059996,26.147175,23.677872,24.151155,27.302946,26.092302,24.27805,22.501524,20.793589,19.654966,20.059656,22.796469,22.5221,22.820475,25.097721,28.599329,23.472097,17.521763,12.041282,9.630281,14.177915,15.388559,20.652975,25.114868,28.777668,36.504528,53.480988,49.30032,42.423996,42.108475,48.415485,46.333725,41.683205,38.46625,37.40308,35.942078,31.2504,26.380386,22.607841,21.36633,24.250612,25.920822,27.460707,29.09662,31.6791,36.67601,31.50762,28.565035,29.741383,33.363026,34.17584,27.316664,24.212887,22.02481,19.459478,16.743246,21.215427,15.282242,9.544542,7.517656,5.641671,4.1360826,2.8980014,2.0063086,1.4164196,0.9602845,0.70649505,0.5007198,0.32924038,0.21263443,0.17490897,0.14061308,0.14061308,0.08916927,0.0,0.0,0.0,0.12003556,0.45613512,0.7305021,0.28465575,0.66191036,1.1694894,1.4267083,1.4198492,1.5124481,1.4232788,1.2072148,2.2600982,4.8837323,8.292743,2.6064866,2.8980014,4.712253,5.9743414,7.006647,12.010415,14.706071,14.441993,12.22648,10.734609,10.319629,9.47595,7.514226,5.6176643,6.824879,6.258997,6.0052075,5.8543057,4.914599,1.605047,1.9342873,1.9582944,2.318401,3.4947495,5.7822843,6.632822,7.3118806,7.1266828,6.2144127,5.535354,5.9571934,6.464772,6.279575,5.9228973,7.2158523,8.275595,7.7371492,6.667118,5.6965446,5.0277753,4.647091,4.712253,5.658819,7.205563,8.368194,9.997248,10.268185,9.578837,8.152129,6.0497923,5.271276,5.007198,4.214963,3.6559403,5.8988905,6.5882373,6.4098988,6.697984,7.363324,6.8900414,6.8797526,7.3358874,7.0718093,6.3790326,7.034084,6.228131,6.228131,6.4544835,6.684266,7.0306544,7.058091,6.8214493,7.0443726,7.6857057,7.9257765,7.750868,7.5759587,7.2192817,7.0478024,7.98065,7.2467184,6.9654922,6.694555,6.4819202,6.869464,7.0958166,5.8680243,5.0140567,4.8425775,4.1429415,4.331569,4.3933015,4.4859004,4.7088237,5.1169443,5.1512403,5.3432975,5.2815647,5.079219,5.3707337,4.9214582,4.537344,4.588788,4.9008803,4.7259717,4.6745276,4.3692946,3.998899,3.7382503,3.7794054,2.9460156,2.5721905,2.4212887,2.4007113,2.5893385,2.4452958,2.2258022,2.1743584,2.253239,2.1091962,2.1915064,1.99602,1.920569,2.0234566,2.0165975,2.369845,2.8088322,2.6819375,2.270387,2.760818,2.4452958,2.4247184,2.8019729,3.117495,2.3424082,1.9171394,2.1812177,2.435007,2.3321195,1.879414,1.6496316,1.670209,1.7971039,1.8759843,1.7456601,1.6804979,1.7662375,1.7662375,1.6427724,1.5638919,1.6530612,1.488441,1.3478279,1.2415106,0.91569984,0.85739684,0.9877212,1.0631721,1.0014396,0.88826317,0.91227025,1.196926,1.3992717,1.3546871,1.0837497,0.9911508,0.9602845,0.88826317,0.7442205,0.5796003,0.6310441,0.6344737,0.61046654,0.5658819,0.490431,0.52472687,0.52472687,0.47328308,0.38754338,0.32924038,0.30866286,0.38754338,0.42869842,0.39097297,0.33266997,0.37039545,0.48014224,0.7133542,1.0288762,1.2758065,1.0700313,1.0871792,1.1797781,1.2860953,1.4369972,1.8485477,2.393852,3.1655092,3.974892,4.341858,4.3590055,4.496189,4.633373,4.8734436,5.5250654,6.560801,7.14726,7.7131424,8.162418,7.846896,7.7885933,8.40249,9.067829,9.431366,9.403929,9.225591,9.798331,10.765475,11.729189,12.264205,10.81006,9.304471,8.752307,9.201583,9.736599,9.084977,9.132992,8.916927,8.604835,9.513676,10.251037,10.731179,10.943813,10.981539,11.008976,11.163307,11.533703,11.585147,11.094715,10.151579,9.829198,10.854645,12.528283,13.821238,13.371962,10.6317215,9.47938,9.770895,10.81006,11.331357,12.205902,12.902108,12.644889,11.760056,11.698323,11.38623,11.159878,11.444533,12.05157,12.199042,13.6086035,14.393978,14.232788,13.354814,12.548861,13.745787,14.256795,14.225929,13.96871,13.992717,15.011304,17.610931,19.099373,18.605513,17.069057,17.03819,18.025911,19.20569,19.95334,19.850452,19.274282,19.94648,19.967058,19.219408,19.342873,19.829874,20.759293,20.766151,19.377169,17.017612,17.87501,18.708399,20.423193,22.796469,24.494114,22.210009,20.954779,20.409475,20.546658,21.630407,21.527521,22.216867,23.184011,24.147726,25.063425,26.373528,25.114868,22.985096,21.417774,21.585823,21.187992,21.77445,22.559826,22.919933,22.36777,0.84024894,0.7339317,0.7305021,0.7613684,0.8093826,0.9294182,1.0254467,0.91227025,0.939707,1.1111864,1.0734608,1.155771,1.2826657,1.4747226,1.7182233,1.9823016,1.6290541,1.5638919,1.4781522,1.3889829,1.6256244,1.8965619,1.9754424,2.194936,2.5961976,2.942586,3.5976372,4.5339146,5.360445,5.5833683,4.6093655,5.7068334,7.233,9.513676,12.229909,14.435134,10.299051,6.3173003,4.245829,3.7279615,2.2806756,1.0014396,0.53158605,0.78194594,1.3684053,1.6187652,1.1866373,0.9362774,0.84367853,0.8711152,0.980862,2.4727325,2.2292318,1.4027013,0.71678376,0.48014224,0.48357183,0.45956472,0.48700142,0.5007198,0.29151493,0.19891608,0.21263443,0.23321195,0.23321195,0.2469303,0.36010668,0.29494452,0.28122616,0.34295875,0.30866286,0.25378948,0.18176813,0.14061308,0.15090185,0.22635277,0.28122616,0.28808534,0.23664154,0.17147937,0.20234565,0.18176813,0.18176813,0.22635277,0.29837412,0.32581082,0.15090185,0.15776102,0.16119061,0.106317215,0.082310095,0.16462019,0.14747226,0.07888051,0.01371835,0.01371835,0.044584636,0.048014224,0.030866288,0.061732575,0.26407823,0.26407823,0.28808534,0.40126175,0.70649505,1.3169615,1.7250825,2.633923,3.4192986,3.799983,3.8479972,4.064061,4.2355404,4.5442033,4.7191124,4.0194764,3.9886103,4.15323,4.1360826,3.782835,3.1620796,4.098357,3.4913201,3.3232703,4.0709205,4.7088237,6.125243,5.4084597,4.5339146,4.190956,3.789694,2.3904223,1.6564908,1.2792361,1.1626302,1.4129901,0.6927767,0.37382504,0.31552204,0.38754338,0.45613512,0.34981793,0.25378948,0.31552204,0.39783216,0.06859175,0.034295876,0.01371835,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.037725464,0.061732575,0.072021335,0.08916927,0.05144381,0.034295876,0.0548734,0.082310095,0.24007112,0.20234565,0.26064864,0.5007198,0.8265306,0.7888051,0.5212973,0.47328308,0.6379033,0.5212973,0.6001778,0.607037,0.65848076,0.77508676,0.91227025,1.4850113,2.0097382,2.843128,3.8891523,4.619654,5.751418,6.931196,8.368194,9.928656,11.122152,12.257345,12.936404,13.831526,15.138199,16.575195,17.724108,18.684393,19.901896,21.812176,24.840502,29.391565,31.987762,34.340458,36.717163,37.962105,37.694595,37.16644,36.00038,34.940636,35.880344,36.73431,36.92294,39.210472,43.600346,47.338596,52.60644,57.93602,67.05872,76.3632,74.88847,51.646156,28.132906,11.924676,5.096367,4.2286816,3.7039545,5.1169443,5.9228973,6.0566516,7.915488,10.998687,12.624311,14.507155,16.602633,17.099922,20.62211,22.395206,24.507832,30.475315,45.246548,38.109577,50.54869,51.241467,40.119312,48.367474,27.02858,22.624989,19.805868,15.522313,19.03421,15.827546,16.19794,17.53891,18.849012,20.718138,22.254593,20.488356,20.95135,23.396646,21.78474,21.578964,21.20171,20.251715,19.233126,19.521212,17.315987,15.54632,15.340545,16.503176,17.504614,19.260563,17.46003,17.734396,19.569225,16.307688,16.2974,14.661487,12.912396,12.703192,15.834405,26.00999,26.946268,25.282919,26.383816,34.340458,30.362139,20.172834,11.530273,9.136421,14.63062,13.680624,23.256033,30.51304,31.593359,31.655092,49.88678,52.52413,49.849052,46.5738,41.827248,39.279064,38.558853,36.89207,35.14984,37.859215,31.09607,25.214327,22.875349,23.571554,23.629858,24.336353,28.914852,31.32928,30.708527,31.356718,24.106571,21.94593,24.058556,27.44356,26.929121,24.802776,24.953678,24.922812,23.324625,19.847023,30.989752,20.426622,10.285333,7.9943686,6.276145,4.383013,3.0420442,2.218943,1.7456601,1.3238207,1.0666018,0.7956643,0.53844523,0.33266997,0.24350071,0.18519773,0.08573969,0.024007112,0.01371835,0.0034295875,0.006859175,0.26750782,0.64819205,0.89169276,0.607037,1.0768905,1.6564908,1.7490896,1.5947582,2.2909644,1.6530612,2.0063086,3.4055803,5.5147767,7.6205435,3.0866287,1.5055889,1.7182233,3.590778,8.008087,9.791472,11.550851,12.092726,11.369082,10.477389,7.613684,8.251588,6.989499,3.9508848,4.7945633,4.249259,6.0052075,7.1026754,5.9914894,2.534465,2.136633,1.3341095,1.6221949,3.2718265,5.3398676,7.932636,7.630832,6.9209075,6.7185616,6.3618846,5.885172,6.307011,6.23499,5.7274113,6.2830043,7.534804,7.8606143,7.1541195,5.8645945,5.020916,4.770556,4.8322887,5.7068334,7.298162,8.934075,9.589127,9.290752,8.378482,7.085528,5.562791,4.602506,3.8891523,3.3644254,3.6010668,5.8165803,7.414768,6.8969,6.7700057,7.531374,7.682276,7.1712675,6.6396813,6.427047,6.560801,6.773435,5.8165803,6.094377,6.375603,6.4544835,7.140401,7.181556,7.0375133,7.233,7.5210853,6.883182,7.500508,7.373613,7.157549,7.4524937,8.80718,7.507367,7.1369715,6.591667,5.8543057,5.98463,6.451054,5.8234396,5.2644167,4.99005,4.2766957,4.280125,4.355576,4.431027,4.5270553,4.7534084,4.931747,5.003768,4.8288593,4.6093655,4.8940215,4.513337,4.1429415,4.1429415,4.3590055,4.1360826,3.806842,3.7108135,3.666229,3.6559403,3.8377085,2.9220085,2.2669573,1.8828435,1.821111,2.177788,2.2463799,2.0646117,1.937717,1.9445761,1.9754424,1.9514352,1.6942163,1.6942163,1.99602,2.2360911,1.8485477,2.085189,2.020027,1.7353712,2.3252604,1.8554068,1.6804979,1.7593783,1.8656956,1.5947582,1.5947582,1.9068506,1.8725548,1.529596,1.6187652,1.5090185,1.6667795,1.8519772,1.9239986,1.8485477,1.8142518,2.0817597,2.1057668,1.8142518,1.5947582,1.587899,1.471293,1.371835,1.2586586,0.9568549,0.96714365,1.0460242,1.1043272,1.0871792,0.96714365,1.0220171,1.4164196,1.587899,1.3855534,1.0700313,1.0082988,0.9328478,0.83681935,0.7442205,0.7339317,0.7888051,0.7510797,0.6859175,0.6310441,0.58645946,0.6310441,0.59674823,0.5178677,0.44584638,0.42869842,0.33609957,0.35324752,0.39783216,0.39783216,0.29494452,0.2503599,0.29151493,0.4664239,0.83681935,1.4815818,1.1934965,1.1111864,1.1832076,1.3478279,1.5227368,1.8142518,2.287535,2.9460156,3.6799474,4.280125,4.0606318,4.280125,4.5682106,4.839148,5.288424,6.3035817,6.917478,7.48336,7.8331776,7.274155,6.992929,7.750868,8.48137,8.803751,9.016385,9.14328,9.623423,10.374502,11.279913,12.188754,10.566559,8.913498,8.155559,8.447074,9.153569,8.937505,9.3764925,9.115844,8.687145,10.497967,11.670886,11.948683,11.369082,10.518545,10.511685,10.840926,11.540562,11.838936,11.670886,11.674315,11.05699,11.413667,12.6586075,13.738928,12.614022,10.635151,9.908078,10.257896,11.266195,12.257345,13.13532,12.871242,12.267634,11.976119,12.483699,11.821788,11.05356,11.070708,12.003556,13.214201,13.245067,13.125031,13.454271,14.201921,14.723219,14.634049,14.7095,14.342535,13.817808,14.321958,16.149927,18.87302,20.083664,19.294859,17.929884,18.420315,19.329155,20.011642,19.932762,18.670673,17.003895,17.655516,17.96761,17.511473,18.094503,19.94648,20.330595,19.634388,18.403166,17.329706,17.960749,18.406595,19.507494,21.321745,23.118849,19.28457,18.320856,18.516342,19.246845,20.94792,21.43835,23.61957,25.032558,24.888515,24.082563,25.142305,25.18346,23.478956,21.273731,21.767591,21.747015,21.767591,21.548098,21.249723,21.493225,0.71678376,0.58302987,0.59674823,0.6379033,0.6962063,0.85396725,1.097468,1.0871792,1.0323058,1.0494537,1.1592005,1.6221949,1.5021594,1.3478279,1.4472859,1.8005334,1.4953002,1.529596,1.4918705,1.430138,1.845118,1.821111,1.7799559,2.0406046,2.6373527,3.2958336,4.0777793,5.579939,6.2212715,5.9400454,6.193835,7.2947326,8.4093485,9.3079,11.005547,15.776102,14.874121,9.283894,4.619654,2.719663,1.6324836,0.864256,0.864256,1.646202,2.411,1.5570327,0.77508676,0.70649505,1.0666018,1.3821237,0.9911508,1.2860953,1.1660597,0.7579388,0.31895164,0.26064864,0.33266997,0.4046913,0.4424168,0.40126175,0.24350071,0.17147937,0.18862732,0.31895164,0.52815646,0.7476501,0.72364295,0.58988905,0.490431,0.4664239,0.4424168,0.31895164,0.216064,0.15090185,0.15090185,0.274367,0.2503599,0.18862732,0.17833854,0.21263443,0.21263443,0.16462019,0.09602845,0.12689474,0.20577525,0.106317215,0.058302987,0.082310095,0.09602845,0.082310095,0.106317215,0.17833854,0.116605975,0.041155048,0.024007112,0.061732575,0.12346515,0.14747226,0.1097468,0.058302987,0.106317215,0.20577525,0.26407823,0.44927597,0.91569984,1.8313997,2.393852,3.3198407,3.6319332,3.3609958,3.5564823,4.057202,3.9165888,4.2938433,5.164959,5.3261495,4.8254294,4.835718,4.5853586,3.9680326,3.5393343,3.1860867,2.8499873,2.4967396,2.2669573,2.486451,3.5599117,4.7808447,5.579939,5.3398676,3.3884325,2.301253,2.1469216,2.3389788,2.1469216,0.71678376,0.48357183,0.31895164,0.39783216,0.7339317,1.1763484,0.89512235,0.6241849,0.86082643,1.1660597,0.15090185,0.09259886,0.048014224,0.024007112,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09259886,0.20920484,0.12346515,0.14747226,0.09602845,0.061732575,0.058302987,0.044584636,0.14404267,0.37725464,0.6893471,0.8505377,0.47328308,0.37382504,0.45270553,0.5418748,0.5693115,0.53501564,0.6790583,0.69963586,0.72364295,0.8505377,1.1454822,1.7559488,2.2841053,3.0043187,3.9611735,4.972902,6.4887795,8.268735,10.007536,11.502836,12.648318,13.725209,14.284232,15.419425,17.343424,19.394318,20.11453,21.054237,22.017952,23.643576,27.405834,30.0912,31.538486,33.164112,35.215004,36.789185,36.044964,34.72457,33.472775,33.781437,37.97925,42.55775,43.31569,42.688076,42.701794,44.982468,54.088024,62.802605,74.43577,82.06317,68.52659,40.794945,20.237995,8.333898,4.448175,5.830299,5.1580997,5.2644167,5.610805,6.3893213,8.515666,11.516555,13.841815,15.302819,15.536031,14.023583,23.043398,28.153484,32.488483,38.14044,46.172535,49.22487,70.419716,66.47569,40.187904,40.42112,24.051697,20.882757,18.313997,14.016724,15.944152,13.296511,13.906977,15.536031,17.569777,21.009653,20.145397,16.897577,15.090185,14.997586,13.337666,10.55284,9.280463,11.015835,13.1593275,9.033533,8.021805,6.660259,5.8543057,6.7391396,10.683165,14.527733,12.411677,12.346515,14.832966,12.878101,13.841815,14.750656,13.817808,13.406258,20.03565,24.77191,30.25925,28.311245,25.162884,41.456852,37.869503,22.827333,11.382801,10.13786,17.240536,12.542002,22.683292,32.24841,35.060673,34.196415,38.723473,37.687737,37.74947,40.376534,41.840965,37.543694,38.949825,37.66716,33.122955,32.563934,23.393215,22.741594,26.411253,29.453297,26.167753,28.67135,34.90977,34.450207,26.634176,20.553518,19.809298,23.221737,22.885637,17.857862,14.160767,14.565458,15.6526375,17.501184,19.12681,18.478617,16.088194,12.432255,9.482809,8.169277,8.378482,4.372724,2.8122618,2.2326615,1.8382589,1.4953002,1.2895249,1.0425946,0.7682276,0.5007198,0.30523327,0.25721905,0.18862732,0.12346515,0.06516216,0.01371835,0.041155048,0.12689474,0.5693115,1.0837497,0.84024894,1.0940384,1.8554068,2.503599,2.7299516,2.5481834,2.085189,3.7725463,6.324159,8.131552,7.2775846,4.7774153,2.5653315,1.9514352,3.1483612,5.3090014,7.4970784,8.158989,8.375052,8.354475,7.4627824,6.48535,4.6848164,3.275256,3.3541365,5.90575,5.4770513,6.368744,6.7974424,6.1629686,5.051782,1.4369972,0.8711152,1.2895249,2.1915064,4.6676683,7.380472,6.1629686,5.0003386,5.312431,5.936616,6.0806584,7.548522,7.0958166,5.051782,5.295283,7.051232,7.7851634,7.2467184,5.9983487,5.3878818,4.8734436,5.2575574,6.252138,7.507367,8.604835,9.129561,8.573969,7.257007,5.6005163,4.1360826,4.170378,4.6676683,4.99005,5.0243454,5.1580997,7.1952744,6.7459984,6.4133286,6.910619,7.034084,6.728851,6.725421,6.608815,6.420188,6.6533995,5.528495,5.5593615,5.6039457,5.6039457,6.591667,7.4696417,7.7714453,7.682276,7.421627,7.2638664,8.337327,7.6445503,6.7357097,6.608815,7.720001,6.927767,6.8385973,6.6568294,6.142391,5.6313825,5.56965,5.0586414,4.8288593,4.8014226,4.105216,3.9337368,4.0023284,4.1360826,4.2183924,4.180667,4.1429415,4.190956,4.1155047,4.016047,4.273266,4.064061,3.782835,3.8274195,4.07435,3.8925817,3.806842,4.0949273,4.187526,3.9371665,3.6319332,2.702515,2.3252604,2.037175,1.7765263,1.862266,2.1434922,2.1126258,1.9514352,1.7902447,1.6942163,1.7662375,1.7113642,1.5776103,1.5055889,1.7250825,1.5913286,1.7319417,2.061182,2.311542,2.0440342,1.7388009,1.7079345,1.7319417,1.6187652,1.1900668,1.1420527,1.2380811,1.3855534,1.5433143,1.7388009,1.5433143,1.4575747,1.4781522,1.6427724,2.0440342,2.1674993,2.3629858,2.393852,2.2052248,1.937717,1.7422304,1.4267083,1.196926,1.1146159,1.1146159,0.881404,0.83338976,0.881404,0.91912943,0.8093826,1.1249046,1.2037852,1.1146159,1.0220171,1.2037852,1.2312219,1.0528834,0.85739684,0.83338976,1.1763484,1.1489118,0.9877212,0.86082643,0.7579388,0.48700142,0.37725464,0.37039545,0.40126175,0.4389872,0.48700142,0.37725464,0.4424168,0.4424168,0.33266997,0.26064864,0.22292319,0.26064864,0.40126175,0.66191036,1.0528834,0.9431366,0.99801,1.138623,1.3272504,1.5707511,1.8999915,2.3492675,2.9048605,3.5461934,4.2423997,4.180667,4.3590055,4.698535,4.9591837,4.715683,5.4976287,6.2144127,6.989499,7.48336,6.8969,6.5059276,7.0032177,7.658269,8.172707,8.697433,8.110974,8.488229,9.438225,10.381361,10.528833,9.345626,8.086967,7.507367,7.881192,9.016385,9.458802,10.419086,10.175586,9.2153015,10.254466,11.976119,12.130451,11.341646,10.521975,10.864933,10.960961,11.427385,11.231899,10.768905,11.856084,10.978109,10.336777,10.635151,11.478829,11.369082,11.002116,10.882081,11.094715,11.842365,13.443983,13.334236,12.46312,11.499407,11.447963,13.656617,14.791811,13.519434,11.650309,10.820349,12.4802685,13.166186,13.776653,14.88098,16.088194,16.050468,15.954441,15.326826,14.654627,14.750656,16.739817,19.435472,20.79016,21.644127,21.640697,19.20912,18.54035,18.855871,19.582945,20.135109,19.929333,17.70696,17.21653,17.916164,18.814716,18.44775,19.754423,19.246845,19.041069,19.490345,19.20912,18.893597,18.135658,18.855871,20.906765,22.079683,19.905325,20.069946,20.423193,20.251715,20.265432,21.20514,22.875349,23.657295,23.009102,21.469217,19.895037,20.344313,21.417774,22.659285,24.552416,22.974806,21.328604,19.709839,18.574646,18.722118,0.607037,0.6207553,0.64476246,0.7099246,0.8093826,0.939707,1.0871792,1.1454822,1.1832076,1.2758065,1.5124481,1.587899,1.6804979,1.6770682,1.6187652,1.728512,1.6084765,1.6873571,1.7147937,1.7182233,2.0165975,2.2841053,2.1332035,2.136633,2.5653315,3.3815732,4.07435,5.1821065,5.4667625,5.1409516,5.8645945,6.4064693,6.8283086,7.589677,10.278474,17.62122,17.021042,10.604284,4.787704,2.1503513,1.4267083,1.4267083,1.5913286,1.6599203,1.5158776,1.1900668,1.1797781,1.2826657,1.2620882,1.0185875,0.58988905,0.7442205,0.58645946,0.44584638,0.47328308,0.6241849,0.58302987,0.4424168,0.31895164,0.2503599,0.20920484,0.20234565,0.33266997,0.48014224,0.59331864,0.6859175,0.69963586,0.66533995,0.6241849,0.59331864,0.53844523,0.4081209,0.23664154,0.14404267,0.20577525,0.44584638,0.32238123,0.23664154,0.1920569,0.18519773,0.22635277,0.31209245,0.39097297,0.36696586,0.2469303,0.12003556,0.1097468,0.13032432,0.14747226,0.14747226,0.14404267,0.1371835,0.07545093,0.041155048,0.06516216,0.1097468,0.10288762,0.116605975,0.14404267,0.20920484,0.37382504,0.5212973,0.5796003,0.6859175,0.91912943,1.3169615,2.0749004,2.9631636,3.5187566,3.8274195,4.5201964,4.7842746,4.746549,4.8322887,5.2575574,6.0223556,5.7068334,5.579939,4.8322887,3.9337368,4.6402316,3.6593697,3.2203827,2.7951138,2.5001693,3.059192,2.386993,3.2375305,4.420738,4.722542,2.8877127,1.8005334,2.095478,2.5824795,2.393852,0.9842916,0.823101,0.5693115,0.5212973,0.8025235,1.371835,1.138623,0.8505377,1.1077567,1.4095604,0.15090185,0.061732575,0.07888051,0.082310095,0.044584636,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.044584636,0.0548734,0.09945804,0.17490897,0.25721905,0.15433143,0.1097468,0.1371835,0.23321195,0.38754338,0.42526886,0.48014224,0.53158605,0.5521636,0.4972902,0.5658819,0.72021335,0.805953,0.83338976,0.9602845,1.1180456,1.1660597,1.1763484,1.2072148,1.3169615,2.0028791,2.7573884,3.5359046,4.3692946,5.353586,6.9346256,9.280463,11.619442,13.495427,14.760944,15.944152,16.897577,18.653526,20.824455,21.61669,22.823904,23.869928,24.250612,24.572994,26.575872,28.695358,30.574772,32.642815,34.56338,35.23901,34.6697,32.389023,30.75654,32.43704,40.39711,43.411716,42.90071,40.836098,40.726353,47.619823,56.265812,66.005844,74.675835,74.36717,51.426662,27.069735,13.670336,7.473071,5.909179,7.610255,6.999788,6.8557453,6.6465406,7.1232533,10.319629,14.184773,14.644339,15.4914465,16.955881,15.707511,22.961088,28.787956,33.69227,38.66174,45.16081,42.24566,51.03912,50.565838,38.576,31.521338,21.177702,20.430052,18.78385,15.9578705,21.891056,13.509145,16.62664,18.78385,16.259674,14.064738,13.656617,10.81006,9.194724,9.736599,10.624862,9.201583,8.735159,15.453721,21.997374,7.4353456,6.9380555,5.8988905,5.813151,7.425057,10.693454,10.789482,9.822338,9.956093,11.47197,12.782072,11.694893,12.171606,12.068718,13.090735,20.803877,19.29143,24.562706,22.823904,19.414894,38.795494,31.34986,21.548098,12.9638405,9.136421,13.557159,14.802099,18.530062,23.873358,29.806545,35.112118,36.32962,29.741383,27.505291,33.486492,43.22995,36.130703,33.387035,32.19011,30.5199,27.155474,22.751883,23.458378,23.406935,21.28059,20.310017,21.805317,23.917942,23.972816,21.87048,20.076805,18.005335,17.233677,15.05246,11.509696,9.410788,9.3936405,9.956093,10.323058,10.463672,11.05699,12.092726,11.650309,10.185875,8.182996,6.142391,3.7211025,2.5207467,1.8519772,1.3649758,1.0323058,0.90198153,0.7579388,0.5796003,0.3806842,0.19548649,0.12689474,0.106317215,0.09259886,0.07545093,0.06516216,0.07888051,0.12689474,0.38754338,0.7373613,0.764798,1.2380811,2.270387,2.726522,2.3492675,1.7662375,3.1209247,4.139512,6.159539,8.419638,8.083538,5.6313825,2.4075704,1.646202,3.7759757,6.444195,9.119273,11.9040985,14.980438,17.137648,15.786391,10.034973,7.6342616,6.608815,6.118384,6.4407654,6.2692857,6.8797526,6.917478,6.125243,5.3570156,1.546744,0.6036074,1.0597426,1.728512,1.728512,3.7725463,3.9200184,4.1017866,4.911169,5.5833683,5.7582774,6.540223,6.094377,5.147811,7.0032177,8.14527,7.9429245,6.7802944,5.501058,5.3981705,5.90232,6.012067,6.9037595,8.460793,9.266746,8.783174,7.8983397,6.550512,5.329579,5.4667625,5.4736214,5.1340923,5.0174866,5.06893,4.6093655,6.245279,6.118384,5.744559,5.785714,6.046363,6.619104,6.893471,6.461343,5.686256,5.7136927,5.0586414,5.0655007,5.329579,5.6005163,5.7994323,6.2487082,6.4407654,6.684266,7.0272245,7.2878733,8.107545,7.490219,6.5950966,6.23499,6.866034,5.9469047,6.046363,6.135532,5.785714,5.164959,4.6676683,4.2869844,4.2081037,4.197815,3.6285036,3.57363,3.6044965,3.6627994,3.690236,3.642222,3.4913201,3.4192986,3.3609958,3.391862,3.7348208,3.8788633,3.7759757,3.6868064,3.673088,3.5976372,3.5221863,3.57363,3.4776018,3.1723683,2.7882545,2.136633,1.9925903,2.095478,2.2155135,2.153781,2.0063086,1.9102802,1.7525192,1.529596,1.3649758,1.4953002,1.587899,1.5638919,1.488441,1.5398848,1.4644338,1.4507155,1.5330256,1.821111,2.5070283,1.9582944,1.670209,1.5227368,1.3238207,0.7990939,1.2792361,1.4644338,1.4747226,1.4164196,1.3992717,1.3203912,1.4918705,1.6324836,1.7182233,1.9823016,2.1743584,2.5619018,2.7299516,2.4830213,1.8519772,1.5090185,1.3066728,1.255229,1.255229,1.0906088,0.9842916,0.8779744,0.8505377,0.91569984,1.039165,1.2312219,1.255229,1.1489118,0.99801,0.9362774,1.371835,1.3615463,1.1489118,0.99801,1.2106444,1.2072148,0.9534253,0.66191036,0.432128,0.28122616,0.25721905,0.26407823,0.29837412,0.34981793,0.37725464,0.42526886,0.4046913,0.35324752,0.31552204,0.31895164,0.3018037,0.2777966,0.33609957,0.52472687,0.85739684,1.1592005,1.2209331,1.2620882,1.3924125,1.6084765,1.937717,2.4075704,2.8328393,3.216953,3.765687,4.1360826,4.4275975,4.557922,4.506478,4.3007026,4.846007,5.7102633,6.310441,6.416758,6.15268,6.094377,6.351596,6.8969,7.5245147,7.8537555,7.8846216,8.399059,9.122703,9.544542,8.930646,8.508806,7.7028537,7.099246,7.2467184,8.663138,9.630281,10.789482,11.489118,11.393089,10.497967,12.151029,13.049581,12.620882,11.694893,12.524854,12.113303,10.597425,9.822338,9.945804,9.451943,8.680285,9.362774,10.652299,12.020704,13.258785,11.64345,12.082437,12.185325,11.537132,11.7086115,11.502836,11.530273,12.22305,13.488567,14.730078,15.367981,14.901558,13.965281,13.440554,14.445422,15.217079,16.540901,18.008764,18.910746,18.20082,18.279701,17.473747,16.726099,16.606062,17.336565,17.71039,20.237995,22.271742,22.456938,20.759293,21.074816,21.074816,21.170843,21.650986,22.673002,19.984205,19.53493,19.360022,18.87302,18.886738,18.924463,17.929884,17.923023,19.065077,19.675543,19.795578,18.584934,17.840714,18.430603,20.296299,20.546658,20.567236,19.524641,18.272842,19.360022,20.330595,21.19485,21.407484,20.968498,20.457489,19.836735,19.641247,20.03222,20.985645,22.28203,22.230585,22.309467,21.43835,19.764713,18.660385,0.5796003,0.6790583,0.67219913,0.70306545,0.8128122,0.9328478,1.0940384,1.1934965,1.2209331,1.2860953,1.6221949,1.670209,1.8965619,1.9274281,1.7662375,1.8005334,1.7559488,1.7079345,1.6942163,1.7490896,1.8862731,2.287535,2.4898806,2.644212,2.8328393,3.0626216,3.4878905,4.523626,4.945465,4.7362604,5.086078,5.1100855,5.669108,6.64997,8.81404,13.786942,13.344524,9.383351,5.144381,2.4247184,1.5844694,1.605047,1.4335675,1.3512574,1.471293,1.7593783,1.8519772,1.4781522,1.0048691,0.6241849,0.33266997,0.36010668,0.34638834,0.4046913,0.5007198,0.45270553,0.41498008,0.29837412,0.23664154,0.26750782,0.34638834,0.42869842,0.48014224,0.4972902,0.51100856,0.5693115,0.5658819,0.5453044,0.5590228,0.5796003,0.51100856,0.4424168,0.37725464,0.37725464,0.44584638,0.5624523,0.42869842,0.34295875,0.29494452,0.28808534,0.32924038,0.42183927,0.48357183,0.4698535,0.37725464,0.2503599,0.15433143,0.2194936,0.30523327,0.33609957,0.31895164,0.2503599,0.116605975,0.044584636,0.06516216,0.11317638,0.12346515,0.17833854,0.23321195,0.3018037,0.45956472,0.85396725,1.0906088,1.2860953,1.4953002,1.7113642,2.5481834,3.7348208,4.6265135,5.3707337,6.9209075,6.5779486,6.557371,5.796003,4.7259717,5.2609873,5.007198,4.763697,4.098357,3.4055803,3.923448,3.192946,2.7333813,2.6407824,2.8534167,3.1415021,2.1915064,2.428148,3.1449318,3.4604537,2.3046827,1.488441,1.786815,2.294394,2.287535,1.2346514,1.2517995,1.097468,0.8505377,0.7339317,1.1351935,1.0563129,0.89512235,1.0220171,1.1283343,0.22635277,0.14404267,0.31895164,0.41840968,0.32581082,0.14404267,0.06516216,0.030866288,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.0548734,0.09602845,0.12689474,0.13375391,0.15433143,0.23321195,0.40126175,0.4046913,0.31895164,0.32581082,0.44584638,0.5453044,0.48357183,0.548734,0.67219913,0.77508676,0.7682276,0.864256,0.7922347,0.8745448,1.1694894,1.4815818,1.4850113,1.4164196,1.4232788,1.5055889,1.5124481,1.8691251,2.5756202,3.3301294,4.2115335,5.658819,7.805741,10.343636,13.330807,16.335125,18.410025,19.78186,21.016512,22.347193,23.626429,24.322634,25.505842,25.996273,26.054577,26.411253,28.242653,28.705647,30.351849,31.974045,33.352737,35.26302,35.359047,31.195528,29.048605,32.11466,40.48628,42.73266,44.13193,44.37543,46.076508,54.77737,60.41218,68.06359,73.03649,67.398254,39.99242,20.21399,11.276484,8.114404,7.4765005,7.9189177,7.1884155,7.3427467,7.534804,8.114404,10.597425,14.04759,14.812388,15.275383,16.12592,16.338554,28.026588,29.470446,30.190659,35.18071,44.907017,38.404522,39.388813,41.209923,39.779785,33.57223,22.251163,25.889956,26.26378,21.44178,25.77335,14.730078,14.815818,15.728088,13.186764,8.940934,8.56025,7.191845,7.3701835,9.0369625,9.544542,8.042382,9.349055,15.014734,19.558937,10.477389,8.447074,5.7754254,4.4104495,5.4633327,9.194724,7.795452,6.7940125,7.023795,8.354475,9.671436,8.388771,12.164746,13.570878,13.639469,21.85676,17.844143,26.472986,24.425522,15.477728,30.50618,26.10945,19.315437,12.936404,10.81006,17.823566,17.857862,17.226818,19.054789,23.69845,28.729654,33.77115,29.076042,26.469557,29.974594,35.81518,28.719366,25.77678,26.466127,27.361248,22.141417,22.035099,22.666143,21.342323,18.488907,17.645227,17.031332,18.310568,19.54179,19.576086,18.073925,18.70154,29.84427,31.84029,22.28546,16.033321,13.742357,10.662587,8.467651,7.7783046,8.1487,10.024684,9.496528,8.443645,7.606825,6.5813785,4.9008803,2.7951138,1.4953002,1.2072148,1.097468,0.64476246,0.4389872,0.31895164,0.24350071,0.28808534,0.082310095,0.034295876,0.058302987,0.13375391,0.28808534,0.2194936,0.6276145,1.2003556,1.5158776,1.039165,1.1043272,1.5673214,1.9685832,2.1503513,2.2498093,3.2958336,3.758828,5.470192,8.351046,10.436234,8.375052,4.2526884,2.7299516,4.5510626,6.5642304,7.6033955,13.032433,19.775002,23.338343,17.830425,11.002116,11.365653,10.861504,8.100685,8.344186,7.157549,7.082098,7.4010496,7.6514096,7.610255,3.0866287,1.1866373,1.1489118,1.9857311,2.4761622,4.383013,4.540774,5.1340923,6.2692857,5.9400454,6.111525,6.4236174,5.9400454,5.796003,9.187865,8.361334,7.1266828,6.193835,5.8543057,5.9880595,5.8645945,6.094377,7.1678376,8.591117,8.899779,7.5519514,7.1129646,6.5950966,6.1046658,6.869464,6.23156,5.4976287,5.2164025,5.188966,4.4516044,5.161529,5.2987127,5.3844523,5.7239814,6.4133286,6.7802944,6.711703,6.3721733,5.9400454,5.6245236,5.6142344,5.4736214,5.5422134,5.785714,5.802862,6.012067,6.3653145,6.790583,7.116394,7.06495,7.425057,6.807731,6.135532,5.892031,6.111525,5.658819,5.9228973,5.8680243,5.2918534,4.8494368,4.2698364,3.8685746,3.6868064,3.5839188,3.2443898,3.2409601,3.1655092,3.0969174,3.1072063,3.2272418,3.1517909,3.1723683,3.223812,3.3198407,3.5564823,3.683377,3.5393343,3.357566,3.292404,3.4055803,3.3781435,3.069481,2.5961976,2.1880767,2.194936,1.7833855,1.6256244,1.7079345,1.920569,2.037175,1.8828435,1.6496316,1.4918705,1.4164196,1.2998136,1.2860953,1.4061309,1.4747226,1.4678634,1.5227368,1.3443983,1.3581166,1.9102802,2.7882545,3.210094,2.1160555,1.4369972,1.138623,1.039165,0.8128122,1.1214751,1.3478279,1.4198492,1.371835,1.3478279,1.4095604,1.5501735,1.728512,1.9239986,2.1434922,2.3561265,2.7059445,2.7230926,2.2806756,1.6221949,1.3443983,1.2963841,1.3066728,1.2380811,1.0014396,0.96371406,0.8779744,0.8676856,0.980862,1.1626302,1.1317638,1.1934965,1.2277923,1.1489118,0.9259886,1.1900668,1.2483698,1.2003556,1.0940384,0.9568549,0.89512235,0.71678376,0.47328308,0.25721905,0.1920569,0.17833854,0.18862732,0.24007112,0.3018037,0.29494452,0.39783216,0.37382504,0.32924038,0.32581082,0.36353627,0.29837412,0.274367,0.31209245,0.42183927,0.607037,0.9294182,1.0666018,1.1626302,1.3306799,1.6633499,1.9857311,2.386993,2.6750782,2.843128,3.069481,3.625074,3.875434,3.9474552,3.9474552,3.9474552,4.262977,5.188966,5.7239814,5.662249,5.6176643,5.7308407,5.90232,6.2727156,6.728851,6.883182,7.3530354,8.128122,8.669997,8.755736,8.491658,7.7542973,7.3393173,7.3221693,7.7920227,8.841476,10.436234,11.55771,12.555719,13.121602,12.260776,12.895248,13.954991,13.749216,12.504276,12.370522,11.821788,10.854645,9.668007,8.580828,8.025234,7.6857057,7.9737906,8.663138,9.935514,12.404818,11.451392,11.489118,11.646879,11.485688,11.002116,11.276484,11.924676,12.850664,14.13676,16.060759,16.588915,16.21852,15.642348,15.37827,15.745236,16.777542,18.20768,19.260563,19.61038,19.360022,18.917604,18.20768,17.339994,16.640358,16.643787,17.521763,19.586374,21.825895,22.978235,21.561817,21.822466,21.146837,20.316875,19.94648,20.488356,19.53836,19.435472,18.831865,17.641798,17.04848,17.04505,16.907866,17.309128,18.265984,19.140528,19.884748,18.986197,18.62266,19.37031,20.207129,18.71183,17.61436,16.832415,16.7844,18.403166,20.090523,20.416334,20.138538,19.816156,19.79901,19.486916,19.065077,18.488907,18.362011,19.963629,20.316875,20.526081,20.056227,18.897026,17.583494,0.6790583,0.77851635,0.75450927,0.805953,0.9602845,1.0631721,1.138623,1.214074,1.2277923,1.2689474,1.6016173,1.728512,1.961724,1.9823016,1.8142518,1.8485477,1.845118,1.762808,1.762808,1.8176813,1.7456601,2.1126258,2.609916,2.8465576,2.784825,2.7230926,3.0111778,3.923448,4.623084,4.773986,4.537344,4.2183924,5.164959,6.310441,7.5210853,9.589127,13.522863,14.177915,11.382801,6.4990683,2.4075704,1.6153357,1.1592005,1.2106444,1.6324836,1.9823016,1.7765263,1.1454822,0.6001778,0.32581082,0.1920569,0.16462019,0.2194936,0.34295875,0.47328308,0.4938606,0.39097297,0.26750782,0.22978236,0.30866286,0.4355576,0.53501564,0.50757897,0.42526886,0.37725464,0.44927597,0.47328308,0.4081209,0.39097297,0.42869842,0.42869842,0.44584638,0.4938606,0.53844523,0.5693115,0.6173257,0.44584638,0.4115505,0.4389872,0.4698535,0.432128,0.5007198,0.52472687,0.5521636,0.5590228,0.432128,0.33952916,0.3806842,0.44584638,0.4629943,0.41498008,0.30866286,0.16462019,0.09945804,0.11317638,0.11317638,0.16804978,0.24007112,0.31895164,0.41840968,0.6001778,1.2758065,1.6153357,1.903421,2.2292318,2.486451,3.1792276,4.636802,5.874883,6.8797526,8.601405,7.0958166,6.2418494,5.051782,3.8308492,4.173808,4.2081037,4.0880685,3.57363,2.9220085,2.9048605,2.836269,2.5070283,2.5481834,2.860276,2.5893385,2.2360911,2.1400626,2.5310357,3.2478194,3.7313912,2.095478,1.862266,2.0131679,1.9411465,1.4507155,1.3169615,1.1489118,0.8848336,0.67219913,0.85396725,0.83338976,0.8128122,0.9774324,1.0528834,0.32238123,0.26407823,0.40126175,0.52815646,0.5178677,0.29494452,0.14404267,0.06516216,0.024007112,0.006859175,0.006859175,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.05144381,0.07888051,0.106317215,0.14061308,0.17833854,0.2469303,0.2194936,0.2469303,0.432128,0.85739684,0.7442205,0.50757897,0.4629943,0.65162164,0.8196714,0.58302987,0.72021335,0.84367853,0.8711152,1.0323058,1.0254467,0.8162418,0.8711152,1.255229,1.670209,1.5193073,1.5090185,1.5536032,1.6187652,1.728512,2.085189,2.6064866,3.450165,4.715683,6.4407654,9.431366,11.8869505,15.175924,19.092514,21.846472,23.324625,24.35007,24.710178,24.662163,24.909094,26.462696,28.163773,28.702217,28.283808,28.623337,28.369547,29.305824,30.122066,30.962317,33.40761,34.055805,29.7551,28.544456,32.886314,39.64603,41.772377,45.270554,47.46892,49.927933,58.460747,61.211277,66.84609,68.279655,58.906593,32.605087,17.165085,10.151579,7.915488,7.5759587,7.0478024,6.2384195,6.708273,7.888051,9.448513,11.324498,13.193623,14.054449,14.260224,14.472859,15.642348,27.392115,25.43382,23.712168,28.829113,40.047295,34.40219,35.043526,37.862644,38.137012,30.547335,20.827885,25.917393,26.52443,20.220848,21.44864,14.935853,12.830087,13.642899,13.732068,7.3255987,6.5127864,6.375603,7.2638664,8.700864,9.379922,7.486789,8.525954,11.406808,13.838386,12.319078,10.052121,6.9071894,4.3178506,3.899441,7.4799304,6.368744,4.7945633,5.15467,6.869464,6.385892,5.5662203,14.538021,17.12393,13.749216,21.428062,17.267973,26.706198,24.682741,13.111313,20.886189,20.104242,15.46744,12.768354,16.074476,27.717926,21.242865,18.265984,16.513464,16.304258,20.570665,25.348082,26.953129,26.34609,24.94339,24.590141,18.71526,18.653526,21.074816,22.69701,20.296299,22.223726,22.926792,21.688711,19.312008,18.115082,16.187653,17.916164,19.233126,18.053349,14.284232,17.511473,31.027477,34.08667,24.590141,19.054789,15.426285,10.580277,7.613684,7.0546613,6.8728933,7.9875093,7.0923867,6.48535,6.5985265,5.98463,5.0243454,3.707384,2.4212887,1.430138,0.8745448,0.432128,0.29837412,0.29837412,0.37382504,0.5796003,1.3375391,1.2517995,1.1832076,1.5981878,2.5824795,1.903421,2.0817597,2.4727325,2.4830213,1.5913286,1.0494537,1.2003556,1.6221949,2.177788,3.0248961,2.7985435,3.4364467,5.0620713,7.6514096,11.015835,10.127572,5.645101,3.1792276,4.331569,6.6739774,5.7822843,12.418536,20.388897,24.007113,18.087645,13.666906,15.151917,14.249936,10.257896,10.076128,7.7611566,7.016936,7.630832,9.153569,10.899229,5.586798,2.5790498,2.0920484,3.350707,4.5922174,5.7994323,5.7719955,6.169828,6.999788,6.5950966,6.5196457,6.708273,6.228131,6.2418494,10.024684,8.937505,7.281014,6.5024977,6.677407,6.5127864,5.662249,5.720552,6.8043017,8.244728,8.611694,6.931196,7.0135064,7.250148,7.116394,7.1678376,6.420188,5.8988905,5.4599032,4.996909,4.482471,4.523626,4.6608095,5.0277753,5.7102633,6.7357097,6.492209,6.2658563,6.2898636,6.3447366,5.73427,5.861165,5.5079174,5.552502,6.029215,6.108095,6.101236,6.5196457,6.8214493,6.869464,6.931196,6.9826403,6.4819202,6.0840883,5.953764,5.73427,5.501058,5.7308407,5.5079174,4.8117113,4.5270553,4.0709205,3.8102717,3.6319332,3.450165,3.2066643,3.0146074,2.8396983,2.784825,2.867135,3.0043187,3.083199,3.2443898,3.3609958,3.3952916,3.3952916,3.3781435,3.1552205,2.959734,2.9322972,3.1140654,2.9460156,2.609916,2.170929,1.8073926,1.8142518,1.6599203,1.5227368,1.4815818,1.5433143,1.6324836,1.5261664,1.3409687,1.3101025,1.4129901,1.3478279,1.3203912,1.3958421,1.4129901,1.3512574,1.3341095,1.1797781,1.3169615,2.136633,3.1552205,2.9974594,1.8691251,1.2826657,1.0528834,1.0151579,1.0117283,1.1180456,1.3203912,1.488441,1.5776103,1.6530612,1.6427724,1.670209,1.8931323,2.2120838,2.2635276,2.4658735,2.8328393,2.7059445,2.0680413,1.5536032,1.3306799,1.313532,1.2758065,1.1351935,0.9294182,0.91569984,0.91912943,0.939707,1.0254467,1.2483698,1.2689474,1.3066728,1.3169615,1.2758065,1.1694894,1.2037852,1.138623,1.0666018,0.96371406,0.6756287,0.5624523,0.47328308,0.33609957,0.18862732,0.16804978,0.16804978,0.1920569,0.22635277,0.2469303,0.24007112,0.3566771,0.37039545,0.33609957,0.30866286,0.36353627,0.28465575,0.2709374,0.30523327,0.36353627,0.41840968,0.64819205,0.8676856,1.0666018,1.2929544,1.646202,1.9137098,2.1983654,2.3904223,2.486451,2.5584722,3.018037,3.3061223,3.3712845,3.357566,3.5942078,3.865145,4.6127954,5.0106273,4.962613,5.099797,5.1821065,5.363875,5.672538,5.9812007,6.012067,6.543653,7.449064,7.953213,7.953213,8.021805,7.267296,7.4181976,7.8434668,8.330468,9.071259,10.573419,11.729189,13.022143,14.225929,14.387119,14.417986,14.750656,14.325387,13.077017,11.938394,10.772334,10.72089,9.640571,7.7131424,7.4456344,7.2707253,7.14726,6.9380555,7.7371492,11.880091,11.825217,11.365653,11.303921,11.393089,10.323058,11.231899,12.696333,13.72178,14.5414505,16.585485,16.756964,16.832415,17.151367,17.532051,17.264544,17.545769,17.847572,18.070496,18.217968,18.37916,17.53548,17.401728,16.849564,15.920145,15.803539,17.415445,18.759844,20.546658,22.19286,21.805317,21.815605,20.721567,18.969048,17.63151,18.430603,18.608942,18.578075,17.785841,16.331696,14.953001,15.289101,16.338554,17.501184,18.478617,19.274282,19.87446,19.929333,20.35803,20.96164,20.430052,17.974468,16.444872,16.221949,17.089634,18.231688,19.006773,18.732407,18.509483,18.800999,19.46291,19.5315,18.550638,17.261114,16.770683,18.554068,18.694681,18.533491,18.163095,17.36057,15.556609,0.8093826,0.86082643,0.8676856,1.0048691,1.2243627,1.2586586,1.2003556,1.1934965,1.196926,1.2689474,1.5638919,1.6942163,1.8416885,1.9308578,1.920569,1.8313997,1.8279701,1.8176813,1.8862731,1.9308578,1.6496316,1.9720128,2.5310357,2.6407824,2.3801336,2.5619018,3.0111778,3.690236,4.523626,5.07236,4.5167665,3.9474552,5.0483527,6.1972647,7.0889573,8.704293,19.994495,25.396095,22.182571,12.5145645,3.4295874,1.6427724,1.0666018,1.1832076,1.471293,1.430138,0.9362774,0.5212973,0.26064864,0.15090185,0.12346515,0.1097468,0.15433143,0.28122616,0.5007198,0.8162418,0.58645946,0.38754338,0.28122616,0.29151493,0.42869842,0.44584638,0.4115505,0.35324752,0.31209245,0.37039545,0.41498008,0.31552204,0.23321195,0.2469303,0.34981793,0.432128,0.4972902,0.5178677,0.53158605,0.64476246,0.45270553,0.48357183,0.58645946,0.6241849,0.48700142,0.5521636,0.59331864,0.6859175,0.75450927,0.58302987,0.548734,0.4938606,0.4698535,0.4629943,0.3806842,0.28465575,0.22292319,0.20920484,0.21263443,0.17833854,0.26750782,0.34981793,0.5007198,0.7305021,0.97400284,1.8142518,2.1572106,2.49331,2.959734,3.3541365,3.7794054,5.363875,6.848886,7.8366075,8.776315,6.48535,4.431027,3.3369887,3.2718265,3.6216443,4.262977,4.266407,3.6079261,2.6887965,2.3424082,2.8499873,2.726522,2.6819375,2.6819375,1.920569,2.3458378,2.335549,2.9940298,4.6882463,7.0272245,3.3747141,2.2326615,1.8279701,1.4404267,1.4232788,1.0082988,0.7579388,0.66191036,0.6790583,0.70649505,0.58645946,0.64819205,1.0323058,1.2929544,0.39440256,0.40126175,0.33266997,0.37039545,0.4698535,0.36010668,0.28808534,0.14404267,0.044584636,0.020577524,0.01371835,0.0034295875,0.006859175,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.11317638,0.16804978,0.20577525,0.22978236,0.24007112,0.59674823,0.53844523,0.4938606,0.71678376,1.2860953,1.0288762,0.6927767,0.6173257,0.85739684,1.1694894,0.8162418,0.9602845,1.039165,0.9945804,1.2895249,1.2895249,1.0940384,1.0563129,1.2655178,1.5638919,1.5021594,1.6359133,1.6393428,1.605047,2.020027,2.486451,2.8259802,3.8891523,5.658819,7.257007,10.834066,13.416546,16.842705,21.02337,23.921373,25.210897,25.571005,25.01884,24.065414,23.715597,26.239773,29.700228,30.814844,29.055466,26.654755,26.548437,26.260351,26.239773,26.870817,28.469006,29.401854,27.553307,28.969725,34.388474,39.25506,42.612625,46.666397,48.923065,50.977386,58.501904,59.53078,64.4831,63.539967,51.721607,28.890844,16.324837,9.458802,6.9792104,6.8626046,6.358455,5.802862,5.8680243,7.6959944,10.576848,11.948683,12.144169,12.490558,13.05301,13.704632,14.147048,20.059656,18.420315,17.909306,22.652426,32.24841,28.712505,33.321873,35.66085,30.633076,18.482046,14.46943,18.849012,19.390888,14.054449,10.971251,12.380811,11.907528,14.863832,17.861292,8.80718,6.7665763,6.783724,7.2364297,7.8503256,9.72288,7.7268605,6.6053853,7.4696417,10.443094,14.647768,10.9369545,8.711152,5.9743414,3.6765177,5.703404,6.4819202,4.434457,4.7019644,6.756287,4.420738,4.108646,15.145059,18.005335,12.617453,18.358582,15.635489,23.218307,21.386908,10.823778,12.600305,12.836946,10.772334,12.644889,20.858751,33.983784,22.299177,19.723558,15.46744,9.626852,13.203912,13.358243,20.60839,22.223726,16.681513,13.660047,9.9801,13.2862215,16.345413,17.37429,20.04251,21.976797,23.43094,23.252604,21.757303,20.731855,18.989626,20.821026,20.913624,17.350283,11.612583,13.817808,16.726099,17.137648,15.824117,17.514904,12.500846,9.030104,7.1061053,6.39961,6.245279,6.5333643,7.157549,7.5725293,7.0546613,4.7191124,4.4550343,4.647091,3.7142432,1.8142518,0.8505377,0.91227025,0.9911508,1.1420527,1.3306799,1.4129901,3.0214665,2.8294096,2.5619018,3.1689389,4.8254294,3.7622573,3.5187566,3.508468,3.3472774,2.8568463,2.5893385,2.6545007,2.7813954,3.117495,4.2218223,2.6853669,3.8857226,5.4153185,6.715132,9.050681,9.369633,5.3570156,2.510458,3.3232703,7.2775846,6.0978065,11.461681,18.0362,22.035099,21.215427,20.073376,18.1288,15.062748,11.976119,11.38623,8.89635,7.438775,7.6685576,9.6645775,12.939834,7.963502,4.0846386,3.1106358,4.540774,5.56965,5.6245236,5.953764,6.108095,6.1904054,6.831738,6.39961,6.708273,6.478491,6.3961806,9.122703,9.345626,7.953213,7.133542,7.2295704,6.756287,5.720552,5.2987127,6.2041235,7.857185,8.419638,7.3084507,7.5931067,7.9463544,7.671987,6.6876955,6.23499,6.060081,5.429037,4.5339146,4.4927597,4.372724,4.437886,4.8185706,5.528495,6.4544835,5.9571934,5.8371577,6.217842,6.6568294,6.135532,5.703404,5.2301207,5.545643,6.385892,6.39961,6.183546,6.5127864,6.5470824,6.3618846,6.975781,6.824879,6.601956,6.495639,6.375603,5.7754254,5.377593,5.295283,5.003768,4.48933,4.290414,3.9886103,3.9371665,3.8479972,3.6216443,3.333559,2.867135,2.633923,2.7230926,2.9974594,3.07634,3.2855449,3.4844608,3.5461934,3.4295874,3.1723683,3.0660512,2.8499873,2.6647894,2.603057,2.6819375,2.318401,2.201795,2.1194851,1.9274281,1.5638919,1.6359133,1.5947582,1.488441,1.3649758,1.2380811,1.1523414,1.1694894,1.2860953,1.430138,1.4644338,1.5330256,1.5090185,1.3684053,1.1626302,1.0048691,1.039165,1.2346514,1.8588364,2.4590142,1.8656956,1.3409687,1.2723769,1.2689474,1.2106444,1.2312219,1.371835,1.5227368,1.7113642,1.903421,2.0131679,1.7971039,1.7833855,2.0508933,2.3595562,2.1743584,2.318401,2.7299516,2.6167753,1.99602,1.6770682,1.4129901,1.2586586,1.1283343,1.0014396,0.91912943,0.89855194,0.99801,1.0323058,1.0323058,1.2483698,1.5810398,1.5433143,1.3821237,1.2929544,1.4164196,1.3924125,1.1694894,0.922559,0.72707254,0.5555932,0.3841138,0.31552204,0.26064864,0.20234565,0.19891608,0.22635277,0.25378948,0.24007112,0.20234565,0.22292319,0.31209245,0.36353627,0.34638834,0.3018037,0.32924038,0.28465575,0.26750782,0.29151493,0.33952916,0.34295875,0.5007198,0.7442205,0.9877212,1.2277923,1.5398848,1.7422304,1.8965619,2.0303159,2.1572106,2.2738166,2.4761622,2.860276,2.9322972,2.7985435,3.1723683,3.566771,3.9783216,4.2046742,4.290414,4.5270553,4.530485,4.835718,5.192395,5.3913116,5.2575574,5.6039457,6.478491,7.0615206,7.1781263,7.291303,7.06495,7.6925645,8.210432,8.450503,9.054111,9.764035,11.05699,12.617453,14.123041,15.241087,15.553179,14.915276,14.164196,13.358243,11.770344,9.897789,9.952662,9.304471,7.840037,7.9600725,7.8503256,7.4765005,6.697984,7.1026754,12.020704,12.620882,12.140739,11.80464,11.540562,9.983529,11.002116,13.313659,14.63062,14.856973,16.060759,16.173935,16.499744,17.394867,18.3723,18.104792,16.894148,15.9578705,15.590904,15.673215,15.680074,14.829536,15.350834,15.505165,15.086755,15.443433,17.12736,18.423744,19.668684,20.889618,21.78474,21.352612,20.440342,18.636377,17.134218,18.69811,18.663815,18.1288,17.099922,15.772673,14.527733,15.134769,17.171944,19.325726,20.814167,21.400625,20.94792,21.589252,22.062536,21.750444,20.697561,19.360022,18.20082,18.108221,18.77699,18.725548,17.079346,16.208231,16.424294,17.600643,19.157675,19.912186,18.310568,16.818697,16.743246,18.224829,17.95732,17.532051,17.089634,16.2974,14.356253,0.7476501,0.8093826,0.91569984,1.1111864,1.2826657,1.1592005,1.2209331,1.1180456,1.0631721,1.196926,1.587899,1.5638919,1.6564908,2.0920484,2.4795918,1.8313997,1.7216529,1.611906,1.6839274,1.786815,1.4198492,2.0063086,2.5550427,2.5310357,2.1983654,2.6236343,3.5050385,4.0880685,4.722542,5.23698,4.945465,3.9063,4.5442033,5.7582774,7.98408,13.183334,27.94085,35.293884,29.189219,13.780083,3.4192986,1.8073926,0.9842916,0.65162164,0.5658819,0.5041494,0.31895164,0.20920484,0.12346515,0.06516216,0.07545093,0.05144381,0.28465575,0.5521636,0.7305021,0.77851635,0.6207553,0.45270553,0.29837412,0.24350071,0.42869842,0.31895164,0.32581082,0.39440256,0.4424168,0.3806842,0.22292319,0.20920484,0.216064,0.216064,0.29151493,0.40126175,0.35324752,0.3841138,0.5453044,0.71678376,0.7305021,0.7407909,0.6859175,0.5727411,0.48700142,0.5624523,0.70649505,0.8711152,0.91227025,0.59674823,0.42526886,0.29837412,0.30523327,0.3806842,0.31895164,0.31895164,0.3566771,0.33266997,0.28808534,0.39783216,0.50757897,0.6893471,1.0563129,1.4987297,1.6942163,2.4247184,2.9220085,3.3301294,3.7553983,4.256118,4.57507,6.293293,7.795452,8.337327,8.056101,7.3839016,5.48734,4.280125,4.1943855,4.197815,5.6005163,5.0174866,3.6936657,2.5619018,2.2429502,2.6956558,2.644212,2.843128,3.1037767,2.2738166,2.8945718,3.1620796,4.602506,7.284444,9.81205,4.0846386,2.0680413,1.3615463,0.86082643,0.7613684,0.7510797,0.764798,0.7613684,0.71678376,0.65505123,0.34981793,0.44927597,0.9568549,1.3101025,0.3806842,0.5658819,0.51100856,0.3566771,0.22635277,0.21263443,0.6276145,0.36696586,0.09259886,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0034295875,0.01371835,0.06516216,0.12346515,0.20920484,0.2777966,0.22978236,1.5707511,1.5330256,1.1592005,0.91912943,0.6859175,1.1146159,1.1489118,1.0940384,1.1077567,1.2037852,1.0940384,1.0666018,1.5021594,2.085189,1.8142518,2.4007113,2.0817597,1.8313997,1.8691251,1.6496316,2.270387,2.1057668,1.7216529,1.6770682,2.534465,2.0337453,2.3286898,3.5873485,5.377593,6.684266,9.72288,13.502286,17.679523,21.551527,24.079134,24.627867,24.326063,23.616138,23.201159,24.03112,27.621897,28.499872,28.359259,27.337242,24.0174,22.710728,20.443771,19.682402,20.683842,21.500084,22.734735,24.94682,29.583622,35.84948,40.695484,48.15484,50.751034,52.20175,55.43928,62.58997,62.408203,67.343376,66.31793,53.77936,29.707087,17.562918,10.398509,7.870903,8.22758,8.299602,8.690575,6.6568294,7.346176,10.288762,9.383351,9.836057,10.662587,13.2690735,15.806969,13.183334,14.904987,16.681513,18.334574,21.61669,30.197517,21.602972,25.27949,25.413242,16.931873,5.4941993,4.773986,12.703192,18.766703,16.719238,4.623084,5.6142344,10.151579,16.78783,20.135109,10.8958,6.159539,4.945465,6.368744,8.916927,10.467101,8.735159,6.8728933,7.1781263,12.586586,26.671902,11.976119,9.39021,7.596536,3.6285036,2.884283,7.267296,5.470192,4.7671266,6.0703697,3.9200184,4.1155047,5.861165,7.953213,9.935514,12.085866,12.233338,21.211998,18.581505,5.888602,6.667118,5.363875,7.442205,11.434244,16.101913,20.4472,16.163645,18.259123,15.6526375,8.114404,6.2727156,8.114404,13.282792,12.566009,6.677407,6.2247014,6.824879,9.674867,12.370522,14.061309,15.426285,17.63494,20.001354,22.186,23.640146,23.588703,23.02968,23.345201,22.216867,19.277712,16.12935,10.744898,8.879202,10.875222,16.403717,24.459818,13.265644,11.859513,9.9801,6.0532217,7.1884155,8.663138,14.003006,15.9750185,12.614022,7.233,6.8043017,4.3178506,2.287535,1.8656956,2.8534167,3.450165,3.6182148,3.7965534,3.9268777,3.4638834,2.1812177,1.6427724,1.2517995,0.881404,0.8711152,1.6153357,2.534465,3.4535947,4.4447455,5.7994323,8.423067,7.459353,6.262427,6.2830043,7.06495,4.856296,5.7411294,6.6876955,6.5985265,6.3173003,5.950334,3.415869,1.786815,3.1037767,8.378482,10.587136,12.099585,17.532051,26.1849,32.042637,30.039757,19.267422,11.657167,11.067279,13.289652,12.569438,9.818909,8.272165,8.838047,10.072699,8.532814,4.3487167,2.1091962,2.5790498,2.702515,2.49331,4.0057583,4.6676683,4.40359,5.662249,5.195825,5.521636,6.1561093,6.8385973,7.5210853,7.267296,6.3138704,5.9469047,6.4133286,6.927767,5.9880595,5.4324665,6.385892,7.956643,7.2467184,7.9429245,8.06296,7.6857057,7.1884155,7.2467184,6.111525,5.2609873,4.619654,4.2355404,4.273266,4.2115335,4.746549,5.360445,5.7582774,5.844017,6.2830043,5.8988905,6.1972647,7.2467184,7.675417,6.2830043,6.0532217,6.584808,7.1198235,6.5470824,6.252138,6.591667,6.701414,6.574519,7.051232,6.341307,6.4407654,6.725421,6.715132,6.042933,5.6656785,5.0106273,4.5647807,4.461893,4.4859004,4.1429415,3.8857226,3.5976372,3.2718265,2.9906003,2.6716487,2.4007113,2.585909,3.1483612,3.5393343,3.8102717,3.7931237,3.666229,3.450165,3.0351849,3.0489032,2.976882,2.6990852,2.3286898,2.2429502,2.085189,1.8416885,1.6427724,1.4918705,1.2963841,1.4541451,1.3409687,1.2620882,1.2998136,1.313532,1.4232788,1.4850113,1.4061309,1.3443983,1.7079345,1.611906,1.4129901,1.2037852,1.039165,0.9294182,1.1008976,1.0528834,1.4198492,1.8416885,0.9602845,1.1214751,1.2895249,1.3306799,1.2826657,1.3443983,1.6496316,1.7971039,1.8828435,1.903421,1.7696671,1.611906,1.7456601,1.9239986,1.9651536,1.7696671,1.8073926,1.9342873,1.9891608,1.9068506,1.7250825,1.3821237,1.039165,0.85739684,0.8711152,0.9911508,0.9431366,1.0048691,1.0528834,1.039165,0.9911508,1.4918705,1.5158776,1.3649758,1.2209331,1.1592005,1.1832076,1.2072148,1.0563129,0.7888051,0.70306545,0.3841138,0.2503599,0.23664154,0.28465575,0.31895164,0.31895164,0.274367,0.2503599,0.26064864,0.26064864,0.22292319,0.28808534,0.37382504,0.40126175,0.30523327,0.26750782,0.23321195,0.24350071,0.30523327,0.36696586,0.47671264,0.6036074,0.6962063,0.8711152,1.4198492,1.6496316,1.7079345,1.7456601,1.821111,1.9068506,1.9925903,2.2155135,2.3081124,2.3149714,2.609916,3.0729103,3.3266997,3.5839188,3.8548563,3.9508848,4.170378,4.7945633,5.1409516,4.9660425,4.4413157,4.8082814,5.686256,6.307011,6.5710897,7.034084,7.023795,7.267296,7.8537555,8.519095,8.652849,8.786603,10.038403,11.149589,11.821788,12.7272,13.7526455,13.505715,13.313659,13.114742,11.427385,10.367643,9.534253,8.930646,8.9100685,10.192734,10.97468,9.174147,8.1041155,8.882631,10.422516,12.154458,12.404818,12.600305,12.778643,11.581717,11.262765,13.656617,14.805529,14.2533655,15.059319,17.134218,15.374841,13.72178,13.927555,15.563468,13.865822,14.448852,14.658057,13.824667,13.275933,12.531713,12.80265,13.46799,14.342535,15.6869335,17.576635,20.001354,21.424633,21.661274,21.880768,19.977346,19.895037,20.382038,20.70099,20.61525,20.395756,18.763273,17.069057,16.393429,17.576635,18.3723,21.150267,24.123718,26.10259,26.503853,24.77191,23.715597,22.587263,21.589252,21.880768,21.342323,19.94648,19.428614,19.689262,18.79757,15.7966795,14.750656,15.055889,16.314548,18.341434,19.805868,18.845583,17.61779,17.357141,18.3723,17.809847,17.384579,16.88043,16.61292,17.4566,0.69963586,0.7510797,0.84024894,0.9877212,1.1214751,1.0871792,1.5090185,1.5536032,1.430138,1.3478279,1.5124481,1.371835,1.5193073,1.7456601,1.845118,1.5981878,1.7250825,1.7319417,1.8039631,1.845118,1.4815818,1.762808,1.9720128,2.270387,2.6887965,3.1380725,3.724532,3.9851806,4.6848164,5.4187484,4.6402316,4.400161,5.1238036,6.6636887,9.80519,16.235666,24.120289,25.224615,18.595222,8.1212635,2.551613,1.4575747,0.8128122,0.53844523,0.4629943,0.33266997,0.20920484,0.17833854,0.15090185,0.14404267,0.28465575,1.0220171,1.0906088,1.097468,1.1420527,0.84024894,0.6036074,0.42183927,0.30523327,0.25721905,0.29151493,0.28122616,0.32238123,0.37039545,0.3841138,0.33266997,0.24350071,0.20234565,0.20577525,0.26407823,0.4355576,0.53501564,0.53158605,0.4938606,0.4698535,0.48357183,0.47671264,0.4355576,0.432128,0.5041494,0.6344737,0.64133286,0.8128122,0.8505377,0.6790583,0.44927597,0.33609957,0.432128,0.66533995,0.8848336,0.83338976,0.58988905,0.548734,0.4629943,0.3806842,0.6790583,0.9534253,1.2449403,1.5021594,1.7216529,1.937717,2.49331,3.100347,3.525616,3.7965534,4.1600895,5.2575574,7.0478024,8.021805,7.671987,6.495639,5.528495,4.979761,5.127233,5.579939,5.2575574,4.7774153,3.765687,3.1895163,3.1620796,2.9631636,2.2429502,2.0303159,2.2360911,2.668219,3.0317552,4.4550343,3.8342788,3.806842,5.0414934,6.258997,3.5016088,2.270387,1.6427724,1.2517995,1.2998136,0.6824879,0.5178677,0.6173257,0.7339317,0.5453044,0.48357183,0.70306545,0.8676856,0.7510797,0.22292319,0.24007112,0.29837412,0.31895164,0.28465575,0.21263443,0.28808534,0.18862732,0.09259886,0.06859175,0.061732575,0.01371835,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.13032432,0.28122616,0.32238123,0.39097297,0.88826317,1.255229,0.91912943,0.71678376,0.85396725,0.89512235,0.9877212,1.5021594,1.6496316,1.3786942,1.3889829,0.84024894,0.83338976,1.3855534,1.8965619,1.1694894,1.0220171,0.9431366,1.0494537,1.2655178,1.3306799,1.5227368,1.5947582,1.9823016,2.5996273,2.8499873,1.9102802,2.6545007,4.033195,5.5422134,7.208993,9.983529,14.123041,18.440891,21.78131,23.02968,24.134007,24.075705,23.828773,24.130577,25.447538,27.837961,28.904564,28.808535,27.361248,24.03112,21.054237,17.686382,15.820687,16.616352,20.512363,24.206028,28.76738,33.788296,38.606865,42.331398,48.364044,50.13714,52.71276,56.61563,57.829704,55.940002,60.381317,58.51905,45.28084,23.142857,13.975569,9.002667,6.8626046,6.2967224,6.166398,6.2247014,6.258997,6.245279,6.166398,6.0154963,7.2467184,9.523964,14.160767,17.580065,11.303921,12.264205,15.87899,17.484037,18.087645,24.374079,28.396984,30.194088,24.710178,13.443983,4.4687524,6.90033,10.048691,15.724659,19.140528,8.906639,7.8949103,8.903209,11.187314,12.950122,11.345076,8.1041155,6.8557453,8.008087,9.757176,8.076678,6.2727156,5.501058,6.3618846,10.600855,21.095392,9.513676,6.210983,4.6127954,2.4487255,1.7730967,5.2164025,6.848886,10.573419,13.564018,6.2418494,6.2898636,8.858624,9.818909,8.851766,9.434795,10.813489,18.828436,17.87158,7.9463544,4.65395,7.2432885,11.201033,12.737488,12.442543,15.29596,14.740367,16.321407,14.479718,9.016385,5.0620713,7.2775846,9.571979,8.505377,6.001778,9.338767,14.095605,14.778092,13.516005,12.205902,12.507706,14.356253,16.033321,17.71039,19.174824,19.819586,16.287111,16.362562,18.20425,20.587814,22.878778,24.593573,24.391226,20.471207,14.5585985,11.910957,7.846896,6.677407,7.1781263,8.076678,8.042382,10.446524,12.840376,13.982429,12.250486,5.645101,6.118384,5.809721,3.923448,1.8931323,3.391862,2.8259802,3.2546785,3.4981792,3.5221863,4.417309,4.139512,4.4516044,3.7451096,2.3767042,2.6750782,3.508468,4.105216,5.5113473,7.8263187,10.216741,10.556271,9.561689,9.283894,9.80519,9.235879,8.522525,7.143831,6.475061,6.632822,6.4990683,5.744559,5.7239814,5.2266912,4.9694724,7.596536,8.663138,10.556271,16.300829,24.542128,29.552755,24.19231,16.650646,13.138749,14.661487,17.04848,15.169065,12.63803,10.693454,10.377932,12.548861,9.935514,6.0635104,4.40359,4.4721823,1.8108221,2.4418662,3.7108135,4.870014,5.768566,6.869464,6.307011,5.720552,6.046363,6.9620624,6.8626046,6.7048435,5.6005163,5.411889,6.1904054,6.193835,6.262427,6.9963584,7.822889,8.05953,6.941485,7.610255,8.512236,9.345626,9.211872,6.636252,5.288424,4.7259717,4.5784993,4.6745276,5.055212,4.7774153,5.0243454,5.302142,5.456474,5.6485305,5.610805,5.442755,6.1801167,7.1952744,6.186976,5.7308407,5.4084597,5.4907694,5.9571934,6.495639,6.478491,6.416758,6.560801,6.7974424,6.660259,6.125243,5.9469047,5.9297566,5.895461,5.6656785,5.579939,4.9694724,4.537344,4.5167665,4.6676683,4.2698364,3.666229,2.884283,2.2292318,2.270387,2.3252604,2.3801336,2.719663,3.316411,3.8342788,3.858286,3.6799474,3.3609958,2.9974594,2.719663,3.0146074,3.2135234,2.9185789,2.2738166,1.9754424,1.9342873,1.6976458,1.5158776,1.4335675,1.2963841,1.2620882,1.1900668,1.2106444,1.2860953,1.2380811,1.2998136,1.2655178,1.155771,1.0906088,1.2826657,1.3101025,1.2483698,1.1797781,1.1351935,1.0666018,1.2072148,1.1934965,1.3615463,1.5330256,1.0357354,1.5158776,1.2655178,1.0117283,1.1111864,1.5638919,1.7113642,1.786815,1.8176813,1.8142518,1.7593783,1.7662375,1.9411465,2.0165975,1.9239986,1.8073926,1.9891608,1.8828435,1.704505,1.5330256,1.3203912,1.2826657,1.0734608,0.86082643,0.7579388,0.8196714,0.8128122,0.7956643,0.9602845,1.1900668,1.0528834,1.2620882,1.3066728,1.2415106,1.1214751,1.0014396,0.89855194,0.85396725,0.75450927,0.6276145,0.64133286,0.36353627,0.23664154,0.23664154,0.2777966,0.23664154,0.23664154,0.25378948,0.26064864,0.25378948,0.28465575,0.2469303,0.274367,0.37382504,0.45613512,0.32924038,0.22292319,0.17833854,0.19548649,0.25721905,0.32924038,0.40126175,0.48357183,0.5555932,0.6859175,1.039165,1.8005334,1.8519772,1.6667795,1.5570327,1.6496316,1.6496316,1.8485477,2.0337453,2.1469216,2.2909644,2.620205,2.983741,3.2786856,3.450165,3.4878905,3.7759757,4.2183924,4.506478,4.513337,4.280125,4.695105,5.096367,5.4804807,5.9469047,6.7048435,6.8866115,7.0135064,7.363324,7.8331776,7.9086285,8.275595,9.132992,9.949233,10.504827,10.871792,12.109874,12.377381,12.545431,12.775213,12.5145645,10.662587,8.680285,7.5862474,7.966932,9.959522,10.1652975,8.683716,8.337327,9.355915,9.373062,10.000677,11.808069,13.934414,15.110763,13.618892,13.282792,14.527733,14.88441,14.201921,14.644339,16.897577,14.935853,13.087306,12.946692,13.392539,13.306799,13.207341,12.946692,12.795791,13.457702,14.208781,14.267084,14.044161,14.027013,14.781522,16.901007,19.260563,20.35803,20.433481,21.503513,21.95279,22.302607,23.506393,24.76505,23.557837,23.708738,22.391777,20.824455,20.087093,21.10568,23.832203,26.400965,27.44013,27.313234,28.115759,27.357819,25.039417,23.976246,25.01884,27.01829,25.817934,23.44123,21.369759,20.128248,19.274282,17.336565,15.409137,14.826107,15.885849,17.864721,18.159666,18.567787,18.506054,18.231688,18.835295,19.552078,17.88873,16.11906,15.522313,16.393429,0.6790583,0.6962063,0.7476501,0.89169276,1.0597426,1.039165,1.2895249,1.4335675,1.5021594,1.529596,1.5604624,1.4095604,1.8005334,1.8656956,1.5433143,1.5604624,1.7936742,1.8313997,1.9137098,1.9925903,1.7422304,1.8313997,1.8862731,2.2566686,2.8534167,3.1380725,3.5393343,4.1017866,5.0003386,5.768566,5.312431,5.809721,7.2364297,9.493098,12.9638405,18.509483,19.384027,15.906426,10.443094,5.130663,1.8588364,0.9602845,0.5693115,0.4389872,0.37725464,0.24350071,0.18519773,0.216064,0.2503599,0.28465575,0.3806842,1.0528834,1.3821237,1.2998136,0.9294182,0.58988905,0.42869842,0.34981793,0.29837412,0.25378948,0.22292319,0.33609957,0.39097297,0.3806842,0.33609957,0.3018037,0.26407823,0.2503599,0.33266997,0.48357183,0.58302987,0.5624523,0.5624523,0.5212973,0.4629943,0.48357183,0.4389872,0.3806842,0.3841138,0.4664239,0.5624523,0.6001778,0.6893471,0.67219913,0.53844523,0.40126175,0.29837412,0.42526886,0.6207553,0.7407909,0.64133286,0.59331864,0.64133286,0.6276145,0.6036074,0.85739684,1.1008976,1.2792361,1.430138,1.6256244,1.961724,2.4315774,2.8225505,3.1380725,3.4776018,4.0263357,5.2026844,6.914048,7.8023114,7.5519514,6.8728933,5.9228973,5.576509,5.336438,4.9077396,4.2046742,3.7211025,3.117495,2.8294096,2.7985435,2.4658735,2.3389788,2.037175,2.1983654,2.9151495,3.7519686,4.3795834,3.2581081,2.7779658,3.4810312,4.033195,3.6010668,3.0729103,2.4041407,1.762808,1.5364552,0.78194594,0.71678376,0.9294182,1.0631721,0.82996017,0.91227025,1.0528834,0.864256,0.39783216,0.1371835,0.15776102,0.2194936,0.25378948,0.23321195,0.17833854,0.15090185,0.116605975,0.08573969,0.06516216,0.048014224,0.024007112,0.020577524,0.020577524,0.020577524,0.0274367,0.0274367,0.020577524,0.01371835,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15433143,0.3018037,0.33609957,0.32924038,0.53158605,0.61046654,0.5418748,1.1043272,1.8588364,1.1489118,1.0734608,1.1351935,1.1832076,1.1900668,1.2517995,0.8711152,1.0220171,1.2758065,1.3855534,1.2826657,1.2586586,1.4404267,1.9411465,2.3321195,1.6187652,2.0989075,2.503599,2.7642474,2.884283,2.9288676,2.7299516,3.6868064,5.2781353,6.914048,7.915488,11.159878,14.946142,18.46147,21.143406,22.69358,23.880217,24.127148,24.476965,25.498983,27.302946,28.835972,28.818823,27.820814,26.150604,23.85964,18.650097,14.887839,13.838386,16.156786,21.901346,28.366117,33.92891,38.349648,41.88555,45.273983,48.71729,50.082264,52.6476,54.94885,50.79219,53.415825,57.9566,53.419254,38.040985,19.294859,12.812939,9.095266,6.9826403,5.754848,5.1169443,4.9831905,5.5147767,5.7411294,5.2609873,4.2286816,5.1100855,7.3393173,11.89038,16.592344,16.13278,14.977009,15.488017,17.607502,20.642687,23.266321,30.362139,31.91917,24.878227,12.3911,3.8102717,10.422516,10.401938,14.205351,20.001354,13.687484,12.30536,8.327039,7.682276,10.30934,10.158438,12.871242,9.702303,7.3701835,7.257007,5.4187484,4.65395,4.822,5.31929,7.98408,17.106783,7.6445503,4.2423997,3.3438478,3.0283258,3.0146074,5.2438393,8.704293,15.350834,19.987637,10.271614,8.416207,9.918367,10.563129,9.355915,8.525954,11.698323,16.074476,14.664916,8.2653055,5.4496145,6.4887795,11.945253,16.62664,18.485476,18.62266,15.117621,15.580616,14.860402,11.163307,6.0703697,7.455923,10.22703,9.688584,7.6445503,12.404818,14.13333,13.111313,13.529722,15.988737,17.511473,14.249936,13.872682,14.928994,16.80155,19.69955,13.924125,12.782072,15.138199,18.28313,17.919594,18.108221,17.154797,13.937843,9.55826,7.363324,6.4064693,6.6431108,13.015285,19.178253,7.514226,8.920357,15.069608,16.88386,13.05301,10.045261,9.592556,7.3084507,4.7979927,3.1723683,3.0386145,4.0949273,4.681387,5.1580997,5.686256,6.210983,6.4407654,4.8734436,3.474172,3.2478194,4.2355404,4.314421,4.664239,6.228131,8.848335,11.249047,12.319078,12.991278,13.29994,12.936404,11.235329,10.251037,8.299602,7.222711,7.284444,7.1884155,5.576509,6.5162163,7.414768,7.39762,7.281014,7.2364297,9.705732,14.79524,20.62554,23.328054,21.04395,19.77843,22.168854,26.033998,24.408375,18.770132,14.407697,11.441104,10.364213,12.05157,9.403929,6.355026,6.5333643,8.045813,3.474172,3.192946,3.4810312,4.105216,5.0414934,6.4407654,5.7582774,5.579939,6.018926,6.742569,6.9552035,6.433906,5.0140567,4.6436615,5.518206,6.0840883,6.7185616,7.5245147,8.097256,8.076678,7.1884155,7.5245147,9.009526,9.956093,9.163857,5.909179,5.003768,4.496189,4.307562,4.331569,4.4516044,4.863155,5.2781353,5.5079174,5.576509,5.7102633,5.425607,5.535354,6.0223556,6.368744,5.5559316,5.2438393,5.1238036,5.4084597,6.0223556,6.6122446,6.7631464,6.550512,6.4098988,6.3824625,6.111525,5.669108,5.4941993,5.4187484,5.3878818,5.48734,5.3501563,4.8151407,4.5201964,4.554492,4.4584637,4.0503426,3.3644254,2.4830213,1.786815,1.9514352,2.2395205,2.609916,2.9871707,3.316411,3.5599117,3.5873485,3.2306714,2.8465576,2.5961976,2.4384367,2.9871707,3.1072063,2.6785078,1.9857311,1.704505,1.6804979,1.4644338,1.2483698,1.1523414,1.2415106,1.2072148,1.1626302,1.1763484,1.2209331,1.1660597,1.1934965,1.1523414,1.1146159,1.1283343,1.2312219,1.138623,1.1832076,1.2415106,1.2620882,1.2826657,1.2415106,1.2209331,1.371835,1.5741806,1.4198492,1.255229,0.9568549,0.89169276,1.1214751,1.4061309,1.611906,1.6153357,1.6496316,1.7490896,1.728512,1.9308578,1.903421,1.762808,1.6221949,1.5604624,1.7936742,1.6942163,1.6359133,1.6599203,1.4781522,1.4095604,1.1660597,0.97057325,0.89855194,0.88826317,0.90198153,0.85739684,0.9842916,1.1934965,1.0871792,1.1317638,1.1694894,1.1111864,0.9774324,0.88826317,0.84024894,0.8196714,0.7305021,0.59331864,0.53501564,0.28808534,0.18862732,0.20234565,0.25721905,0.23321195,0.26750782,0.30866286,0.29151493,0.2469303,0.29837412,0.2709374,0.25721905,0.36010668,0.5007198,0.41840968,0.28808534,0.18862732,0.15433143,0.19548649,0.274367,0.33609957,0.44584638,0.53501564,0.6173257,0.7990939,1.2963841,1.4438564,1.4129901,1.371835,1.4781522,1.5981878,1.7765263,1.937717,2.0817597,2.2841053,2.4624438,2.7230926,2.9871707,3.1963756,3.316411,3.5564823,3.882293,4.1600895,4.2869844,4.1772375,4.5167665,4.770556,5.0106273,5.442755,6.4133286,7.0032177,7.2467184,7.394191,7.534804,7.6033955,7.846896,8.549961,9.407358,10.124143,10.4533825,11.249047,11.465111,11.753197,12.195613,12.291641,10.336777,8.611694,7.740579,7.915488,8.89635,8.875772,8.368194,8.9100685,10.446524,11.334786,11.080997,10.847785,11.609154,12.908967,12.874671,13.457702,14.544881,15.165636,14.949572,14.147048,14.493437,13.54687,13.533153,14.38369,13.7526455,13.697772,13.323947,13.015285,13.173045,14.2190695,14.366542,14.79524,14.733508,14.020154,13.101024,14.342535,17.017612,18.725548,19.239986,20.519222,22.847912,24.322634,25.159454,25.166313,23.753323,23.952238,23.509823,22.727877,22.350622,23.561266,26.136887,27.073164,26.754211,26.133457,26.743923,26.253492,24.209457,23.78076,25.228045,25.917393,25.20061,24.284908,23.074265,21.644127,20.244854,17.62808,15.3302555,14.723219,15.837835,17.38115,18.04649,18.396307,18.197392,17.929884,18.79414,19.78186,18.547209,16.925014,15.985307,16.03675,0.67219913,0.6893471,0.7476501,0.90198153,1.0940384,1.155771,1.2106444,1.3238207,1.4541451,1.5604624,1.5844694,1.4850113,1.9480057,1.9823016,1.546744,1.546744,1.7147937,1.7971039,1.8588364,1.8897027,1.7971039,1.9720128,2.0303159,2.3286898,2.8088322,2.976882,3.4947495,4.3007026,5.56965,6.7871537,6.7459984,7.81603,9.506817,12.445972,16.266533,19.644676,14.973578,9.373062,5.453044,3.4707425,1.3032433,0.5761707,0.35324752,0.34981793,0.39783216,0.45270553,0.47671264,0.5144381,0.4938606,0.44584638,0.51100856,0.94999576,1.4095604,1.2689474,0.64476246,0.40126175,0.29837412,0.28465575,0.29151493,0.2777966,0.2469303,0.39440256,0.432128,0.39440256,0.35324752,0.4115505,0.44927597,0.45270553,0.50757897,0.59331864,0.6001778,0.58645946,0.58988905,0.5521636,0.48357183,0.4698535,0.4424168,0.4081209,0.38754338,0.38754338,0.4081209,0.45613512,0.5178677,0.53501564,0.50757897,0.5007198,0.4938606,0.607037,0.67219913,0.6379033,0.5693115,0.70306545,0.86082643,0.980862,1.0700313,1.1866373,1.2209331,1.2517995,1.3821237,1.6324836,1.9514352,2.2223728,2.428148,2.6785078,3.0523329,3.6147852,4.513337,6.0737996,6.90033,6.7700057,6.6225333,6.1801167,5.7136927,5.137522,4.3795834,3.3747141,3.1517909,2.8534167,2.5893385,2.2978237,1.7525192,1.9823016,2.1572106,2.4007113,2.74367,3.1346428,3.2375305,2.5790498,2.435007,3.000889,3.3884325,4.0194764,3.9337368,3.391862,2.6990852,2.201795,1.5776103,1.4575747,1.5913286,1.6324836,1.1214751,1.0906088,1.0871792,0.8265306,0.3841138,0.19891608,0.16462019,0.18519773,0.20577525,0.1920569,0.14747226,0.1097468,0.10288762,0.1097468,0.12003556,0.1097468,0.26064864,0.31895164,0.35324752,0.41498008,0.5144381,0.4081209,0.2503599,0.13375391,0.082310095,0.058302987,0.0274367,0.010288762,0.006859175,0.0034295875,0.0,0.2194936,0.2709374,0.25721905,0.1920569,0.0,0.09602845,0.29151493,0.37382504,0.31209245,0.26407823,0.33952916,0.48357183,1.1146159,1.7902447,1.2037852,1.0014396,0.9774324,1.1077567,1.2826657,1.2929544,1.0117283,1.1249046,1.1626302,1.1180456,1.4404267,1.6290541,1.6873571,2.170929,2.7162333,2.037175,2.411,3.0077481,3.018037,2.6236343,3.0043187,3.6319332,4.6402316,6.183546,7.864044,8.721441,12.548861,16.156786,18.95876,20.941061,22.655855,23.760181,24.751333,25.865948,27.230925,28.84969,29.662502,28.733084,26.723345,24.11343,21.191422,15.899568,13.262215,13.920695,17.71039,23.643576,31.305275,36.871494,40.47942,43.099625,46.54636,46.868744,48.11368,50.2366,51.06999,46.340588,55.182064,57.839993,49.327755,32.543354,18.272842,13.954991,10.477389,7.716572,5.7377,4.8185706,4.290414,4.372724,4.7362604,4.6745276,3.117495,3.806842,5.73427,9.89436,15.477728,19.881319,17.737827,17.182234,20.927343,27.035439,28.911423,32.121517,30.68109,22.652426,10.8958,3.0523329,14.321958,11.46854,13.557159,21.04395,15.80011,15.758954,8.292743,4.763697,7.140401,8.011517,13.920695,11.111863,6.8591747,4.5339146,3.6044965,4.2252517,4.6127954,4.5819287,5.8474464,11.993267,7.589677,4.616225,3.782835,4.7362604,6.077229,8.522525,13.186764,19.435472,23.170294,16.825556,12.075578,10.14129,9.5033865,9.136421,8.501947,11.907528,14.424845,13.042721,9.163857,8.594546,9.054111,12.5145645,17.04848,20.330595,19.634388,18.1288,16.462019,14.55174,11.965831,7.8949103,8.155559,11.458252,11.526843,9.743458,15.138199,13.989287,12.504276,13.416546,16.191082,17.017612,13.485138,13.22106,13.55373,14.068168,16.575195,13.265644,12.476839,14.928994,17.171944,11.578287,10.151579,8.831187,8.7283,8.796892,5.8200097,6.385892,7.486789,14.020154,19.8676,7.9086285,8.621983,14.225929,14.46257,10.666017,15.772673,15.501736,10.662587,7.4284863,6.5299344,3.2546785,5.130663,5.456474,6.0086374,7.085528,7.4799304,7.747438,5.658819,4.3178506,4.629943,5.2781353,5.219832,5.7582774,7.016936,8.8929205,11.06042,13.238208,14.160767,13.701202,12.253916,10.748327,9.438225,8.423067,8.2653055,8.666568,8.457363,7.4970784,8.241299,9.506817,10.038403,8.525954,8.1384115,9.918367,13.838386,17.78927,17.590355,18.506054,21.503513,27.481285,32.17982,26.19176,20.334024,15.515453,12.154458,10.635151,11.30735,9.534253,8.786603,10.360784,11.5645685,5.689686,3.6765177,2.9563043,3.508468,4.6573796,5.0826488,4.8117113,6.0086374,7.349606,8.165848,8.412778,6.684266,5.284994,4.8734436,5.504488,6.6465406,7.5416627,7.9600725,7.8674736,7.4627824,7.160979,7.56224,8.676856,9.31133,8.604835,6.018926,5.2301207,4.4996185,4.262977,4.3658648,4.057202,4.7945633,5.40503,5.5902276,5.5113473,5.7891436,5.456474,5.576509,5.65539,5.5662203,5.545643,5.360445,5.3844523,5.761707,6.358455,6.7459984,6.9826403,6.8214493,6.759717,6.725421,6.094377,5.2781353,5.0140567,4.9248877,4.9591837,5.363875,5.099797,4.6745276,4.461893,4.431027,4.1292233,3.649081,2.9288676,2.1743584,1.7147937,2.0028791,2.4007113,2.8259802,3.0420442,3.0351849,3.0351849,2.9563043,2.603057,2.3835633,2.3629858,2.2806756,2.784825,2.7230926,2.318401,1.821111,1.5398848,1.4027013,1.2723769,1.1523414,1.1043272,1.2723769,1.2003556,1.1249046,1.0871792,1.097468,1.1660597,1.138623,1.1077567,1.1592005,1.255229,1.2346514,1.255229,1.3341095,1.3238207,1.2620882,1.3615463,1.2312219,1.3169615,1.3889829,1.3752645,1.3752645,0.94999576,0.8196714,0.88826317,1.0460242,1.155771,1.430138,1.4987297,1.546744,1.6256244,1.6770682,1.7593783,1.6599203,1.6530612,1.7113642,1.5055889,1.4987297,1.4610043,1.5707511,1.7696671,1.7319417,1.5261664,1.2346514,1.0837497,1.0597426,0.91912943,0.9568549,0.94656616,0.9842916,1.0494537,0.9774324,0.9842916,1.0460242,1.0117283,0.8711152,0.764798,0.84024894,0.805953,0.6824879,0.5144381,0.36353627,0.20577525,0.14061308,0.18176813,0.26750782,0.28808534,0.30523327,0.36353627,0.33609957,0.2469303,0.29151493,0.29151493,0.26064864,0.3566771,0.5144381,0.4664239,0.32924038,0.20577525,0.14404267,0.15433143,0.2194936,0.2503599,0.37382504,0.4972902,0.58302987,0.6790583,0.84024894,1.0151579,1.1489118,1.2380811,1.3375391,1.5707511,1.7079345,1.8005334,1.9171394,2.1332035,2.2909644,2.5070283,2.7951138,3.1037767,3.3369887,3.3198407,3.4810312,3.6936657,3.8548563,3.8720043,4.139512,4.496189,4.791134,5.178677,6.0875177,7.0272245,7.431916,7.5416627,7.56567,7.6616983,7.7371492,8.419638,9.328478,10.024684,10.024684,9.877212,9.97667,10.491108,11.177026,11.375941,9.798331,8.796892,8.292743,8.179566,8.333898,8.152129,7.9943686,8.858624,10.55284,11.705182,11.46854,9.575408,8.707723,9.571979,10.916377,12.151029,13.090735,14.225929,14.932424,13.4645605,13.128461,13.231348,14.339106,15.580616,14.634049,14.514014,14.579176,14.479718,14.411126,15.103903,13.937843,14.30138,14.479718,13.725209,12.253916,12.823228,15.436573,17.593784,18.53692,19.288,21.314886,23.681301,24.703318,24.10314,22.988525,23.184011,23.012531,22.624989,22.583834,23.842491,25.787067,26.150604,25.416672,24.151155,23.009102,23.053686,22.340332,22.36434,23.043398,22.748453,23.132568,23.201159,22.755312,21.819035,20.649546,17.895588,15.820687,15.138199,15.820687,17.099922,18.214539,18.485476,18.427174,18.584934,19.53493,19.895037,19.298288,18.20768,17.2131,17.021042,0.66191036,0.72364295,0.8471081,0.99801,1.1660597,1.371835,1.430138,1.4335675,1.4335675,1.4644338,1.5193073,1.5261664,1.8691251,1.9480057,1.6976458,1.611906,1.5536032,1.7079345,1.7422304,1.6290541,1.6496316,2.0234566,2.153781,2.3801336,2.7162333,2.8705647,3.8205605,4.5510626,6.046363,7.846896,8.06296,9.201583,10.504827,13.409687,17.075916,18.37916,11.115293,5.7891436,3.1552205,2.369845,1.0185875,0.50757897,0.28465575,0.2777966,0.4389872,0.7373613,0.84024894,0.8779744,0.77851635,0.64819205,0.7510797,1.097468,1.3615463,1.1317638,0.5624523,0.3806842,0.26064864,0.25721905,0.30866286,0.34638834,0.30523327,0.3841138,0.4081209,0.39783216,0.41840968,0.5453044,0.6276145,0.6379033,0.59674823,0.5521636,0.5796003,0.72707254,0.7133542,0.61389613,0.4972902,0.42869842,0.4629943,0.44584638,0.38754338,0.33266997,0.34638834,0.39783216,0.5212973,0.6241849,0.70649505,0.84024894,1.0425946,1.1523414,1.0700313,0.90541106,0.9602845,1.1694894,1.371835,1.7696671,2.1743584,1.9823016,1.5741806,1.4095604,1.4987297,1.728512,1.8485477,1.8965619,2.1057668,2.3801336,2.6887965,3.0489032,3.6182148,4.839148,5.4941993,5.3707337,5.284994,5.453044,5.2301207,4.979761,4.5784993,3.40901,3.093488,2.7230926,2.3664153,1.9651536,1.3375391,1.1934965,1.8931323,2.2600982,2.054323,1.9857311,2.428148,2.9563043,3.542764,4.0434837,4.184097,4.712253,4.540774,4.0709205,3.549623,3.083199,2.7779658,2.3492675,2.2155135,2.136633,1.2175035,0.8848336,0.78537554,0.8676856,0.91227025,0.5144381,0.20234565,0.1371835,0.16119061,0.17490897,0.12346515,0.09602845,0.12003556,0.18862732,0.26407823,0.28808534,0.82996017,0.9842916,1.0460242,1.2072148,1.5364552,0.9534253,0.58988905,0.3841138,0.26750782,0.15776102,0.08573969,0.041155048,0.020577524,0.01371835,0.0,0.4424168,0.5418748,0.5144381,0.3806842,0.0,0.0,0.34295875,0.5041494,0.40126175,0.41498008,0.45270553,0.59331864,0.59674823,0.5727411,0.96371406,0.8196714,1.2723769,1.670209,1.762808,1.6976458,1.1180456,0.94656616,0.9568549,1.0734608,1.3649758,1.670209,1.5193073,1.8005334,2.6167753,3.2615378,2.4624438,2.8122618,2.9254382,2.668219,3.1723683,4.3007026,5.164959,6.392751,8.032094,9.537683,13.437123,17.144508,20.097382,22.103691,23.338343,24.380938,26.147175,27.975145,29.449867,30.396433,30.564484,29.34012,26.44212,22.076254,16.914726,13.821238,13.646329,16.228807,20.855322,26.243204,32.563934,36.689728,39.433395,41.834106,45.14709,42.928146,44.152508,45.164238,44.852146,44.64637,57.335842,56.087475,44.107925,28.246082,18.989626,15.758954,11.869802,8.22758,5.579939,4.513337,3.6044965,3.0900583,3.2272418,3.4433057,2.3424082,3.5804894,6.121814,9.73317,14.102464,18.821575,17.010754,18.313997,24.02083,32.00834,36.748028,37.114994,30.279827,19.648108,9.033533,2.644212,17.110212,13.704632,15.182784,22.415783,14.38369,16.595774,8.611694,2.8259802,3.3781435,6.1629686,10.323058,9.736599,6.6225333,3.5118976,3.2409601,4.5784993,4.633373,4.386442,4.863155,7.157549,8.937505,7.6514096,6.0875177,6.1629686,8.9100685,13.80066,19.54179,22.62156,22.624989,22.261452,16.37971,10.4705305,7.534804,7.7885933,8.659708,11.413667,13.461131,12.4802685,10.000677,11.38966,13.910407,13.516005,13.413116,14.651197,16.13278,23.019392,18.687822,13.557159,11.537132,9.997248,9.434795,11.358793,11.688034,11.290202,15.978448,14.620332,14.260224,14.023583,13.2690735,11.585147,11.441104,13.46799,13.289652,10.820349,10.254466,12.905538,16.194511,18.293419,16.770683,8.567109,8.110974,7.466212,9.582268,12.089295,7.3187394,9.126132,8.237869,8.663138,10.360784,9.266746,9.8429165,9.757176,7.1369715,6.807731,20.296299,20.498644,14.616901,11.55771,11.214751,4.479041,5.8680243,5.5113473,5.5079174,6.543653,7.8983397,7.953213,7.5279446,7.14726,6.831738,6.077229,6.2555676,7.040943,7.8606143,8.889491,11.032983,13.63604,13.077017,11.022695,9.187865,9.321619,7.9292064,8.162418,9.126132,10.021255,10.134431,11.331357,11.667457,12.130451,12.363663,10.666017,10.621432,10.477389,12.360233,14.894698,13.210771,14.490007,18.348293,23.725885,26.833092,21.139977,19.469769,17.027903,14.400838,12.325937,11.674315,10.401938,12.171606,13.999576,13.13189,7.0375133,3.9886103,2.620205,3.525616,5.2335505,4.214963,4.695105,6.7631464,8.961512,10.244178,9.997248,7.257007,6.2727156,6.0635104,6.2864337,7.2535777,8.309891,8.385342,7.623973,6.708273,6.8557453,7.373613,7.6274023,7.939495,7.905199,6.39961,5.353586,4.57507,4.4859004,4.7431192,4.249259,4.57164,5.219832,5.4153185,5.267846,5.761707,5.5079174,5.381023,5.164959,5.0655007,5.693115,5.720552,5.778855,6.159539,6.6876955,6.7459984,7.082098,6.842027,7.0478024,7.449064,6.550512,5.0620713,4.554492,4.4275975,4.513337,5.055212,4.846007,4.6093655,4.40702,4.201245,3.8685746,3.3266997,2.534465,1.961724,1.8416885,2.1812177,2.5310357,2.7779658,2.750529,2.5310357,2.4487255,2.2292318,2.0817597,2.1332035,2.287535,2.218943,2.4418662,2.2120838,1.9548649,1.786815,1.5364552,1.2380811,1.1900668,1.2312219,1.2929544,1.4129901,1.2415106,1.08032,0.9534253,0.9328478,1.1523414,1.1489118,1.1111864,1.2243627,1.4095604,1.313532,1.4918705,1.5055889,1.3615463,1.1797781,1.1934965,1.2243627,1.4061309,1.2826657,0.9534253,1.0734608,0.91227025,0.91569984,0.89855194,0.8711152,1.0254467,1.3341095,1.5536032,1.5981878,1.5604624,1.7079345,1.4541451,1.4267083,1.7113642,1.99602,1.587899,1.3101025,1.3203912,1.4850113,1.6804979,1.8073926,1.5776103,1.3101025,1.2003556,1.1660597,0.8711152,0.9328478,0.96714365,0.9602845,0.90884066,0.83338976,0.84024894,0.91227025,0.91227025,0.8196714,0.71678376,0.83338976,0.75450927,0.58302987,0.3806842,0.18862732,0.15776102,0.13032432,0.18519773,0.30523327,0.37382504,0.31552204,0.4115505,0.4115505,0.30866286,0.33952916,0.34981793,0.31552204,0.3841138,0.5178677,0.48700142,0.36010668,0.2469303,0.17147937,0.14747226,0.17490897,0.16119061,0.26064864,0.38754338,0.50757897,0.64133286,0.71678376,0.7990939,0.94656616,1.1317638,1.2380811,1.4918705,1.5707511,1.646202,1.7730967,1.8691251,2.1057668,2.3561265,2.6819375,3.0523329,3.3369887,2.9974594,2.9871707,3.117495,3.2615378,3.3644254,3.6387923,4.1360826,4.633373,5.130663,5.8337283,6.7802944,7.3187394,7.6376915,7.864044,8.049242,8.018375,8.539673,9.321619,9.832627,9.273604,8.385342,8.491658,9.325048,10.281903,10.429376,9.379922,8.97866,8.7283,8.48137,8.436785,8.014946,7.48336,7.922347,9.167287,9.80862,10.117283,8.608265,7.4799304,7.8023114,9.4862385,10.6488695,11.314209,12.4802685,13.653188,12.826657,13.543441,14.291091,15.258235,15.96816,15.271953,15.594335,15.909856,15.693792,15.179354,15.364552,13.4645605,13.152468,13.197053,13.05301,12.843805,12.919256,14.733508,16.578627,17.669235,18.142517,18.259123,20.224277,21.589252,21.482935,20.649546,21.050808,20.735287,20.306587,20.340883,21.397196,23.19773,24.27805,24.02426,22.306036,19.469769,20.296299,20.539799,20.412905,20.272291,20.61868,21.723007,21.462358,20.7833,20.248285,20.028791,18.296848,16.88729,16.167076,16.37285,17.593784,18.969048,19.486916,19.836735,20.412905,21.342323,20.759293,20.334024,19.459478,18.44432,18.516342,0.6241849,0.7339317,0.9362774,1.0768905,1.1763484,1.4198492,1.6256244,1.605047,1.5364552,1.4815818,1.371835,1.5913286,1.9411465,1.9342873,1.7079345,2.0131679,1.6839274,1.8485477,1.8931323,1.7079345,1.7079345,1.9274281,2.020027,2.3389788,2.7985435,2.884283,4.4584637,4.9351764,5.813151,7.1849856,7.720001,7.8537555,8.721441,9.966381,11.31078,12.542002,7.0375133,3.4638834,1.8759843,1.6187652,1.313532,0.90884066,0.50757897,0.25721905,0.23664154,0.45613512,0.5796003,0.7373613,0.86082643,0.9568549,1.1283343,1.4472859,1.3512574,1.0288762,0.65162164,0.3806842,0.22292319,0.274367,0.40126175,0.45270553,0.24350071,0.25721905,0.34295875,0.42183927,0.4355576,0.34981793,0.32581082,0.36696586,0.42869842,0.5418748,0.823101,1.1283343,0.9842916,0.6756287,0.45613512,0.5658819,0.6379033,0.5178677,0.45270553,0.50757897,0.5796003,0.7888051,0.94999576,1.1249046,1.3409687,1.5707511,2.0097382,2.0749004,1.8142518,1.5090185,1.6942163,2.095478,2.287535,3.3369887,4.5819287,3.6319332,2.411,1.7936742,1.5433143,1.4575747,1.371835,1.5193073,1.8691251,2.1915064,2.452155,2.7916842,3.2443898,3.6696587,4.197815,4.650521,4.5167665,4.431027,5.381023,5.521636,4.4584637,3.2512488,2.8945718,2.452155,1.9857311,1.5673214,1.2517995,1.0185875,0.7613684,0.9294182,1.7559488,3.2203827,4.1600895,5.528495,6.7322803,7.1026754,5.90575,5.967482,4.8288593,3.6387923,3.0077481,3.0214665,3.2649672,2.510458,2.1091962,2.0714707,1.0837497,0.5453044,0.5041494,1.3409687,2.2498093,1.2346514,0.30866286,0.06859175,0.06859175,0.07545093,0.07545093,0.07545093,0.16804978,0.30866286,0.44584638,0.5178677,1.7147937,1.9239986,1.879414,2.0886188,2.8088322,0.96371406,0.65162164,0.72364295,0.61046654,0.30523327,0.18176813,0.09602845,0.041155048,0.01371835,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.548734,0.7339317,0.47671264,0.548734,0.24350071,0.45956472,0.4355576,0.18176813,0.48700142,0.9877212,1.5707511,1.9514352,2.1126258,2.318401,1.0871792,0.6036074,0.48700142,0.6310441,1.2037852,1.961724,2.4624438,3.292404,4.8014226,7.0958166,3.8377085,3.1689389,3.9200184,4.602506,3.4192986,4.945465,5.353586,6.3481665,8.303031,10.268185,13.114742,16.506605,20.975357,25.19375,25.999702,27.062874,28.482723,30.447878,32.457615,33.325302,32.99606,31.521338,27.491573,21.297739,15.121051,14.057879,16.520323,20.893047,26.328943,32.776566,35.132694,35.115547,36.528538,39.81408,42.08447,39.48484,40.517147,38.565712,35.39677,41.168766,51.728466,47.05394,35.18071,23.578413,19.133669,15.055889,10.88894,7.373613,4.804852,3.0351849,2.5481834,2.2326615,2.3321195,2.5619018,2.136633,4.5167665,9.705732,11.118723,9.568549,13.289652,11.032983,11.924676,17.820137,27.289227,35.612835,47.599243,38.082138,22.354052,9.80862,3.9371665,16.80155,20.320305,22.559826,22.673002,10.878652,14.579176,9.030104,4.166949,3.9680326,6.468202,6.7494283,5.2472687,4.5270553,4.9008803,4.4241676,4.523626,4.6573796,4.6573796,5.2644167,8.131552,9.657719,12.850664,10.611144,5.1409516,7.936065,17.394867,24.11686,24.147726,19.565796,18.478617,17.96418,11.684605,7.1129646,6.81802,8.453933,13.1421795,10.878652,7.857185,7.191845,8.9100685,13.011855,13.313659,10.597425,8.697433,14.496866,27.460707,21.290878,14.099034,12.72034,12.696333,11.89038,9.921797,10.103564,12.133881,12.085866,10.851214,13.152468,16.026463,17.333136,15.745236,10.731179,13.71492,13.831526,9.2153015,7.0203657,12.706621,25.571005,24.77191,11.30049,7.98065,7.8949103,7.4970784,8.498518,11.691463,16.952452,19.881319,11.238758,7.3701835,10.621432,9.352485,8.608265,7.0306544,5.9640527,9.249598,23.238884,19.600092,14.781522,14.13676,14.891269,6.1629686,8.323608,7.1712675,5.3398676,5.0655007,8.179566,8.213862,9.167287,9.815479,9.3593445,7.431916,6.2830043,6.245279,7.3187394,9.297611,11.763485,14.634049,13.327377,10.964391,10.031544,12.373952,9.993818,9.592556,9.506817,9.709162,11.794352,14.699212,15.875561,15.405707,13.656617,11.276484,11.348505,9.56512,7.4044795,6.3138704,7.706283,6.924337,10.501397,11.465111,10.497967,15.916716,18.45461,20.680412,19.668684,15.87213,13.138749,9.561689,10.569988,11.780633,10.686595,6.684266,5.4016004,3.7725463,3.9303071,5.56965,5.936616,6.5813785,6.451054,7.39762,9.009526,8.604835,7.4936485,6.9346256,6.910619,7.0478024,6.608815,7.9875093,8.045813,7.682276,7.346176,7.06495,6.368744,6.9654922,7.1095347,6.2418494,4.9591837,4.166949,4.461893,4.5784993,4.249259,4.2115335,3.8685746,4.4241676,5.096367,5.4941993,5.6142344,5.470192,5.1855364,4.8014226,4.6436615,5.3398676,5.0243454,5.2918534,6.385892,7.431916,6.4544835,7.1026754,6.018926,5.645101,6.40304,6.684266,4.914599,4.297273,4.139512,4.105216,4.2252517,4.482471,4.629943,4.496189,4.125794,3.782835,3.4535947,2.5927682,2.0680413,2.061182,2.061182,2.095478,2.2052248,2.194936,2.0337453,1.862266,1.99602,2.0749004,2.16064,2.218943,2.1194851,2.2052248,1.7971039,1.5055889,1.5364552,1.6942163,1.3752645,1.214074,1.1729189,1.2655178,1.5707511,1.4507155,1.1523414,0.8779744,0.7613684,0.8848336,1.2037852,1.1729189,1.3066728,1.6530612,1.8005334,1.3238207,1.2037852,1.2723769,1.255229,0.77851635,1.2792361,1.138623,0.881404,0.9294182,1.587899,1.1729189,0.91227025,0.78537554,0.82996017,1.1592005,1.5741806,1.7696671,1.8245405,1.8554068,2.0131679,1.7696671,1.5981878,1.4953002,1.4027013,1.2209331,1.3443983,1.4541451,1.5227368,1.5501735,1.587899,1.7079345,1.5364552,1.3924125,1.2895249,0.94656616,0.9945804,1.0082988,1.0425946,1.0768905,0.9911508,0.881404,0.7613684,0.72021335,0.7888051,0.9602845,0.8505377,0.8505377,0.66876954,0.32238123,0.15090185,0.18862732,0.17833854,0.20920484,0.31552204,0.47328308,0.36353627,0.490431,0.5693115,0.5453044,0.59674823,0.51100856,0.4424168,0.4664239,0.5624523,0.61046654,0.548734,0.38754338,0.23664154,0.15090185,0.1371835,0.12346515,0.18519773,0.23664154,0.32238123,0.64133286,0.77508676,0.72707254,0.805953,1.0563129,1.2517995,1.4953002,1.5090185,1.7250825,2.0749004,2.0131679,2.2326615,2.3149714,2.5070283,2.8122618,3.0214665,2.6304936,2.651071,2.867135,3.0351849,2.8980014,3.3026927,3.642222,4.2526884,5.127233,5.919468,6.2487082,6.9654922,7.73372,8.354475,8.759167,8.601405,8.378482,8.786603,9.469091,9.016385,8.820899,8.947794,9.839486,10.834066,10.161868,9.355915,9.191295,9.136421,8.851766,8.179566,7.4456344,6.924337,6.5779486,6.8900414,8.879202,8.868914,9.122703,9.321619,9.595985,10.511685,11.135871,12.144169,12.199042,11.705182,12.80265,14.04759,15.3302555,16.506605,17.075916,16.173935,17.151367,15.426285,13.756075,13.365103,13.96185,13.107883,12.161317,11.777204,12.442543,14.479718,12.905538,13.173045,13.848674,14.846684,17.412016,16.811838,15.920145,15.361122,14.949572,13.704632,14.778092,15.46744,15.498305,15.340545,16.221949,18.687822,19.77843,20.443771,20.899906,20.62897,21.44864,19.884748,18.927893,19.713268,21.544668,21.558388,20.893047,19.696121,18.564358,18.54035,17.929884,17.254255,17.62122,18.910746,19.792149,22.172283,22.583834,21.980227,21.70929,23.5304,22.70044,22.089973,20.745575,18.95533,18.235117,0.61389613,0.7442205,0.91227025,1.0871792,1.2449403,1.3821237,1.2758065,1.3238207,1.4678634,1.5673214,1.3992717,1.821111,1.9445761,1.7319417,1.4678634,1.7319417,1.7147937,1.8039631,1.8348293,1.8588364,2.16064,2.0474637,1.9823016,2.2326615,2.726522,3.0660512,4.396731,4.73969,5.003768,5.3741636,5.3158607,5.305572,5.6142344,6.4887795,7.939495,9.760606,7.2535777,4.4413157,2.6647894,2.1400626,1.9720128,2.0165975,1.6976458,1.2826657,0.922559,0.66533995,0.4355576,0.3806842,0.48357183,0.70306545,0.97057325,1.3272504,1.1249046,0.7339317,0.38754338,0.19891608,0.22635277,0.3806842,0.4972902,0.51100856,0.48700142,0.89169276,0.8471081,0.61046654,0.39097297,0.36353627,0.4081209,0.42869842,0.4698535,0.53501564,0.59331864,0.77165717,0.77851635,0.6756287,0.5555932,0.52815646,0.47328308,0.44927597,0.4389872,0.50757897,0.7888051,1.7971039,2.3904223,3.100347,3.625074,2.8396983,2.2635276,1.8554068,1.5090185,1.214074,1.0357354,1.3684053,1.7216529,2.177788,2.5001693,2.1057668,1.3924125,1.0494537,0.9602845,1.0014396,1.0425946,1.3375391,1.6907866,2.2498093,2.9391565,3.4776018,3.7622573,4.1360826,4.434457,4.513337,4.2595477,5.1409516,6.324159,6.444195,5.271276,3.7005248,2.9391565,2.5584722,2.1880767,1.7319417,1.3855534,1.0357354,0.939707,1.2003556,2.0508933,3.8171308,6.3207297,8.021805,8.1212635,7.1026754,6.7357097,5.381023,4.3624353,3.5530527,2.9563043,2.702515,3.2409601,2.8396983,2.2909644,1.8245405,1.1214751,0.64133286,0.52472687,0.9842916,1.5570327,1.1008976,0.26064864,0.05144381,0.044584636,0.041155048,0.041155048,0.048014224,0.08573969,0.13375391,0.21263443,0.37382504,0.97400284,1.5090185,1.4198492,0.90884066,0.91569984,0.4389872,0.3806842,0.42869842,0.4115505,0.28122616,0.14061308,0.06516216,0.0274367,0.01371835,0.0,0.0034295875,0.0,0.0,0.030866288,0.15776102,0.70649505,0.5041494,0.29151493,0.30523327,0.28122616,0.5041494,0.72021335,0.6036074,0.4698535,1.2929544,1.7353712,1.9068506,1.9514352,1.7936742,1.1729189,0.72021335,1.2380811,2.020027,2.5996273,2.74367,2.9048605,3.8205605,4.280125,3.8960114,3.1037767,2.5996273,2.7128036,3.5290456,4.6436615,5.188966,5.6005163,7.716572,8.680285,8.718011,11.122152,13.214201,16.510035,20.797018,25.18003,28.074602,29.988314,33.126385,34.902912,34.868614,34.728004,33.705986,30.053474,25.52985,20.824455,15.536031,17.158226,21.736725,27.086882,31.555634,34.00779,34.343887,36.905792,40.249638,42.146202,39.580868,39.687187,38.84694,35.38991,34.35761,47.503216,55.075745,47.931915,37.24189,28.92514,23.664154,18.667244,13.594885,9.441654,6.557371,4.6608095,4.297273,4.125794,3.858286,3.625074,3.9783216,5.65539,8.841476,8.992378,6.944915,8.920357,8.076678,8.327039,12.339656,19.37374,25.286348,41.268227,35.99352,21.880768,9.9869585,10.0041065,15.769243,13.999576,14.441993,18.248835,17.971039,23.01596,13.814379,5.4633327,3.9268777,6.018926,6.3481665,5.7274113,4.729401,3.9097297,3.8137012,4.3521466,5.518206,6.4819202,6.9346256,7.1061053,11.924676,18.296848,17.29884,9.97324,7.349606,11.585147,20.574095,24.85079,21.829325,15.830976,16.695232,13.766364,10.110424,8.450503,11.201033,13.485138,14.013294,11.777204,8.460793,8.436785,7.9943686,9.352485,9.530824,10.422516,18.766703,20.766151,17.947031,16.973028,17.319416,11.279913,9.644,8.110974,7.14726,7.9463544,12.425395,17.600643,19.202261,19.771572,19.322296,15.343974,11.965831,11.71547,11.046701,8.824328,6.334448,14.476289,15.247946,12.363663,8.968371,7.6376915,6.8111606,6.492209,7.8846216,10.744898,13.38911,16.228807,14.009865,13.234778,14.891269,14.4317045,14.30138,13.821238,11.880091,11.101575,17.857862,14.363112,16.921585,20.093952,18.800999,8.323608,12.020704,10.984968,8.601405,7.267296,8.399059,10.340206,10.38479,9.8429165,9.712592,10.652299,9.956093,8.539673,8.237869,9.424506,11.019264,10.069269,10.065839,10.491108,10.618003,9.506817,8.824328,9.383351,10.659158,12.46998,14.956431,15.645778,15.29939,14.79867,14.448852,13.972139,12.795791,10.882081,7.997798,5.8371577,7.997798,7.6651278,9.362774,11.441104,12.919256,13.485138,10.518545,9.777754,9.108984,7.936065,7.291303,9.788043,11.900668,10.871792,7.610255,6.684266,6.81802,5.360445,4.5784993,5.1992545,6.375603,7.764586,8.213862,8.755736,9.139851,7.8503256,7.14726,7.233,7.425057,7.438775,7.3530354,6.279575,6.6293926,6.711703,6.4064693,7.15069,7.099246,6.8728933,6.4887795,5.8645945,4.835718,4.4241676,4.9831905,4.722542,3.9303071,4.9694724,4.7534084,4.931747,5.1855364,5.336438,5.3227196,5.3913116,5.144381,4.979761,4.955754,4.791134,5.23698,6.142391,6.6636887,6.6739774,6.773435,6.989499,6.258997,5.9469047,6.1972647,5.950334,4.7191124,4.2869844,4.1326528,4.0949273,4.372724,4.5819287,4.3349986,3.7862647,3.357566,3.7485392,3.758828,2.8396983,2.2120838,2.201795,2.2292318,2.0714707,2.1846473,2.1469216,1.9411465,1.9480057,2.0131679,2.2566686,2.352697,2.2086544,1.9754424,1.9137098,1.7525192,1.5433143,1.3581166,1.2895249,1.4129901,1.2723769,1.097468,1.0288762,1.1214751,1.1832076,1.1832076,1.0700313,0.90884066,0.8848336,1.0837497,1.2449403,1.214074,1.0940384,1.2517995,1.255229,1.0563129,0.9328478,1.0151579,1.2895249,1.2723769,1.0117283,0.8196714,0.8676856,1.196926,0.89855194,0.78537554,0.89512235,1.2072148,1.6359133,1.4541451,1.488441,1.6599203,1.8485477,1.879414,1.5090185,1.3066728,1.1934965,1.155771,1.2449403,1.5536032,1.5433143,1.5673214,1.6393428,1.4404267,1.3855534,1.2072148,1.0185875,0.8711152,0.7613684,0.881404,0.91569984,0.89512235,0.84367853,0.8093826,0.7579388,0.65162164,0.6310441,0.67219913,0.6207553,0.75450927,0.96714365,0.82996017,0.3841138,0.16462019,0.2709374,0.29837412,0.32924038,0.38754338,0.44927597,0.4938606,0.58302987,0.64476246,0.67219913,0.6927767,0.6173257,0.6036074,0.6241849,0.6379033,0.59674823,0.7407909,0.50757897,0.2469303,0.12346515,0.11317638,0.12003556,0.15776102,0.17147937,0.21263443,0.42183927,0.5555932,0.52815646,0.6036074,0.8471081,1.1420527,1.4815818,1.5433143,1.6907866,1.9480057,2.0131679,1.9685832,2.1023371,2.3424082,2.5961976,2.7642474,2.510458,2.5310357,2.6750782,2.7711067,2.6064866,3.1072063,3.8514268,4.633373,5.3158607,5.8474464,5.8645945,6.3824625,7.051232,7.6514096,8.110974,8.683716,8.735159,8.855195,9.187865,9.421077,10.319629,11.084427,11.382801,11.187314,10.762046,9.6817255,8.7317295,8.460793,8.834618,9.2153015,7.857185,6.835168,6.293293,6.4304767,7.500508,7.9189177,8.39563,9.033533,9.537683,9.23245,10.401938,11.499407,12.902108,14.55174,15.964729,15.920145,16.307688,15.889278,15.12448,16.173935,16.242527,14.291091,12.788932,12.607163,13.008426,13.101024,12.840376,13.176475,13.972139,13.978998,14.291091,14.424845,13.87954,13.265644,14.335675,14.400838,14.5243025,14.123041,13.179905,12.236768,14.356253,15.525743,16.177364,16.684942,17.367432,18.12537,19.12681,19.819586,20.220848,20.910194,22.127699,21.311457,20.831314,21.19485,21.033659,22.755312,23.657295,22.882208,21.013083,20.090523,18.667244,17.638369,17.53891,18.804428,21.743584,24.418663,25.27606,24.3535,22.594122,21.843042,22.46037,23.266321,23.249174,22.19286,20.663265,0.6379033,0.7956643,1.0014396,1.1832076,1.3306799,1.4815818,1.2998136,1.2449403,1.3272504,1.4198492,1.2312219,1.4781522,1.4850113,1.3306799,1.2209331,1.5090185,1.6564908,1.8759843,1.9137098,1.8691251,2.1812177,2.2806756,2.0474637,2.1160555,2.651071,3.333559,4.2081037,4.3933015,4.5510626,4.8940215,5.1992545,5.429037,5.7377,6.385892,7.548522,9.301042,8.790032,6.914048,4.887162,3.5976372,3.6387923,3.5187566,2.843128,2.037175,1.3443983,0.8265306,0.4355576,0.31209245,0.41840968,0.64476246,0.78537554,1.0837497,1.2243627,0.8745448,0.2709374,0.216064,0.31209245,0.4081209,0.5212973,0.64133286,0.72364295,0.939707,0.8128122,0.5727411,0.39440256,0.4115505,0.42869842,0.42869842,0.48357183,0.5727411,0.58988905,0.58302987,0.53844523,0.5041494,0.48700142,0.4629943,0.58988905,0.66876954,0.70649505,0.7956643,1.1043272,1.8005334,2.0303159,2.3629858,2.6990852,2.270387,1.7833855,1.4095604,1.1763484,1.0528834,0.91569984,1.3855534,1.8313997,2.1332035,2.1983654,1.9720128,1.4164196,1.2243627,1.2483698,1.3169615,1.2449403,1.4953002,1.920569,2.5447538,3.1895163,3.4535947,3.9543142,4.437886,4.664239,4.633373,4.5819287,5.336438,6.0978065,5.8645945,4.5510626,2.9734523,2.5173173,2.3424082,2.0646117,1.6187652,1.2723769,1.2449403,1.4061309,1.7113642,2.417859,4.0846386,7.191845,8.419638,7.8983397,6.375603,5.212973,4.1463714,3.3987212,2.6716487,2.061182,2.0646117,3.2683969,3.8274195,3.4707425,2.4624438,1.6153357,0.939707,0.61389613,0.66876954,0.8505377,0.6207553,0.22635277,0.09945804,0.06516216,0.037725464,0.030866288,0.034295876,0.072021335,0.14747226,0.23321195,0.26407823,0.50757897,0.7888051,0.70649505,0.34638834,0.28808534,0.19548649,0.23664154,0.32924038,0.4081209,0.44927597,0.28122616,0.14747226,0.06516216,0.0274367,0.010288762,0.0034295875,0.006859175,0.006859175,0.017147938,0.07888051,0.5007198,0.28808534,0.17833854,0.36010668,0.48014224,0.8196714,1.0700313,1.1763484,1.1900668,1.2929544,1.3992717,1.4987297,1.6599203,1.7696671,1.5158776,1.5021594,2.2258022,2.8877127,3.1826572,3.3198407,3.882293,4.0606318,3.865145,3.4844608,3.2683969,3.6559403,4.190956,4.7842746,5.754848,7.8091707,9.379922,10.47396,11.358793,12.404818,14.085316,16.311117,18.560926,21.93221,26.178041,29.710516,31.881445,34.933777,36.453087,35.767166,33.963203,32.495342,30.327843,26.68219,22.182571,18.845583,21.959648,25.145735,28.839401,32.58451,35.012657,36.665718,40.5583,44.09078,45.380302,43.277966,42.015877,37.43052,34.84461,39.601448,57.051186,57.819416,49.334614,42.430855,39.48141,34.41591,27.309805,21.246294,16.45173,12.55229,8.580828,6.975781,6.3173003,5.5833683,5.5593615,8.824328,7.3530354,9.331907,9.071259,6.677407,8.038953,7.9086285,7.829748,13.022143,22.36434,28.400414,31.075493,24.593573,14.267084,7.5039372,13.790371,14.874121,14.832966,15.391989,16.619781,16.942162,20.093952,16.026463,9.935514,5.892031,6.848886,7.3427467,6.5162163,5.3844523,4.506478,3.9646032,4.3692946,5.0655007,11.046701,16.811838,6.375603,10.240748,16.846134,17.274832,11.348505,7.630832,10.233889,17.192522,21.942501,21.973368,18.849012,19.915615,18.663815,15.590904,12.648318,13.224489,13.9481325,14.099034,12.569438,10.295622,10.247607,10.299051,11.962401,13.13532,14.846684,21.28402,19.065077,17.367432,16.012743,13.903547,9.002667,8.464222,9.678296,8.447074,6.252138,10.268185,19.342873,18.6158,15.782962,14.472859,14.246507,10.333347,9.866923,9.935514,9.177576,7.747438,11.907528,10.556271,8.934075,8.56368,7.2432885,6.7494283,7.5039372,8.995808,11.046701,13.807519,15.563468,14.277372,12.926115,12.600305,12.4974165,15.436573,15.285671,12.912396,11.629731,17.195951,13.375391,15.71437,17.065628,14.661487,10.082987,14.96672,14.596324,11.444533,8.429926,8.9100685,11.578287,12.63803,11.893809,10.360784,10.268185,11.022695,10.374502,9.438225,8.772884,8.381912,8.923786,10.374502,11.067279,10.676306,10.233889,10.4705305,10.659158,11.790922,13.786942,15.481158,17.278261,16.952452,16.945591,17.408587,16.187653,13.231348,10.840926,8.683716,7.2604365,7.915488,7.1095347,8.361334,10.871792,13.365103,14.085316,11.821788,10.076128,9.331907,8.865483,6.7357097,9.088407,10.669447,10.484249,9.002667,8.155559,8.045813,7.500508,6.9037595,6.790583,7.840037,8.375052,9.1981535,9.657719,9.253027,7.658269,7.208993,7.2158523,7.1232533,6.9380555,7.2158523,6.3310184,6.6396813,6.776865,6.550512,6.941485,7.205563,7.1095347,6.783724,6.1046658,4.722542,4.787704,5.271276,4.931747,4.2252517,5.312431,5.305572,5.425607,5.5079174,5.5250654,5.579939,5.627953,5.254128,5.1238036,5.2026844,4.7362604,4.822,5.6176643,5.970912,5.9126086,6.660259,6.9380555,6.217842,5.7651367,5.8165803,5.5833683,4.839148,4.8597255,4.8254294,4.5510626,4.5099077,4.331569,3.9611735,3.3952916,2.9185789,3.0900583,3.3609958,2.9460156,2.4624438,2.2463799,2.3561265,2.061182,1.9857311,1.9308578,1.8725548,1.9857311,2.0440342,2.1880767,2.1640697,1.9514352,1.7559488,1.5844694,1.4335675,1.3409687,1.2929544,1.2449403,1.2072148,1.0871792,0.96714365,0.9328478,1.08032,1.138623,1.0460242,0.9911508,1.0151579,1.0117283,1.214074,1.2072148,0.9877212,0.7476501,0.8848336,0.9328478,0.77165717,0.7305021,0.9294182,1.255229,1.0940384,0.9945804,0.90198153,0.84367853,0.9431366,0.83681935,0.88826317,1.0494537,1.2655178,1.4541451,1.2037852,1.2380811,1.4953002,1.7490896,1.5810398,1.2723769,1.2277923,1.2003556,1.1797781,1.3992717,1.5981878,1.4095604,1.3238207,1.3924125,1.2312219,1.1832076,1.0494537,0.89512235,0.78537554,0.78194594,0.7922347,0.8128122,0.7956643,0.7407909,0.71678376,0.65162164,0.59331864,0.6241849,0.70649505,0.66191036,0.82996017,1.0082988,0.8848336,0.5212973,0.34295875,0.48014224,0.6036074,0.64476246,0.6036074,0.5521636,0.5796003,0.61389613,0.66191036,0.72707254,0.7990939,0.7922347,0.7922347,0.7510797,0.67219913,0.6036074,0.6962063,0.4938606,0.2503599,0.116605975,0.12346515,0.09945804,0.116605975,0.13375391,0.17490897,0.32924038,0.3841138,0.44584638,0.5796003,0.78194594,1.0048691,1.4129901,1.5536032,1.7319417,1.9925903,2.095478,2.0097382,2.061182,2.2120838,2.393852,2.5070283,2.4487255,2.6579304,2.7916842,2.750529,2.6613598,3.069481,3.7691166,4.588788,5.302142,5.6176643,5.658819,6.018926,6.4819202,6.9380555,7.3564653,7.846896,8.344186,8.855195,9.407358,10.014396,11.187314,12.404818,13.004995,12.867812,12.394529,11.324498,10.010965,9.23245,9.153569,9.338767,8.594546,8.110974,7.6514096,7.3290286,7.623973,8.141841,8.639131,9.328478,9.757176,8.81061,10.034973,10.676306,11.736049,13.512574,15.611482,15.477728,14.774663,13.9309845,13.646329,14.88441,14.167625,12.576297,11.63659,11.605724,11.454823,11.893809,12.075578,12.373952,12.788932,12.950122,13.72178,14.472859,14.232788,13.258785,13.025573,12.9707,13.296511,13.395968,13.210771,13.207341,15.206791,17.151367,18.612371,19.346302,19.28457,19.174824,19.29143,19.198832,19.017063,19.425184,19.819586,19.270851,19.459478,20.416334,20.512363,23.012531,23.928232,23.1943,21.654415,21.064526,20.148827,19.486916,19.257133,20.087093,23.063976,24.94682,25.910534,25.869379,24.888515,23.180582,23.643576,25.351511,27.056015,27.615038,25.985985,0.66876954,0.7990939,1.0117283,1.1420527,1.1900668,1.2998136,1.1763484,1.0768905,1.0700313,1.0906088,0.94999576,1.0185875,1.0185875,1.0048691,1.0631721,1.3169615,1.5981878,1.9342873,2.0680413,2.0577524,2.2738166,2.428148,2.2566686,2.2566686,2.6887965,3.5633414,3.9886103,4.280125,4.6402316,5.206114,6.0532217,6.3721733,6.574519,6.9552035,7.7611566,9.2153015,10.131001,9.280463,7.3873315,5.597087,5.48734,4.695105,3.415869,2.2120838,1.3478279,0.7956643,0.42526886,0.29837412,0.34295875,0.44927597,0.45956472,0.65505123,0.9602845,0.77165717,0.24350071,0.29494452,0.47328308,0.4664239,0.5144381,0.6756287,0.83338976,0.8128122,0.6173257,0.42526886,0.33952916,0.3806842,0.36010668,0.35324752,0.38754338,0.45956472,0.53501564,0.51100856,0.44584638,0.45956472,0.5590228,0.6276145,0.881404,0.90884066,0.86082643,0.8676856,1.0254467,1.2243627,1.155771,1.1523414,1.2792361,1.3443983,1.2758065,1.1283343,1.0460242,1.08032,1.1763484,1.5227368,1.9171394,2.1263442,2.1023371,1.978872,1.5707511,1.5055889,1.5638919,1.5913286,1.4575747,1.6736387,2.2635276,2.8980014,3.3609958,3.5461934,4.2526884,4.616225,4.7774153,4.852866,4.945465,5.020916,4.979761,4.341858,3.1689389,2.0886188,2.1057668,2.2909644,2.1880767,1.8348293,1.7662375,1.978872,2.277246,2.767677,3.4467354,4.2218223,6.6122446,7.2432885,6.5127864,4.98662,3.3678548,3.2581081,2.7779658,2.020027,1.3615463,1.4815818,2.651071,3.6970954,3.7965534,2.9803114,2.1503513,1.2792361,0.8162418,0.61046654,0.53844523,0.48014224,0.4081209,0.28122616,0.15776102,0.082310095,0.08573969,0.09945804,0.12689474,0.18519773,0.23664154,0.18862732,0.2469303,0.29151493,0.24350071,0.14404267,0.14061308,0.08916927,0.12689474,0.216064,0.33609957,0.47328308,0.5007198,0.5041494,0.34981793,0.11317638,0.058302987,0.0274367,0.017147938,0.010288762,0.0,0.0,0.216064,0.18519773,0.20234565,0.3566771,0.53501564,0.85739684,1.0597426,1.3066728,1.488441,1.2072148,1.1866373,1.3649758,1.5158776,1.6016173,1.786815,1.9480057,2.8328393,3.2272418,3.1483612,3.8445675,4.5682106,4.0880685,3.957744,4.523626,4.90431,5.086078,5.967482,6.6876955,7.4936485,9.72631,11.118723,12.394529,14.455711,17.154797,19.277712,20.12139,20.95135,23.557837,27.618467,30.701668,32.793716,35.18071,36.08612,34.878906,32.039207,30.993181,30.015749,27.954567,25.3618,24.51469,27.865398,29.10348,30.557625,33.157253,36.453087,39.74549,43.782112,46.837875,48.343464,48.8922,45.442036,38.23647,37.47853,46.175964,60.141247,54.551018,47.80845,44.31027,43.010456,37.42709,31.072062,26.496992,22.134558,17.312557,12.260776,9.177576,7.3839016,6.4304767,6.8866115,10.340206,8.886061,9.517105,8.772884,6.999788,8.344186,9.122703,9.06097,14.79867,25.005123,30.396433,22.213438,13.900118,6.9517736,4.746549,12.545431,12.264205,16.46545,19.082224,17.971039,14.922135,17.61779,17.017612,13.474849,8.824328,6.385892,6.392751,6.48535,7.274155,7.7028537,5.038064,4.4275975,4.547633,10.39508,16.37971,6.3207297,7.7028537,11.4033785,12.682614,10.690024,8.460793,10.233889,15.179354,18.989626,20.827885,23.35206,23.897366,23.039968,20.436913,17.106783,15.426285,14.390549,14.527733,13.193623,10.72432,10.460241,10.765475,12.096155,13.234778,15.525743,22.865059,19.939621,17.63151,14.918706,12.445972,12.528283,10.0041065,11.550851,10.1481495,6.166398,7.363324,14.79867,13.670336,11.492548,11.338216,11.828648,9.071259,9.033533,9.849775,10.2921915,9.757176,10.371073,9.716022,8.724871,7.8194594,6.8866115,8.056101,12.041282,16.434584,18.488907,15.148488,14.006435,13.310229,12.878101,11.842365,8.663138,14.188204,15.54632,14.150477,12.782072,15.584045,11.989838,12.617453,12.88839,12.034423,13.111313,18.145947,17.027903,13.214201,9.928656,10.161868,14.435134,16.208231,15.282242,12.72034,10.844356,11.513125,11.177026,9.966381,8.471081,7.7440085,9.431366,11.163307,12.05157,12.22305,12.830087,12.878101,12.55229,13.516005,15.580616,16.715809,18.986197,18.756414,19.071936,20.03908,18.835295,14.894698,11.526843,9.225591,8.045813,7.5759587,7.6033955,8.652849,10.834066,13.327377,14.363112,14.644339,13.766364,13.193623,12.490558,9.321619,10.117283,10.563129,10.734609,10.600855,10.041832,9.551401,9.445084,8.995808,8.4264965,8.920357,8.947794,9.647429,9.719451,8.707723,6.9963584,7.0032177,7.06838,6.9860697,6.917478,7.4010496,6.636252,6.5985265,6.667118,6.6876955,6.948344,7.363324,7.1266828,6.6122446,5.9160385,4.839148,4.856296,5.099797,4.9694724,4.73969,5.552502,5.7102633,5.885172,5.7102633,5.394741,5.7479887,5.90575,5.48734,5.435896,5.610805,4.804852,4.5956473,5.2575574,5.6142344,5.669108,6.584808,6.7185616,6.0737996,5.7651367,5.919468,5.689686,5.1409516,5.353586,5.363875,4.9523244,4.633373,4.064061,3.6799474,3.192946,2.6887965,2.6476414,2.9460156,3.0386145,2.843128,2.5138876,2.452155,2.153781,1.8313997,1.7010754,1.7765263,1.8828435,1.9102802,1.9685832,1.8554068,1.5981878,1.4541451,1.3615463,1.2003556,1.155771,1.2277923,1.2312219,0.94999576,0.8471081,0.8162418,0.83338976,0.94656616,0.980862,0.84367853,0.84367853,0.9842916,0.9534253,0.9911508,0.89512235,0.6962063,0.52815646,0.6173257,0.64476246,0.607037,0.6790583,0.8745448,1.0357354,0.8676856,0.9294182,0.96714365,0.91227025,0.89512235,0.9911508,1.0940384,1.1146159,1.0871792,1.1729189,1.1214751,1.155771,1.3649758,1.5810398,1.371835,1.1489118,1.155771,1.2483698,1.3821237,1.605047,1.6496316,1.3203912,1.138623,1.2003556,1.1866373,1.1214751,1.0254467,0.9328478,0.8711152,0.8711152,0.75450927,0.6927767,0.6379033,0.6036074,0.64476246,0.58302987,0.5658819,0.6310441,0.7442205,0.7956643,1.2277923,1.214074,0.9842916,0.7373613,0.65848076,0.71678376,0.7510797,0.7339317,0.6756287,0.61389613,0.61046654,0.6241849,0.66191036,0.7305021,0.82996017,0.8162418,0.7682276,0.6927767,0.6241849,0.6276145,0.70306545,0.5178677,0.26750782,0.10288762,0.11317638,0.07888051,0.08916927,0.1097468,0.16119061,0.30523327,0.28122616,0.35324752,0.47328308,0.6173257,0.7956643,1.2003556,1.4027013,1.646202,1.937717,2.0303159,2.0303159,2.0131679,2.0920484,2.2326615,2.2395205,2.4315774,2.8568463,2.9871707,2.8156912,2.8568463,3.1826572,3.7794054,4.5682106,5.295283,5.5387836,5.6793966,5.8645945,6.042933,6.228131,6.495639,6.9689217,7.7440085,8.625413,9.523964,10.449953,11.519984,12.836946,13.869251,14.263655,13.838386,12.768354,11.616013,10.645439,9.9698105,9.55826,9.469091,9.39021,8.98209,8.399059,8.275595,8.920357,9.266746,9.616563,9.791472,9.098696,9.825768,9.935514,10.233889,11.218181,13.070158,12.864383,12.05843,11.862943,12.432255,12.843805,11.962401,11.341646,11.276484,11.341646,10.38479,10.947243,10.840926,10.854645,11.372512,12.373952,12.860953,14.366542,14.911846,13.924125,12.229909,12.271064,12.603734,12.991278,13.399398,13.982429,16.21166,18.416885,20.135109,21.153696,21.517231,21.187992,20.591244,19.637817,18.478617,17.494326,16.935303,16.564907,17.415445,19.068506,19.62753,20.594673,20.76958,20.27572,19.5315,19.267422,19.277712,19.349733,19.668684,20.673553,23.046827,25.306927,26.315224,26.479845,25.900244,24.377508,24.696459,26.123167,28.715937,31.226395,31.120077,0.65162164,0.7339317,0.91569984,0.9945804,0.939707,0.90541106,0.8196714,0.7613684,0.72364295,0.6962063,0.64133286,0.66191036,0.7099246,0.7990939,0.9431366,1.1317638,1.6221949,2.0063086,2.2566686,2.3767042,2.4212887,2.352697,2.4418662,2.5241764,2.74367,3.5564823,3.724532,4.262977,4.887162,5.6039457,6.7185616,7.0032177,6.9689217,7.0375133,7.5107965,8.543102,10.357354,10.443094,9.030104,7.099246,6.3618846,4.9660425,3.3061223,1.9582944,1.1523414,0.7442205,0.4664239,0.32581082,0.22978236,0.15090185,0.11317638,0.18519773,0.33609957,0.33952916,0.26750782,0.4664239,0.6344737,0.53844523,0.53501564,0.72364295,0.939707,0.7339317,0.5007198,0.37382504,0.36696586,0.3806842,0.31209245,0.32924038,0.33952916,0.34295875,0.42869842,0.52472687,0.52472687,0.6001778,0.77851635,0.94999576,1.0768905,0.939707,0.75450927,0.65162164,0.64819205,0.64819205,0.5796003,0.5590228,0.6344737,0.8025235,0.99801,1.0494537,1.0700313,1.1626302,1.4335675,1.5330256,1.728512,1.7490896,1.6084765,1.6187652,1.4335675,1.488441,1.529596,1.488441,1.4918705,1.8691251,2.6750782,3.4398763,3.957744,4.2869844,4.846007,4.7499785,4.636802,4.7259717,4.8185706,4.15323,3.426158,2.6476414,1.9720128,1.6839274,2.037175,2.5961976,2.8122618,2.7882545,3.2889743,3.3781435,3.642222,4.431027,5.1512403,4.266407,5.219832,5.3913116,4.705394,3.4707425,2.3595562,2.9117198,2.5756202,1.8245405,1.1489118,1.0597426,1.5227368,2.3252604,2.8465576,2.819121,2.318401,1.5638919,1.1489118,0.85739684,0.67219913,0.77851635,0.7682276,0.5453044,0.3018037,0.15433143,0.15776102,0.1920569,0.1920569,0.17147937,0.15090185,0.1371835,0.12346515,0.15090185,0.14747226,0.10288762,0.07545093,0.061732575,0.0548734,0.08573969,0.17147937,0.32581082,0.6379033,0.881404,0.72364295,0.29151493,0.17490897,0.082310095,0.037725464,0.01371835,0.0034295875,0.0,0.1371835,0.20577525,0.2469303,0.29837412,0.4081209,0.64476246,0.7682276,1.0425946,1.3889829,1.3924125,1.4781522,1.7388009,1.6393428,1.3238207,1.6084765,1.9582944,2.952875,3.3026927,3.2443898,4.5510626,4.9351764,4.413879,4.866585,6.118384,5.9297566,5.813151,6.807731,7.9189177,8.872343,10.110424,11.173596,14.38369,17.724108,20.491785,23.321196,22.230585,22.450079,25.02227,28.993732,31.435598,33.116096,34.75201,34.776016,32.797146,29.576763,29.624777,28.92514,28.76395,29.624777,31.209246,34.41248,34.714283,34.50508,35.39334,38.212463,41.22364,44.255398,46.65954,48.744728,51.773052,47.2117,39.4917,39.16246,46.347446,50.751034,43.689514,40.383392,37.862644,34.16212,28.318104,25.485264,24.048267,21.136547,16.561478,12.80608,9.541112,6.869464,6.0978065,7.040943,8.035523,9.599416,8.964942,7.6616983,7.143831,8.796892,9.949233,10.254466,14.918706,22.559826,25.19718,15.87899,7.9086285,3.2718265,3.117495,7.7680154,8.30646,15.278812,20.183123,19.438902,14.390549,18.413456,17.79613,15.37827,11.739478,5.192395,4.266407,5.5593615,8.659708,10.827208,7.010077,5.2644167,5.3570156,5.9297566,6.3207297,6.591667,6.5950966,7.016936,8.244728,9.55826,9.105555,9.825768,13.642899,17.864721,21.674994,26.112879,27.1006,25.797358,23.098272,19.9602,17.422304,15.097044,15.594335,13.594885,9.338767,8.604835,7.7542973,8.934075,9.983529,12.833516,23.499533,21.939072,18.646667,15.515453,14.832966,19.263992,14.771234,13.615462,11.842365,8.419638,5.24041,8.172707,9.547972,11.821788,13.512574,9.218731,9.0644,8.961512,9.9869585,11.605724,11.677745,11.550851,10.515115,8.495089,6.7219915,7.7268605,9.901219,15.8138275,23.36921,26.215767,13.759505,10.350495,12.271064,14.88098,14.260224,7.2192817,12.147599,15.337115,15.618341,13.615462,11.753197,9.568549,10.405369,12.068718,13.841815,16.486027,19.812727,17.669235,14.472859,12.576297,12.257345,18.523201,19.823015,18.581505,16.496315,14.55174,12.826657,11.746337,10.621432,9.554831,9.451943,10.528833,11.372512,13.145609,15.237658,15.275383,15.076467,15.309678,16.609491,18.3723,18.78042,20.258574,20.165974,20.423193,21.342323,21.637268,17.895588,13.663476,10.39508,8.704293,8.368194,9.928656,10.858074,12.6586075,14.71636,14.287662,15.340545,15.357693,15.3302555,14.901558,12.367092,12.432255,12.181894,11.746337,11.489118,12.010415,11.4754,11.1393,10.295622,9.266746,9.403929,9.692014,9.836057,9.321619,8.052671,6.355026,6.6396813,6.9037595,7.2535777,7.671987,8.008087,6.680836,6.183546,6.0978065,6.3001523,6.9552035,7.5725293,6.8763227,5.844017,5.1409516,5.130663,4.7602673,4.8185706,4.9934793,5.2575574,5.8988905,5.9983487,6.1629686,5.720552,5.086078,5.754848,6.23499,5.977771,6.0052075,6.108095,4.863155,4.629943,5.284994,5.658819,5.669108,6.3035817,6.2144127,5.8371577,5.895461,6.2418494,5.878313,5.3741636,5.425607,5.394741,5.0757895,4.7019644,3.9783216,3.590778,3.1243541,2.633923,2.6236343,2.8396983,3.1552205,3.2203827,2.942586,2.5241764,2.2738166,1.7936742,1.5810398,1.670209,1.6530612,1.6016173,1.6633499,1.5638919,1.2998136,1.1454822,1.2106444,1.1249046,1.097468,1.1489118,1.1249046,0.8196714,0.72364295,0.7510797,0.7990939,0.7407909,0.71678376,0.65162164,0.6927767,0.7956643,0.72707254,0.50757897,0.47328308,0.44927597,0.4081209,0.45956472,0.6310441,0.71678376,0.7990939,0.88826317,0.9328478,0.8196714,0.89512235,0.9842916,0.99801,0.9431366,1.1489118,1.2243627,1.0940384,0.91912943,1.097468,1.2072148,1.1797781,1.2517995,1.3992717,1.3341095,1.1351935,1.0940384,1.313532,1.670209,1.8039631,1.704505,1.3306799,1.1111864,1.1660597,1.3101025,1.2175035,1.0940384,1.0048691,0.97057325,0.94999576,0.7888051,0.6001778,0.45613512,0.42183927,0.5418748,0.5521636,0.5693115,0.6344737,0.7510797,0.89512235,1.6187652,1.4781522,1.1351935,0.9431366,0.9259886,0.881404,0.6893471,0.58302987,0.6036074,0.6001778,0.6241849,0.6344737,0.65162164,0.6927767,0.7888051,0.7373613,0.64133286,0.5555932,0.52815646,0.6173257,0.78194594,0.58988905,0.29837412,0.08916927,0.06859175,0.058302987,0.072021335,0.08573969,0.13032432,0.2777966,0.24007112,0.25378948,0.29151493,0.36696586,0.5453044,0.86082643,1.0871792,1.4027013,1.7490896,1.8348293,2.0028791,1.920569,1.961724,2.1263442,2.0234566,2.3904223,2.9494452,3.0969174,2.901431,3.083199,3.4055803,3.9783216,4.6779575,5.3090014,5.56965,5.8062916,5.895461,5.8337283,5.703404,5.6965446,6.3035817,7.085528,8.001227,9.0644,10.350495,11.372512,12.583157,13.858963,14.767803,14.586036,13.450842,12.624311,11.89038,11.1393,10.367643,10.254466,10.017825,9.5205345,8.958082,8.851766,9.609704,9.619993,9.499957,9.537683,9.668007,9.602845,9.421077,9.345626,9.613133,10.484249,9.956093,9.932085,10.528833,11.266195,11.067279,10.55284,10.912948,11.581717,11.766914,10.419086,10.981539,10.251037,10.031544,10.998687,12.699762,12.579727,14.335675,15.237658,14.201921,11.766914,12.401388,12.9638405,13.38225,13.862392,14.918706,17.21996,19.133669,20.567236,21.736725,23.180582,23.012531,22.076254,20.53637,18.53692,16.21166,15.285671,15.114192,16.153357,17.717249,17.977898,16.39,16.067617,16.0539,15.916716,15.721229,16.194511,16.88386,17.95732,19.459478,21.318316,24.651875,25.975695,26.044287,25.61559,25.464687,26.126596,26.239773,28.112328,31.58307,34.052376,0.5178677,0.6276145,0.8471081,1.0185875,1.039165,0.8711152,0.5761707,0.42869842,0.40126175,0.42183927,0.39783216,0.4081209,0.42869842,0.5144381,0.6790583,0.90198153,1.7902447,2.2600982,2.452155,2.4075704,2.0920484,1.9445761,2.1915064,2.3801336,2.5070283,3.0043187,3.275256,3.690236,4.3349986,5.2026844,6.1801167,6.924337,7.0923867,7.0306544,7.0272245,7.3084507,9.163857,9.829198,8.700864,6.39961,4.7774153,3.8960114,2.7882545,1.8725548,1.3443983,1.1592005,0.84367853,0.58988905,0.36353627,0.17490897,0.07545093,0.05144381,0.044584636,0.09602845,0.31895164,0.9294182,0.65162164,0.4698535,0.67219913,1.1489118,1.4027013,0.72021335,0.5590228,0.69963586,0.8711152,0.7476501,0.53844523,0.6344737,0.7373613,0.7099246,0.5658819,0.6001778,0.6756287,0.75450927,0.8505377,1.0220171,0.7407909,0.5796003,0.4938606,0.5007198,0.67219913,0.8162418,0.6344737,0.52472687,0.59674823,0.65505123,0.75450927,0.8711152,0.9431366,0.9842916,1.0666018,1.5673214,1.4815818,1.2380811,1.0940384,1.1283343,1.0425946,1.196926,1.2209331,1.1626302,1.4815818,2.3972816,3.357566,4.6402316,5.8508763,5.936616,5.703404,4.9420357,4.081209,3.525616,3.6456516,2.6579304,2.0646117,1.7936742,1.7936742,2.0131679,2.5138876,3.1620796,3.865145,4.681387,5.830299,5.3878818,5.579939,6.5470824,6.975781,4.1189346,4.448175,4.15666,3.5153272,2.836269,2.4555845,2.5413244,2.1229146,1.5124481,0.9602845,0.65505123,0.8745448,1.2415106,1.6256244,1.8554068,1.7079345,1.7319417,1.611906,1.2758065,0.9259886,1.0220171,1.0220171,0.7305021,0.4046913,0.19548649,0.12346515,0.13375391,0.1371835,0.12003556,0.08916927,0.07545093,0.09945804,0.116605975,0.12346515,0.11317638,0.07545093,0.15090185,0.15776102,0.14061308,0.15433143,0.29151493,0.47328308,0.6276145,0.67219913,0.5761707,0.3806842,0.17490897,0.07545093,0.034295876,0.01371835,0.0,0.0,0.06516216,0.24007112,0.48357183,0.64133286,0.5555932,0.8162418,1.3306799,1.8176813,1.8313997,1.8313997,2.0680413,1.862266,1.4129901,1.8142518,2.8294096,3.117495,3.474172,4.170378,4.99005,5.2575574,5.1683884,5.3090014,5.5147767,4.866585,5.610805,5.8543057,6.842027,8.388771,8.865483,15.395418,19.490345,20.584383,19.672113,19.318867,20.063087,22.316326,25.838512,29.823692,32.91375,33.548225,34.144974,33.469345,30.969175,26.795366,27.611609,28.990303,30.93488,33.50364,36.789185,41.281944,41.81696,40.81552,39.80036,39.3991,38.726902,39.622025,41.100178,43.178505,46.88932,42.82526,35.647133,31.072062,29.59391,26.507282,27.495003,24.572994,19.490345,14.486577,12.315649,11.519984,10.618003,9.006097,7.226141,6.958633,6.7494283,5.2987127,5.0655007,6.351596,7.2775846,8.889491,8.460793,7.4353456,7.3084507,9.626852,8.2481575,9.239308,12.9638405,16.808409,15.199932,9.290752,4.5819287,2.4624438,3.0557625,5.2026844,5.6073756,10.38479,14.345964,15.121051,13.169616,16.304258,19.041069,18.355152,13.697772,6.9723516,5.861165,4.715683,5.2644167,7.4970784,9.657719,8.498518,9.033533,8.416207,6.5539417,6.1046658,8.4093485,10.871792,11.262765,9.654288,8.423067,8.604835,9.575408,18.756414,30.252392,24.85765,30.17694,28.047167,23.581844,19.77843,17.532051,16.798119,14.493437,10.72775,7.2878733,7.630832,7.130112,9.904649,11.866373,13.989287,22.340332,24.61072,22.11055,17.741257,14.867262,17.333136,22.131128,18.735836,16.554619,15.347404,5.2026844,9.170717,14.363112,19.185112,19.630959,9.294182,8.865483,8.282454,9.400499,11.97269,13.656617,13.4474125,10.329918,7.534804,7.5210853,11.962401,10.288762,8.690575,11.523414,14.640909,5.3878818,6.0566516,12.22305,16.091625,15.0456,11.626302,10.333347,11.996697,12.253916,10.288762,8.834618,9.493098,13.166186,15.8138275,16.362562,16.691803,15.5085945,16.29397,17.014183,16.602633,14.970149,20.560377,20.666695,19.603521,19.678972,21.19485,15.738377,14.246507,13.958421,12.977559,10.268185,11.842365,12.000127,14.390549,17.62808,15.275383,17.165085,20.303158,22.03167,21.28402,18.584934,20.697561,22.141417,22.251163,21.819035,23.101702,20.220848,16.6335,13.937843,12.79922,12.9707,13.310229,15.062748,17.912735,19.853882,17.182234,14.335675,11.667457,12.168177,14.4317045,12.648318,12.4802685,13.049581,13.677195,14.099034,14.466,13.646329,13.231348,11.595435,9.541112,10.285333,10.504827,10.072699,9.599416,9.054111,7.795452,7.016936,6.7665763,7.442205,8.423067,8.056101,6.944915,6.228131,5.6793966,5.442755,6.025785,7.160979,6.824879,5.5902276,4.5442033,5.2644167,5.164959,5.360445,5.5387836,5.7651367,6.48535,6.0566516,5.9880595,5.778855,5.5593615,6.0737996,6.9037595,6.992929,6.800872,6.3173003,5.0346346,4.2526884,4.616225,4.928317,4.839148,4.852866,5.425607,5.3398676,5.377593,5.5833683,5.2781353,5.1580997,5.055212,5.0414934,5.007198,4.65395,4.15323,3.690236,3.2272418,2.8088322,2.5619018,3.0043187,3.2581081,3.3026927,3.0866287,2.5481834,2.170929,1.7902447,1.6256244,1.6187652,1.4335675,1.2620882,1.3032433,1.3203912,1.2037852,0.9602845,0.90198153,1.0048691,1.1249046,1.1489118,0.9911508,0.980862,0.8745448,0.9362774,1.1077567,1.0220171,0.70649505,0.5144381,0.44927597,0.50757897,0.70306545,0.53158605,0.4424168,0.4046913,0.42526886,0.53501564,1.0940384,1.1523414,1.1214751,1.1660597,1.1900668,1.2517995,1.2106444,1.0666018,0.881404,0.8093826,0.85739684,1.0254467,1.1351935,1.1729189,1.2826657,1.1489118,1.0494537,1.1180456,1.2963841,1.3581166,1.1489118,1.2826657,1.6290541,1.961724,1.937717,1.5844694,1.2929544,1.1043272,1.0906088,1.3581166,1.4918705,1.196926,0.9534253,0.9259886,0.9602845,0.89855194,0.64819205,0.42183927,0.33266997,0.3806842,0.5418748,0.6173257,0.6893471,0.8093826,0.9911508,1.2003556,1.3169615,1.2175035,0.9602845,0.77851635,0.8505377,0.65848076,0.59331864,0.6859175,0.6241849,0.69963586,0.66191036,0.61389613,0.6310441,0.77851635,0.8505377,0.8711152,0.7305021,0.50757897,0.45613512,0.70306545,0.5796003,0.31895164,0.09259886,0.030866288,0.030866288,0.041155048,0.044584636,0.06859175,0.16804978,0.216064,0.28465575,0.3018037,0.29151493,0.34981793,0.51100856,0.7407909,1.1454822,1.6016173,1.786815,2.1880767,1.8862731,1.8073926,2.0714707,1.9994495,2.2292318,2.7470996,3.0283258,3.059192,3.3266997,3.6799474,4.1635194,4.695105,5.1409516,5.3261495,5.7754254,6.0806584,6.0566516,5.720552,5.295283,5.4907694,6.125243,6.8214493,7.689135,9.338767,10.779194,12.109874,13.574307,14.805529,14.832966,13.7938,12.610593,12.133881,12.22305,11.732618,10.683165,10.038403,9.383351,8.851766,9.108984,9.523964,8.988949,8.786603,9.266746,9.825768,9.253027,9.163857,9.421077,9.959522,10.789482,10.347065,10.604284,10.367643,9.918367,11.015835,10.748327,10.882081,11.334786,11.787492,11.688034,11.96926,11.5645685,11.245617,11.756626,13.807519,12.96727,13.773223,13.852104,12.867812,12.511135,13.817808,15.042171,15.683503,16.46888,19.363451,19.044498,20.834743,22.20658,22.508383,22.9508,22.985096,21.52066,19.603521,17.847572,16.417435,16.088194,15.96816,15.964729,15.817257,15.121051,13.924125,14.5414505,14.774663,14.29452,14.647768,14.270514,14.870691,15.573756,16.314548,17.854433,19.757853,22.038528,24.332924,26.709627,29.662502,30.530188,29.254381,28.472435,29.803116,33.84317,0.42183927,0.490431,0.61389613,0.6927767,0.67219913,0.5418748,0.4424168,0.39783216,0.39097297,0.4046913,0.4081209,0.4389872,0.4972902,0.7442205,1.0734608,1.1077567,1.5090185,2.335549,2.620205,2.318401,2.2738166,2.3321195,2.3801336,2.3458378,2.3218307,2.5790498,3.0214665,3.590778,4.3521466,5.2335505,6.0326443,7.157549,7.6342616,7.548522,7.1849856,7.016936,6.958633,7.298162,7.301592,6.40304,4.214963,3.1792276,2.428148,1.937717,1.6873571,1.6599203,1.3443983,0.980862,0.6379033,0.3566771,0.16119061,0.09945804,0.07545093,0.09945804,0.22635277,0.5521636,0.4972902,0.41498008,0.53501564,0.85396725,1.1592005,0.64133286,0.5007198,0.53844523,0.61046654,0.6241849,0.65162164,0.67219913,0.7476501,0.8265306,0.7613684,0.7682276,0.71678376,0.64476246,0.6036074,0.66876954,0.58302987,0.5521636,0.52815646,0.5041494,0.5007198,0.4424168,0.3841138,0.39440256,0.4972902,0.65505123,0.83338976,0.922559,0.9774324,1.0288762,1.1043272,1.2346514,1.3546871,1.3992717,1.3684053,1.3375391,1.5536032,1.7388009,2.0028791,2.4212887,3.0317552,3.799983,4.681387,5.610805,6.279575,6.1321025,5.254128,4.1463714,3.309552,2.8328393,2.3904223,1.879414,1.8519772,2.2360911,2.9974594,4.125794,4.695105,5.2266912,5.641671,5.953764,6.279575,6.15268,6.416758,6.684266,6.217842,3.9474552,3.8205605,3.3541365,2.942586,2.651071,2.2120838,1.9171394,1.4541451,1.0288762,0.7579388,0.66876954,0.8093826,1.0323058,1.2998136,1.4404267,1.1489118,1.0563129,0.823101,0.5658819,0.40126175,0.44927597,0.4698535,0.37039545,0.25378948,0.18176813,0.19548649,0.23664154,0.23321195,0.18862732,0.12689474,0.07545093,0.09945804,0.20234565,0.22292319,0.13375391,0.041155048,0.044584636,0.037725464,0.034295876,0.048014224,0.09602845,0.15090185,0.18519773,0.20577525,0.20920484,0.19891608,0.1097468,0.0548734,0.020577524,0.0034295875,0.0,0.0,0.041155048,0.24007112,0.47671264,0.42183927,0.864256,1.0460242,1.4507155,1.9685832,1.903421,1.6221949,1.5913286,1.471293,1.7388009,3.6970954,3.069481,3.40901,3.9783216,4.6779575,6.0635104,5.4941993,5.113515,4.554492,4.48933,6.625963,5.857735,7.3290286,9.774324,11.4754,10.281903,13.238208,16.153357,16.86671,15.837835,16.156786,18.217968,23.280039,27.741934,30.732533,34.08667,35.90092,36.075832,34.686848,32.11123,29.041746,31.497332,32.42675,33.970062,37.495678,43.610634,47.770725,49.440933,50.034252,49.677574,47.235706,44.845287,43.7341,44.22453,46.71098,51.663307,50.809338,44.553772,36.878353,29.316114,20.913624,18.173384,14.033872,10.744898,9.153569,8.687145,6.4407654,4.705394,3.875434,3.8171308,3.882293,3.3026927,3.6044965,4.266407,5.1992545,6.742569,8.488229,8.488229,8.176137,8.570539,10.275044,8.086967,6.7494283,9.578837,14.020154,11.657167,7.9086285,4.557922,2.7985435,2.8156912,3.8102717,5.5902276,8.525954,9.80519,9.033533,8.213862,8.820899,9.383351,9.026674,7.716572,6.252138,6.773435,5.3878818,4.962613,6.7665763,10.487679,8.762596,9.177576,11.622872,14.088745,12.668896,12.593445,10.295622,8.951223,8.916927,7.716572,9.177576,11.132441,18.399736,25.670462,17.521763,19.19197,17.583494,14.321958,11.105004,9.709162,10.820349,13.639469,14.448852,12.449403,9.764035,11.382801,12.312219,15.254805,18.835295,17.566347,20.227707,19.164536,16.904436,15.107333,14.575747,17.741257,19.795578,25.811075,28.60619,8.755736,20.097382,20.718138,21.407484,23.19773,17.350283,10.367643,8.755736,11.63659,14.977009,11.595435,8.690575,11.482259,11.900668,8.663138,7.274155,7.4799304,13.54687,24.422092,29.130917,6.8145905,6.684266,8.81747,9.89093,9.499957,10.175586,11.077567,11.495977,11.447963,11.365653,12.082437,12.127021,14.435134,15.896138,15.902997,16.352274,18.927893,20.680412,22.182571,22.70044,20.2037,27.241213,27.724785,25.090862,21.795029,19.315437,17.724108,16.619781,16.431154,16.503176,15.103903,14.589465,14.3974085,15.155347,15.937293,14.273943,16.39,18.259123,19.871029,21.35947,22.978235,21.644127,22.175713,23.406935,24.061985,22.748453,21.380049,18.262554,16.153357,15.614912,14.997586,15.162207,16.780972,19.243416,21.596113,22.576975,17.171944,14.4145565,13.7526455,13.954991,13.101024,15.96816,15.364552,14.79524,15.175924,14.819247,14.246507,13.817808,12.63117,11.197603,11.444533,10.209882,8.98209,8.114404,7.3393173,5.7582774,5.5250654,5.6245236,6.358455,7.2158523,6.8591747,6.1904054,6.217842,6.6396813,6.848886,5.9434752,6.7940125,6.5539417,5.4770513,4.506478,5.2644167,6.3961806,6.1732574,6.2041235,6.852316,7.2295704,6.2247014,5.6176643,5.3844523,5.48734,5.8543057,6.5470824,6.893471,6.7048435,5.9400454,4.7191124,4.756838,5.1580997,5.3741636,5.3227196,5.363875,5.4016004,5.4667625,5.3090014,4.9660425,4.7671266,5.103226,5.188966,5.0620713,4.787704,4.434457,3.9131594,3.4810312,2.9803114,2.527606,2.5378947,2.8911421,3.0077481,2.9288676,2.7299516,2.534465,1.9823016,1.6324836,1.3752645,1.1797781,1.1043272,1.0494537,0.96714365,0.94999576,1.0014396,1.0220171,0.84367853,0.91227025,1.0220171,1.0837497,1.0906088,1.1249046,0.939707,0.9911508,1.214074,1.0117283,0.6344737,0.53158605,0.61046654,0.72707254,0.6893471,0.65505123,0.53501564,0.44927597,0.51100856,0.8162418,1.2003556,1.0906088,0.922559,0.89169276,0.94656616,1.1626302,1.3032433,1.2929544,1.2209331,1.3341095,1.0117283,0.939707,1.0288762,1.1729189,1.2449403,1.2483698,1.214074,1.2620882,1.3958421,1.5158776,1.3958421,1.1626302,1.1832076,1.4369972,1.5090185,1.2449403,1.255229,1.2380811,1.1592005,1.2620882,1.1489118,1.0563129,0.99801,0.96714365,0.9259886,0.805953,0.7133542,0.65848076,0.66533995,0.77165717,0.8025235,0.7373613,0.75450927,0.8848336,1.0288762,1.039165,1.2243627,1.255229,1.0425946,0.75450927,0.8676856,0.77851635,0.77165717,0.84367853,0.72364295,0.805953,0.8162418,0.7956643,0.805953,0.91227025,1.0254467,1.1043272,1.1283343,1.0323058,0.6893471,0.6001778,0.6001778,0.48700142,0.24007112,0.041155048,0.024007112,0.020577524,0.030866288,0.058302987,0.106317215,0.25378948,0.25721905,0.23664154,0.2469303,0.29151493,0.37039545,0.58302987,0.84367853,1.138623,1.5158776,1.8999915,1.7902447,1.7422304,1.8725548,1.8759843,2.1674993,2.6545007,2.9254382,2.9974594,3.3129816,3.6868064,4.029765,4.4516044,4.852866,4.897451,5.439326,5.778855,5.8234396,5.586798,5.195825,5.147811,5.435896,5.9160385,6.6122446,7.716572,9.184435,10.851214,12.30193,13.234778,13.4645605,12.857523,12.085866,11.72233,11.736049,11.502836,10.998687,10.48082,10.131001,10.39508,11.989838,11.605724,10.347065,10.127572,10.916377,10.765475,11.238758,10.209882,9.932085,10.947243,12.082437,10.628291,9.465661,9.283894,10.319629,12.346515,11.47197,10.31277,9.89093,10.14129,9.904649,10.967821,11.4033785,11.338216,11.266195,12.037852,12.651748,13.564018,13.605173,13.087306,13.807519,14.273943,14.774663,16.160215,18.28313,19.984205,20.21399,20.845032,21.20514,21.527521,22.923363,21.544668,19.997925,18.756414,17.689812,16.077906,16.21509,14.997586,13.660047,12.795791,12.373952,12.264205,11.773774,11.413667,11.581717,12.562579,14.205351,16.012743,17.117071,17.775553,19.390888,21.647556,24.36036,26.003132,26.02714,24.840502,26.949697,28.318104,28.822252,29.268099,31.415022,0.34295875,0.36696586,0.4046913,0.4355576,0.4355576,0.40126175,0.39783216,0.8093826,1.1489118,1.2586586,1.3443983,1.2003556,1.0082988,1.0871792,1.4164196,1.646202,2.16064,2.784825,2.7916842,2.294394,2.2463799,2.2909644,2.4555845,2.5173173,2.4795918,2.5619018,2.8019729,3.3712845,4.3007026,5.456474,6.526505,7.205563,7.0752387,6.495639,5.878313,5.6793966,5.422178,5.98463,6.667118,6.6225333,4.870014,2.668219,1.8554068,1.8382589,2.020027,1.8142518,1.4438564,1.0460242,0.69963586,0.44927597,0.3018037,0.18519773,0.1371835,0.1920569,0.34638834,0.5693115,0.6036074,0.5212973,0.53501564,0.6756287,0.7956643,0.47328308,0.4698535,0.5624523,0.64133286,0.6962063,0.7956643,0.84024894,1.0151579,1.2209331,1.0837497,0.9877212,0.91569984,0.7682276,0.6001778,0.6173257,0.5418748,0.5007198,0.5007198,0.5041494,0.4115505,0.32581082,0.3806842,0.5555932,0.7339317,0.6824879,0.8711152,1.0528834,1.2586586,1.4644338,1.5913286,1.5741806,1.5227368,1.5193073,1.605047,1.7456601,2.0165975,2.2635276,2.5893385,3.0729103,3.7553983,4.417309,5.1992545,5.90232,6.121814,5.254128,4.2526884,3.40901,2.8054025,2.4212887,2.1572106,2.1640697,2.6922262,3.5393343,4.5819287,5.7891436,6.3447366,6.475061,6.4304767,6.262427,5.8062916,5.65539,5.3570156,5.2026844,4.914599,3.642222,3.1689389,2.7951138,2.411,2.0131679,1.6942163,1.3924125,0.91912943,0.5658819,0.41840968,0.36010668,0.4664239,0.6241849,0.864256,1.0768905,0.9877212,0.7922347,0.548734,0.42869842,0.48014224,0.6241849,0.5693115,0.4938606,0.4081209,0.33952916,0.32238123,0.30523327,0.28465575,0.24350071,0.18519773,0.13032432,0.14747226,0.21263443,0.20920484,0.13032432,0.058302987,0.037725464,0.041155048,0.05144381,0.06516216,0.072021335,0.06859175,0.061732575,0.061732575,0.07545093,0.08916927,0.06516216,0.06516216,0.0548734,0.030866288,0.010288762,0.0034295875,0.01371835,0.17147937,0.39440256,0.40126175,0.939707,0.84024894,1.0494537,1.6976458,2.0886188,1.5193073,2.0303159,2.393852,2.5790498,3.7348208,3.875434,4.098357,4.4584637,4.835718,4.90431,5.120374,4.434457,3.7142432,3.7931237,5.453044,5.5662203,8.217292,10.439664,11.334786,12.082437,13.917266,15.193072,16.496315,17.919594,19.044498,21.085104,24.909094,28.647345,31.895163,35.722584,37.859215,38.15759,36.943516,34.937206,33.25328,34.693707,35.705437,37.259037,40.685196,47.671265,55.12376,61.62283,65.6766,65.98869,61.461636,57.075195,52.54471,49.512955,49.656998,54.70535,55.813107,50.997967,42.24566,31.91917,22.748453,18.86959,15.395418,12.346515,9.743458,7.589677,4.962613,3.0146074,2.1983654,2.2326615,2.1229146,2.8294096,3.4947495,3.758828,3.9680326,5.195825,6.64997,7.8983397,8.724871,9.431366,10.847785,9.174147,8.018375,11.331357,16.88043,16.256245,9.897789,5.099797,2.651071,2.3801336,3.1620796,4.9420357,6.48535,6.866034,6.3893213,6.5985265,5.5113473,5.3501563,5.130663,5.0414934,6.447624,7.3393173,5.926327,4.996909,6.2247014,10.155008,8.471081,9.39707,10.851214,11.430815,10.39508,10.257896,9.685155,10.017825,10.64201,8.985519,10.408798,12.751206,19.562366,25.76992,17.700102,22.11055,18.550638,14.280802,12.445972,12.044711,10.381361,12.812939,17.322845,20.838173,19.226267,14.863832,12.55229,15.313108,20.724997,20.930773,18.602083,18.025911,17.95732,17.230247,14.781522,16.331696,21.174273,27.374968,28.959436,15.885849,19.997925,17.87158,18.578075,22.659285,22.137987,11.629731,9.956093,12.535142,14.942713,12.936404,15.306249,13.461131,12.202472,12.555719,11.770344,15.772673,21.225718,22.60441,17.518333,6.694555,6.6225333,7.610255,9.030104,10.504827,11.907528,15.704081,15.604623,15.151917,15.666355,16.269962,12.411677,15.4742985,17.70696,16.571766,14.764374,20.066517,21.846472,22.789608,23.959099,24.754763,28.551315,28.616478,28.002583,27.162333,23.952238,22.494663,21.081675,20.526081,20.639257,20.237995,18.79757,18.70154,18.927893,19.006773,19.003344,19.432043,19.521212,20.334024,22.186,24.627867,22.18943,22.11055,22.961088,23.022821,20.296299,20.083664,18.512913,17.662374,17.878439,17.765263,16.935303,19.682402,22.347193,23.225166,22.590693,17.981327,16.20137,14.788382,13.694343,15.29253,18.169954,16.839275,15.717799,15.913286,15.237658,15.165636,14.260224,13.1421795,12.367092,12.439114,10.868362,9.746887,8.433355,6.708273,4.791134,4.8185706,5.4187484,6.166398,6.6876955,6.6636887,6.1458206,6.5642304,7.1266828,7.2604365,6.6053853,6.8969,6.2555676,5.6245236,5.4599032,5.7308407,6.7631464,6.883182,6.6533995,6.420188,6.3173003,5.8817425,5.3090014,5.212973,5.6039457,5.8817425,6.210983,6.776865,6.684266,5.885172,5.1512403,5.1169443,5.0620713,5.0449233,5.144381,5.4667625,5.2575574,5.2918534,5.099797,4.6573796,4.355576,4.9248877,4.887162,4.8151407,4.7499785,4.2046742,3.6285036,3.1655092,2.7333813,2.4315774,2.534465,2.9734523,2.9185789,2.6819375,2.486451,2.452155,1.9480057,1.5810398,1.2758065,1.0631721,1.0494537,1.0837497,1.039165,0.9362774,0.86082643,0.94656616,0.85739684,0.88826317,1.0082988,1.1283343,1.0940384,1.1008976,0.94656616,0.9259886,1.0288762,0.9534253,0.8471081,0.7442205,0.65162164,0.5624523,0.45613512,0.59674823,0.607037,0.6001778,0.72364295,1.1592005,1.3752645,1.1866373,1.0151579,0.9911508,0.94999576,1.0528834,1.255229,1.3169615,1.2655178,1.4095604,1.2449403,1.1317638,1.2723769,1.4918705,1.2449403,1.2380811,1.3169615,1.3889829,1.4610043,1.6496316,1.4541451,1.2963841,1.2346514,1.2517995,1.2380811,1.2449403,1.3203912,1.3478279,1.2723769,1.1077567,0.922559,0.864256,0.86082643,0.8745448,0.91569984,0.91912943,0.91912943,0.89169276,0.84024894,0.7888051,0.8162418,0.8265306,0.8848336,0.99801,1.1111864,1.155771,1.1832076,1.2277923,1.214074,0.9842916,0.9328478,0.83338976,0.7922347,0.7990939,0.7373613,0.9259886,0.9774324,0.922559,0.86082643,0.97400284,0.9431366,0.980862,1.0734608,1.1111864,0.8848336,0.6927767,0.64476246,0.50757897,0.2469303,0.044584636,0.020577524,0.0274367,0.044584636,0.072021335,0.1097468,0.22978236,0.20920484,0.19891608,0.22635277,0.2194936,0.216064,0.32924038,0.50757897,0.7579388,1.155771,1.6016173,1.6427724,1.6530612,1.7662375,1.8999915,2.1846473,2.4761622,2.627064,2.7093742,3.018037,3.433017,4.040054,4.547633,4.7842746,4.671098,5.0277753,5.40503,5.56965,5.470192,5.23698,5.2301207,5.312431,5.562791,6.025785,6.7322803,7.8434668,9.383351,10.738038,11.605724,11.996697,11.670886,11.324498,11.22161,11.293632,11.149589,11.482259,11.598865,11.526843,11.650309,12.6929035,12.171606,10.645439,10.1481495,10.933525,11.506266,11.650309,11.125582,11.05356,11.821788,13.073587,11.664027,11.084427,11.211322,11.674315,11.88352,11.399949,10.820349,10.587136,10.5597,10.028113,10.100135,10.868362,11.441104,11.543991,11.533703,12.041282,12.490558,12.696333,12.864383,13.588025,14.791811,14.983868,16.074476,18.255693,19.994495,20.652975,20.587814,20.364891,20.364891,20.776442,19.065077,17.995045,17.593784,17.28169,15.899568,15.422854,14.040731,12.593445,11.835506,12.421966,11.818358,11.005547,11.032983,11.941824,12.754636,14.688923,16.04361,16.606062,17.014183,18.766703,22.453508,25.831654,27.42641,26.709627,24.130577,24.840502,26.35981,27.982004,29.199507,29.710516,0.31209245,0.31552204,0.32581082,0.4389872,0.7682276,1.4267083,1.7833855,2.3046827,2.469303,2.294394,2.3389788,2.07833,1.728512,1.6153357,1.8382589,2.2978237,3.0077481,3.3129816,3.069481,2.4898806,2.1194851,2.0063086,2.1812177,2.294394,2.2429502,2.1983654,2.386993,2.9734523,3.9028704,5.079219,6.358455,6.6053853,6.23156,5.6142344,5.1992545,5.4976287,5.453044,5.8474464,6.4236174,6.5024977,4.972902,2.194936,1.488441,1.6839274,1.9651536,1.8485477,1.4232788,1.0048691,0.6893471,0.4972902,0.37382504,0.28122616,0.29837412,0.39783216,0.5521636,0.7133542,0.6276145,0.5212973,0.5521636,0.6927767,0.7305021,0.45956472,0.45270553,0.5453044,0.6276145,0.66533995,0.82996017,0.94999576,1.1077567,1.2517995,1.2003556,1.1008976,1.1008976,0.980862,0.764798,0.72707254,0.70649505,0.6790583,0.66876954,0.64476246,0.4972902,0.4664239,0.548734,0.7407909,0.9362774,0.90884066,1.1214751,1.4027013,1.6393428,1.8073926,1.9514352,1.8828435,1.6599203,1.6221949,1.8245405,2.037175,2.4452958,2.877424,3.2478194,3.6319332,4.2766957,5.0140567,5.7479887,6.0497923,5.638242,4.3761535,3.3850029,2.843128,2.5619018,2.4144297,2.3389788,2.8739944,3.5633414,4.5339146,5.5662203,6.1321025,6.262427,5.830299,5.4187484,5.086078,4.3658648,4.290414,3.8377085,3.7519686,3.8617156,3.1106358,2.5173173,2.0817597,1.7079345,1.3752645,1.138623,0.8745448,0.52815646,0.3018037,0.23664154,0.21263443,0.34981793,0.5727411,0.805953,0.96371406,0.9328478,0.7133542,0.5212973,0.5212973,0.7305021,1.0220171,0.82996017,0.65848076,0.4972902,0.36353627,0.30523327,0.30866286,0.33952916,0.36010668,0.33609957,0.26064864,0.24350071,0.22635277,0.17833854,0.106317215,0.05144381,0.048014224,0.061732575,0.06859175,0.06859175,0.06859175,0.041155048,0.030866288,0.030866288,0.041155048,0.041155048,0.041155048,0.072021335,0.07888051,0.05144381,0.01371835,0.0034295875,0.0,0.07545093,0.2194936,0.33609957,0.66191036,0.5418748,0.70306545,1.2723769,1.762808,1.3478279,2.0920484,2.5310357,2.5310357,3.3026927,4.1600895,4.5682106,4.671098,4.5613513,4.262977,5.038064,4.5819287,4.0709205,4.232111,5.3330083,6.9654922,9.983529,12.30193,13.886399,16.763824,16.108772,16.064188,16.842705,18.276272,19.826445,22.11398,25.351511,29.309254,33.4179,36.76175,38.30506,38.881233,38.291344,36.868065,35.482513,35.537384,36.134132,37.365356,40.177616,46.371452,53.38153,61.51994,66.33508,65.83779,60.52536,56.090904,50.4801,46.29943,45.36315,48.669277,49.69129,45.249977,36.826912,27.261791,20.735287,18.392878,16.739817,14.287662,10.88551,7.7131424,5.254128,3.3952916,2.277246,1.7833855,1.5330256,2.633923,3.3541365,3.4021509,3.2581081,4.15323,5.439326,7.2775846,8.669997,9.530824,10.683165,9.770895,9.746887,13.347955,19.696121,24.326063,14.167625,6.560801,2.8225505,2.620205,3.974892,5.0655007,5.796003,6.0532217,5.9880595,6.036074,4.5201964,4.5853586,4.9831905,5.6519604,7.723431,9.352485,7.98408,7.1712675,8.553391,11.866373,10.189304,9.89436,9.884071,9.97324,10.8958,9.126132,9.517105,10.343636,10.5597,9.794902,11.262765,12.860953,21.160555,29.683079,18.883308,27.68363,24.377508,18.866161,16.671225,18.948471,14.417986,12.548861,17.336565,25.18003,24.878227,17.04848,12.130451,13.05301,18.437462,22.580404,17.71039,17.55263,18.962189,19.37374,16.7844,16.894148,20.141968,23.547548,24.699888,21.740154,17.943602,14.7197895,15.940722,20.443771,22.021381,13.728639,11.430815,12.154458,13.704632,14.668345,18.296848,14.308239,16.420864,22.350622,13.828096,15.436573,18.468328,15.035312,7.0478024,6.2075534,7.3873315,10.659158,12.099585,12.2093315,15.923574,23.393215,23.10856,20.714708,19.421753,20.008213,14.956431,17.545769,19.823015,18.338005,14.140189,20.244854,22.196291,22.20315,22.546108,25.61559,25.420103,24.730755,26.02371,28.637054,28.76738,27.77966,26.03057,24.411804,23.36578,22.851341,21.825895,22.055677,22.004232,21.674994,22.60441,22.731306,21.873909,21.606401,22.408924,23.681301,21.969936,22.666143,22.830763,21.242865,18.36887,18.650097,19.03078,19.236557,19.29143,19.521212,19.408035,22.635277,24.377508,23.509823,22.60098,18.386019,16.571766,15.073037,14.531162,18.344864,18.838724,17.415445,16.407146,16.112202,14.784951,15.920145,15.0250225,13.797231,13.162757,13.282792,11.976119,10.964391,9.139851,6.701414,5.1580997,4.972902,5.5079174,6.060081,6.3824625,6.711703,6.416758,7.140401,7.5690994,7.3118806,6.90033,6.8111606,6.0737996,5.8200097,6.1904054,6.324159,6.9380555,7.1849856,6.7665763,5.8405876,5.003768,5.137522,4.976331,5.212973,5.8817425,6.3447366,6.228131,6.5367937,6.444195,5.8817425,5.5490727,5.446185,4.99005,4.6882463,4.804852,5.3741636,5.2644167,5.178677,4.8905916,4.4413157,4.1463714,4.602506,4.5956473,4.636802,4.6848164,4.15666,3.4878905,2.8225505,2.3561265,2.2600982,2.6853669,3.1140654,2.9734523,2.6133456,2.3252604,2.3424082,1.9239986,1.5741806,1.3066728,1.1454822,1.0940384,1.1077567,1.0940384,0.9911508,0.85739684,0.8471081,0.922559,0.90884066,0.980862,1.1249046,1.155771,1.1420527,0.980862,0.881404,0.8745448,0.805953,0.8848336,0.8265306,0.6893471,0.548734,0.48700142,0.67219913,0.7510797,0.85396725,1.0631721,1.4267083,1.529596,1.2998136,1.1111864,1.08032,1.0768905,1.1008976,1.2689474,1.3478279,1.313532,1.3615463,1.3649758,1.2929544,1.4129901,1.5810398,1.2209331,1.2483698,1.371835,1.4987297,1.5913286,1.6770682,1.4335675,1.4404267,1.4335675,1.3272504,1.2072148,1.3169615,1.3615463,1.3924125,1.3443983,1.039165,0.8711152,0.78194594,0.7407909,0.75450927,0.89855194,1.039165,1.0734608,1.0151579,0.89169276,0.72021335,0.7922347,0.90198153,0.9774324,1.0185875,1.1111864,1.1832076,1.1592005,1.1797781,1.2175035,1.0666018,0.939707,0.8745448,0.8471081,0.84367853,0.8676856,0.9534253,0.9568549,0.91912943,0.89169276,0.9362774,0.9602845,0.9774324,1.0734608,1.1694894,1.0323058,0.8711152,0.8676856,0.71678376,0.37725464,0.07545093,0.037725464,0.030866288,0.044584636,0.072021335,0.10288762,0.16119061,0.15776102,0.16462019,0.18176813,0.13375391,0.106317215,0.14061308,0.25721905,0.4629943,0.7613684,1.2037852,1.3992717,1.4953002,1.6256244,1.8999915,2.0920484,2.201795,2.2738166,2.417859,2.8294096,3.2546785,3.8685746,4.3109913,4.4413157,4.341858,4.619654,5.0003386,5.223262,5.2301207,5.1683884,5.2164025,5.271276,5.4084597,5.6965446,6.1629686,6.852316,8.06639,9.235879,10.086417,10.679735,10.652299,10.576848,10.700313,11.022695,11.286773,11.712041,12.380811,12.545431,12.212761,12.144169,12.000127,10.816919,10.285333,10.868362,11.787492,11.297061,11.283342,11.640019,12.401388,13.732068,12.641459,12.490558,12.483699,12.017275,10.662587,10.803201,11.032983,11.2250395,11.0981455,10.230459,9.170717,10.034973,11.262765,11.873232,11.447963,11.451392,11.835506,12.271064,12.566009,12.63803,14.195063,14.407697,15.254805,17.147938,18.934752,20.27572,20.484926,20.258574,19.977346,19.696121,17.881868,17.312557,17.388008,17.267973,15.861842,15.011304,14.1299,13.474849,13.485138,14.774663,13.862392,13.138749,13.279363,14.016724,14.150477,15.539461,16.462019,16.386568,15.844694,16.438013,19.775002,23.883648,26.675331,26.881107,24.082563,22.868488,22.991955,24.655304,27.083452,28.537598,0.32238123,0.36010668,0.47328308,0.94656616,1.903421,3.309552,3.9714622,4.2081037,3.858286,3.2649672,3.2443898,3.018037,2.5070283,2.1332035,2.1434922,2.6236343,3.4364467,3.590778,3.3198407,2.767677,1.9857311,1.6839274,1.670209,1.6667795,1.5810398,1.4987297,1.8245405,2.4761622,3.2958336,4.232111,5.346727,5.48734,5.48734,5.3844523,5.528495,6.5779486,6.5985265,6.3207297,6.2898636,6.142391,4.616225,2.0303159,1.4198492,1.4095604,1.4164196,1.6290541,1.3512574,0.9774324,0.7133542,0.58302987,0.4355576,0.4355576,0.52815646,0.64133286,0.7510797,0.881404,0.6310441,0.5521636,0.6790583,0.88826317,0.91912943,0.71678376,0.66876954,0.66533995,0.64133286,0.58988905,0.8025235,0.9328478,0.94656616,0.91912943,1.039165,1.0631721,1.2106444,1.196926,1.0048691,0.881404,0.96371406,1.0288762,1.0700313,1.0323058,0.8196714,0.89512235,0.9534253,1.0837497,1.2758065,1.4404267,1.6427724,1.8999915,2.0097382,2.020027,2.2429502,2.1297739,1.7765263,1.6873571,1.9068506,2.0303159,2.651071,3.3232703,3.7965534,4.139512,4.7362604,5.7308407,6.5642304,6.5367937,5.552502,4.1292233,3.1243541,2.6990852,2.6716487,2.784825,2.6990852,3.415869,3.841138,4.5956473,5.377593,4.9591837,4.4721823,3.7691166,3.292404,3.0626216,2.644212,2.767677,2.6476414,2.7813954,2.959734,2.2566686,1.7662375,1.196926,0.90884066,0.8676856,0.65162164,0.4081209,0.28808534,0.25378948,0.28122616,0.34981793,0.5453044,0.85396725,1.0357354,1.0151579,0.8711152,0.6756287,0.6001778,0.6756287,0.91912943,1.3443983,1.0220171,0.72364295,0.47671264,0.31895164,0.2709374,0.3806842,0.5041494,0.5693115,0.53844523,0.40126175,0.33609957,0.2503599,0.15433143,0.06859175,0.017147938,0.041155048,0.058302987,0.05144381,0.030866288,0.030866288,0.006859175,0.0034295875,0.017147938,0.030866288,0.024007112,0.024007112,0.0548734,0.06516216,0.044584636,0.020577524,0.0274367,0.0274367,0.041155048,0.08573969,0.18862732,0.274367,0.5212973,0.9431366,1.3478279,1.3306799,1.4747226,1.8862731,1.9102802,1.9891608,3.6696587,3.9063,4.537344,4.57507,4.1772375,4.629943,5.4804807,5.442755,5.254128,5.562791,6.9689217,9.499957,12.572867,15.844694,19.013634,21.815605,18.931322,19.054789,18.506054,17.223389,18.739265,20.742146,24.621008,29.978024,35.046955,36.710304,36.902363,37.262466,37.224743,36.432507,34.75201,34.127827,33.397324,33.67855,35.650562,39.539715,41.443134,46.079937,48.12054,45.97362,41.796383,39.501987,36.81319,35.846046,36.49081,36.429077,35.91121,31.219534,24.068846,17.20967,14.424845,15.285671,15.073037,13.310229,10.463672,7.939495,5.7068334,4.0606318,2.7368107,1.7833855,1.5364552,1.7765263,2.417859,2.6956558,2.8122618,3.940596,5.055212,6.464772,7.8023114,8.838047,9.465661,8.858624,10.80663,15.29596,22.12084,30.890295,18.149376,8.110974,3.4192986,3.7382503,5.7479887,6.3961806,7.291303,7.7440085,7.5245147,6.869464,5.442755,6.186976,7.140401,7.795452,9.102125,12.020704,12.075578,13.642899,16.660936,16.606062,14.836395,11.71547,11.122152,13.502286,15.875561,11.351934,9.945804,9.246168,8.700864,9.609704,10.991828,13.694343,24.428951,34.474213,19.692692,29.08633,27.50872,21.726437,18.471758,24.43238,20.735287,14.225929,15.782962,23.458378,22.484375,17.21653,12.408247,11.650309,15.093615,19.480057,17.233677,17.473747,18.962189,20.069946,18.763273,18.485476,17.648657,18.317427,20.731855,23.321196,18.12194,15.745236,15.594335,16.61292,17.29884,15.501736,12.343085,11.091286,12.445972,14.538021,16.417435,16.050468,22.563255,28.777668,11.207891,8.093826,9.043822,9.712592,8.81747,8.124693,11.667457,15.899568,15.237658,12.79922,20.395756,30.85257,31.181808,27.025148,23.266321,24.010542,21.211998,21.630407,22.930222,22.374628,16.818697,20.62897,22.44322,21.585823,20.083664,22.676432,20.443771,19.816156,21.53438,25.20061,29.271528,30.053474,28.709076,26.370098,24.380938,24.267761,23.245745,23.506393,23.125708,22.141417,22.570116,24.140865,23.636717,22.820475,22.511812,22.570116,22.161995,23.310905,22.748453,20.189981,18.327715,18.550638,20.378609,21.067955,20.248285,19.912186,21.554956,24.675882,25.070284,22.899355,22.683292,17.912735,15.498305,14.860402,16.245956,20.714708,18.79757,17.62465,16.859852,15.889278,13.834956,16.475739,16.139639,14.71636,13.601744,13.684054,12.908967,11.753197,9.541112,6.9792104,6.1458206,5.610805,5.6793966,5.970912,6.279575,6.6053853,6.5127864,7.490219,7.915488,7.31531,6.3790326,6.23156,6.166398,6.2247014,6.4236174,6.742569,7.06495,6.869464,6.3790326,5.579939,4.2252517,4.5099077,4.9008803,5.4804807,6.2144127,6.9380555,6.6122446,6.3378778,6.111525,5.90232,5.641671,5.5833683,5.0620713,4.6676683,4.729401,5.288424,5.446185,5.2815647,4.8425775,4.3521466,4.201245,4.2835546,4.4241676,4.4927597,4.386442,4.029765,3.3987212,2.5996273,2.1194851,2.2326615,2.9665933,3.1895163,3.0729103,2.6990852,2.3046827,2.2806756,1.8588364,1.5364552,1.3478279,1.255229,1.1592005,1.0597426,1.0048691,0.9877212,0.96371406,0.85396725,1.0117283,0.97057325,0.9774324,1.1214751,1.3272504,1.2826657,1.0494537,0.939707,0.9294182,0.65162164,0.6893471,0.70306545,0.71678376,0.7407909,0.764798,0.89169276,0.9945804,1.2003556,1.4644338,1.5913286,1.5947582,1.371835,1.1351935,1.0563129,1.2483698,1.2758065,1.3752645,1.4541451,1.4610043,1.3786942,1.3306799,1.2723769,1.313532,1.3821237,1.2243627,1.3889829,1.4507155,1.5707511,1.7113642,1.6187652,1.3924125,1.471293,1.5364552,1.4644338,1.3101025,1.3203912,1.3341095,1.3375391,1.2620882,1.0048691,0.88826317,0.8093826,0.77165717,0.7990939,0.9328478,1.0768905,1.0837497,0.99801,0.8745448,0.78194594,0.8471081,0.9431366,0.9774324,0.980862,1.08032,1.1283343,1.1866373,1.2380811,1.214074,0.99801,0.89512235,0.91569984,0.9328478,0.9294182,0.99801,0.90884066,0.8676856,0.89855194,0.94999576,0.85739684,1.0837497,1.1317638,1.2037852,1.2929544,1.1729189,1.0528834,1.1729189,1.0734608,0.66191036,0.21263443,0.13032432,0.061732575,0.034295876,0.0548734,0.07888051,0.08573969,0.106317215,0.12003556,0.106317215,0.0548734,0.0548734,0.061732575,0.12346515,0.2503599,0.4046913,0.7613684,1.0837497,1.2860953,1.4369972,1.7525192,1.8588364,1.9068506,2.0063086,2.253239,2.726522,3.1312134,3.4638834,3.6868064,3.8137012,3.8857226,4.15323,4.479041,4.73969,4.8905916,4.98662,5.007198,5.0929375,5.2335505,5.453044,5.802862,6.217842,7.0752387,7.956643,8.707723,9.448513,9.81205,9.839486,10.028113,10.6145735,11.598865,11.55428,12.55229,12.946692,12.298501,11.38623,11.561139,11.129011,10.9369545,11.255906,11.797781,11.101575,11.087856,11.578287,12.46312,13.694343,12.867812,12.528283,11.986408,10.967821,9.613133,10.175586,10.768905,11.235329,11.262765,10.360784,9.067829,9.80519,11.235329,12.212761,11.80121,11.238758,11.667457,12.147599,12.195613,11.794352,12.936404,13.402828,14.373401,15.995596,17.388008,19.089085,20.080235,20.272291,19.987637,19.95677,18.235117,17.87501,17.820137,17.29198,15.786391,15.446862,15.282242,15.590904,16.410576,17.521763,17.04505,16.62664,16.2974,15.971589,15.446862,16.266533,17.302269,17.182234,15.841265,14.520873,14.980438,18.79071,23.043398,25.464687,24.408375,22.12427,20.27572,20.491785,23.02968,26.77822,0.33609957,0.4698535,0.9534253,2.2463799,3.882293,4.4550343,4.3590055,4.5339146,4.5270553,4.3795834,4.623084,4.513337,3.2855449,2.194936,1.7936742,1.9548649,2.942586,3.2615378,3.1517909,2.719663,1.937717,1.546744,1.3581166,1.2243627,1.1454822,1.2655178,1.4369972,2.0920484,3.0351849,3.9543142,4.4550343,4.5647807,4.7842746,5.0346346,5.5662203,6.958633,7.0546613,6.3310184,6.0669403,6.2898636,5.751418,2.8705647,1.4198492,0.764798,0.5418748,0.64133286,1.1043272,0.9842916,0.82996017,0.8162418,0.71678376,0.75450927,0.6790583,0.71678376,0.90541106,1.1146159,1.0768905,1.1420527,1.2037852,1.1489118,0.8711152,1.2346514,1.5570327,1.5090185,1.138623,0.8711152,0.96714365,0.864256,0.8093826,0.84367853,0.7922347,0.96371406,1.2723769,1.3821237,1.2243627,0.9911508,1.0048691,1.2003556,1.5227368,1.7353712,1.4198492,1.6393428,1.786815,2.1160555,2.4795918,2.318401,2.3081124,2.277246,2.3081124,2.534465,3.1586502,2.9871707,2.194936,1.646202,1.5913286,1.6633499,2.2258022,2.9871707,3.6456516,4.173808,4.822,6.090947,7.2775846,7.7680154,7.0478024,4.715683,3.7519686,3.3644254,3.3026927,3.3609958,3.3712845,3.2375305,3.2958336,3.649081,3.82399,2.760818,2.2360911,2.2978237,2.2429502,1.9857311,2.061182,2.1332035,1.903421,1.5501735,1.2072148,0.9602845,0.71678376,0.51100856,0.3806842,0.31209245,0.21263443,0.16462019,0.18176813,0.25378948,0.37382504,0.53501564,0.71678376,0.864256,0.90198153,0.86082643,0.8848336,0.6276145,0.764798,0.89512235,1.0117283,1.5261664,1.1832076,0.8505377,0.65505123,0.6241849,0.6859175,0.83338976,0.91569984,0.82996017,0.61046654,0.42869842,0.34295875,0.18176813,0.072021335,0.041155048,0.030866288,0.041155048,0.06516216,0.058302987,0.030866288,0.030866288,0.006859175,0.017147938,0.030866288,0.024007112,0.0,0.0,0.010288762,0.01371835,0.020577524,0.044584636,0.13032432,0.14404267,0.20577525,0.274367,0.15090185,0.3841138,1.1660597,2.253239,2.9665933,2.1983654,2.819121,2.9220085,2.6956558,3.1312134,6.012067,4.180667,4.0434837,4.3349986,4.4104495,4.2252517,5.98463,5.3330083,5.2301207,6.495639,7.8126,9.815479,14.387119,18.571217,20.556948,19.713268,21.94936,25.26234,25.34122,23.050257,24.428951,22.426073,24.61072,30.365568,36.185577,35.66085,34.08667,32.84173,32.694256,33.273857,33.06465,32.34444,29.539038,28.410702,29.35727,29.419,27.076593,26.040857,24.69303,22.813616,21.592682,21.836184,25.68761,31.325851,35.012657,31.082352,29.569902,26.479845,21.225718,15.683503,14.205351,17.830425,16.338554,12.922686,9.626852,7.3564653,4.9248877,3.5942078,2.534465,1.5638919,1.1592005,1.0734608,0.7888051,0.764798,1.5364552,3.707384,3.8171308,4.5510626,6.118384,7.6616983,7.233,6.1458206,12.236768,21.397196,29.154922,30.670801,17.802988,7.747438,3.865145,5.2609873,6.773435,8.399059,11.111863,12.178465,11.592006,12.068718,9.335337,10.710602,10.39508,7.98065,8.467651,11.97269,17.562918,26.949697,33.68541,23.163433,21.671564,16.750105,15.614912,18.193962,17.1205,13.495427,10.813489,9.4862385,9.3764925,9.781183,9.122703,21.297739,32.900032,35.14641,23.880217,23.917942,19.384027,14.771234,14.339106,22.12427,26.006561,20.066517,17.250826,18.893597,14.695783,14.438563,14.610043,16.400288,18.159666,15.426285,18.550638,18.399736,17.960749,18.238546,18.248835,20.237995,18.327715,17.364002,18.560926,19.500635,19.819586,21.006224,16.46545,8.875772,10.192734,13.512574,11.451392,10.467101,11.718901,11.046701,22.20315,24.682741,18.646667,10.13786,11.063849,16.78783,13.780083,13.680624,17.744686,16.828985,23.310905,17.12393,12.130451,14.472859,22.566685,32.32043,35.383053,34.4845,32.23812,31.126936,29.491022,28.441568,29.816833,31.061773,25.252052,22.237446,21.575535,19.922474,17.62122,18.708399,17.854433,19.963629,21.599543,21.94936,22.827333,24.535269,25.20061,24.77534,25.111439,29.967735,24.85422,24.003683,23.485815,21.973368,20.752434,22.93708,23.647005,24.068846,24.830214,25.999702,25.464687,22.288889,20.265432,20.268862,20.29287,20.426622,22.035099,22.77589,21.839613,19.973917,20.522652,25.008553,26.737064,23.502962,17.593784,14.003006,13.365103,14.870691,17.54234,20.2037,19.932762,18.612371,17.103354,15.690363,14.054449,17.250826,17.20967,15.494876,13.622321,13.059869,12.939834,11.763485,9.647429,7.3050213,6.0737996,5.888602,6.1629686,6.5779486,6.7631464,6.2864337,5.8234396,6.831738,7.6376915,7.233,5.2781353,5.2301207,6.7185616,7.3839016,6.852316,6.728851,6.742569,5.802862,5.2472687,5.2026844,4.5922174,4.887162,5.720552,6.2555676,6.4133286,6.852316,7.034084,6.584808,6.262427,6.1561093,5.693115,5.1066556,4.8322887,4.945465,5.2781353,5.3878818,5.5833683,5.528495,5.1752477,4.7019644,4.530485,4.2526884,4.125794,3.9611735,3.642222,3.1277838,2.9940298,2.6750782,2.6819375,3.0146074,3.1723683,3.07634,3.0248961,2.860276,2.585909,2.3664153,1.7799559,1.3855534,1.1900668,1.1729189,1.2826657,1.0734608,0.939707,0.9534253,1.0631721,1.097468,1.0494537,1.0837497,1.1934965,1.3649758,1.5707511,1.3409687,1.0906088,1.1317638,1.2517995,0.70306545,0.59331864,0.5453044,0.59674823,0.70649505,0.77851635,0.97400284,1.3066728,1.6359133,1.8245405,1.7388009,1.5570327,1.4472859,1.2517995,1.1008976,1.4198492,1.3203912,1.4541451,1.5741806,1.587899,1.5261664,1.2312219,1.0768905,1.138623,1.3341095,1.4198492,1.7593783,1.6804979,1.5844694,1.5913286,1.5570327,1.3615463,1.4027013,1.4164196,1.3203912,1.2346514,1.2483698,1.2689474,1.1523414,0.91912943,0.7476501,0.7099246,0.77508676,1.0254467,1.2998136,1.1900668,1.08032,0.980862,0.88826317,0.8779744,1.097468,0.9877212,0.8779744,0.91569984,1.0940384,1.2517995,1.3478279,1.371835,1.605047,1.8039631,1.2037852,0.9362774,0.91569984,0.82996017,0.66876954,0.71678376,0.9602845,1.1317638,1.155771,1.039165,0.8711152,0.96714365,1.0288762,1.1008976,1.2209331,1.4027013,1.1489118,1.2106444,1.1797781,0.922559,0.5796003,0.4081209,0.1920569,0.06859175,0.06859175,0.09259886,0.06859175,0.061732575,0.0548734,0.041155048,0.030866288,0.030866288,0.030866288,0.048014224,0.09945804,0.19891608,0.4664239,0.8093826,1.1146159,1.313532,1.371835,1.6187652,1.7525192,1.978872,2.2498093,2.2738166,2.6887965,3.0317552,3.2546785,3.3952916,3.5564823,3.433017,3.642222,4.098357,4.619654,4.914599,4.9248877,4.846007,4.914599,5.164959,5.446185,5.874883,6.375603,6.869464,7.3598948,7.936065,8.776315,8.858624,8.841476,9.328478,10.878652,11.135871,12.555719,13.282792,12.730629,11.581717,11.032983,11.197603,11.427385,11.616013,12.175035,12.116733,11.979549,11.773774,11.71547,12.253916,11.787492,11.88352,11.125582,9.736599,9.551401,10.2236,11.032983,11.684605,12.006986,11.948683,11.729189,11.928105,12.507706,13.193623,13.474849,11.777204,10.840926,10.796341,11.393089,11.979549,13.101024,13.9481325,14.946142,16.095055,16.997036,17.192522,18.056778,18.605513,18.674105,18.907316,18.259123,17.748116,16.96617,15.981877,15.333686,16.37285,16.496315,16.818697,17.412016,17.302269,17.401728,17.470318,16.726099,15.470869,15.107333,16.071047,17.144508,18.108221,18.341434,16.815268,13.214201,13.677195,17.04162,22.172283,27.985434,26.140316,22.69358,20.083664,19.795578,22.384918,0.432128,2.2566686,2.877424,2.983741,3.316411,4.650521,5.137522,5.857735,5.977771,5.5902276,5.6965446,4.746549,3.0043187,1.8656956,1.7422304,2.037175,1.8862731,1.8691251,1.7730967,1.6804979,1.9754424,1.7593783,1.6736387,1.5330256,1.3786942,1.4610043,1.6530612,1.7559488,2.311542,3.175798,3.5393343,3.8171308,4.15666,4.262977,4.256118,4.698535,5.099797,4.4721823,3.789694,3.7622573,4.835718,3.4981792,2.1332035,1.0837497,0.50757897,0.37382504,0.45613512,0.48014224,0.5658819,0.7476501,0.97400284,1.3924125,1.5604624,1.5776103,1.6564908,2.1263442,2.4041407,2.3767042,2.0131679,1.4335675,0.91912943,1.3032433,1.5844694,1.7559488,1.7182233,1.2860953,1.1660597,1.1626302,1.0837497,0.91912943,0.82996017,1.0700313,1.1660597,1.1832076,1.2277923,1.4438564,1.9239986,2.3389788,2.6613598,2.8122618,2.6407824,2.760818,3.192946,3.6525106,3.8891523,3.6627994,2.860276,2.2052248,2.085189,2.3732746,2.452155,2.5721905,2.2052248,1.879414,1.9137098,2.3972816,3.4844608,4.7088237,5.689686,6.3481665,6.8969,7.0718093,7.130112,6.8283086,6.1732574,5.422178,4.2252517,3.6079261,3.3061223,3.0797696,2.750529,2.3904223,2.2600982,2.2326615,2.153781,1.8348293,1.5810398,1.7250825,1.5741806,1.1111864,0.99801,1.08032,1.0528834,0.91912943,0.7373613,0.6207553,0.48357183,0.4424168,0.4938606,0.5624523,0.4938606,0.33952916,0.37039545,0.41840968,0.4629943,0.6310441,0.65848076,0.61389613,0.5555932,0.53501564,0.5693115,0.5761707,0.64476246,0.8196714,1.0768905,1.3546871,1.08032,0.7305021,0.53501564,0.5796003,0.7956643,1.0597426,1.039165,0.8505377,0.6379033,0.5624523,0.52472687,0.37039545,0.29151493,0.28122616,0.15090185,0.116605975,0.07545093,0.05144381,0.05144381,0.030866288,0.024007112,0.034295876,0.0274367,0.0034295875,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.010288762,0.0274367,0.037725464,0.05144381,0.06859175,0.041155048,0.09945804,1.6633499,3.3301294,4.3521466,4.6265135,6.958633,6.2247014,5.9400454,7.034084,7.8537555,6.7357097,7.840037,8.419638,7.997798,8.351046,9.026674,8.258447,8.440215,10.052121,11.694893,15.4914465,17.703531,18.886738,19.397747,19.384027,16.70552,20.697561,26.294647,31.517908,37.464813,34.182697,31.140654,30.327843,31.572783,32.522778,31.222963,30.324413,30.567913,31.730543,32.625664,31.58307,26.966846,24.182022,24.84736,26.795366,24.617579,23.887077,21.997374,19.401176,19.62753,22.076254,31.202387,41.353966,47.101955,43.24024,43.483738,38.277626,27.772799,17.185663,16.780972,71.592636,43.199085,11.924676,6.368744,3.3747141,1.9994495,1.6599203,1.3546871,0.881404,0.82996017,0.6173257,0.52472687,0.94999576,1.6187652,1.5844694,2.1640697,4.0537724,5.288424,5.394741,5.377593,3.7725463,9.860064,17.758404,24.17859,28.438139,14.417986,6.228131,4.9351764,7.949784,9.033533,8.128122,11.461681,13.015285,11.574858,10.703742,11.80464,17.370861,19.641247,16.170506,9.822338,11.71547,15.169065,19.517782,21.112541,13.323947,16.852993,16.818697,15.395418,14.195063,14.2533655,13.838386,12.120162,11.55428,11.931535,10.39165,8.580828,13.145609,18.331144,22.391777,27.577312,23.434372,22.583834,21.078245,19.089085,20.879328,20.738716,19.102802,16.53747,13.152468,8.591117,8.354475,13.653188,18.547209,19.490345,15.340545,17.96761,19.881319,19.226267,17.20967,18.091074,19.19197,19.723558,21.12283,22.765602,21.980227,19.78529,20.838173,16.588915,8.388771,7.4696417,11.962401,12.655178,14.448852,17.778982,18.591793,29.68994,21.006224,16.180794,18.36544,10.220171,10.007536,11.286773,12.946692,14.085316,14.009865,11.118723,10.830637,14.085316,21.829325,35.029808,27.625326,31.977474,38.137012,39.96841,35.1567,31.655092,31.699677,33.126385,32.769707,26.462696,19.490345,17.717249,18.135658,18.732407,18.46147,16.592344,19.19197,22.11055,23.417223,23.389786,20.721567,21.187992,23.753323,26.7645,27.94085,30.982893,29.43272,27.131466,25.711617,24.61072,24.909094,24.60729,23.962528,23.52697,24.134007,23.976246,21.764162,20.893047,21.716148,21.513802,21.335464,22.978235,23.612709,22.223726,19.596663,19.987637,24.202599,25.752771,22.312897,15.700651,17.326277,17.237106,17.909306,19.263992,18.653526,16.273392,17.494326,18.02934,17.051908,17.20281,18.574646,17.497755,15.978448,14.596324,12.511135,12.349944,12.734058,11.406808,8.498518,6.5127864,6.0737996,6.1561093,6.3173003,6.464772,6.848886,7.058091,6.9552035,6.601956,5.909179,4.619654,4.7362604,6.6053853,7.421627,6.725421,6.385892,7.3358874,6.7048435,5.8405876,5.302142,4.835718,4.7671266,5.593657,6.4407654,6.7185616,6.0806584,6.869464,6.8145905,6.228131,5.6039457,5.6176643,5.1580997,5.003768,5.209543,5.576509,5.6656785,6.1732574,5.953764,5.3673043,4.8117113,4.6916757,4.125794,3.9303071,3.8034124,3.6044965,3.3369887,3.2409601,2.867135,2.7642474,2.9940298,3.1243541,2.8705647,2.7951138,2.6304936,2.2463799,1.6564908,1.5021594,1.3821237,1.2209331,1.1592005,1.5638919,1.4541451,1.2929544,1.1420527,1.0837497,1.2072148,1.0631721,1.1660597,1.471293,1.7936742,1.8142518,1.2826657,0.89512235,0.8025235,0.939707,1.0425946,0.7682276,0.6276145,0.65505123,0.805953,0.9842916,1.4335675,1.845118,1.9994495,1.8656956,1.605047,1.3341095,1.2175035,1.1694894,1.1729189,1.2860953,1.255229,1.3306799,1.4781522,1.5776103,1.4267083,1.1454822,1.1900668,1.3581166,1.4781522,1.4061309,1.6221949,1.6633499,1.646202,1.6187652,1.5810398,1.3375391,1.138623,1.0631721,1.039165,0.85739684,0.88826317,0.9534253,0.9534253,0.89855194,0.89512235,0.7613684,0.89512235,1.2620882,1.6427724,1.6290541,1.2449403,1.0631721,0.9945804,0.980862,0.9774324,0.9362774,1.1146159,1.3443983,1.4747226,1.3615463,1.3512574,1.3546871,1.4747226,1.5707511,1.2655178,0.9294182,0.78194594,0.7990939,0.89169276,0.89855194,0.9602845,0.94999576,1.039165,1.1214751,0.83338976,0.94999576,0.8471081,0.7682276,0.89855194,1.3546871,1.1489118,1.2003556,1.3752645,1.3409687,0.5796003,0.67219913,0.4698535,0.22635277,0.07545093,0.041155048,0.048014224,0.072021335,0.09259886,0.09259886,0.030866288,0.020577524,0.017147938,0.0274367,0.05144381,0.09945804,0.24350071,0.4629943,0.7510797,1.0734608,1.3992717,1.5913286,1.7593783,1.9308578,2.085189,2.1400626,2.4075704,2.603057,2.7711067,2.8945718,2.9082901,3.0386145,3.4433057,3.9543142,4.4104495,4.6436615,4.715683,4.664239,4.7431192,4.99005,5.24041,5.4907694,5.830299,6.138962,6.4544835,6.9689217,7.6857057,7.9189177,7.9463544,8.14527,9.012956,10.22703,12.97413,14.613472,14.417986,13.584596,12.22305,11.893809,12.133881,12.367092,11.88352,11.938394,12.061859,12.30193,12.538571,12.459691,12.277924,11.873232,11.008976,10.076128,10.076128,10.463672,9.993818,10.038403,10.882081,11.739478,10.906088,11.4376745,12.178465,12.977559,14.695783,12.596875,11.516555,11.499407,12.0309925,12.037852,12.380811,12.771784,14.057879,15.693792,15.728088,15.395418,15.666355,16.19794,16.407146,15.4742985,16.263103,16.414005,15.484588,14.164196,14.249936,14.973578,16.314548,17.2131,17.343424,17.096493,17.134218,15.8138275,14.706071,14.565458,15.313108,15.741806,18.313997,19.768143,19.53836,19.768143,19.010202,18.550638,19.058218,20.958208,24.4461,30.667372,31.377296,29.35384,27.18291,27.230925,3.07634,3.9028704,3.1895163,2.3389788,2.2806756,3.4638834,3.5564823,4.040054,4.016047,3.4227283,3.018037,2.4452958,1.5913286,1.2037852,1.4369972,1.8313997,1.6770682,1.4507155,1.1660597,0.980862,1.2072148,1.3272504,1.4815818,1.6290541,1.728512,1.7593783,2.1126258,2.1263442,2.201795,2.4418662,2.633923,3.0523329,3.5599117,3.882293,4.1360826,4.839148,4.90431,4.0606318,3.4981792,3.9303071,5.6073756,4.1772375,2.609916,1.3649758,0.64133286,0.34295875,0.37382504,0.41840968,0.548734,0.8093826,1.2037852,1.3649758,1.5433143,1.8519772,2.3218307,2.901431,2.7059445,2.201795,1.5604624,0.9877212,0.7305021,1.2072148,1.4095604,1.5158776,1.5810398,1.5090185,1.5570327,1.670209,1.8759843,2.1194851,2.277246,2.16064,1.903421,1.728512,1.8142518,2.287535,2.7711067,3.0797696,3.1209247,2.9151495,2.6064866,2.6236343,2.7642474,2.877424,2.8259802,2.486451,1.9754424,1.5330256,1.3889829,1.529596,1.6976458,2.1846473,2.7711067,3.1792276,3.2786856,3.083199,4.0023284,4.4756117,4.8837323,5.3330083,5.6656785,6.807731,7.1541195,6.917478,6.420188,6.094377,5.8474464,5.2918534,4.448175,3.508468,2.8122618,2.1572106,1.728512,1.4747226,1.3478279,1.2998136,1.1111864,1.0597426,0.89169276,0.6241849,0.53158605,0.6310441,0.6824879,0.7133542,0.70649505,0.59674823,0.5624523,0.66876954,0.7922347,0.85739684,0.8471081,0.6207553,0.53844523,0.490431,0.45613512,0.48357183,0.44927597,0.36353627,0.3566771,0.4629943,0.6173257,0.78537554,0.9568549,1.1626302,1.2723769,1.0014396,0.70649505,0.52815646,0.53501564,0.6893471,0.8505377,0.939707,0.939707,0.8505377,0.8128122,1.1180456,1.0631721,0.6893471,0.4046913,0.29494452,0.1371835,0.082310095,0.044584636,0.030866288,0.034295876,0.030866288,0.030866288,0.0274367,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.19891608,0.939707,2.2635276,4.715683,7.507367,9.661148,9.983529,11.461681,13.070158,14.682064,15.690363,14.997586,14.623761,16.2974,16.184223,14.273943,14.373401,14.225929,14.870691,17.086205,19.908754,20.61868,23.468666,23.091412,21.685282,20.35803,19.147387,17.826996,20.62554,26.160892,32.522778,37.293335,38.685745,37.526546,35.16699,32.82801,31.627655,30.732533,29.978024,30.7634,32.848587,34.35761,30.904013,27.004572,24.720467,24.480396,25.094292,23.067406,21.750444,20.738716,20.62554,23.005672,29.079472,45.72326,62.34304,71.46917,68.77351,62.367046,47.29058,29.854559,17.261114,17.607502,57.562195,35.489372,10.861504,5.1100855,1.5844694,0.7373613,0.64133286,0.6207553,0.4664239,0.44584638,0.4424168,0.5007198,0.8265306,1.2037852,0.97057325,1.8485477,3.1792276,3.9303071,4.040054,4.417309,2.9563043,6.7528577,11.132441,14.13333,16.499744,8.375052,5.4667625,6.5230756,9.246168,10.302481,12.874671,15.662926,15.789821,13.430264,11.825217,10.028113,13.474849,16.667795,17.61779,17.844143,15.971589,18.279701,22.175713,23.396646,15.999025,18.516342,17.689812,16.304258,15.340545,13.992717,13.073587,12.267634,11.8115,11.382801,10.096705,10.281903,13.437123,17.21996,23.681301,39.25163,25.142305,23.725885,25.629307,24.483826,16.925014,15.477728,16.21509,13.581166,7.939495,5.5833683,6.9552035,11.736049,15.539461,16.654078,16.060759,15.656067,16.585485,16.115631,14.510585,15.038741,18.862732,21.764162,22.378057,21.397196,21.582394,20.848463,19.137098,15.367981,10.518545,7.613684,12.061859,15.724659,16.513464,15.055889,14.7095,20.632399,19.305147,17.357141,15.782962,9.956093,14.870691,13.234778,9.97324,8.865483,12.545431,12.4802685,10.645439,13.704632,23.492674,37.00182,28.215216,32.948048,39.96498,41.453423,33.00635,29.981453,30.02604,30.626217,30.0912,27.532728,20.745575,17.847572,16.311117,15.470869,16.516893,17.021042,17.816708,18.749556,19.69955,20.563807,18.019053,20.889618,24.312346,26.147175,27.004572,29.33669,28.712505,27.76937,27.450418,26.983994,26.689049,26.404394,25.680752,24.795918,24.747904,24.055126,23.396646,22.556396,21.921923,22.470657,24.161444,25.306927,24.10314,21.095392,19.198832,20.176264,23.382927,24.343212,22.007662,18.742695,18.605513,18.499195,18.523201,18.04992,15.728088,12.905538,16.146498,18.389448,17.837284,17.991615,18.348293,16.945591,15.426285,14.30138,12.932974,12.308789,11.790922,10.628291,8.820899,7.1266828,6.8145905,6.958633,6.9963584,6.790583,6.6396813,7.085528,6.989499,5.9228973,4.65395,5.1409516,5.9297566,6.941485,7.0923867,6.574519,6.852316,7.706283,7.116394,6.217842,5.6519604,5.576509,5.5250654,6.1458206,7.116394,7.6514096,6.475061,7.1952744,6.9689217,6.2144127,5.545643,5.7822843,5.5387836,5.422178,5.576509,5.8543057,5.802862,6.101236,5.8200097,5.23698,4.650521,4.3624353,4.0503426,3.9680326,3.7279615,3.2958336,2.983741,3.07634,2.8122618,2.5241764,2.428148,2.644212,2.6236343,2.5447538,2.452155,2.2360911,1.6256244,1.5193073,1.4781522,1.3889829,1.3409687,1.6427724,1.4987297,1.3855534,1.2655178,1.1729189,1.2072148,1.1900668,1.5261664,1.6873571,1.5638919,1.4747226,1.2072148,1.0254467,0.9945804,1.0700313,1.0837497,0.96371406,0.9294182,0.9431366,1.0563129,1.4027013,1.8725548,1.9514352,1.7936742,1.5810398,1.5158776,1.4129901,1.3032433,1.2860953,1.3306799,1.2895249,1.430138,1.4781522,1.4610043,1.3924125,1.3032433,1.3169615,1.3238207,1.3478279,1.3958421,1.4678634,1.6290541,1.8073926,1.7490896,1.529596,1.5604624,1.2895249,1.1317638,1.0906088,1.0734608,0.90884066,0.90198153,0.84367853,0.78537554,0.7510797,0.72021335,0.78194594,0.9568549,1.1523414,1.2758065,1.2449403,1.1077567,1.0940384,1.1489118,1.196926,1.1283343,1.1763484,1.2175035,1.3581166,1.5124481,1.3786942,1.2483698,1.2895249,1.3615463,1.3512574,1.1626302,0.91227025,0.805953,0.8196714,0.8848336,0.89169276,0.9842916,1.0357354,1.0768905,1.0460242,0.77851635,0.7682276,0.7579388,0.6790583,0.66876954,1.0768905,0.9911508,0.9877212,1.1489118,1.2449403,0.7442205,0.881404,0.6824879,0.39097297,0.16462019,0.08573969,0.048014224,0.041155048,0.05144381,0.05144381,0.020577524,0.024007112,0.020577524,0.020577524,0.034295876,0.048014224,0.106317215,0.26064864,0.4972902,0.805953,1.1763484,1.313532,1.5364552,1.7833855,1.961724,1.9411465,2.1434922,2.277246,2.3835633,2.4624438,2.4898806,2.7162333,3.0351849,3.4398763,3.8788633,4.266407,4.396731,4.5030484,4.6848164,4.931747,5.1340923,5.3330083,5.552502,5.693115,5.7479887,5.830299,6.2658563,6.6739774,6.9963584,7.284444,7.7028537,8.615124,11.218181,13.522863,14.610043,14.651197,13.982429,13.392539,12.908967,12.593445,12.55229,12.63803,12.065289,11.746337,11.770344,11.413667,11.89038,11.688034,11.008976,10.367643,10.583707,11.303921,10.316199,9.513676,9.56512,9.904649,9.72631,10.199594,10.645439,11.22161,12.902108,11.818358,11.149589,11.201033,11.660598,11.605724,11.825217,12.092726,12.703192,13.21763,12.452832,11.732618,11.585147,11.712041,11.825217,11.616013,11.979549,12.6586075,12.723769,12.397959,13.063298,13.512574,14.3974085,14.88098,15.073037,16.03675,15.453721,14.96672,14.874121,15.12448,15.3302555,16.208231,18.056778,19.342873,20.28601,22.823904,25.20061,25.951689,25.591581,24.93996,25.097721,30.605639,35.26302,36.213013,33.68884,31.024048,4.822,3.6559403,2.2566686,1.5433143,1.8245405,2.8156912,2.2258022,2.311542,2.2498093,1.7182233,0.89512235,0.7613684,0.67219913,0.78537554,1.0734608,1.3169615,1.3786942,1.2346514,0.9294182,0.607037,0.53501564,0.72364295,0.94999576,1.2758065,1.6187652,1.7765263,2.2120838,2.2155135,2.1091962,2.1023371,2.3218307,2.551613,3.1826572,3.8857226,4.681387,5.9400454,5.751418,4.602506,3.8308492,4.108646,5.4153185,3.9543142,2.6236343,1.6221949,0.980862,0.5555932,0.64476246,0.7922347,1.1077567,1.546744,1.9102802,1.8279701,1.9891608,2.5996273,3.590778,4.616225,3.9611735,2.5790498,1.3101025,0.6379033,0.6859175,1.0906088,1.0768905,1.0460242,1.1660597,1.3546871,1.5158776,1.7319417,2.0680413,2.503599,2.935727,3.0866287,3.1312134,3.093488,3.0386145,3.100347,3.175798,3.2649672,3.0420442,2.5241764,2.0817597,2.0337453,1.9480057,1.9102802,1.9137098,1.845118,1.8965619,1.937717,2.0028791,2.1229146,2.3389788,2.8877127,3.5873485,4.1429415,4.290414,3.782835,3.8857226,3.5873485,3.4878905,3.7005248,3.8720043,5.0655007,5.5079174,5.4736214,5.4016004,5.888602,7.2947326,6.7871537,5.4324665,4.0537724,3.223812,2.411,1.7113642,1.2723769,1.08032,0.9774324,0.7922347,0.65505123,0.5624523,0.5041494,0.4698535,0.5761707,0.66191036,0.805953,0.922559,0.7510797,0.70306545,0.8128122,0.980862,1.1146159,1.1043272,0.84024894,0.6859175,0.61046654,0.5521636,0.4081209,0.37039545,0.3841138,0.42869842,0.5041494,0.6241849,0.8162418,1.2175035,1.6016173,1.6564908,0.96371406,0.6173257,0.6379033,0.8128122,0.9328478,0.7956643,1.0460242,1.2620882,1.4198492,1.5776103,1.879414,1.4644338,0.8505377,0.4081209,0.22635277,0.09945804,0.0548734,0.034295876,0.030866288,0.037725464,0.030866288,0.030866288,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12003556,0.764798,2.2223728,4.6882463,7.2604365,10.285333,12.915827,14.527733,14.71636,14.939283,16.414005,19.421753,22.662714,23.280039,24.957108,24.957108,23.149715,21.064526,21.904776,22.412354,24.456388,27.200058,28.808535,26.44212,27.254932,26.10945,25.087433,24.566135,23.221737,24.418663,26.02028,29.144634,32.924038,34.51537,37.543694,38.483402,37.49225,35.057243,31.970613,29.566473,28.396984,30.046616,33.376743,34.532516,30.701668,27.388685,25.711617,25.090862,23.238884,21.421204,20.35803,20.323736,21.637268,24.672453,32.210686,48.13426,63.828053,73.45148,73.95905,64.69574,45.867302,26.826233,14.757515,14.668345,26.987423,17.864721,7.5759587,3.6147852,0.70649505,0.34981793,0.39097297,0.5144381,0.548734,0.45613512,0.4938606,0.6824879,0.8162418,0.9842916,1.5501735,2.4590142,3.2615378,3.625074,3.6799474,4.0091877,2.6064866,4.029765,5.8371577,7.222711,9.002667,7.675417,8.947794,10.48082,11.622872,13.395968,16.431154,18.324286,17.943602,15.71437,13.6086035,9.678296,9.825768,12.185325,16.077906,22.017952,20.028791,23.931662,27.93399,28.372976,23.746464,23.242313,21.04052,20.255144,20.409475,17.429163,15.7795315,14.5585985,13.138749,11.413667,9.784613,10.768905,12.960411,16.232237,22.823904,37.365356,22.868488,22.484375,26.078583,25.632736,15.241087,13.581166,12.648318,9.421077,4.9934793,4.5682106,12.044711,15.271953,16.112202,16.146498,16.688372,13.903547,13.797231,14.177915,14.29452,14.860402,17.885298,21.081675,21.37319,19.288,18.982767,19.54522,16.760393,14.603184,13.341095,9.571979,11.399949,15.13134,15.525743,12.332796,10.2921915,12.641459,17.027903,17.775553,15.090185,15.069608,15.21022,11.739478,8.450503,7.953213,11.64345,18.221397,15.117621,14.918706,21.894485,32.015198,31.140654,35.90778,39.934116,38.73376,29.710516,29.18236,29.052036,29.717375,30.5199,29.779108,23.509823,19.936192,17.521763,15.844694,15.577187,14.894698,13.893259,13.817808,14.778092,15.734947,16.832415,19.473198,21.602972,22.998814,25.27263,27.6802,27.539587,27.824244,29.052036,29.285248,28.17406,27.313234,26.34609,25.553856,25.821363,25.066854,24.898806,23.821915,22.511812,23.818485,25.289778,24.957108,22.817045,20.262003,20.076805,21.369759,22.53582,21.832754,19.843594,19.476627,18.344864,17.905876,17.470318,16.650646,15.313108,12.771784,15.234227,17.71382,18.70497,20.169403,20.814167,19.03764,16.636929,14.743796,13.80066,13.155897,11.458252,9.949233,8.97523,7.9909387,7.64798,7.7714453,7.795452,7.5519514,7.2878733,7.0718093,6.56766,5.3741636,4.3692946,5.693115,6.6705475,6.941485,6.8763227,6.9380555,7.682276,7.589677,7.016936,6.492209,6.200694,5.970912,6.186976,6.680836,7.6376915,8.327039,7.099246,7.4970784,7.0546613,6.279575,5.7274113,5.98463,5.857735,5.7479887,5.8508763,6.0635104,5.960623,5.919468,5.5593615,5.0483527,4.523626,4.0949273,3.875434,3.6799474,3.3266997,2.9151495,2.8259802,2.9254382,2.784825,2.3835633,2.0131679,2.2806756,2.428148,2.3835633,2.352697,2.2806756,1.8416885,1.6633499,1.6393428,1.5913286,1.5158776,1.5810398,1.3889829,1.3478279,1.3101025,1.2312219,1.1900668,1.2860953,1.7388009,1.8073926,1.430138,1.2175035,1.2792361,1.3889829,1.471293,1.4061309,1.0460242,0.9568549,0.9877212,1.0906088,1.3169615,1.7936742,2.136633,1.9548649,1.605047,1.3478279,1.3581166,1.4061309,1.3375391,1.3032433,1.3272504,1.3306799,1.5741806,1.5741806,1.4438564,1.2929544,1.2106444,1.3786942,1.4164196,1.3684053,1.3786942,1.6804979,1.7971039,1.903421,1.762808,1.488441,1.546744,1.2723769,1.1523414,1.1214751,1.1180456,1.0940384,0.9294182,0.77851635,0.6756287,0.61046654,0.53158605,0.75450927,0.90884066,0.97400284,0.9568549,0.922559,0.8128122,0.91912943,1.1180456,1.2655178,1.196926,1.3375391,1.3341095,1.3821237,1.488441,1.4575747,1.2243627,1.2175035,1.2620882,1.2415106,1.1249046,0.8779744,0.7305021,0.71678376,0.77165717,0.7373613,0.86082643,0.90884066,0.91227025,0.88826317,0.8196714,0.6824879,0.7682276,0.7133542,0.5624523,0.77851635,0.84024894,0.7956643,0.922559,1.097468,0.78194594,0.8162418,0.7442205,0.5727411,0.36696586,0.28122616,0.14404267,0.061732575,0.024007112,0.01371835,0.01371835,0.0274367,0.024007112,0.024007112,0.030866288,0.024007112,0.0548734,0.14404267,0.29151493,0.5178677,0.8505377,1.039165,1.2998136,1.5810398,1.7730967,1.7079345,1.9102802,1.9925903,2.0440342,2.1194851,2.2155135,2.4144297,2.6304936,2.9288676,3.3198407,3.74168,3.899441,4.1635194,4.4447455,4.6779575,4.8151407,5.137522,5.2575574,5.2747054,5.23698,5.137522,5.1992545,5.689686,6.101236,6.276145,6.3961806,6.8969,8.618553,10.786053,12.740917,13.924125,14.438563,13.985858,13.107883,12.452832,12.80265,12.847235,12.161317,11.574858,11.321068,11.022695,11.640019,11.753197,11.297061,10.563129,10.206452,10.374502,9.589127,8.766026,8.309891,8.128122,8.711152,9.1810055,9.499957,9.798331,10.364213,10.604284,10.748327,10.933525,11.153018,11.269625,11.55428,11.667457,11.427385,10.796341,9.873782,9.273604,8.97523,8.834618,8.927217,9.544542,9.054111,9.626852,10.209882,10.556271,11.211322,12.370522,13.207341,13.54687,13.985858,15.87899,15.6697855,16.13278,16.897577,17.463459,17.189093,17.775553,18.241976,18.766703,19.871029,22.408924,26.10945,28.986874,29.954018,29.17893,28.105469,30.705097,35.49623,37.759758,36.33648,33.630535,4.170378,1.9171394,1.0768905,1.3306799,2.277246,3.4467354,2.1846473,1.903421,1.8965619,1.6290541,0.72707254,0.65505123,0.6927767,0.8128122,0.9294182,0.90541106,0.9602845,1.0460242,0.91569984,0.607037,0.44927597,0.35324752,0.39783216,0.64133286,1.0288762,1.3992717,1.7662375,1.7936742,1.8485477,2.1160555,2.5756202,2.335549,2.9940298,3.9886103,5.103226,6.4579134,6.252138,5.0586414,3.9611735,3.57363,4.0537724,3.2272418,2.6750782,2.2463799,1.8142518,1.2517995,1.4918705,1.845118,2.417859,2.9871707,3.0146074,2.9048605,3.3266997,4.0503426,4.9214582,5.844017,5.096367,3.199805,1.5021594,0.7133542,0.9259886,1.0666018,0.84367853,0.82996017,1.0597426,1.039165,1.155771,1.3786942,1.5947582,1.8519772,2.3767042,3.2375305,4.4104495,5.206114,5.1580997,4.0263357,3.2375305,3.0111778,2.6545007,2.054323,1.6359133,1.5981878,1.5364552,1.6804979,2.1160555,2.8054025,3.0797696,3.2786856,3.426158,3.5564823,3.724532,4.012617,3.9611735,3.9474552,4.0057583,3.8137012,3.1792276,2.6922262,2.510458,2.585909,2.668219,2.6853669,2.6579304,2.668219,3.1415021,4.8322887,7.6651278,7.222711,5.579939,4.0606318,3.2443898,2.6133456,1.8416885,1.2758065,0.980862,0.7579388,0.6207553,0.6241849,0.65505123,0.65505123,0.607037,0.65848076,0.7442205,0.9431366,1.1351935,0.9842916,0.90884066,0.91227025,1.0631721,1.2483698,1.1694894,0.922559,0.78537554,0.7305021,0.6893471,0.53844523,0.5727411,0.67219913,0.6790583,0.58302987,0.53844523,0.69963586,1.3341095,1.937717,2.0508933,1.255229,0.8711152,0.99801,1.1763484,1.1317638,0.78194594,1.6016173,2.0440342,2.3595562,2.5550427,2.4075704,1.4575747,0.7442205,0.33952916,0.18862732,0.12003556,0.10288762,0.08916927,0.10288762,0.12003556,0.0548734,0.034295876,0.024007112,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.3566771,1.9754424,4.187526,7.010077,11.146159,13.677195,15.927004,16.383139,15.532601,15.875561,15.110763,15.031882,19.071936,26.298077,31.418451,35.173847,32.03235,28.290667,27.320093,29.556185,31.140654,33.73685,35.115547,33.637394,28.235794,26.908543,26.298077,27.481285,29.467016,29.209797,30.804554,31.720255,32.766277,33.702557,33.242992,33.712845,34.542805,35.57854,35.58197,32.203827,27.51215,25.824793,28.420992,32.67025,32.049496,30.022608,26.496992,24.874798,24.627867,21.301168,19.881319,19.696121,19.637817,19.905325,21.980227,28.139765,35.540813,43.178505,49.667286,53.216908,46.88932,33.781437,20.186552,11.173596,10.590566,7.891481,5.1100855,3.018037,1.6324836,0.2194936,0.51100856,0.7476501,0.94999576,1.0357354,0.8162418,0.61389613,0.84367853,0.89169276,1.0357354,2.4487255,3.2581081,4.383013,4.770556,4.3452873,3.9851806,2.651071,2.6236343,3.8445675,6.060081,8.80718,10.786053,13.128461,14.030442,14.037301,16.023033,15.87213,17.7927,19.123379,18.313997,14.953001,11.609154,10.213311,11.005547,14.095605,19.473198,21.44521,28.215216,31.497332,30.286688,30.876575,28.643915,26.620459,26.846811,27.772799,24.27462,22.518671,19.805868,16.588915,13.310229,10.381361,9.990388,9.578837,11.245617,15.693792,22.258022,16.87357,19.243416,22.035099,21.160555,15.803539,15.971589,10.9198065,6.90033,5.768566,4.972902,17.432592,21.390337,20.591244,18.265984,17.141079,13.735497,13.327377,14.335675,15.566897,16.204802,15.385129,17.422304,18.8593,18.28313,16.328266,16.225378,14.445422,14.376831,15.261664,12.21619,9.942374,11.091286,12.836946,12.922686,9.688584,12.8197975,16.273392,17.995045,18.519772,20.965069,9.156999,8.944365,11.039842,11.866373,13.560589,21.729866,20.385468,18.259123,19.847023,25.426962,33.325302,37.845497,37.56427,33.397324,28.599329,30.430729,30.331272,31.92603,34.340458,32.19354,26.407824,23.581844,22.36434,21.057667,17.62808,11.650309,9.239308,9.822338,11.502836,11.084427,16.29397,16.19794,16.496315,18.975908,21.52066,26.232914,27.659622,28.10204,28.784527,29.875137,29.508171,28.01973,26.167753,25.073713,26.246634,25.910534,25.046278,24.044838,23.68473,25.125158,23.540688,21.808746,20.351171,19.87446,21.37319,22.165424,20.779871,18.358582,16.39,16.691803,17.343424,16.71238,16.002455,15.981877,17.000465,15.46744,15.247946,16.907866,20.255144,24.339783,25.711617,23.221737,19.312008,15.927004,14.493437,14.325387,12.147599,10.155008,9.211872,8.875772,8.443645,8.368194,8.375052,8.419638,8.687145,7.1129646,5.7308407,4.99005,5.055212,5.7891436,6.4990683,6.6396813,6.831738,7.377043,8.255017,7.3187394,7.006647,7.0306544,6.9552035,6.166398,6.5367937,7.016936,7.891481,8.577398,7.658269,7.7680154,7.2192817,6.492209,6.012067,6.1149545,5.970912,5.9126086,6.018926,6.2041235,6.23156,5.953764,5.4804807,5.0243454,4.633373,4.180667,3.8377085,3.3747141,2.959734,2.7916842,3.093488,2.9322972,2.7882545,2.4487255,2.07833,2.194936,2.3732746,2.4555845,2.4384367,2.3046827,2.037175,1.821111,1.7799559,1.7182233,1.5707511,1.4404267,1.2415106,1.2655178,1.2998136,1.2723769,1.2449403,1.3272504,1.646202,1.7765263,1.5981878,1.2929544,1.4267083,1.7113642,1.8485477,1.6599203,1.0906088,0.85739684,0.83681935,1.0666018,1.488441,1.9823016,2.1229146,1.9137098,1.5844694,1.2998136,1.1729189,1.2655178,1.2826657,1.2620882,1.2723769,1.4369972,1.6359133,1.5364552,1.3924125,1.2860953,1.1454822,1.2792361,1.4404267,1.4644338,1.471293,1.862266,1.9480057,1.8519772,1.6667795,1.5090185,1.5193073,1.2895249,1.138623,1.0597426,1.0494537,1.1146159,0.8093826,0.6756287,0.59674823,0.5178677,0.45613512,0.66876954,0.7613684,0.8162418,0.86082643,0.85396725,0.58988905,0.72364295,1.0048691,1.2106444,1.1180456,1.3272504,1.471293,1.5055889,1.471293,1.5158776,1.2517995,1.1420527,1.1249046,1.138623,1.1351935,0.8265306,0.5658819,0.53844523,0.65848076,0.5555932,0.6344737,0.58645946,0.59674823,0.72364295,0.91227025,0.7407909,0.8162418,0.77508676,0.58988905,0.5624523,0.7339317,0.66876954,0.78194594,0.97400284,0.6344737,0.5453044,0.64133286,0.65505123,0.5453044,0.4938606,0.29494452,0.14747226,0.061732575,0.024007112,0.01371835,0.0274367,0.030866288,0.030866288,0.024007112,0.017147938,0.05144381,0.082310095,0.1371835,0.26064864,0.52815646,0.8196714,1.0940384,1.3375391,1.5124481,1.5330256,1.7730967,1.8108221,1.821111,1.8897027,2.0097382,2.1434922,2.3218307,2.5756202,2.8808534,3.1689389,3.2889743,3.5942078,3.9200184,4.170378,4.2938433,4.729401,4.8288593,4.866585,4.938606,4.9523244,4.7088237,5.0620713,5.2506986,5.1066556,5.0346346,5.3981705,6.142391,7.4353456,9.187865,11.046701,12.620882,12.785502,12.312219,11.89038,12.120162,12.130451,12.034423,11.832077,11.629731,11.646879,11.979549,12.1921835,11.897239,11.008976,9.72631,8.625413,8.207003,7.9120584,7.56224,7.380472,8.2310095,8.868914,9.273604,9.304471,8.697433,9.561689,10.353925,10.751757,10.837497,11.115293,11.324498,11.204462,10.556271,9.56512,8.80718,8.711152,8.48137,8.31675,8.491658,9.362774,8.64942,8.608265,8.868914,9.211872,9.551401,11.616013,13.070158,13.924125,14.747226,16.660936,17.641798,18.28313,19.123379,19.963629,19.87446,19.44576,18.845583,18.478617,18.728977,19.949911,23.1943,27.491573,30.646793,31.751122,31.17838,31.898594,33.863747,35.407063,35.863197,35.527096,1.5707511,1.2312219,1.2723769,1.9514352,3.2546785,4.914599,2.8980014,2.037175,1.786815,1.6187652,1.0082988,0.89855194,0.9259886,1.1077567,1.3443983,1.4198492,1.2963841,1.2929544,1.2277923,1.0837497,1.0220171,0.5453044,0.29151493,0.28465575,0.48357183,0.77851635,1.0460242,1.371835,1.6804979,2.0646117,2.7470996,2.1743584,2.7333813,3.6147852,4.3349986,4.7602673,4.3692946,3.8685746,3.5770597,3.5770597,3.724532,3.7485392,4.0023284,4.0366244,3.6559403,2.8980014,3.5702004,4.0674906,4.4996185,4.6265135,3.8445675,3.6868064,5.0483527,5.597087,4.5270553,2.5481834,1.9754424,1.5021594,1.1592005,1.0460242,1.3272504,1.2037852,1.1660597,1.5810398,2.0063086,1.1763484,1.3101025,1.3341095,1.430138,1.6564908,1.937717,2.5241764,5.188966,7.8503256,8.615124,5.7822843,3.5118976,2.6716487,2.2669573,1.879414,1.6496316,1.6976458,1.6804979,1.9308578,2.7573884,4.4413157,4.2081037,3.590778,2.884283,2.527606,3.1140654,3.1380725,2.8225505,2.369845,1.9582944,1.7388009,1.8725548,1.7696671,1.6976458,1.704505,1.6187652,1.5673214,1.3821237,1.4129901,2.0714707,3.8308492,6.478491,6.4819202,4.8597255,2.8156912,1.7559488,1.8142518,1.371835,0.8848336,0.61046654,0.61046654,0.61046654,0.7922347,0.9328478,0.91227025,0.71678376,0.58302987,0.5761707,0.7476501,1.0357354,1.2655178,1.4267083,1.4267083,1.3306799,1.1797781,1.0220171,0.91227025,0.764798,0.6207553,0.5727411,0.7922347,1.0631721,0.97400284,0.8093826,0.7099246,0.6859175,0.9568549,1.5981878,2.0817597,2.061182,1.3889829,1.0357354,1.1111864,1.0940384,0.9534253,1.1592005,2.4795918,2.7162333,2.6716487,2.5653315,2.0303159,0.9911508,0.4389872,0.26750782,0.29151493,0.22978236,0.25378948,0.23321195,0.28122616,0.33609957,0.15090185,0.0548734,0.041155048,0.034295876,0.01371835,0.01371835,0.0034295875,0.0,0.01371835,0.041155048,0.09259886,1.786815,8.666568,13.334236,14.747226,18.187103,18.296848,16.78783,13.450842,10.213311,11.1393,8.831187,13.502286,20.954779,29.707087,41.000717,43.03789,38.404522,34.052376,33.119526,34.926918,34.693707,36.84406,37.471672,35.42421,32.286137,29.028028,27.18977,27.505291,28.818823,28.060884,26.52443,26.448978,27.865398,29.960876,31.082352,31.473324,32.056355,33.34245,33.963203,30.653652,27.213776,26.160892,29.120626,32.683968,28.410702,26.582733,23.36921,21.939072,22.144846,20.508932,19.86074,19.003344,17.055338,15.2033615,16.695232,20.845032,23.262892,25.622448,28.047167,29.144634,23.324625,18.231688,13.543441,10.652299,12.665466,5.0346346,2.1126258,1.2689474,0.89169276,0.36696586,1.3306799,1.5536032,1.5913286,1.5261664,0.9774324,0.53844523,0.5555932,0.5796003,0.83681935,2.2292318,3.2032347,5.381023,6.5779486,6.0223556,4.3624353,4.046913,3.2889743,4.7842746,7.658269,7.4765005,6.636252,7.449064,9.767465,11.931535,10.772334,11.530273,16.177364,21.163984,22.44665,15.501736,11.866373,11.423956,12.034423,12.977559,14.970149,20.045938,26.260351,29.281818,29.792826,33.476204,33.34245,32.24841,33.352737,35.43107,32.865738,29.803116,26.308365,21.390337,15.9613,12.847235,11.273054,8.224151,7.3701835,10.220171,16.12935,13.869251,15.117621,15.05246,13.227919,13.581166,21.112541,14.819247,10.669447,11.444533,6.742569,8.916927,17.936743,20.899906,17.117071,18.142517,14.932424,13.488567,12.867812,12.175035,10.590566,10.981539,13.649758,16.098484,17.20624,17.243965,15.083325,12.792361,13.049581,15.011304,14.328816,10.041832,9.575408,12.260776,14.692352,10.72775,17.744686,23.801336,23.547548,17.816708,13.642899,9.15014,17.034761,19.346302,15.772673,23.61957,18.945042,20.148827,20.86904,20.543228,24.415234,31.579641,35.112118,31.92603,26.586163,31.294985,31.380726,31.318993,32.92061,34.611397,31.449318,29.17893,30.029469,28.949148,25.512701,23.924803,14.404267,9.462232,9.47938,11.571428,9.582268,14.246507,14.4317045,15.573756,17.652086,15.199932,17.652086,26.85367,27.793377,21.304598,24.061985,31.068632,31.631084,28.414133,24.991404,25.831654,25.015411,23.667583,23.35549,24.19574,24.85765,20.155685,19.70641,19.325726,18.44432,20.080235,19.44576,16.348843,14.870691,15.522313,15.227368,16.667795,16.688372,15.848124,15.158776,16.098484,17.21996,16.523752,18.255693,23.060547,27.954567,28.27009,24.909094,20.063087,15.848124,14.29795,14.335675,12.175035,10.182446,9.338767,9.2153015,9.400499,9.105555,8.875772,8.89635,9.016385,6.2212715,4.928317,5.0620713,5.813151,5.6313825,6.6431108,6.8866115,6.6053853,6.509357,7.7680154,7.8263187,8.320179,8.453933,7.997798,7.2775846,7.1198235,7.4936485,8.285883,8.951223,8.498518,8.522525,7.7611566,6.917478,6.3721733,6.1629686,5.970912,6.121814,6.262427,6.341307,6.6225333,6.3035817,5.7754254,5.3570156,5.07236,4.6676683,4.57164,4.2252517,3.7382503,3.3644254,3.508468,2.9494452,2.568761,2.5138876,2.5721905,2.1812177,2.534465,2.935727,2.8945718,2.4418662,2.136633,1.9274281,1.7662375,1.6393428,1.5021594,1.2826657,1.1111864,1.1866373,1.3169615,1.4027013,1.4644338,1.4267083,1.3821237,1.5227368,1.7216529,1.5261664,1.3546871,1.5124481,1.6187652,1.5158776,1.2963841,1.1146159,1.0048691,1.1626302,1.5398848,1.845118,1.7730967,1.5981878,1.4335675,1.3066728,1.1592005,1.2826657,1.4404267,1.5433143,1.6084765,1.7559488,1.7799559,1.546744,1.3032433,1.1454822,1.0220171,1.255229,1.4027013,1.4541451,1.4575747,1.5570327,1.6907866,1.6599203,1.5638919,1.4575747,1.371835,1.2895249,1.2209331,1.0940384,0.89512235,0.6859175,0.5761707,0.5212973,0.4664239,0.41840968,0.4424168,0.5418748,0.5727411,0.58645946,0.58645946,0.548734,0.7442205,1.0117283,1.2586586,1.3478279,1.1283343,1.3478279,1.5055889,1.4678634,1.2963841,1.2346514,1.0906088,1.0151579,0.8711152,0.7339317,0.91569984,0.7339317,0.5761707,0.5693115,0.64133286,0.5178677,0.5693115,0.5796003,0.5727411,0.6207553,0.84024894,0.764798,0.7476501,0.78537554,0.7579388,0.42869842,0.59674823,0.4664239,0.44927597,0.5727411,0.48700142,0.42869842,0.42183927,0.39783216,0.36010668,0.39783216,0.33609957,0.26407823,0.16804978,0.06516216,0.01371835,0.0274367,0.041155048,0.034295876,0.017147938,0.030866288,0.041155048,0.0548734,0.08573969,0.15090185,0.26064864,0.5041494,0.7922347,1.0425946,1.2620882,1.5570327,1.8382589,1.9342873,1.8931323,1.8005334,1.8005334,1.9480057,2.1126258,2.3252604,2.568761,2.7779658,2.7539587,2.867135,3.1895163,3.6216443,3.8925817,4.0263357,4.3349986,4.6676683,4.880303,4.804852,4.5613513,4.4104495,4.3109913,4.2183924,4.057202,4.170378,4.4241676,4.7602673,5.2609873,6.166398,8.460793,9.719451,10.343636,10.64201,10.847785,10.957532,10.8958,11.122152,11.660598,12.099585,12.771784,12.782072,12.662037,12.421966,11.581717,10.323058,9.3764925,8.553391,7.939495,7.905199,8.501947,9.273604,9.462232,9.074688,8.879202,8.759167,9.047252,9.736599,10.504827,10.710602,10.539123,10.360784,10.172156,9.661148,8.210432,8.368194,8.213862,7.9943686,8.093826,9.033533,9.424506,9.026674,8.995808,9.626852,10.347065,10.991828,12.188754,13.701202,15.29596,16.722668,17.761833,18.176813,18.567787,19.054789,19.288,18.907316,17.916164,17.429163,18.44775,21.86705,25.053137,28.009441,31.391014,33.754,31.555634,31.312134,32.797146,34.889194,36.748028,37.811203,1.1454822,1.2998136,1.5193073,1.8416885,2.253239,2.702515,1.5604624,1.1489118,1.2758065,1.5707511,1.5090185,1.4164196,1.3101025,1.3169615,1.4164196,1.430138,1.5638919,1.5433143,1.3546871,1.0906088,0.9602845,0.58302987,0.32238123,0.22635277,0.29837412,0.47328308,0.70306545,0.980862,1.2517995,1.4850113,1.6599203,1.6804979,2.4144297,2.9563043,3.1860867,3.758828,5.7719955,6.5299344,6.831738,7.130112,7.517656,6.848886,6.1321025,5.363875,4.7499785,4.705394,7.3873315,8.790032,8.652849,7.181556,5.055212,3.3712845,3.8377085,3.99204,2.867135,0.9842916,0.6379033,0.84367853,0.99801,0.89512235,0.71678376,0.94656616,1.3032433,1.9171394,2.4795918,2.2258022,2.5721905,2.2841053,2.1297739,2.3252604,2.534465,2.8568463,3.8377085,5.096367,5.7891436,4.5853586,2.8156912,2.1263442,2.0063086,2.1983654,2.6990852,2.9220085,2.651071,2.5996273,2.8499873,2.867135,2.469303,2.1846473,2.0714707,2.1469216,2.3801336,2.1983654,1.8348293,1.5913286,1.5193073,1.3992717,1.4815818,1.4404267,1.3238207,1.1729189,1.0185875,0.97057325,0.9534253,1.4953002,2.867135,5.0620713,6.842027,6.461343,4.605936,2.4247184,1.5090185,1.2895249,1.1694894,0.9328478,0.6173257,0.548734,0.490431,0.5624523,0.6207553,0.61389613,0.59674823,0.48014224,0.4424168,0.48014224,0.58302987,0.71678376,0.7476501,0.764798,0.7510797,0.70649505,0.64476246,0.5624523,0.48357183,0.42869842,0.4629943,0.6824879,0.89512235,0.7305021,0.5555932,0.5727411,0.83338976,1.3272504,1.5810398,1.7696671,1.9651536,2.1332035,1.7319417,1.1729189,0.9534253,1.3684053,2.503599,3.6044965,3.7965534,3.192946,2.1503513,1.2723769,0.59674823,0.274367,0.17147937,0.23664154,0.4972902,1.039165,1.097468,1.1592005,1.2037852,0.6790583,0.19891608,0.20577525,0.28122616,0.24350071,0.12346515,0.11317638,0.08916927,0.106317215,0.15433143,0.16462019,3.7176728,12.151029,15.529172,12.662037,11.0981455,9.294182,6.0154963,5.874883,7.7783046,4.938606,7.3393173,15.100473,23.166862,29.158352,33.42133,36.943516,34.467354,33.33216,35.194427,36.024387,34.367897,33.26014,30.75997,27.875687,28.565035,26.994284,24.720467,23.434372,23.091412,21.884197,23.160004,25.670462,27.906553,29.425861,30.84914,32.481625,33.9975,34.230713,32.711407,29.67965,28.372976,29.731094,32.39931,33.65454,29.412142,24.291767,23.105131,23.825344,24.010542,20.814167,16.640358,13.591455,13.22106,15.097044,16.79126,20.755863,21.167414,21.517231,22.230585,20.673553,16.530611,14.201921,14.476289,17.816708,24.37065,8.567109,3.865145,2.8088322,1.6942163,0.5727411,0.77508676,0.77165717,0.8093826,0.8848336,0.7442205,0.607037,0.490431,0.40126175,0.548734,1.3238207,2.5070283,5.7582774,7.764586,6.9792104,3.6182148,4.650521,4.6265135,5.353586,7.7028537,11.602294,7.8503256,7.0375133,6.7974424,6.3790326,6.636252,9.325048,11.777204,15.323397,17.412016,11.609154,10.5597,12.109874,16.667795,21.86705,22.597551,24.442669,30.26611,36.09984,39.6769,40.42455,40.932125,40.277077,36.40164,31.367006,31.353289,31.66881,29.460155,25.955118,21.719578,16.643787,15.899568,13.262215,10.607714,10.261326,15.018164,27.896265,20.814167,12.593445,10.635151,10.9198065,17.933313,12.3533745,7.085528,6.262427,5.2438393,11.976119,16.811838,16.55119,13.231348,14.140189,12.850664,10.834066,9.9869585,10.268185,9.685155,10.446524,14.939283,16.259674,13.646329,12.483699,12.370522,11.094715,10.97468,12.000127,11.825217,10.381361,11.262765,11.849225,11.255906,10.323058,28.211786,23.657295,15.96816,12.751206,9.89436,9.921797,13.262215,23.334913,32.91718,24.158014,16.688372,18.578075,21.335464,21.839613,22.340332,29.611057,34.83089,34.51194,30.461596,29.792826,28.60962,29.85113,32.19354,33.66826,31.66881,30.128925,29.525318,27.707638,24.52841,21.839613,17.785841,13.570878,12.487128,14.102464,14.270514,15.388559,14.572317,15.086755,16.232237,13.317088,16.554619,26.205479,31.367006,30.365568,30.75311,25.20061,23.729315,25.296637,27.035439,24.233465,23.406935,22.642136,22.724447,22.312897,17.923023,18.02934,20.052797,20.426622,18.30028,15.553179,15.590904,16.918156,19.322296,21.44521,20.76958,18.900457,17.171944,16.489456,16.21852,14.181344,13.029003,15.285671,22.570116,33.047504,41.41913,33.122955,24.151155,18.550638,16.396858,13.773223,14.123041,12.668896,10.912948,9.89093,10.168727,10.2921915,10.131001,9.06097,7.641121,7.6274023,7.0958166,6.420188,6.3138704,6.3618846,5.007198,5.8543057,6.0154963,5.8165803,5.8165803,6.790583,6.9209075,7.6616983,8.114404,7.956643,7.4627824,7.1266828,7.507367,8.179566,8.738589,8.803751,8.505377,7.5759587,6.9380555,6.866034,6.9689217,6.334448,6.3035817,6.509357,6.742569,6.9654922,6.958633,6.5024977,6.135532,5.98463,5.768566,4.938606,4.2046742,3.5702004,3.1277838,3.059192,2.8877127,3.083199,3.0111778,2.6785078,2.719663,2.7882545,2.9288676,2.6819375,2.1503513,2.0028791,2.0577524,1.8519772,1.6942163,1.6016173,1.2929544,1.1832076,1.2860953,1.4335675,1.4953002,1.3924125,1.5501735,1.9411465,2.1023371,1.8588364,1.3306799,1.2860953,1.2415106,1.1523414,1.0597426,1.1146159,1.1077567,0.980862,1.0425946,1.3375391,1.6496316,1.5673214,1.529596,1.5570327,1.5947582,1.5261664,1.4335675,1.6496316,1.879414,1.9857311,1.9754424,1.9685832,1.7662375,1.5536032,1.3992717,1.2792361,1.3341095,1.2998136,1.3272504,1.3924125,1.3238207,1.6256244,1.6564908,1.5741806,1.5330256,1.6907866,1.1934965,1.155771,1.2106444,1.1523414,0.9568549,0.9534253,0.7407909,0.607037,0.6207553,0.6241849,0.59674823,0.66533995,0.65162164,0.5624523,0.58645946,0.9774324,1.097468,1.1832076,1.2689474,1.1660597,1.2963841,1.313532,1.2586586,1.1694894,1.0906088,0.90541106,0.8711152,0.8676856,0.805953,0.64819205,0.70649505,0.58988905,0.51100856,0.48700142,0.33609957,0.32581082,0.39783216,0.39440256,0.36696586,0.5590228,0.5624523,0.4972902,0.50757897,0.53844523,0.35324752,0.47671264,0.39097297,0.34295875,0.4081209,0.48700142,0.5727411,0.5590228,0.48700142,0.41498008,0.432128,0.33266997,0.26750782,0.23321195,0.18519773,0.041155048,0.024007112,0.0274367,0.030866288,0.024007112,0.017147938,0.020577524,0.037725464,0.058302987,0.08916927,0.15090185,0.4424168,0.65505123,0.89855194,1.196926,1.5193073,1.6530612,1.7216529,1.7525192,1.8039631,1.9582944,1.9102802,2.0268862,2.1846473,2.3561265,2.5927682,2.5584722,2.5378947,2.719663,3.0626216,3.292404,3.4467354,3.9063,4.40702,4.763697,4.856296,4.7088237,4.383013,4.0606318,3.8514268,3.789694,3.8891523,3.9611735,4.105216,4.3487167,4.6265135,5.4084597,6.166398,6.9380555,7.5245147,7.466212,7.7714453,8.388771,9.012956,9.784613,11.2593355,12.72034,12.644889,11.664027,10.604284,10.494537,10.381361,10.021255,9.561689,9.1810055,9.074688,9.595985,9.578837,9.462232,9.235879,8.453933,8.378482,8.477941,8.772884,9.194724,9.589127,9.448513,9.349055,9.249598,8.903209,7.829748,7.4044795,7.06838,7.0478024,7.3187394,7.6033955,8.06296,8.790032,9.72288,10.744898,11.688034,11.38623,11.499407,12.151029,13.341095,14.904987,16.53747,17.257685,17.110212,16.39,15.6252,15.316538,14.5585985,14.092175,14.774663,17.607502,22.638706,27.169191,30.605639,32.43361,32.23812,34.885765,36.00381,37.550552,39.594585,40.32509,1.0288762,1.1763484,1.1660597,1.3992717,1.8142518,1.8588364,1.3341095,1.3752645,1.587899,1.7147937,1.6427724,1.7696671,1.6221949,1.3752645,1.1900668,1.2037852,1.2620882,1.2517995,1.1317638,0.9294182,0.7442205,0.48700142,0.31895164,0.23321195,0.23664154,0.36010668,0.5007198,0.6790583,0.922559,1.1592005,1.2243627,1.4369972,2.2120838,2.7299516,2.952875,3.6387923,5.3501563,5.521636,5.5730796,6.1766872,7.2878733,5.9983487,5.0346346,4.7328305,5.120374,5.9434752,7.613684,8.200144,7.455923,5.597087,3.3129816,1.9411465,1.7971039,1.7079345,1.1660597,0.31895164,0.64133286,1.155771,1.4027013,1.3512574,1.3786942,1.8073926,1.5741806,1.4747226,1.7593783,2.1469216,2.901431,2.877424,2.6819375,2.633923,2.7402403,2.9665933,3.3541365,3.9783216,4.496189,4.149801,3.5564823,3.1140654,2.819121,2.7711067,3.2066643,3.2203827,2.7985435,2.5790498,2.5001693,1.8039631,1.6633499,1.862266,2.1263442,2.287535,2.2806756,1.879414,1.3821237,1.1111864,1.1077567,1.1214751,1.1866373,1.0906088,0.9877212,0.97057325,1.0631721,0.881404,1.3066728,2.9665933,5.254128,6.324159,5.4770513,4.664239,3.4981792,2.0817597,1.0185875,0.7922347,0.84367853,0.85396725,0.7510797,0.70649505,0.5178677,0.45613512,0.44584638,0.44927597,0.47328308,0.45956472,0.490431,0.53501564,0.5693115,0.607037,0.6207553,0.6344737,0.61046654,0.5555932,0.5041494,0.45956472,0.42526886,0.40126175,0.432128,0.6001778,0.66533995,0.6001778,0.5727411,0.66191036,0.86082643,1.1592005,1.2483698,1.546744,2.2223728,3.1792276,2.7573884,1.6530612,1.0425946,1.3855534,2.4452958,4.506478,4.931747,3.6696587,1.6839274,0.94656616,0.5658819,0.33952916,0.26407823,0.36010668,0.66533995,1.937717,2.0646117,1.8348293,1.9754424,3.1415021,1.728512,0.7613684,0.64476246,0.94999576,0.40126175,0.42526886,0.70649505,1.1763484,1.6804979,1.9514352,3.3815732,6.81802,7.81603,5.9400454,4.7534084,3.9303071,2.7162333,3.3129816,4.98662,4.064061,6.2144127,8.621983,11.825217,15.944152,20.69413,31.51105,29.573332,28.650774,31.490473,29.827122,28.108898,27.35096,25.745913,23.815056,24.43924,23.10856,22.655855,23.225166,24.11686,23.801336,25.001692,26.174612,27.885975,30.077482,32.09065,33.242992,35.863197,36.80633,35.407063,33.479633,31.415022,33.122955,35.75002,36.796043,34.120964,28.036877,26.164322,25.498983,23.76361,19.397747,15.193072,12.466551,11.835506,13.516005,17.319416,21.969936,22.930222,21.740154,19.37031,16.21166,11.447963,10.9198065,13.718349,17.748116,19.716698,8.073249,5.0586414,3.566771,1.2346514,0.432128,0.58302987,1.1077567,1.0425946,0.4698535,0.5212973,0.4698535,0.45613512,0.40126175,0.40126175,0.72364295,2.2258022,5.312431,7.675417,7.4765005,3.340418,4.262977,5.164959,6.252138,7.7542973,9.932085,7.466212,7.205563,7.016936,6.447624,6.7357097,9.0369625,10.508256,12.181894,13.495427,12.291641,10.593996,11.825217,16.561478,22.494663,24.442669,26.747353,30.235243,33.74714,39.279064,51.982258,56.95173,54.283512,44.433735,32.683968,29.154922,27.77966,26.93598,26.040857,24.140865,19.929333,18.108221,16.684942,16.695232,16.907866,13.786942,23.376068,22.77932,16.88386,10.80663,9.887501,27.697348,29.394995,20.28944,10.8958,16.942162,16.167076,14.421415,12.953552,12.291641,12.240198,13.361672,10.666017,8.988949,10.1652975,13.011855,10.30591,13.512574,13.807519,10.079557,8.930646,9.2153015,8.64256,8.793462,9.743458,10.072699,9.877212,11.684605,11.866373,10.587136,11.814929,22.096832,16.650646,13.440554,16.067617,13.780083,11.674315,12.017275,19.301718,26.894825,17.031332,19.308577,21.606401,22.395206,21.942501,22.340332,25.19718,29.809975,31.161232,28.523878,25.4544,28.897703,29.645353,29.923151,30.358707,29.974594,26.723345,24.44953,22.981665,21.626978,19.164536,16.084764,12.212761,11.286773,13.735497,16.678083,17.04162,16.780972,15.999025,13.88983,8.738589,13.917266,19.37031,24.843931,30.218096,35.520237,29.902573,26.219196,25.680752,26.260351,22.679861,21.925352,20.351171,19.672113,19.12681,15.4742985,16.438013,17.765263,17.477179,15.62863,14.308239,14.29795,16.016174,19.397747,22.991955,23.959099,22.131128,19.613811,16.925014,14.064738,10.487679,13.190193,25.128588,41.24765,52.664745,46.686974,28.92857,18.907316,16.12249,16.726099,13.533153,13.066729,12.3533745,11.303921,10.463672,11.008976,11.14273,10.2236,9.081548,8.385342,8.64256,8.31332,7.1952744,6.4407654,6.1321025,5.2815647,5.65539,5.425607,5.2266912,5.4667625,6.3173003,6.447624,7.301592,7.8537555,7.781734,7.442205,7.394191,8.038953,8.779744,9.153569,8.834618,8.484799,7.671987,7.2707253,7.394191,7.4010496,6.4133286,6.5470824,6.728851,6.6636887,6.8111606,7.1987042,6.8626046,6.3001523,5.8234396,5.521636,4.846007,4.383013,3.9097297,3.4433057,3.2546785,3.4535947,3.673088,3.3541365,2.750529,2.9185789,2.8088322,2.4898806,2.1983654,2.037175,1.978872,2.085189,1.9308578,1.670209,1.4335675,1.3169615,1.3203912,1.5193073,1.611906,1.5227368,1.3924125,1.4232788,1.670209,1.7490896,1.5433143,1.2175035,1.2037852,1.1660597,1.1111864,1.0871792,1.196926,1.2929544,1.1283343,1.0494537,1.1866373,1.4815818,1.5947582,1.7182233,1.728512,1.6427724,1.6187652,1.3821237,1.3992717,1.6564908,1.9823016,2.020027,2.037175,1.8588364,1.6427724,1.4335675,1.1763484,1.2346514,1.1317638,1.1866373,1.4164196,1.5330256,1.4129901,1.3341095,1.2895249,1.2723769,1.3032433,0.9534253,0.96371406,1.138623,1.2655178,1.1146159,1.0666018,0.823101,0.64476246,0.607037,0.607037,0.5761707,0.6276145,0.6276145,0.607037,0.7613684,1.039165,1.1180456,1.2037852,1.3169615,1.2929544,1.2792361,1.2449403,1.138623,0.9911508,0.9328478,0.7442205,0.7305021,0.84024894,0.91227025,0.6893471,0.78194594,0.6344737,0.5521636,0.58302987,0.52815646,0.30523327,0.30866286,0.29837412,0.2503599,0.36010668,0.37725464,0.36353627,0.39440256,0.41840968,0.28122616,0.33952916,0.30866286,0.28465575,0.3566771,0.58988905,0.7922347,0.764798,0.6310441,0.5007198,0.4698535,0.42526886,0.40126175,0.37725464,0.31895164,0.14747226,0.0548734,0.0274367,0.020577524,0.020577524,0.024007112,0.010288762,0.024007112,0.041155048,0.06859175,0.13032432,0.31895164,0.490431,0.6893471,0.9294182,1.2003556,1.4198492,1.5021594,1.5090185,1.5570327,1.8348293,1.7353712,1.862266,2.0577524,2.2223728,2.318401,2.6064866,2.5653315,2.5790498,2.7402403,2.8396983,3.0351849,3.3712845,3.858286,4.355576,4.5922174,4.7259717,4.461893,3.9646032,3.5118976,3.4776018,3.5290456,3.6216443,3.7931237,4.0263357,4.2046742,4.513337,4.7431192,5.055212,5.329579,5.147811,5.305572,5.562791,5.9571934,6.680836,8.052671,9.078118,9.6645775,9.6645775,9.355915,9.482809,9.534253,9.294182,8.968371,8.64942,8.30646,8.22758,8.080108,8.22758,8.536243,8.347616,8.601405,8.436785,8.354475,8.443645,8.3922,8.237869,8.14527,8.086967,7.9120584,7.3530354,6.461343,6.118384,6.427047,7.0958166,7.421627,7.9257765,8.783174,9.246168,9.3593445,9.928656,9.633711,9.613133,9.997248,10.960961,12.72034,14.774663,14.860402,14.592895,14.668345,14.856973,14.496866,14.157337,14.198492,15.079896,17.364002,22.666143,27.090311,30.42044,32.93776,35.403633,39.152172,41.669487,43.082478,43.603775,43.528324,1.039165,1.1934965,1.1043272,1.3032433,1.7182233,1.6633499,1.529596,1.6804979,1.8108221,1.8039631,1.7456601,2.0131679,1.937717,1.5844694,1.2003556,1.2003556,1.1146159,1.0425946,0.97400284,0.88826317,0.7682276,0.66533995,0.59331864,0.4629943,0.32238123,0.36010668,0.40126175,0.4698535,0.61389613,0.7990939,0.90198153,1.155771,1.7182233,2.0646117,2.2052248,2.702515,3.3644254,3.1072063,3.0660512,3.673088,4.650521,3.9886103,3.758828,4.5030484,5.8062916,6.310441,5.895461,5.284994,4.2766957,2.901431,1.4027013,0.7476501,0.45270553,0.32238123,0.23664154,0.16119061,0.69963586,1.2312219,1.5570327,1.7079345,1.9651536,2.1332035,1.5433143,1.1111864,1.2586586,1.9411465,2.5927682,2.8568463,2.9906003,3.1346428,3.3266997,3.532475,3.9131594,4.5956473,5.2987127,5.3090014,4.911169,4.3178506,3.7142432,3.3061223,3.3369887,3.4467354,3.216953,2.9220085,2.510458,1.5913286,1.7079345,2.061182,2.3252604,2.3389788,2.07833,1.6770682,1.2483698,1.0151579,1.0220171,1.138623,1.1008976,0.9328478,0.7922347,0.764798,0.8745448,0.8196714,1.8279701,3.9714622,6.0703697,5.6999745,3.8377085,2.976882,2.4795918,1.879414,0.89855194,0.59331864,0.6790583,0.8162418,0.8505377,0.7922347,0.5624523,0.4424168,0.40126175,0.4115505,0.45613512,0.6173257,0.7373613,0.864256,0.9534253,0.85739684,0.7305021,0.6379033,0.5658819,0.5212973,0.51100856,0.45956472,0.45613512,0.48700142,0.5624523,0.71678376,1.0014396,1.0494537,1.0082988,0.9774324,1.0117283,1.1832076,1.2826657,1.7079345,2.5961976,3.858286,3.3369887,1.9857311,1.1866373,1.4472859,2.4075704,4.945465,5.171818,3.5187566,1.3169615,0.7922347,0.6379033,0.53844523,0.58988905,0.7990939,1.0871792,2.3081124,2.369845,1.9171394,1.978872,3.9474552,3.590778,1.920569,1.1420527,1.3958421,0.7476501,0.8196714,1.3615463,2.1812177,2.952875,3.2135234,3.340418,3.6627994,3.9165888,3.7142432,2.527606,2.527606,2.3972816,2.5173173,3.0797696,4.1155047,4.8254294,5.435896,6.108095,8.165848,14.078457,25.19032,24.624437,23.890507,26.551867,28.198069,24.120289,20.803877,19.552078,20.61525,23.173723,21.70929,21.897917,23.03311,24.35007,25.046278,25.94483,25.248623,25.896814,28.417562,30.93145,33.551655,38.785206,41.99873,42.15306,41.799812,39.611736,40.56516,42.4823,43.024174,39.694046,33.57566,30.825132,27.968287,23.69159,18.852442,15.059319,12.603734,11.784062,13.474849,19.150816,22.813616,25.162884,23.238884,17.71039,12.871242,7.6342616,8.14527,10.840926,12.617453,10.837497,5.288424,3.789694,3.0283258,1.8348293,1.1660597,0.5693115,1.1214751,1.0871792,0.3841138,0.5761707,0.38754338,0.4664239,0.5007198,0.45613512,0.58988905,1.7353712,4.2081037,7.0752387,8.1487,3.9954693,3.865145,5.8405876,8.766026,10.875222,9.774324,6.5470824,6.584808,7.2878733,7.366754,6.8454566,9.194724,10.179015,10.655728,11.077567,11.499407,10.093276,10.762046,14.500296,19.37031,20.512363,22.480946,27.299517,31.528198,37.550552,53.577015,63.467945,64.802055,57.27068,44.430305,33.712845,26.785078,24.922812,25.138876,25.204039,23.633287,19.871029,18.03277,19.675543,21.349182,14.606613,17.758404,20.76958,18.180243,12.089295,12.164746,30.029469,37.931236,30.825132,18.132229,23.69845,18.21111,13.687484,11.550851,11.543991,11.746337,14.273943,10.7757635,9.606275,13.015285,17.161655,12.442543,12.250486,10.799771,7.5553813,7.2192817,7.7097125,7.1541195,7.016936,7.6925645,8.512236,9.006097,10.868362,12.267634,12.826657,13.615462,15.422854,14.081886,16.897577,22.165424,19.178253,21.150267,24.027689,26.040857,24.85422,17.53891,23.61957,23.516682,21.53781,20.817596,23.317764,22.748453,25.93111,27.378397,25.673891,23.482386,28.897703,27.85511,27.01486,28.026588,27.52587,24.236895,20.896477,19.404606,19.109661,16.815268,14.191633,11.825217,11.489118,13.491997,16.647217,18.811287,19.387459,18.04992,14.575747,8.834618,10.772334,12.30193,16.208231,22.758743,29.68994,29.881996,29.058895,27.625326,25.19375,20.598103,20.36832,18.718689,18.091074,18.063637,15.361122,14.856973,15.789821,16.026463,15.326826,15.333686,15.5085945,16.431154,18.862732,22.244305,24.68617,22.597551,19.11309,15.319967,12.751206,13.368532,26.160892,45.445465,59.61309,60.02121,41.007576,22.055677,13.406258,12.977559,15.734947,13.690913,13.488567,12.05843,11.084427,11.077567,11.399949,11.177026,10.237319,9.705732,9.630281,8.995808,8.848335,7.48336,6.5333643,6.351596,6.0326443,5.967482,5.768566,6.0497923,6.7048435,6.9037595,6.756287,7.250148,7.610255,7.596536,7.473071,7.658269,8.501947,9.277034,9.537683,9.126132,9.22216,8.680285,8.272165,8.172707,7.936065,6.8454566,6.883182,6.914048,6.6225333,6.5367937,7.099246,6.824879,6.1492505,5.501058,5.271276,4.9831905,4.6608095,4.2389703,3.8342788,3.7451096,4.0674906,4.184097,3.7725463,3.1072063,3.07634,2.7916842,2.311542,2.0646117,2.0680413,1.9480057,2.0680413,1.9651536,1.6804979,1.371835,1.3341095,1.3375391,1.5536032,1.5810398,1.430138,1.488441,1.4575747,1.430138,1.3752645,1.2895249,1.1763484,1.0837497,1.1214751,1.1660597,1.1729189,1.1489118,1.2380811,1.0700313,0.9259886,0.97400284,1.2689474,1.587899,1.728512,1.7319417,1.6633499,1.6221949,1.4232788,1.3409687,1.4438564,1.7216529,2.0577524,2.0303159,1.8245405,1.6187652,1.430138,1.1180456,1.1694894,1.1832076,1.3101025,1.5604624,1.8005334,1.3443983,1.214074,1.1626302,1.08032,0.99801,1.0048691,0.939707,0.9877212,1.138623,1.1626302,1.1077567,0.89512235,0.72021335,0.66191036,0.6927767,0.6276145,0.6962063,0.7956643,0.881404,0.96714365,1.1146159,1.1866373,1.2689474,1.3546871,1.371835,1.2209331,1.1694894,1.0117283,0.78537554,0.7579388,0.6824879,0.66533995,0.78537554,0.90198153,0.66533995,0.72021335,0.61046654,0.5555932,0.6001778,0.607037,0.3566771,0.31895164,0.29151493,0.24007112,0.28122616,0.28465575,0.30523327,0.34981793,0.3806842,0.31209245,0.31552204,0.29837412,0.28122616,0.32581082,0.4972902,0.6207553,0.6276145,0.5658819,0.490431,0.48700142,0.58988905,0.61389613,0.5727411,0.4664239,0.28122616,0.116605975,0.044584636,0.020577524,0.017147938,0.030866288,0.006859175,0.010288762,0.024007112,0.048014224,0.09945804,0.18176813,0.31895164,0.48357183,0.66191036,0.84367853,1.0837497,1.196926,1.2312219,1.3101025,1.6221949,1.6016173,1.7422304,1.9171394,2.0337453,2.037175,2.393852,2.3835633,2.3458378,2.4041407,2.4795918,2.760818,2.952875,3.2718265,3.690236,3.9474552,4.372724,4.3795834,3.9303071,3.3198407,3.175798,3.2066643,3.2649672,3.433017,3.7142432,4.0537724,4.2286816,4.15323,4.0434837,3.974892,3.8788633,3.99204,4.0606318,4.245829,4.6745276,5.446185,5.8645945,6.540223,7.082098,7.3427467,7.4181976,7.4181976,7.39762,7.373613,7.301592,7.06838,6.701414,6.4887795,6.660259,7.1541195,7.589677,7.8537555,7.716572,7.5931067,7.486789,6.9963584,6.708273,6.6225333,6.48535,6.279575,6.228131,5.768566,5.586798,5.9571934,6.6739774,7.0546613,7.5039372,8.045813,8.131552,7.870903,8.05953,8.021805,8.296172,8.694004,9.335337,10.624862,12.284782,12.401388,12.689473,13.649758,14.5585985,14.486577,14.764374,15.206791,15.9578705,17.497755,22.234016,26.538147,29.731094,32.334152,36.044964,41.06588,44.690956,46.364594,46.6321,47.16369,1.097468,1.3169615,1.3924125,1.5330256,1.6942163,1.5810398,1.6530612,1.6530612,1.6942163,1.8005334,1.920569,2.1503513,2.1503513,1.862266,1.488441,1.4781522,1.3512574,1.2003556,1.097468,1.0563129,1.0254467,1.0460242,1.0220171,0.8128122,0.5178677,0.4698535,0.41840968,0.37725464,0.36696586,0.4115505,0.5521636,0.7990939,1.0563129,1.138623,1.097468,1.2312219,1.2209331,1.3684053,1.7113642,2.0577524,2.0165975,2.668219,3.532475,4.914599,6.111525,5.435896,3.7142432,2.5721905,1.7765263,1.1694894,0.6893471,0.3806842,0.216064,0.15090185,0.16462019,0.24350071,0.53844523,0.90884066,1.3272504,1.6976458,1.8656956,1.5981878,1.3032433,1.2415106,1.4644338,1.821111,1.9823016,2.294394,2.8396983,3.4981792,3.9371665,4.2526884,4.846007,5.895461,6.992929,7.1266828,6.118384,5.164959,4.355576,3.799983,3.6079261,4.341858,4.4721823,4.0777793,3.2821152,2.2429502,2.3767042,2.4658735,2.3904223,2.1023371,1.6256244,1.4472859,1.3203912,1.2689474,1.2929544,1.371835,1.1694894,0.9431366,0.71678376,0.5178677,0.3841138,0.764798,2.2841053,3.9371665,4.7088237,3.57363,2.7128036,2.2566686,2.2395205,2.2669573,1.529596,0.7922347,0.7099246,0.8128122,0.84024894,0.72707254,0.5658819,0.47671264,0.4389872,0.45270553,0.53501564,0.83338976,0.97400284,1.155771,1.3101025,1.1180456,0.8128122,0.59674823,0.4972902,0.5007198,0.5590228,0.5624523,0.64476246,0.77508676,0.94656616,1.1626302,1.7730967,1.7971039,1.5810398,1.3821237,1.3649758,1.5947582,1.7593783,2.1194851,2.8122618,3.8514268,3.1860867,1.9720128,1.4061309,1.8931323,3.0454736,5.2644167,4.9248877,3.1312134,1.214074,0.7305021,0.6893471,0.75450927,0.9945804,1.3443983,1.5913286,2.085189,1.9994495,1.5227368,1.3169615,2.5138876,4.3521466,2.8568463,1.5090185,1.3889829,1.2106444,1.3443983,1.9308578,2.7162333,3.340418,3.333559,4.0194764,5.0003386,6.0635104,6.2555676,3.858286,3.3678548,2.386993,1.9925903,2.527606,3.590778,3.8925817,8.1212635,10.110424,10.117283,14.812388,19.185112,21.654415,21.956219,23.211449,31.92603,23.101702,15.909856,13.965281,17.367432,22.683292,21.897917,21.369759,21.551527,22.412354,23.44809,25.02227,23.77733,23.537258,25.526419,28.383266,33.390465,41.3231,47.29401,50.37035,53.587303,54.19091,54.22521,53.995426,51.838215,44.114784,37.64658,35.033237,31.078922,24.977686,20.316875,16.095055,13.039291,12.823228,15.954441,21.757303,21.829325,24.09971,22.196291,15.614912,9.72288,5.0003386,6.351596,7.514226,6.23156,4.2595477,2.1503513,1.0151579,2.6750782,5.4839106,4.307562,1.1866373,0.9945804,1.0906088,0.71678376,0.9842916,0.4664239,0.48014224,0.59674823,0.6790583,0.90541106,1.2998136,3.0043187,6.0635104,8.23444,5.020916,3.8445675,6.711703,11.348505,14.599753,12.428825,6.2692857,5.662249,6.701414,6.9723516,5.5559316,8.4264965,9.259886,9.400499,9.263316,8.320179,8.738589,9.331907,12.000127,15.302819,14.472859,14.5585985,22.549538,29.552755,34.302734,43.195656,54.966,66.060715,70.03903,63.893215,48.058807,33.359596,26.987423,25.351511,26.033998,27.807095,22.86163,19.078794,19.068506,20.560377,16.417435,17.099922,17.655516,16.657507,15.45715,18.169954,26.77136,36.792614,34.529087,22.930222,21.592682,17.147938,15.450292,13.066729,10.295622,11.156448,14.205351,10.48082,10.611144,16.077906,19.185112,15.9921665,12.517994,8.944365,6.3618846,6.776865,9.472521,8.364764,6.9620624,7.0546613,8.707723,9.283894,10.353925,13.173045,16.112202,14.651197,14.942713,18.763273,23.465237,26.215767,24.0174,40.626892,51.30663,46.944195,32.35473,26.301506,25.85223,22.61813,20.018501,20.131678,23.677872,23.749893,25.913963,26.19176,24.35693,23.94195,26.815945,24.761621,24.566135,26.558725,24.641586,23.52354,20.656404,18.763273,17.87501,15.343974,13.63604,13.344524,13.759505,14.496866,15.501736,20.303158,20.255144,18.331144,15.851553,12.4802685,8.3922,8.419638,10.302481,12.847235,15.947581,21.53095,27.254932,28.400414,24.43238,19.017063,18.883308,17.861292,17.998474,18.44432,15.433144,13.265644,15.21022,16.973028,17.117071,17.027903,17.881868,17.70696,18.149376,19.888178,22.624989,19.473198,15.405707,12.932974,14.695783,23.454948,45.706112,63.656574,65.313065,49.941654,28.081463,15.721229,10.093276,10.854645,14.291091,13.313659,14.568888,12.3911,11.235329,11.880091,11.423956,10.408798,10.422516,10.477389,9.836057,7.997798,9.3079,7.8126,6.807731,7.0889573,6.9552035,6.591667,6.9037595,8.004657,9.088407,8.423067,7.9086285,7.7542973,7.7440085,7.747438,7.7028537,8.011517,8.81404,9.493098,9.815479,9.928656,10.593996,10.39165,9.856634,9.242738,8.549961,7.6205435,7.298162,7.0889573,6.776865,6.4236174,6.7665763,6.468202,5.936616,5.5147767,5.4976287,5.521636,5.0174866,4.479041,4.245829,4.4859004,4.557922,4.513337,4.149801,3.5599117,3.1517909,2.784825,2.4761622,2.287535,2.1640697,1.9308578,2.020027,1.9137098,1.704505,1.471293,1.3066728,1.2346514,1.4027013,1.4164196,1.3203912,1.605047,1.5981878,1.430138,1.2929544,1.2312219,1.155771,0.9774324,1.039165,1.1351935,1.1249046,0.9431366,0.922559,0.7956643,0.72364295,0.8162418,1.1351935,1.4781522,1.471293,1.5364552,1.6839274,1.4815818,1.4369972,1.6496316,1.6221949,1.5021594,2.0749004,1.9445761,1.6770682,1.5261664,1.4644338,1.1832076,1.1797781,1.3409687,1.5090185,1.6359133,1.7971039,1.3924125,1.3203912,1.2312219,1.0563129,0.9911508,1.2483698,1.097468,0.9568549,0.980862,1.0597426,1.1111864,1.0220171,0.90884066,0.85739684,0.9328478,0.78194594,0.90198153,1.138623,1.2963841,1.1454822,1.255229,1.3478279,1.3889829,1.3752645,1.3409687,1.0940384,1.0082988,0.8505377,0.64133286,0.64819205,0.7407909,0.6962063,0.71678376,0.7613684,0.5418748,0.5555932,0.53501564,0.4972902,0.45956472,0.45613512,0.37382504,0.37382504,0.34981793,0.29494452,0.29837412,0.30523327,0.31209245,0.33952916,0.3806842,0.39783216,0.4081209,0.3806842,0.34981793,0.32238123,0.29151493,0.20920484,0.25378948,0.31209245,0.3566771,0.432128,0.6756287,0.7682276,0.7510797,0.64819205,0.45270553,0.23664154,0.10288762,0.037725464,0.020577524,0.030866288,0.010288762,0.0034295875,0.006859175,0.017147938,0.041155048,0.07545093,0.17147937,0.31552204,0.4698535,0.58302987,0.72364295,0.8676856,0.9842916,1.1283343,1.4061309,1.5090185,1.646202,1.7353712,1.7662375,1.7902447,1.903421,1.9068506,1.9308578,2.0268862,2.16064,2.49331,2.6476414,2.784825,2.959734,3.1312134,3.6593697,3.9714622,3.789694,3.2649672,2.9665933,2.9871707,2.935727,3.0146074,3.3026927,3.7622573,3.8274195,3.7348208,3.5221863,3.3198407,3.333559,3.549623,3.841138,4.0503426,4.180667,4.40702,4.5647807,4.6916757,4.8254294,4.931747,4.8837323,4.791134,5.079219,5.411889,5.638242,5.785714,5.6210938,5.295283,5.1992545,5.4839106,6.0532217,5.9880595,6.060081,6.15268,6.0737996,5.545643,5.0414934,4.9934793,4.787704,4.465323,4.7191124,5.219832,5.2609873,5.48734,5.9914894,6.3173003,6.677407,6.9346256,7.1198235,7.2158523,7.1678376,7.2878733,7.8777623,8.378482,8.683716,9.156999,9.877212,10.690024,11.753197,12.953552,13.906977,14.538021,15.436573,15.944152,16.101913,16.674654,20.183123,24.45296,27.60132,29.796255,33.26014,40.31823,45.356293,48.55953,50.438942,51.824497,1.2209331,1.1489118,1.2655178,1.4061309,1.4335675,1.2517995,1.4095604,1.4781522,1.6290541,1.8691251,2.0303159,2.1160555,1.9514352,1.7319417,1.611906,1.7079345,1.7216529,1.670209,1.5227368,1.3066728,1.097468,1.0494537,1.039165,0.90198153,0.7133542,0.7613684,0.6036074,0.45613512,0.34981793,0.33266997,0.4424168,0.6001778,0.88826317,1.1763484,1.3786942,1.4644338,1.4541451,2.2086544,3.0077481,3.275256,2.5790498,2.9460156,3.7794054,4.0880685,3.6285036,2.884283,2.3835633,2.1469216,1.8965619,1.5330256,1.1283343,0.66533995,0.36696586,0.26407823,0.31895164,0.42869842,0.9259886,1.0631721,1.2689474,1.4987297,1.2037852,1.1934965,1.4747226,1.845118,1.9445761,1.2346514,1.4438564,1.5776103,1.920569,2.4967396,3.083199,3.8377085,4.650521,5.6519604,6.601956,6.883182,6.478491,5.8371577,5.0757895,4.557922,4.914599,6.5367937,6.6053853,5.878313,4.7945633,3.4638834,3.3061223,3.0283258,2.4795918,1.786815,1.3581166,1.3821237,1.5707511,1.704505,1.6667795,1.4335675,1.1420527,0.85739684,0.6310441,0.4698535,0.33609957,1.1660597,2.819121,3.5633414,3.1106358,2.609916,2.2052248,2.335549,3.199805,4.029765,3.0660512,1.3341095,0.71678376,0.65162164,0.7133542,0.64133286,0.5178677,0.4972902,0.48014224,0.47328308,0.59674823,0.764798,0.78194594,0.805953,0.8471081,0.7613684,0.66533995,0.5590228,0.4972902,0.4972902,0.53501564,0.88826317,1.2415106,1.4850113,1.6770682,2.0303159,2.1023371,1.8005334,1.5810398,1.6187652,1.8142518,2.095478,2.1469216,2.2326615,2.5447538,3.2032347,2.5070283,1.786815,1.9137098,2.9734523,4.2423997,6.355026,5.967482,3.9097297,1.5604624,0.84024894,0.7407909,0.864256,1.138623,1.4198492,1.4815818,1.7593783,1.6942163,1.2620882,0.85396725,1.2826657,2.16064,1.704505,1.2037852,1.2963841,1.9685832,2.201795,2.633923,3.018037,3.234101,3.2958336,3.6970954,4.4413157,4.9831905,4.979761,4.273266,2.7093742,1.8245405,2.0028791,2.9940298,3.9200184,5.470192,10.436234,12.823228,12.284782,14.1299,17.439453,23.821915,24.744474,22.60098,30.732533,18.245405,15.570327,15.422854,14.908417,15.518884,17.545769,18.005335,19.987637,23.091412,23.420652,26.411253,26.26378,25.913963,27.10403,30.34842,32.91375,39.460835,46.72813,54.78423,67.01414,74.32602,74.18541,69.7681,61.327885,46.203403,37.975822,36.40507,33.52765,27.6802,23.468666,18.46147,14.867262,15.601193,19.87789,23.225166,17.754974,15.573756,14.016724,11.55428,7.781734,3.8034124,6.715132,7.517656,4.029765,0.91569984,0.8196714,0.5658819,5.9914894,13.831526,11.718901,3.5290456,2.5138876,2.5378947,1.5604624,1.6324836,0.65505123,0.39440256,0.5453044,0.9294182,1.4815818,2.07833,2.6476414,4.064061,5.5833683,4.835718,3.9954693,6.989499,9.606275,10.902658,13.200482,7.9257765,6.773435,6.5470824,5.693115,4.2869844,5.446185,6.8626046,6.8214493,5.90232,6.989499,7.7714453,8.165848,9.321619,11.406808,13.642899,13.2862215,17.024471,18.70497,20.19684,31.404732,38.349648,55.988014,73.173676,80.602165,70.80041,48.178844,34.09353,27.374968,26.905113,31.617367,28.465576,23.815056,19.901896,17.309128,14.953001,16.064188,19.435472,22.43979,24.494114,27.069735,41.9953,51.6976,42.530315,22.436361,20.934202,14.332246,18.4649,17.53891,9.925226,8.179566,12.586586,10.611144,9.829198,12.703192,16.585485,17.367432,14.184773,9.589127,6.0223556,5.813151,15.62863,14.033872,10.7586155,10.786053,14.373401,13.251926,13.190193,14.856973,16.578627,14.359683,18.104792,25.011982,26.43869,24.151155,30.303835,67.902405,87.1664,69.980736,33.318443,29.26467,21.647556,21.236006,22.847912,23.2869,21.345753,26.730206,29.292107,28.163773,24.552416,21.743584,22.391777,23.787619,23.873358,22.371199,20.7833,21.002794,21.20514,19.984205,17.394867,14.953001,12.562579,12.202472,13.810948,16.002455,16.0539,21.10568,16.7844,11.266195,8.868914,10.041832,8.296172,8.608265,8.786603,8.303031,8.31675,12.943263,20.882757,24.507832,22.642136,20.553518,17.940172,16.071047,15.539461,15.481158,13.564018,12.161317,15.217079,16.54776,15.553179,17.2131,18.787281,16.139639,14.352823,15.217079,17.243965,14.911846,12.871242,14.112752,20.673553,33.6614,50.922516,55.2095,48.30231,33.987213,18.080786,10.000677,9.637141,13.004995,15.206791,10.422516,12.339656,13.704632,13.985858,13.13189,11.581717,9.626852,10.412228,9.716022,7.3873315,7.3393173,11.941824,8.98209,6.5882373,7.2604365,7.857185,7.2124224,7.9292064,9.331907,10.460241,10.069269,9.705732,9.294182,9.023245,8.790032,8.179566,8.899779,9.400499,9.887501,10.48082,11.201033,11.592006,11.787492,11.47197,10.456812,8.697433,8.100685,7.720001,7.3290286,6.910619,6.667118,6.3378778,5.9812007,5.871454,5.950334,5.830299,6.0840883,5.4976287,4.98662,5.0483527,5.768566,5.144381,4.6127954,4.033195,3.3850029,2.760818,2.6887965,2.4590142,2.270387,2.1743584,2.0920484,1.8965619,1.728512,1.5981878,1.4541451,1.1592005,1.196926,1.4438564,1.529596,1.4472859,1.5570327,1.3238207,1.2380811,1.1832076,1.1214751,1.0837497,1.0117283,0.94656616,0.9568549,1.0048691,0.9294182,0.72364295,0.66191036,0.7888051,1.0734608,1.4027013,1.4164196,1.2003556,1.3169615,1.5398848,0.8711152,0.89512235,2.0268862,2.3801336,1.8073926,1.8931323,1.7319417,1.4644338,1.4164196,1.488441,1.1592005,1.1351935,1.1008976,1.1317638,1.2106444,1.2346514,1.2106444,1.1694894,1.0940384,1.0048691,0.9294182,1.039165,1.1592005,1.313532,1.3032433,0.71678376,0.9362774,1.2106444,1.2243627,1.0425946,1.1283343,0.9568549,1.08032,1.3306799,1.4850113,1.2655178,1.3752645,1.587899,1.6427724,1.4747226,1.2037852,0.89855194,0.7510797,0.6962063,0.70649505,0.7922347,0.91569984,0.7888051,0.65505123,0.6173257,0.64133286,0.6036074,0.5590228,0.45956472,0.34638834,0.33609957,0.31209245,0.36010668,0.39097297,0.37382504,0.33609957,0.4081209,0.41840968,0.38754338,0.34638834,0.33609957,0.48357183,0.5178677,0.51100856,0.48357183,0.4115505,0.3018037,0.22978236,0.18519773,0.17833854,0.21263443,0.39783216,0.6344737,0.82996017,0.89169276,0.7339317,0.48700142,0.24350071,0.08573969,0.030866288,0.030866288,0.030866288,0.020577524,0.010288762,0.0034295875,0.01371835,0.041155048,0.09259886,0.17833854,0.29151493,0.4115505,0.58302987,0.71678376,0.8025235,0.90541106,1.1763484,1.2963841,1.4095604,1.4644338,1.4850113,1.5707511,1.5947582,1.5090185,1.5844694,1.7936742,1.8313997,2.0268862,2.2498093,2.4212887,2.534465,2.6545007,2.8637056,3.1449318,3.2821152,3.199805,2.9288676,2.8945718,2.8465576,2.9220085,3.1277838,3.3712845,3.40901,3.4467354,3.3644254,3.1483612,2.867135,2.976882,3.1620796,3.4227283,3.7108135,3.9063,4.1155047,4.266407,4.2835546,4.197815,4.149801,3.5530527,3.6216443,3.7279615,3.7005248,3.8445675,3.8925817,3.7691166,3.8308492,4.1360826,4.4413157,4.2698364,4.1429415,4.249259,4.482471,4.4721823,3.8102717,3.8102717,3.8617156,3.789694,3.875434,4.3761535,4.4927597,4.8905916,5.645101,6.2555676,6.7459984,7.1129646,7.15069,6.852316,6.4236174,6.5813785,7.2638664,7.8537555,8.268735,8.927217,9.342196,9.949233,10.820349,12.037852,13.687484,15.127911,16.239098,16.62321,16.331696,15.868701,17.103354,19.94648,23.259462,26.606739,30.25925,39.364803,49.331184,57.126637,60.68655,58.930603,0.96371406,0.91227025,0.89512235,0.84024894,0.7956643,0.9328478,1.1523414,1.2826657,1.4815818,1.6942163,1.6873571,1.7353712,1.5638919,1.3855534,1.3512574,1.5261664,1.8897027,2.0063086,1.9514352,1.7559488,1.3924125,1.1660597,1.0734608,0.91227025,0.7373613,0.8848336,0.89169276,0.7099246,0.5007198,0.37039545,0.3806842,0.53158605,0.6962063,0.94656616,1.255229,1.5261664,1.3855534,1.7319417,2.0337453,2.1572106,2.3595562,3.4878905,3.5804894,3.1312134,2.5927682,2.3972816,2.2841053,2.2429502,2.1880767,2.0886188,1.9582944,1.7593783,1.3786942,1.0700313,0.94656616,0.9877212,1.3443983,1.6599203,1.7765263,1.7216529,1.7319417,1.5124481,1.728512,1.7182233,1.3443983,0.96714365,1.1454822,1.2723769,1.4472859,1.6942163,1.9480057,2.5961976,3.309552,4.280125,5.2026844,5.2575574,4.866585,4.0366244,3.3850029,3.3609958,4.2423997,5.8371577,7.9086285,8.471081,7.034084,4.5990767,3.4638834,2.4452958,1.7490896,1.3821237,1.1489118,1.371835,1.5193073,1.4644338,1.2483698,1.1043272,0.91912943,0.66876954,0.6207553,0.72707254,0.65162164,1.2277923,1.9548649,2.2669573,2.1126258,1.961724,2.4007113,2.9700227,3.625074,3.8342788,2.6167753,1.3203912,0.939707,0.85396725,0.7442205,0.59331864,0.5178677,0.51100856,0.5555932,0.65162164,0.8025235,0.7682276,0.72364295,0.7099246,0.7442205,0.83681935,0.6790583,0.6310441,0.7476501,0.9259886,0.9259886,1.4335675,2.07833,2.4761622,2.5996273,2.750529,2.6750782,2.2052248,1.7079345,1.7593783,3.1449318,3.7965534,3.5770597,3.1552205,2.7779658,2.2635276,1.6359133,1.3855534,1.9171394,3.1689389,4.5853586,6.3618846,5.2575574,3.1689389,1.4507155,0.8745448,1.0906088,1.0700313,1.1008976,1.3272504,1.7593783,1.8073926,1.6153357,1.2415106,0.9431366,1.1832076,1.6804979,1.7456601,1.9754424,2.5241764,3.0660512,2.4007113,2.3732746,2.6956558,3.175798,3.7348208,4.029765,4.0846386,4.0057583,3.8548563,3.673088,3.4878905,3.6868064,4.0606318,4.3007026,4.0057583,4.5990767,5.6656785,6.444195,7.6685576,11.55428,16.317978,25.488693,32.74913,35.93865,37.07727,34.443348,29.566473,24.154585,20.21399,20.069946,24.69303,26.905113,28.575323,29.741383,28.585611,28.547886,26.119738,26.016851,28.417562,28.969725,32.889744,39.666607,48.669277,61.722286,83.10233,99.74955,103.07282,96.889275,82.44728,58.409306,45.95304,37.197304,32.022057,28.60619,23.406935,18.79414,15.79325,15.110763,17.346853,23.01596,14.472859,10.628291,10.412228,10.861504,7.099246,3.2443898,3.525616,3.5461934,2.1126258,1.2449403,1.587899,0.9877212,5.535354,13.509145,15.391989,11.38966,7.346176,3.9165888,1.8828435,2.1332035,0.7956643,0.58988905,1.097468,1.7353712,1.7353712,2.5310357,2.6236343,3.457024,4.887162,5.178677,3.9851806,5.0174866,7.0306544,9.211872,11.183885,7.6788464,8.31332,8.796892,7.373613,4.835718,4.756838,5.9297566,6.7048435,6.866034,7.610255,8.556821,9.342196,10.357354,11.794352,13.615462,16.698662,22.072824,23.338343,21.208569,23.516682,29.868277,37.464813,47.225418,56.406425,58.5945,56.883137,46.690403,36.871494,32.557076,35.118977,32.625664,26.877676,25.581293,27.615038,23.022821,18.6158,22.789608,27.704208,29.782537,29.741383,40.805233,48.844185,44.14908,30.993181,27.635616,15.748666,16.527182,15.199932,8.742019,5.885172,13.776653,14.805529,14.404267,15.45715,18.28313,18.838724,14.832966,10.734609,10.179015,15.9578705,16.750105,12.329367,10.676306,13.015285,13.80066,14.140189,16.417435,16.599203,14.956431,16.0539,22.69358,25.303495,26.77822,29.374416,34.734863,61.62283,68.814674,53.096874,29.724234,32.42675,27.93399,26.538147,24.77191,22.213438,21.493225,24.61072,27.217207,25.876238,21.757303,20.62211,20.680412,21.678423,22.549538,22.52553,21.12283,23.852781,23.314335,22.000803,20.272291,16.345413,12.936404,13.282792,15.518884,17.343424,16.016174,16.510035,15.676644,13.361672,10.923236,11.235329,12.9981365,15.7966795,15.512024,11.485688,6.5470824,10.48082,15.830976,20.090523,21.383478,18.4649,17.62122,17.833855,16.602633,14.054449,12.919256,14.520873,16.849564,17.545769,16.732958,17.017612,17.144508,15.587475,14.376831,14.2533655,14.678635,13.989287,13.481709,16.890718,24.586712,33.551655,39.309933,39.99585,35.568253,25.965406,11.125582,5.885172,6.012067,9.373062,13.241637,14.315098,13.087306,12.88496,13.327377,13.032433,9.616563,8.659708,9.047252,9.280463,8.961512,8.81747,8.906639,7.654839,6.4579134,6.2212715,7.3564653,9.678296,8.656279,8.381912,9.884071,11.146159,10.583707,9.997248,9.606275,9.47595,9.5205345,9.880642,10.172156,10.419086,10.621432,10.786053,10.628291,11.348505,11.379372,10.261326,8.659708,7.956643,7.39762,7.1952744,7.205563,6.910619,6.23156,5.844017,5.7239814,5.686256,5.3878818,5.65539,5.693115,5.562791,5.4153185,5.4976287,4.8288593,4.262977,3.7176728,3.1483612,2.5550427,2.4795918,2.2806756,2.1263442,2.0989075,2.201795,2.1023371,1.6290541,1.2655178,1.1866373,1.2449403,1.3409687,1.5055889,1.5741806,1.5330256,1.5433143,1.430138,1.3512574,1.3786942,1.4232788,1.2312219,1.1866373,1.0494537,0.9774324,1.0151579,1.0768905,0.77165717,0.8848336,0.96714365,0.97057325,1.2209331,1.1249046,1.0425946,1.2415106,1.4918705,1.0666018,1.8313997,2.0886188,1.9480057,1.6873571,1.7319417,1.5741806,1.2758065,1.2483698,1.4027013,1.1592005,0.90198153,0.8093826,0.8093826,0.8779744,1.0288762,1.0528834,1.2792361,1.4095604,1.371835,1.3101025,1.2826657,0.9945804,0.84367853,0.82996017,0.5453044,0.65848076,0.8128122,0.7990939,0.6790583,0.7613684,0.83681935,0.89512235,1.1249046,1.4267083,1.3992717,1.5193073,1.7182233,1.6770682,1.3992717,1.2312219,0.9259886,0.84024894,0.8265306,0.7682276,0.61046654,0.6241849,0.64819205,0.64133286,0.6001778,0.5693115,0.4629943,0.45956472,0.4389872,0.39440256,0.42183927,0.42526886,0.5178677,0.5144381,0.4046913,0.34638834,0.39097297,0.3806842,0.37725464,0.38754338,0.33609957,0.4046913,0.50757897,0.5727411,0.5624523,0.51100856,0.4081209,0.32238123,0.26750782,0.23321195,0.20234565,0.22978236,0.39783216,0.64819205,0.86082643,0.8676856,0.7407909,0.5453044,0.3018037,0.082310095,0.041155048,0.024007112,0.024007112,0.020577524,0.01371835,0.01371835,0.030866288,0.041155048,0.08573969,0.15433143,0.216064,0.3566771,0.5658819,0.7579388,0.89512235,0.980862,1.0528834,1.0871792,1.097468,1.1420527,1.3169615,1.5536032,1.728512,1.879414,1.9823016,1.9411465,1.8931323,1.99602,2.1812177,2.3801336,2.5207467,2.5721905,2.702515,2.8980014,3.069481,3.0626216,2.976882,3.0660512,3.1792276,3.2272418,3.175798,3.1826572,3.2855449,3.2821152,3.1312134,2.9665933,2.9494452,2.959734,3.0351849,3.1243541,3.1243541,3.3026927,3.5873485,3.7279615,3.649081,3.4433057,3.069481,3.0489032,3.0454736,2.9700227,2.9906003,3.3438478,3.2203827,3.1963756,3.3781435,3.391862,3.1037767,2.983741,3.083199,3.2958336,3.3609958,2.8294096,2.5893385,2.5927682,2.7368107,2.8637056,3.4604537,3.6525106,3.9371665,4.465323,5.0346346,5.5833683,6.0086374,6.090947,5.8234396,5.435896,5.2438393,5.394741,5.7274113,6.125243,6.509357,7.1781263,7.671987,8.848335,10.871792,13.224489,14.781522,16.221949,17.147938,17.545769,17.785841,18.588364,20.11796,21.976797,23.650434,24.497543,29.785967,43.950165,64.26018,85.37615,99.33114,0.59674823,0.6379033,0.6036074,0.5693115,0.6001778,0.7613684,0.864256,0.90198153,1.0288762,1.2758065,1.5570327,1.6016173,1.3306799,1.1043272,1.1523414,1.5536032,1.9239986,2.1194851,2.201795,2.1400626,1.7936742,1.4164196,1.0837497,0.85396725,0.77851635,0.90541106,1.0220171,0.9362774,0.7579388,0.5796003,0.4938606,0.6344737,0.7682276,0.90884066,1.1008976,1.430138,1.670209,1.8382589,1.9651536,2.1229146,2.4418662,3.5393343,3.5153272,2.9665933,2.5310357,2.8877127,3.1243541,2.767677,2.435007,2.369845,2.4795918,2.5996273,2.8019729,2.8534167,2.7230926,2.5927682,2.9322972,2.9220085,2.527606,2.0234566,1.9994495,1.9068506,1.9514352,1.862266,1.5810398,1.2586586,1.039165,1.1489118,1.2998136,1.3821237,1.471293,1.7696671,2.054323,2.5756202,3.2375305,3.5873485,3.8205605,3.0351849,2.411,2.527606,3.340418,5.703404,8.920357,10.353925,9.047252,5.7068334,3.865145,2.3732746,1.3821237,0.91569984,0.88826317,1.1866373,1.371835,1.313532,1.1317638,1.214074,1.1077567,0.89512235,0.764798,0.823101,1.1077567,1.8245405,2.0508933,2.0406046,2.0028791,2.1126258,2.5310357,2.6853669,2.6956558,2.5927682,2.3389788,1.2620882,0.75450927,0.64133286,0.8025235,1.1763484,0.89512235,0.77851635,0.75450927,0.764798,0.7613684,0.6344737,0.6207553,0.7407909,0.881404,0.78194594,0.6036074,0.6241849,0.91227025,1.3478279,1.5981878,2.1263442,2.726522,3.083199,3.1277838,3.0111778,2.6750782,2.2806756,2.177788,2.5310357,3.3129816,4.2046742,4.0674906,3.4398763,2.6373527,1.7353712,1.3375391,1.4267083,2.054323,3.0214665,3.8720043,4.530485,3.590778,2.3801336,1.5776103,1.2243627,1.2449403,1.2106444,1.214074,1.430138,2.1160555,2.3081124,2.3561265,2.369845,2.486451,2.8705647,2.8122618,2.7745364,3.117495,3.6182148,3.4776018,2.784825,2.6236343,3.1209247,4.0366244,4.7328305,4.3795834,4.5510626,4.6436615,4.434457,4.1017866,4.232111,4.0057583,3.8308492,3.7519686,3.4604537,4.0194764,4.0263357,4.0949273,5.0174866,7.7714453,11.622872,19.70641,28.043737,34.148403,37.046402,35.211575,30.561054,29.00402,31.58993,34.51194,36.878353,34.878906,31.898594,29.34012,26.627317,25.927681,23.924803,27.251501,33.157253,29.51503,34.367897,38.431957,45.407738,59.325005,84.55648,108.40583,119.57256,114.70255,95.78495,70.16936,54.85282,41.875263,34.0901,29.813404,22.813616,18.399736,15.594335,13.951562,14.692352,20.683842,12.288212,10.549411,11.317638,10.871792,5.9400454,2.301253,2.3252604,2.7128036,1.99602,0.548734,0.86082643,0.8471081,4.681387,12.079007,18.307138,14.181344,10.81006,6.5985265,2.5001693,2.0097382,0.83338976,0.5796003,0.9294182,1.5158776,1.937717,3.0729103,2.7162333,3.1140654,4.479041,5.0003386,4.338428,5.885172,7.6857057,9.0644,10.635151,9.585697,9.616563,9.14328,7.795452,6.4407654,8.690575,7.3598948,6.0703697,6.2487082,7.1266828,8.275595,10.034973,12.072148,13.992717,15.3302555,18.584934,25.999702,29.936869,28.26666,24.336353,30.399864,31.284697,34.64226,41.110466,44.32742,53.182613,52.80536,46.65268,39.24477,36.16157,32.15238,26.150604,25.1183,28.520449,28.33525,20.886189,21.321745,24.60729,27.11089,26.582733,37.125286,49.986237,51.529552,40.921837,30.135784,17.652086,15.285671,12.651748,7.3873315,5.144381,16.47231,17.881868,16.012743,14.987297,16.400288,15.906426,13.694343,11.941824,11.993267,14.356253,11.718901,11.523414,12.003556,11.914387,10.535692,10.64201,12.017275,12.651748,13.54687,18.71183,20.889618,22.134558,24.422092,29.59391,39.385384,50.342915,45.099075,33.802013,25.835083,29.813404,25.426962,22.007662,20.639257,22.186,27.316664,27.786518,27.18634,24.78563,21.061096,17.665806,17.778982,18.276272,19.980776,21.969936,21.61326,22.089973,21.20171,21.249723,21.28059,17.04848,14.640909,16.304258,18.080786,17.580065,13.975569,13.906977,15.563468,15.6252,13.670336,12.157887,14.435134,17.95046,17.981327,13.615462,7.7680154,10.511685,13.790371,16.438013,17.470318,16.105343,16.098484,16.53404,16.163645,14.695783,12.775213,14.435134,16.96617,16.431154,13.262215,12.260776,13.516005,15.470869,15.6697855,13.814379,11.766914,11.122152,12.555719,17.446312,24.43238,29.439579,30.821703,29.494452,24.298628,15.721229,5.90575,3.3987212,4.15323,7.1884155,10.906088,13.101024,11.269625,11.595435,12.21619,11.489118,7.98065,8.210432,9.633711,10.659158,10.367643,8.525954,6.8900414,6.8557453,7.4524937,7.881192,7.5245147,8.56025,9.122703,9.335337,10.110424,13.1421795,11.478829,10.535692,10.618003,11.043272,10.168727,9.97667,10.209882,10.460241,10.542552,10.515115,10.494537,10.9198065,11.019264,10.412228,9.091836,8.110974,7.459353,7.1095347,6.910619,6.5985265,6.1801167,5.754848,5.6656785,5.8234396,5.6999745,5.7068334,5.8337283,5.8200097,5.56965,5.164959,4.5990767,4.0503426,3.5153272,3.0489032,2.7402403,2.469303,2.0749004,1.8519772,1.8759843,1.9994495,1.8588364,1.6564908,1.4472859,1.313532,1.3581166,1.4027013,1.5433143,1.5261664,1.4404267,1.7147937,1.4918705,1.5124481,1.5536032,1.4918705,1.3032433,1.4335675,1.3272504,1.2998136,1.4541451,1.6633499,1.1797781,1.5124481,1.5810398,1.2758065,1.4507155,0.75450927,0.9602845,1.4095604,1.5570327,0.94999576,2.633923,2.4075704,1.8313997,1.529596,1.2003556,1.2380811,1.0151579,0.99801,1.1934965,1.1420527,0.7579388,0.67219913,0.64133286,0.65505123,0.94999576,0.90541106,0.90198153,1.1283343,1.3684053,1.039165,0.91912943,0.6173257,0.47671264,0.4938606,0.32924038,0.45956472,0.5761707,0.607037,0.5761707,0.58988905,0.8128122,0.8745448,1.0563129,1.313532,1.2895249,1.3066728,1.4267083,1.3958421,1.2243627,1.1729189,0.8505377,0.7099246,0.69963586,0.7305021,0.66533995,0.6241849,0.607037,0.59331864,0.58302987,0.58645946,0.4698535,0.4389872,0.4355576,0.4355576,0.4424168,0.41840968,0.45270553,0.48014224,0.45270553,0.34295875,0.37725464,0.37725464,0.36353627,0.34981793,0.32581082,0.39097297,0.52815646,0.69963586,0.823101,0.7442205,0.6310441,0.47328308,0.3566771,0.30523327,0.26407823,0.18519773,0.2503599,0.39440256,0.5555932,0.67219913,0.70649505,0.7510797,0.58988905,0.26750782,0.09945804,0.0548734,0.034295876,0.024007112,0.01371835,0.006859175,0.010288762,0.017147938,0.041155048,0.08573969,0.15090185,0.23321195,0.37382504,0.548734,0.71678376,0.8128122,0.8505377,0.823101,0.8471081,0.97057325,1.1592005,1.4027013,1.6084765,1.7250825,1.7799559,1.8862731,1.7833855,1.7593783,1.8656956,2.054323,2.194936,2.411,2.469303,2.5481834,2.7059445,2.867135,2.9185789,2.9460156,3.0077481,3.0969174,3.1380725,3.2683969,3.316411,3.2546785,3.1655092,3.2375305,3.0489032,2.9185789,2.843128,2.8019729,2.7470996,2.8499873,2.9322972,2.9117198,2.7951138,2.6613598,2.6647894,2.7916842,2.8088322,2.6579304,2.4487255,2.7642474,2.6647894,2.5173173,2.486451,2.5413244,2.2978237,2.0749004,2.0817597,2.2600982,2.287535,1.879414,1.7593783,1.937717,2.2806756,2.5070283,2.9391565,3.0420442,3.192946,3.525616,3.923448,4.2595477,4.5201964,4.715683,4.8425775,4.866585,4.602506,4.5990767,4.856296,5.2918534,5.7479887,6.64997,7.7577267,9.349055,11.406808,13.612033,14.685493,15.446862,15.861842,16.307688,17.576635,20.03222,21.527521,22.247734,22.330044,21.884197,25.18689,34.899483,51.574135,73.92476,98.8167,0.52472687,0.5144381,0.47671264,0.4698535,0.52472687,0.67219913,0.66533995,0.7407909,0.89855194,1.1420527,1.4472859,1.4129901,1.1146159,0.9431366,1.1111864,1.6393428,2.020027,2.270387,2.417859,2.411,2.1057668,1.5364552,1.0597426,0.823101,0.84367853,1.0288762,1.2517995,1.2517995,1.08032,0.8505377,0.72707254,0.91912943,1.0528834,1.1351935,1.2998136,1.8039631,2.3595562,2.5481834,2.702515,2.9220085,3.093488,3.99204,4.0023284,3.5530527,3.2306714,3.7725463,3.7313912,3.216953,2.8808534,2.9185789,3.093488,3.590778,4.6093655,5.223262,5.103226,4.5030484,5.15467,4.3692946,3.0146074,1.8965619,1.786815,1.8965619,1.8485477,1.7936742,1.7353712,1.5193073,1.3375391,1.4095604,1.4164196,1.3101025,1.313532,1.4472859,1.5227368,1.6804979,2.0131679,2.551613,3.292404,2.5619018,1.9857311,2.2738166,3.2203827,5.6313825,9.050681,10.840926,9.705732,5.6828265,3.5050385,2.6853669,1.9514352,1.0357354,0.6756287,0.9328478,1.0940384,1.0288762,0.8779744,1.0425946,0.97400284,0.89855194,0.83681935,0.8848336,1.1934965,1.7936742,1.8313997,1.6907866,1.6633499,1.9480057,2.5996273,2.4967396,2.054323,1.7216529,1.9480057,1.0734608,0.51100856,0.40126175,0.71678376,1.2483698,0.96371406,0.8128122,0.7579388,0.7579388,0.78194594,0.84367853,0.84024894,0.8505377,0.823101,0.5624523,0.432128,0.6241849,1.1351935,1.762808,2.1194851,2.311542,2.7368107,3.07634,3.1552205,2.9391565,2.386993,2.0303159,2.2429502,2.8705647,3.234101,3.7759757,3.6044965,3.1689389,2.7402403,2.4144297,2.2498093,2.294394,2.7333813,3.5153272,4.341858,4.0949273,3.0214665,2.2463799,2.0268862,1.7422304,1.4575747,1.3889829,1.4987297,1.8588364,2.651071,3.1380725,3.1037767,2.8980014,2.7642474,2.877424,2.6545007,2.5447538,2.7882545,3.1483612,2.9117198,2.6785078,2.7162333,3.1346428,3.74168,4.0674906,3.8720043,4.40359,4.791134,4.629943,4.0229063,4.0880685,3.666229,3.4055803,3.391862,3.1312134,3.6868064,3.6456516,3.6079261,4.012617,5.1512403,7.2947326,12.984418,20.172834,27.611609,34.865185,35.25959,32.24155,33.16754,38.24333,40.56173,40.023285,36.470234,32.25184,28.883986,27.066305,26.569014,25.51956,29.621347,35.42764,30.33813,35.190998,36.281605,39.306503,49.821617,73.23541,94.91726,114.17097,116.5511,99.77356,73.72927,58.94432,46.930473,38.857227,32.85888,24.010542,19.823015,17.322845,15.011304,14.4145565,20.080235,11.71547,10.206452,10.422516,9.174147,5.192395,1.7525192,2.294394,3.4433057,3.1655092,0.77508676,0.4389872,0.53844523,5.662249,14.376831,19.239986,14.891269,14.061309,9.767465,2.8054025,1.7662375,0.805953,0.5624523,0.7682276,1.155771,1.4850113,3.0626216,2.8294096,3.0900583,4.2115335,4.6436615,5.206114,8.694004,9.517105,7.881192,9.788043,10.213311,9.568549,8.608265,7.8126,7.3839016,9.410788,6.9346256,4.90431,5.212973,6.711703,8.368194,9.791472,11.650309,13.660047,14.55174,15.158776,20.78673,25.375517,26.34952,24.617579,30.242102,28.76052,30.375856,36.861206,41.57346,52.45554,57.69252,54.37611,45.112793,38.027267,33.877464,27.76594,24.987974,26.613598,29.463587,25.27263,23.28347,24.77534,28.27352,29.542467,38.126724,52.21547,59.328434,54.19091,38.723473,24.161444,16.756964,11.612583,7.4284863,6.495639,18.95533,19.092514,16.187653,14.784951,14.685493,13.622321,14.490007,16.482597,16.918156,11.2250395,11.283342,12.456262,12.329367,10.827208,10.199594,9.499957,9.55826,10.412228,12.370522,15.999025,16.479168,18.173384,21.849901,29.76539,45.661526,40.088448,30.269539,25.495554,26.582733,25.859089,21.726437,18.139088,18.37916,22.61127,27.896265,28.307816,25.821363,24.202599,23.475527,19.936192,17.933313,16.942162,17.665806,19.421753,20.135109,18.725548,18.44432,19.603521,20.28258,16.355703,15.889278,18.152807,18.835295,17.04162,15.278812,15.1862135,16.177364,16.736387,16.098484,14.249936,15.656067,17.96761,17.017612,12.579727,8.375052,9.716022,12.590015,14.675205,15.090185,14.417986,14.767803,14.774663,14.839825,14.490007,12.360233,13.570878,15.313108,14.126471,10.563129,9.167287,11.094715,14.081886,14.942713,13.176475,10.960961,9.187865,10.854645,14.956431,19.53836,21.688711,22.083115,20.148827,14.959861,8.344186,4.8734436,3.0797696,3.5153272,5.3741636,7.723431,9.506817,8.375052,9.139851,10.065839,9.650859,6.625963,7.846896,10.007536,11.149589,10.30934,7.507367,5.785714,7.3839016,9.554831,10.254466,8.158989,8.097256,9.510246,9.860064,9.705732,12.71691,11.043272,10.419086,11.1393,11.897239,9.80862,9.770895,10.199594,10.185875,9.746887,9.832627,10.158438,10.182446,10.251037,10.113853,8.920357,7.966932,7.514226,7.164408,6.7528577,6.3653145,6.159539,5.7377,5.672538,5.9812007,6.1286726,6.0703697,6.0737996,5.953764,5.576509,4.863155,4.2423997,3.6113555,3.1037767,2.8156912,2.8328393,2.726522,2.3081124,1.9068506,1.7182233,1.8108221,1.7833855,1.7730967,1.704505,1.6187652,1.6564908,1.6359133,1.7456601,1.7250825,1.6393428,1.8725548,1.961724,1.978872,1.9102802,1.7662375,1.5776103,1.8313997,1.6770682,1.646202,1.8691251,2.07833,1.6290541,2.061182,2.054323,1.5433143,1.704505,0.99801,1.0254467,1.6359133,2.1674993,1.4369972,4.0434837,2.819121,1.5570327,1.3958421,0.8265306,0.89169276,0.77165717,0.7956643,0.96714365,0.9568549,0.64476246,0.65505123,0.58645946,0.45613512,0.69963586,0.6001778,0.490431,0.70649505,1.0254467,0.65848076,0.66191036,0.4355576,0.32581082,0.36010668,0.2503599,0.3566771,0.42869842,0.47671264,0.5144381,0.5761707,0.7407909,0.83338976,0.9842916,1.1454822,1.097468,1.2106444,1.2346514,1.1146159,0.94999576,0.97057325,0.75450927,0.6241849,0.6036074,0.66191036,0.72707254,0.72021335,0.61046654,0.548734,0.5658819,0.5693115,0.5521636,0.5212973,0.48357183,0.44927597,0.4424168,0.39783216,0.3806842,0.41498008,0.45270553,0.35324752,0.3806842,0.37382504,0.34981793,0.33266997,0.34981793,0.41498008,0.5212973,0.69963586,0.8676856,0.85396725,0.8196714,0.6859175,0.5212973,0.39097297,0.35324752,0.21263443,0.1920569,0.22292319,0.28808534,0.4081209,0.53158605,0.7476501,0.7339317,0.45956472,0.20577525,0.09602845,0.044584636,0.0274367,0.017147938,0.006859175,0.006859175,0.010288762,0.024007112,0.05144381,0.09945804,0.15433143,0.22292319,0.33952916,0.5007198,0.65848076,0.7133542,0.7099246,0.7613684,0.8779744,0.9842916,1.2037852,1.3821237,1.5055889,1.6084765,1.786815,1.7216529,1.6290541,1.6633499,1.8245405,1.9685832,2.2360911,2.3046827,2.3629858,2.49331,2.6853669,2.7230926,2.7162333,2.7470996,2.843128,2.952875,3.1312134,3.0969174,2.976882,2.9082901,3.0351849,2.8499873,2.7230926,2.651071,2.5927682,2.4967396,2.5070283,2.4144297,2.277246,2.1846473,2.2292318,2.3732746,2.4624438,2.4590142,2.3218307,2.0131679,2.1572106,2.0920484,1.9445761,1.8485477,1.961724,1.8691251,1.6873571,1.6564908,1.762808,1.7353712,1.5844694,1.6016173,1.7833855,2.0508933,2.253239,2.411,2.428148,2.5173173,2.7230926,2.9288676,3.1552205,3.3884325,3.6765177,4.040054,4.4584637,4.6676683,5.0003386,5.4839106,5.9812007,6.2075534,6.7700057,7.8263187,9.575408,12.082437,15.282242,15.88242,15.453721,14.908417,14.980438,16.242527,19.243416,21.500084,22.60441,22.69358,22.456938,24.837072,30.403294,40.5,56.20065,78.32835,0.7339317,0.6207553,0.5761707,0.5178677,0.48014224,0.6207553,0.59674823,0.823101,1.0837497,1.2483698,1.2620882,1.1351935,0.9602845,0.9911508,1.2963841,1.7662375,2.194936,2.4658735,2.5721905,2.4761622,2.1126258,1.4918705,1.0700313,0.85396725,0.881404,1.2072148,1.5124481,1.5193073,1.3238207,1.08032,1.0048691,1.2449403,1.371835,1.4850113,1.7319417,2.311542,2.8945718,3.2032347,3.4947495,3.8479972,4.184097,5.137522,5.079219,4.6265135,4.297273,4.530485,3.875434,3.625074,3.7451096,4.064061,4.2869844,5.48734,7.473071,8.450503,7.8503256,6.324159,6.9723516,5.2987127,3.0317552,1.4610043,1.4438564,1.6496316,1.7182233,1.8073926,1.9068506,1.8279701,2.095478,2.085189,1.8485477,1.546744,1.4404267,1.5158776,1.5947582,1.6290541,1.7422304,2.2360911,3.0729103,2.4590142,1.9720128,2.3664153,3.566771,5.346727,8.196714,9.757176,8.64599,4.4584637,2.5207467,3.1072063,3.1449318,1.8279701,0.6310441,0.7613684,0.84367853,0.72707254,0.5178677,0.58302987,0.6173257,0.70306545,0.8128122,0.89855194,0.90884066,1.1729189,1.2449403,1.1626302,1.1283343,1.4987297,2.527606,2.4761622,2.0028791,1.5776103,1.4815818,0.8779744,0.51100856,0.42183927,0.5624523,0.7613684,0.7682276,0.6859175,0.6893471,0.8196714,1.0117283,1.3066728,1.2689474,0.9911508,0.6241849,0.36696586,0.42183927,0.90198153,1.6564908,2.3389788,2.4075704,2.1194851,2.3972816,2.7539587,2.8808534,2.644212,1.9857311,1.6667795,1.9651536,2.7333813,3.4192986,3.4124396,3.0420442,2.9734523,3.3952916,4.029765,3.9714622,3.8137012,4.15666,5.0586414,6.060081,5.3878818,3.858286,2.8568463,2.603057,2.1674993,1.7696671,1.8485477,2.3629858,3.216953,4.2698364,5.0243454,4.5853586,3.4673128,2.2258022,1.4541451,1.4027013,1.5536032,1.9754424,2.5070283,2.7573884,2.6750782,2.726522,2.6545007,2.4624438,2.4144297,3.1106358,3.8891523,4.3521466,4.266407,3.5599117,3.3609958,3.2272418,3.433017,3.7382503,3.3781435,3.724532,3.7759757,3.82399,4.0263357,4.3795834,5.813151,10.456812,16.640358,23.647005,31.699677,34.896053,33.50364,33.987213,36.74117,36.09641,33.291004,31.730543,30.818274,30.5199,31.32928,30.85257,30.691378,32.365017,34.035225,30.475315,33.284145,33.42476,33.232704,37.437378,53.162037,65.71776,90.2736,103.25459,94.72178,68.358536,56.252094,48.689854,43.185364,37.07727,27.532728,23.581844,21.03709,18.139088,16.317978,20.186552,12.919256,9.335337,7.8537555,7.0546613,5.689686,2.218943,4.2835546,5.950334,5.0140567,3.0043187,1.0185875,1.1111864,9.15014,20.124819,18.149376,15.018164,15.484588,11.063849,2.8808534,1.6839274,0.9259886,0.77508676,0.94999576,1.0734608,0.65848076,2.503599,2.7779658,3.1243541,3.8548563,3.9543142,5.4770513,10.271614,9.966381,5.744559,8.330468,8.652849,8.299602,7.970361,7.750868,7.1129646,5.8543057,4.32128,3.6525106,4.434457,6.691125,8.954653,9.609704,10.511685,11.893809,12.380811,9.613133,9.97324,12.154458,15.505165,20.011642,26.335802,25.337791,28.499872,37.67059,45.06478,53.052288,57.85028,54.849392,45.833008,38.97726,36.195866,30.34499,25.828222,24.747904,26.911972,29.333261,28.410702,30.701668,36.477093,39.72148,43.50432,55.137478,67.91612,72.16538,55.236935,34.395332,21.462358,13.63261,9.410788,8.625413,19.709839,18.581505,16.414005,16.763824,15.594335,14.284232,18.060207,22.546108,22.330044,10.981539,14.832966,13.461131,11.540562,11.2593355,12.315649,12.271064,12.367092,12.168177,11.406808,10.007536,12.668896,16.969599,22.43979,31.034336,47.13625,33.09895,27.457277,27.817385,28.818823,22.144846,20.587814,18.972477,20.045938,22.666143,21.819035,24.36036,23.238884,23.598991,25.872808,25.76992,22.000803,17.899017,15.649208,15.944152,17.95389,16.45516,17.003895,18.025911,17.830425,14.586036,15.46058,17.158226,17.20281,16.37285,18.69811,17.984756,16.732958,16.80155,17.576635,15.971589,16.70552,16.979887,14.280802,9.657719,7.716572,7.8023114,11.252477,14.112752,14.623761,13.234778,13.605173,13.21763,12.9638405,12.792361,11.688034,12.566009,12.332796,11.334786,10.079557,9.235879,10.357354,11.331357,11.849225,12.085866,12.696333,10.155008,9.945804,10.971251,12.199042,12.648318,13.248496,11.650309,8.529384,6.0052075,7.6445503,4.835718,3.8891523,3.875434,4.417309,5.65539,5.686256,6.23156,7.682276,8.652849,6.0086374,7.301592,9.427936,10.271614,9.242738,7.2535777,6.0806584,9.006097,11.667457,11.760056,9.0369625,9.6645775,10.340206,9.908078,9.016385,10.127572,9.760606,9.863494,10.909517,11.64345,9.081548,9.431366,10.2921915,9.757176,8.299602,8.772884,9.431366,9.194724,9.235879,9.47938,8.615124,7.922347,7.7371492,7.4936485,6.999788,6.464772,6.3138704,6.001778,5.9469047,6.2041235,6.4544835,6.540223,6.368744,5.9743414,5.3570156,4.496189,3.758828,3.1037767,2.7059445,2.6236343,2.784825,3.0283258,2.7813954,2.2566686,1.7902447,1.8519772,2.037175,1.9514352,1.8828435,1.9548649,2.1229146,2.0337453,2.0474637,2.0646117,2.054323,2.0337453,2.5584722,2.486451,2.3218307,2.2360911,2.0646117,2.2498093,1.9823016,1.8588364,2.0097382,2.0817597,1.9685832,2.4247184,2.2395205,1.6290541,2.218943,1.9308578,1.488441,2.0131679,3.0248961,2.435007,5.693115,3.2992632,1.3101025,1.3752645,0.7613684,0.7442205,0.67219913,0.6790583,0.7373613,0.65162164,0.5761707,0.77851635,0.66191036,0.28808534,0.39097297,0.28808534,0.2709374,0.4081209,0.5761707,0.4355576,0.6962063,0.5144381,0.36353627,0.37382504,0.31552204,0.31552204,0.32924038,0.36010668,0.4389872,0.6310441,0.66191036,0.7407909,0.90198153,1.0528834,0.9842916,1.2758065,1.2312219,0.97057325,0.7099246,0.7579388,0.71678376,0.6790583,0.64476246,0.64133286,0.7305021,0.764798,0.6241849,0.5521636,0.58645946,0.5453044,0.64819205,0.66191036,0.59331864,0.5007198,0.51100856,0.4424168,0.40126175,0.40126175,0.42526886,0.4081209,0.41840968,0.38754338,0.37039545,0.39097297,0.432128,0.4629943,0.5007198,0.5727411,0.6824879,0.7922347,0.8848336,0.8711152,0.70649505,0.47671264,0.4046913,0.25378948,0.19548649,0.17833854,0.18519773,0.22978236,0.33609957,0.5727411,0.6790583,0.5727411,0.34295875,0.14061308,0.06516216,0.048014224,0.044584636,0.024007112,0.020577524,0.01371835,0.020577524,0.034295876,0.041155048,0.09602845,0.1371835,0.19891608,0.30866286,0.48700142,0.59674823,0.6859175,0.7510797,0.77851635,0.7613684,0.980862,1.138623,1.3272504,1.5330256,1.6256244,1.6599203,1.5981878,1.6153357,1.7525192,1.920569,2.0749004,2.1915064,2.3046827,2.428148,2.568761,2.486451,2.527606,2.5619018,2.5653315,2.6167753,2.6922262,2.6236343,2.5138876,2.435007,2.428148,2.369845,2.3424082,2.3424082,2.3321195,2.2155135,2.201795,2.136633,2.0680413,2.0680413,2.2223728,2.2155135,2.0440342,1.9308578,1.8759843,1.6599203,1.6633499,1.6427724,1.6084765,1.5981878,1.6839274,1.6907866,1.670209,1.6804979,1.7113642,1.6770682,1.7971039,1.8588364,1.8691251,1.8588364,1.8828435,1.8588364,1.8656956,1.9857311,2.1812177,2.3081124,2.5207467,2.8294096,3.1209247,3.450165,4.0263357,4.8288593,5.586798,6.310441,6.790583,6.601956,6.619104,7.0272245,8.879202,12.713481,18.54378,19.336014,17.278261,15.237658,14.373401,14.160767,15.9613,19.023922,21.753874,23.592133,25.049707,27.254932,32.097507,39.200184,48.55267,60.52536,0.8093826,0.91912943,0.9362774,0.8162418,0.6310441,0.59674823,0.6310441,0.805953,0.939707,0.980862,0.9911508,1.0048691,1.097468,1.3684053,1.7559488,2.061182,2.3046827,2.4487255,2.435007,2.1846473,1.587899,1.4644338,1.2312219,0.939707,0.7922347,1.1592005,1.4027013,1.3443983,1.2243627,1.1763484,1.2346514,1.3101025,1.4095604,1.587899,1.7490896,1.6633499,2.0920484,2.4727325,2.9494452,3.7451096,5.171818,6.660259,6.40304,5.693115,5.1512403,4.698535,4.2595477,4.57164,5.212973,5.9228973,6.6053853,9.39021,12.751206,13.440554,11.046701,7.9943686,6.848886,4.7842746,2.6990852,1.4541451,1.9068506,1.9685832,2.469303,2.9871707,3.2066643,2.9151495,3.2306714,3.0626216,2.7642474,2.4795918,2.136633,1.6839274,1.3992717,1.3169615,1.529596,2.1503513,2.8122618,2.6716487,2.270387,2.1263442,2.760818,4.8254294,6.7494283,7.4456344,6.2658563,3.0077481,2.201795,3.2546785,3.7794054,2.8294096,0.89855194,0.864256,0.9568549,0.83338976,0.5453044,0.53501564,0.94999576,0.99801,0.85739684,0.7133542,0.7613684,1.2037852,1.4850113,1.5638919,1.5947582,1.937717,2.1469216,1.7593783,1.4953002,1.4918705,1.2963841,1.0288762,0.99801,0.881404,0.6893471,0.7613684,1.08032,1.039165,1.1214751,1.3786942,1.4644338,1.3684053,1.2963841,1.1077567,0.8162418,0.61046654,1.0871792,1.8828435,2.8225505,3.3952916,2.760818,2.4452958,2.7230926,2.942586,2.7813954,2.2429502,1.5364552,1.6153357,2.218943,3.0900583,3.981751,4.4721823,4.1155047,4.0606318,4.616225,5.2644167,5.055212,5.2506986,6.3001523,7.490219,6.927767,5.802862,4.698535,3.6936657,2.8259802,2.1057668,2.020027,2.9700227,4.5853586,6.5642304,8.652849,9.554831,9.047252,7.1198235,4.482471,2.5790498,2.3595562,3.0557625,4.482471,5.919468,6.1046658,4.664239,3.450165,2.6990852,2.609916,3.340418,4.1943855,4.931747,5.267846,5.096367,4.4859004,3.4981792,2.9391565,3.117495,3.7691166,4.07435,4.4413157,4.8254294,4.6127954,4.0846386,4.4413157,8.200144,15.868701,22.889067,26.472986,25.619019,20.028791,18.430603,22.964518,31.0069,35.1567,29.089762,26.236343,27.693918,31.524769,32.7457,31.538486,33.1744,33.963203,32.488483,29.631636,26.630747,29.741383,30.540476,28.407272,30.5199,39.038994,64.212166,83.10919,82.80053,60.36417,48.55953,43.329407,41.66263,39.580868,32.135235,28.204927,23.797907,20.148827,17.501184,15.121051,15.693792,12.579727,10.175586,9.496528,8.179566,4.1635194,10.820349,12.243628,6.8591747,7.4456344,2.2086544,4.249259,14.243076,23.935091,16.160215,14.5585985,10.672876,6.5813785,3.5153272,1.8313997,1.5501735,1.488441,1.4472859,1.2209331,0.61046654,2.0749004,2.3149714,2.6476414,3.07634,2.2600982,2.7951138,5.171818,5.967482,5.4153185,7.414768,6.5367937,7.1781263,7.7268605,7.394191,6.210983,3.7691166,3.0660512,3.1963756,4.0880685,6.5299344,8.824328,11.97269,14.30481,15.237658,15.275383,12.13731,8.652849,8.4264965,10.844356,11.063849,22.28203,20.60839,22.210009,29.401854,30.670801,36.285034,41.041874,40.050724,34.618256,32.227833,29.052036,25.008553,22.422644,22.052248,23.101702,25.800787,27.909983,35.75002,46.323437,47.362602,45.48319,60.868317,83.36298,95.60318,73.057076,42.492588,28.424421,20.073376,12.860953,8.3922,17.425734,17.412016,18.139088,21.256582,20.29287,17.401728,22.371199,23.232025,17.514904,12.253916,10.398509,10.353925,11.794352,12.88839,10.299051,15.306249,17.53548,15.093615,10.618003,11.276484,12.092726,22.95423,30.454737,30.75311,29.556185,27.834532,28.68507,26.647894,21.325174,17.394867,21.925352,22.086544,21.805317,21.318316,17.182234,20.258574,23.050257,22.642136,20.958208,24.778769,27.42984,18.248835,12.531713,14.973578,19.69955,17.672665,17.20281,16.609491,15.172495,13.121602,12.706621,13.107883,14.699212,16.55119,16.403717,15.6697855,15.909856,17.37429,17.87501,12.771784,14.640909,14.356253,12.260776,9.523964,8.131552,7.5210853,9.9869585,12.247057,12.662037,11.245617,11.149589,10.583707,10.590566,11.2250395,11.5645685,11.029553,9.174147,8.525954,9.270175,9.246168,9.050681,8.738589,8.98209,10.765475,15.3817,15.076467,12.22648,9.400499,7.6788464,6.6533995,7.997798,6.958633,6.4887795,7.9257765,11.002116,7.949784,5.4016004,3.6868064,2.9322972,3.0660512,4.3007026,4.9934793,7.250148,9.623423,7.0958166,6.48535,8.601405,9.774324,9.352485,9.719451,8.827758,10.463672,11.63659,11.207891,9.901219,11.784062,12.46312,11.705182,10.14129,9.263316,9.959522,9.784613,10.326488,11.108434,9.582268,8.690575,10.096705,9.328478,6.831738,7.98065,8.968371,8.3922,8.447074,9.517105,10.179015,9.349055,8.865483,8.272165,7.4765005,6.7459984,6.975781,6.9346256,6.910619,6.9552035,6.883182,6.869464,6.492209,5.7102633,4.6916757,3.799983,3.3952916,3.2032347,3.117495,3.0626216,2.9906003,2.843128,2.633923,2.369845,2.170929,2.2429502,2.3389788,2.1812177,2.1091962,2.2566686,2.5619018,2.3081124,2.1229146,2.0268862,2.0817597,2.411,2.253239,2.2223728,2.3081124,2.4418662,2.503599,2.369845,2.1160555,1.9137098,1.8245405,1.8005334,2.2155135,2.867135,2.417859,1.7182233,3.8308492,3.0248961,2.7573884,2.8945718,3.093488,2.8396983,6.0840883,3.974892,1.9308578,1.5776103,0.7476501,1.0666018,0.8711152,0.58302987,0.432128,0.45613512,0.65162164,1.1214751,0.9259886,0.28122616,0.548734,0.42869842,0.2503599,0.28808534,0.45956472,0.34981793,0.6790583,0.5796003,0.41498008,0.34981793,0.34981793,0.26407823,0.2709374,0.34638834,0.45956472,0.59674823,0.7888051,0.7305021,0.94999576,1.3272504,1.0837497,1.1214751,1.0940384,0.939707,0.7682276,0.85396725,0.84367853,0.77508676,0.7510797,0.77851635,0.77851635,0.65505123,0.6173257,0.65162164,0.71678376,0.71678376,0.7407909,0.764798,0.75450927,0.7305021,0.77851635,0.59674823,0.4938606,0.4698535,0.4938606,0.5178677,0.5178677,0.5007198,0.51100856,0.5555932,0.5796003,0.53158605,0.5178677,0.5418748,0.61046654,0.7339317,0.7922347,0.84367853,0.75450927,0.52815646,0.31895164,0.2469303,0.20234565,0.18862732,0.1920569,0.16804978,0.216064,0.39440256,0.53501564,0.5624523,0.48700142,0.2194936,0.13375391,0.12346515,0.1097468,0.061732575,0.037725464,0.01371835,0.01371835,0.030866288,0.030866288,0.0548734,0.08916927,0.09945804,0.12346515,0.24350071,0.40126175,0.52472687,0.59674823,0.6173257,0.5796003,0.6893471,0.8265306,1.039165,1.2483698,1.2346514,1.4918705,1.5844694,1.6256244,1.7113642,1.9068506,2.1400626,2.2326615,2.1846473,2.1194851,2.287535,2.3629858,2.4247184,2.4247184,2.3835633,2.3972816,2.3458378,2.335549,2.3149714,2.270387,2.1983654,2.0989075,2.0028791,1.9171394,1.862266,1.862266,2.0440342,2.218943,2.3389788,2.393852,2.3801336,2.2086544,1.8999915,1.6770682,1.587899,1.5261664,1.587899,1.611906,1.611906,1.6221949,1.7079345,1.5021594,1.4404267,1.471293,1.5330256,1.5570327,1.6187652,1.7525192,1.7765263,1.6633499,1.5398848,1.6633499,1.7319417,1.9137098,2.2326615,2.5619018,2.4658735,2.4967396,2.6922262,3.0351849,3.4638834,3.865145,4.197815,4.48933,4.722542,4.8082814,5.3330083,6.0223556,8.718011,14.476289,23.557837,25.913963,21.45893,16.61292,13.732068,11.108434,11.852654,14.750656,18.550638,22.69358,27.282368,30.200947,35.040096,42.57147,53.762215,69.77839,0.65162164,0.5144381,0.6344737,0.764798,0.8162418,0.84024894,0.85739684,0.7990939,0.77165717,0.805953,0.85739684,1.0254467,1.255229,1.5433143,1.8931323,2.3149714,2.5207467,2.4418662,2.2635276,2.0131679,1.5501735,1.2243627,1.1523414,1.1077567,1.0425946,1.0871792,1.4267083,1.5055889,1.3478279,1.1454822,1.2346514,1.4747226,1.4987297,1.4815818,1.4369972,1.2346514,1.3786942,1.8519772,2.2738166,2.6956558,3.5873485,4.822,4.65395,4.2081037,4.081209,4.3349986,4.431027,5.051782,5.435896,5.809721,7.4010496,11.979549,15.158776,15.175924,12.21962,8.433355,6.1046658,4.1635194,2.8054025,2.1674993,2.335549,3.2443898,4.016047,4.314421,4.0503426,3.3781435,3.1209247,3.1963756,3.093488,2.6579304,2.0989075,1.8519772,1.879414,2.1434922,2.4830213,2.627064,3.1209247,2.6785078,2.1743584,2.0749004,2.4452958,3.3266997,4.2252517,4.249259,3.3541365,2.3218307,2.4452958,3.625074,3.9028704,2.7711067,1.1934965,0.7956643,0.7373613,0.65162164,0.5041494,0.6207553,0.9774324,1.0460242,1.1797781,1.4610043,1.7147937,1.646202,1.5261664,1.488441,1.6153357,1.937717,1.8313997,1.5055889,1.3409687,1.3203912,1.0288762,1.3855534,1.4953002,1.2449403,0.7476501,0.37382504,0.72021335,1.3306799,1.6839274,1.6667795,1.587899,1.6633499,1.6907866,1.5604624,1.2998136,1.0734608,1.3649758,2.0131679,2.609916,2.9665933,3.1037767,3.7039545,3.426158,2.7779658,2.0817597,1.4850113,1.3341095,1.5398848,2.1434922,3.018037,3.8617156,3.4021509,2.9563043,2.942586,3.2855449,3.433017,3.508468,3.6799474,4.012617,4.3624353,4.3761535,4.2389703,3.5702004,2.9254382,2.651071,2.8980014,4.07435,6.684266,10.216741,14.160767,18.025911,18.224829,16.359133,12.641459,8.30646,5.579939,5.4976287,6.9517736,8.834618,10.024684,9.386781,7.507367,6.0086374,5.1512403,4.835718,4.6127954,4.4104495,4.180667,4.046913,3.8720043,3.2409601,2.7985435,3.0214665,3.625074,4.3452873,4.9523244,5.662249,6.276145,6.451054,6.1321025,5.586798,6.9826403,11.777204,18.533491,23.880217,22.508383,24.404943,25.10458,28.033447,33.08866,36.634853,29.892284,24.806206,24.000254,27.124607,30.85257,32.282707,36.00038,38.006687,35.90092,28.877127,29.59391,30.231813,31.17152,31.66538,29.820263,31.205816,42.07075,55.401554,62.308746,52.04056,41.933567,39.766068,44.114784,48.707,42.413708,34.460495,26.34266,23.640146,24.332924,18.818146,17.089634,15.782962,11.63659,5.90575,4.383013,2.9048605,9.253027,14.143619,14.057879,11.266195,4.0194764,8.587687,19.342873,26.35638,15.426285,18.12537,12.116733,5.874883,3.175798,3.1140654,2.2669573,2.07833,2.177788,2.1674993,1.6359133,1.8313997,1.8485477,2.2155135,2.5927682,1.7456601,2.6064866,6.8283086,7.857185,5.8543057,7.7097125,5.2575574,6.1286726,7.1541195,7.0786686,6.540223,5.90575,4.746549,3.7211025,3.415869,4.3349986,6.7940125,11.770344,16.341984,18.975908,19.521212,14.46943,14.225929,14.1299,14.109323,18.70497,25.752771,29.635065,33.92205,37.879795,36.49081,36.511387,39.128162,40.266785,38.353077,34.289017,27.618467,23.44809,22.004232,22.155134,21.417774,21.743584,23.94195,32.17982,40.853245,34.59425,38.89838,59.578793,83.671646,96.323395,80.79765,53.405537,35.221863,22.258022,12.912396,7.9772205,12.919256,14.805529,16.180794,18.03277,19.792149,16.568336,16.410576,16.393429,14.891269,11.592006,11.05699,12.902108,15.004445,15.241087,11.519984,14.3974085,14.249936,14.2362175,15.29253,16.146498,18.156237,26.112879,27.52587,24.408375,33.280716,34.33017,30.368998,26.304935,23.636717,20.457489,19.70641,19.233126,19.665255,21.342323,24.322634,27.01829,27.004572,24.891945,21.325174,16.993607,15.337115,11.773774,12.668896,17.895588,20.821026,18.190533,16.221949,14.634049,13.443983,12.977559,12.932974,13.841815,15.518884,17.233677,17.720678,16.335125,15.553179,16.324837,17.545769,16.067617,17.806417,17.103354,14.507155,11.2593355,9.280463,9.342196,9.6645775,9.901219,9.777754,9.084977,9.956093,10.487679,11.118723,11.746337,11.736049,12.919256,11.698323,10.717461,10.600855,9.942374,8.272165,7.7440085,8.186425,9.880642,13.536582,15.450292,12.641459,8.944365,6.4716315,5.6039457,6.135532,7.5450926,8.165848,7.81603,7.81603,5.593657,4.7774153,4.331569,3.957744,4.091498,3.8685746,4.976331,6.9792104,8.529384,7.3530354,8.958082,7.7714453,7.2124224,8.659708,11.427385,11.808069,11.012405,10.666017,11.286773,12.295071,12.788932,12.339656,11.170166,9.633711,8.186425,8.776315,9.301042,9.208443,8.584257,8.141841,7.377043,7.966932,8.615124,8.594546,7.747438,8.934075,8.827758,9.0369625,9.781183,9.932085,9.191295,8.423067,8.076678,8.028665,7.599966,7.449064,7.3427467,7.298162,7.2535777,7.051232,6.3481665,5.4667625,4.4756117,3.642222,3.433017,3.4604537,3.3541365,3.3541365,3.532475,3.7725463,3.3438478,3.000889,2.7059445,2.4967396,2.510458,2.5001693,2.3081124,2.3424082,2.568761,2.503599,2.510458,2.503599,2.4967396,2.5413244,2.702515,2.633923,2.6613598,2.620205,2.6133456,3.0283258,2.884283,2.4658735,2.1469216,1.99602,1.7765263,2.4144297,3.2718265,3.1826572,2.9734523,5.4667625,5.830299,6.5024977,9.146709,11.4205265,6.9620624,8.423067,4.6745276,2.2292318,2.301253,0.7956643,0.78194594,0.6001778,0.41498008,0.37725464,0.6173257,0.48014224,0.70649505,0.6173257,0.26064864,0.40126175,0.39783216,0.24350071,0.2194936,0.33952916,0.33952916,0.6893471,0.66533995,0.45613512,0.2709374,0.33952916,0.22292319,0.29494452,0.45270553,0.5761707,0.53501564,0.9534253,1.0014396,1.039165,1.138623,1.0700313,0.84367853,0.88826317,0.91227025,0.8265306,0.7579388,0.8025235,0.91227025,0.97057325,0.90884066,0.70649505,0.64133286,0.6756287,0.7305021,0.8093826,0.9842916,1.0871792,1.1043272,0.9534253,0.7339317,0.70649505,0.64819205,0.59331864,0.5693115,0.59331864,0.6790583,0.75450927,0.7133542,0.6859175,0.6893471,0.6173257,0.607037,0.6173257,0.6241849,0.6276145,0.67219913,0.64476246,0.72707254,0.6824879,0.490431,0.33266997,0.26064864,0.22978236,0.2194936,0.216064,0.1920569,0.2503599,0.30523327,0.37382504,0.45956472,0.5624523,0.37039545,0.26750782,0.22292319,0.1920569,0.12346515,0.08916927,0.048014224,0.0274367,0.030866288,0.030866288,0.044584636,0.061732575,0.07545093,0.08916927,0.13375391,0.216064,0.3018037,0.37725464,0.42183927,0.432128,0.4938606,0.6036074,0.75450927,0.91912943,1.0528834,1.2689474,1.3649758,1.4232788,1.4918705,1.5913286,1.821111,2.0337453,2.1469216,2.153781,2.1297739,2.0680413,2.1194851,2.1915064,2.253239,2.335549,2.2360911,2.2498093,2.2806756,2.2498093,2.0886188,2.0097382,1.99602,2.0131679,2.0234566,1.99602,1.9823016,2.1674993,2.2258022,2.1057668,2.0268862,1.903421,1.7971039,1.704505,1.6359133,1.6221949,1.704505,1.7319417,1.7250825,1.7250825,1.8313997,1.6324836,1.546744,1.5364552,1.5638919,1.5673214,1.670209,1.7182233,1.670209,1.5604624,1.5158776,1.7456601,1.9514352,2.1880767,2.4555845,2.6990852,2.5721905,2.551613,2.633923,2.7573884,2.7916842,2.884283,3.2066643,3.4227283,3.4673128,3.5599117,3.882293,4.616225,7.2192817,12.336226,19.78872,19.829874,13.828096,9.191295,8.241299,8.203573,9.5033865,11.962401,15.529172,20.179693,25.889956,29.611057,34.364468,40.592598,49.85934,64.87064,1.0048691,0.84367853,0.9602845,1.0323058,1.0151579,1.1008976,1.0837497,1.0117283,0.9602845,1.0014396,1.1729189,1.313532,1.605047,1.8382589,2.0234566,2.3801336,2.5378947,2.3972816,2.1674993,1.8931323,1.4232788,1.0357354,0.9602845,0.9877212,1.0288762,1.0940384,1.3752645,1.4987297,1.4953002,1.4198492,1.3546871,1.5330256,1.5638919,1.5398848,1.4678634,1.2586586,1.3101025,1.529596,1.7662375,2.153781,3.1072063,4.0434837,3.7622573,3.3850029,3.5050385,4.187526,4.5956473,5.360445,5.3227196,4.715683,5.164959,9.89436,11.670886,11.269625,9.599416,7.7131424,5.754848,4.1360826,3.0317552,2.6236343,3.100347,4.173808,5.003768,5.5147767,5.446185,4.3624353,3.2581081,2.836269,2.6579304,2.4384367,2.0268862,1.6633499,1.6942163,2.1674993,2.8739944,3.350707,3.2032347,2.5824795,2.1194851,2.095478,2.428148,2.568761,2.719663,2.6990852,2.5378947,2.4727325,2.5481834,3.0386145,3.0797696,2.4384367,1.5124481,0.9602845,0.89169276,0.85739684,0.77851635,0.97057325,1.2106444,1.1180456,1.0597426,1.2346514,1.6873571,1.903421,1.7696671,1.6976458,1.862266,2.2292318,1.99602,1.7765263,1.5810398,1.3512574,0.9602845,1.3992717,1.4129901,1.1317638,0.77165717,0.64133286,1.039165,1.4404267,1.9102802,2.2258022,1.8931323,1.546744,1.5158776,1.5055889,1.4781522,1.646202,1.8485477,2.2292318,2.585909,2.9700227,3.666229,4.5099077,4.4550343,3.7382503,2.7299516,1.937717,2.2326615,2.061182,1.9548649,2.136633,2.5207467,2.287535,2.0714707,2.3904223,3.0420442,3.093488,3.1826572,3.3609958,3.57363,4.07435,5.4153185,5.802862,5.212973,4.90431,5.3878818,6.447624,9.746887,15.367981,23.087982,30.811415,34.577103,30.969175,24.308916,17.665806,12.902108,10.690024,11.482259,13.227919,14.167625,13.519434,11.499407,9.9698105,9.067829,8.1487,6.9620624,5.6348124,4.7362604,4.396731,4.5442033,4.8117113,4.557922,4.90431,7.3221693,9.304471,9.671436,8.570539,9.331907,9.647429,9.788043,9.781183,9.407358,9.071259,11.612583,16.907866,22.78275,25.015411,25.4544,29.206367,32.9309,34.36104,32.306713,30.26611,24.476965,22.035099,24.723896,29.01774,30.475315,31.809423,33.122955,32.714836,27.083452,26.469557,30.629646,34.25472,33.325302,25.114868,29.196077,32.138664,36.535397,40.887543,39.622025,32.965195,33.380177,42.300533,54.355534,57.3427,49.927933,37.101276,29.456726,27.861969,23.461807,21.95279,18.564358,12.178465,5.295283,4.029765,2.4967396,7.7783046,14.188204,16.29054,8.889491,4.763697,11.365653,19.61038,22.470657,15.014734,13.821238,9.0644,4.4413157,2.3252604,3.7794054,2.6887965,3.357566,3.9131594,3.6010668,2.7882545,2.3458378,1.8348293,1.6770682,1.8176813,1.7182233,2.9665933,6.6568294,7.623973,6.0566516,7.4799304,4.482471,7.7920227,9.016385,7.239859,9.030104,9.39707,6.684266,4.383013,3.7279615,3.6936657,7.8777623,13.896688,16.695232,15.937293,16.016174,13.488567,12.737488,11.893809,13.876111,26.380386,27.882545,34.127827,41.161907,46.70069,50.143997,51.70103,52.335506,49.979378,44.72868,38.843506,28.26666,23.420652,23.074265,24.240324,22.186,20.063087,20.097382,24.94682,30.24896,24.638157,34.51194,58.899734,76.17457,78.50326,71.83957,54.05716,37.605427,23.221737,12.754636,9.174147,13.011855,14.006435,15.241087,17.55263,19.54179,17.007324,17.590355,17.20624,15.12448,13.965281,13.001566,14.778092,16.901007,16.414005,9.767465,11.845795,13.80066,15.738377,17.604073,19.20569,22.083115,21.472647,24.267761,33.291004,47.30087,34.41248,28.582182,27.26522,26.195189,19.36688,14.874121,16.345413,18.310568,20.004784,25.365229,35.58197,36.00381,30.382715,21.674994,12.05157,10.635151,11.262765,14.490007,18.787281,20.526081,17.604073,15.004445,13.114742,12.202472,12.445972,13.080446,15.13134,17.528622,19.198832,19.085653,16.105343,14.466,14.544881,15.954441,17.532051,19.754423,19.44576,16.47231,12.243628,9.73317,9.496528,8.656279,8.213862,8.443645,8.875772,10.556271,11.519984,12.3911,12.9809885,12.284782,13.039291,13.498857,13.015285,11.900668,11.423956,8.889491,7.874333,7.7714453,8.460793,10.31277,12.689473,12.082437,10.63858,9.506817,8.848335,7.9600725,8.368194,8.652849,8.165848,6.999788,5.439326,4.290414,3.9371665,4.2286816,4.496189,4.0194764,4.32128,5.171818,6.310441,7.4524937,8.786603,7.010077,6.852316,9.595985,13.073587,11.739478,11.273054,11.115293,11.211322,11.979549,11.96926,10.14129,8.529384,8.2481575,9.458802,8.738589,9.23245,9.208443,8.303031,7.517656,8.351046,9.002667,9.465661,9.379922,8.028665,7.966932,9.777754,10.635151,9.609704,7.658269,7.64798,8.81404,8.752307,7.3050213,6.5779486,6.392751,6.2487082,6.40304,6.7219915,6.6739774,5.970912,5.0140567,4.0949273,3.4878905,3.4433057,3.590778,3.8514268,4.0023284,4.07435,4.3349986,4.0674906,3.6044965,3.210094,2.959734,2.7711067,2.7402403,2.4418662,2.428148,2.6476414,2.4590142,2.6956558,2.7882545,2.7573884,2.6990852,2.7779658,2.49331,2.7402403,2.836269,2.7745364,3.223812,3.508468,3.2889743,2.7813954,2.318401,2.3561265,2.5310357,3.1380725,3.1792276,3.1209247,4.8940215,6.711703,10.88894,20.306587,29.148064,22.916504,18.3723,9.163857,3.2821152,2.5756202,2.750529,2.335549,1.1763484,0.37039545,0.25378948,0.40126175,0.33952916,0.5727411,0.58988905,0.3566771,0.31209245,0.33609957,0.24007112,0.18519773,0.216064,0.26407823,0.48357183,0.58988905,0.490431,0.29837412,0.35324752,0.20920484,0.29151493,0.48014224,0.6241849,0.5453044,0.9431366,1.0048691,1.0014396,1.0494537,1.1420527,0.91569984,0.91227025,0.9362774,0.89855194,0.823101,0.9294182,1.0117283,0.9774324,0.8265306,0.65848076,0.77851635,0.96714365,1.0837497,1.1454822,1.3272504,1.1729189,1.0254467,0.8745448,0.7442205,0.6962063,0.61389613,0.58302987,0.6036074,0.67219913,0.7990939,0.88826317,0.8505377,0.823101,0.84367853,0.8265306,0.9362774,0.9294182,0.8471081,0.7442205,0.66533995,0.6824879,0.75450927,0.69963586,0.5212973,0.41840968,0.33609957,0.274367,0.24007112,0.22635277,0.216064,0.29837412,0.30866286,0.33609957,0.4081209,0.4972902,0.37725464,0.3018037,0.28465575,0.28808534,0.20234565,0.16462019,0.11317638,0.072021335,0.044584636,0.020577524,0.034295876,0.044584636,0.06859175,0.09602845,0.106317215,0.116605975,0.16804978,0.22635277,0.26750782,0.26750782,0.31895164,0.39440256,0.50757897,0.65162164,0.823101,1.0185875,1.0768905,1.1214751,1.2106444,1.371835,1.5913286,1.821111,1.9994495,2.0749004,2.0097382,1.961724,1.9480057,1.9308578,1.9720128,2.2086544,2.1880767,2.16064,2.1469216,2.1194851,2.0337453,2.0028791,2.0131679,2.0234566,2.0063086,1.9480057,1.9514352,2.0234566,2.0749004,2.0920484,2.1023371,2.0063086,2.0165975,1.9925903,1.9342873,1.9857311,1.961724,1.9480057,1.8931323,1.8142518,1.8073926,1.7490896,1.6976458,1.6736387,1.6873571,1.7182233,1.7765263,1.7902447,1.7353712,1.6496316,1.6496316,1.670209,1.8279701,1.9823016,2.0989075,2.2360911,2.1674993,2.1469216,2.2155135,2.3664153,2.5241764,2.6545007,3.0557625,3.350707,3.433017,3.4776018,3.724532,3.9474552,5.178677,7.4284863,9.6817255,9.019815,6.4064693,4.822,5.188966,6.3790326,8.704293,11.406808,14.54831,18.005335,21.44178,24.415234,27.464136,31.867727,38.65145,48.576675,1.430138,1.5364552,1.6770682,1.4507155,1.0323058,1.1694894,1.1454822,1.0563129,1.0117283,1.0734608,1.2586586,1.4095604,1.7456601,2.0131679,2.1880767,2.4658735,2.49331,2.3046827,2.0646117,1.7833855,1.3306799,1.0323058,0.90541106,0.8848336,0.9602845,1.1626302,1.3615463,1.5981878,1.762808,1.8073926,1.7388009,1.7456601,1.7079345,1.6256244,1.4953002,1.2929544,1.3889829,1.5193073,1.7971039,2.527606,4.2218223,4.5990767,4.0537724,3.4878905,3.4364467,4.046913,4.6093655,5.3330083,4.914599,3.5804894,3.07634,6.5299344,7.6616983,7.363324,6.6568294,6.691125,5.439326,4.4275975,3.690236,3.4364467,4.064061,5.6210938,6.9071894,8.011517,8.23444,6.0840883,3.6182148,2.4727325,2.1915064,2.3081124,2.3561265,1.9274281,2.061182,2.5550427,3.1449318,3.4981792,2.7916842,2.1469216,1.8588364,1.961724,2.2292318,2.1434922,2.0680413,2.194936,2.4727325,2.6064866,2.551613,2.5070283,2.4761622,2.3458378,1.8862731,1.5021594,1.4987297,1.605047,1.704505,1.862266,1.9308578,1.6427724,1.3032433,1.1900668,1.5364552,1.9754424,1.9137098,1.8656956,2.0337453,2.335549,2.1057668,1.9342873,1.6839274,1.3169615,0.8745448,1.1043272,1.097468,1.0528834,1.08032,1.214074,1.3101025,1.3478279,1.8245405,2.3972816,1.8691251,1.1729189,1.0460242,1.155771,1.3649758,1.7456601,2.0440342,2.2841053,2.4247184,2.633923,3.2855449,3.7519686,3.9371665,3.7382503,3.2032347,2.5653315,2.5447538,2.037175,1.6016173,1.5638919,2.020027,1.821111,1.762808,2.3972816,3.690236,5.0483527,5.3878818,5.23698,5.456474,6.368744,7.7748747,8.2481575,8.738589,9.781183,11.667457,14.455711,22.919933,33.002922,42.6675,48.648697,46.46405,38.42167,28.386696,20.742146,17.175373,16.647217,19.740705,21.921923,21.434921,18.471758,15.155347,13.773223,12.662037,11.084427,8.971801,6.914048,5.754848,5.3844523,5.6142344,5.960623,5.6348124,6.1801167,8.89635,11.22161,11.88352,10.875222,12.034423,12.511135,12.878101,13.368532,13.893259,12.47341,13.588025,16.931873,21.578964,25.968836,23.86307,28.534168,32.26556,31.552204,27.124607,27.52587,23.465237,20.927343,22.306036,26.390675,28.160343,26.918833,27.09374,28.520449,26.455837,26.075153,33.09895,37.968964,35.50652,24.888515,33.050934,31.891733,29.456726,29.76196,32.78343,28.702217,30.855999,41.25794,57.09577,70.73867,72.77585,59.760563,45.966763,37.9038,34.289017,32.200397,24.737614,15.117621,7.2158523,5.5422134,5.212973,7.133542,11.667457,14.606613,7.181556,4.588788,10.175586,16.266533,17.641798,11.540562,9.1810055,5.7582774,3.0660512,2.194936,3.5118976,2.620205,4.3624353,5.3158607,4.4413157,3.093488,2.4658735,1.8691251,1.4369972,1.2826657,1.4815818,3.7519686,7.7920227,9.47938,8.594546,8.81747,5.305572,7.517656,8.244728,6.9209075,9.626852,9.80862,9.277034,8.004657,6.358455,5.113515,10.981539,18.067066,18.509483,13.564018,13.622321,11.838936,9.544542,7.8091707,10.521975,24.35693,21.747015,27.323523,36.459946,45.9599,54.050297,59.03006,60.885468,58.738544,53.63875,48.583534,34.858326,26.898254,25.228045,26.798796,24.957108,21.10568,20.580954,22.000803,22.727877,18.855871,29.563044,51.718178,60.45334,54.19434,54.664196,47.595814,34.028366,20.906765,12.864383,12.205902,14.280802,13.780083,13.989287,15.656067,16.969599,17.847572,19.898466,18.763273,15.179354,14.977009,14.061309,15.412566,16.46888,15.083325,9.534253,11.321068,14.699212,18.238546,21.606401,25.59501,21.753874,18.982767,30.0912,50.147427,56.488735,31.401302,24.380938,25.10115,24.6896,15.748666,11.324498,16.53747,20.21056,20.03565,22.594122,42.204502,45.939323,37.23846,22.813616,12.662037,11.153018,13.375391,16.19794,17.830425,17.816708,18.166525,14.757515,12.229909,12.22648,13.419975,13.708061,15.590904,17.724108,18.9519,18.296848,16.12592,13.934414,13.423406,15.1862135,18.70497,22.830763,22.391777,18.578075,13.29994,9.177576,10.477389,9.462232,8.508806,8.841476,10.535692,12.099585,12.977559,13.958421,14.664916,13.54687,12.768354,13.701202,14.064738,13.289652,12.511135,9.458802,7.9943686,7.534804,7.716572,8.388771,9.767465,10.439664,11.080997,11.626302,11.283342,9.829198,8.368194,7.421627,6.7974424,5.6039457,5.2575574,4.1017866,3.5942078,4.0194764,4.4721823,4.2389703,3.9063,3.875434,4.647091,6.835168,7.3050213,6.5470824,7.39762,10.302481,13.317088,10.158438,10.041832,10.731179,11.173596,11.489118,10.429376,8.639131,7.7748747,8.378482,9.904649,9.026674,9.184435,9.534253,9.235879,7.449064,9.6817255,11.485688,12.257345,12.075578,11.701753,10.185875,11.132441,10.984968,9.078118,7.630832,8.155559,10.48082,10.679735,8.22758,5.9983487,6.2247014,6.447624,6.7528577,7.0478024,7.051232,5.007198,4.1155047,3.642222,3.3952916,3.74168,3.9303071,4.431027,4.7979927,4.8905916,4.9008803,4.835718,4.3281393,3.8514268,3.4707425,2.819121,2.5961976,2.3801336,2.3286898,2.428148,2.5138876,2.884283,3.1277838,3.1277838,2.9974594,3.0523329,2.3286898,2.510458,2.6853669,2.5961976,2.6476414,3.3301294,3.2512488,2.7779658,2.4144297,2.8122618,2.5310357,3.1655092,3.4913201,3.4227283,4.0229063,6.23499,11.478829,24.819925,38.833218,33.613388,25.145735,13.519434,4.9077396,1.9137098,3.5359046,4.4756117,2.3321195,0.5418748,0.2469303,0.29151493,0.35324752,0.4972902,0.490431,0.33609957,0.23321195,0.28465575,0.22635277,0.16119061,0.14061308,0.17147937,0.28122616,0.4664239,0.48014224,0.34638834,0.34638834,0.26407823,0.29837412,0.42526886,0.5453044,0.4972902,0.7476501,0.90884066,1.0323058,1.138623,1.2277923,1.0768905,1.0597426,1.0494537,0.9945804,0.9294182,0.9431366,0.9534253,0.89512235,0.7888051,0.7339317,0.86082643,1.0837497,1.2209331,1.2517995,1.3032433,1.0837497,0.88826317,0.78194594,0.7442205,0.66533995,0.5727411,0.61046654,0.6893471,0.78537554,0.91569984,0.980862,0.9568549,0.96714365,1.0185875,1.0151579,1.1763484,1.1626302,1.0631721,0.91227025,0.70649505,0.72021335,0.72707254,0.65848076,0.52815646,0.45956472,0.37382504,0.32581082,0.2777966,0.23664154,0.23664154,0.31895164,0.33952916,0.3806842,0.45613512,0.53844523,0.41498008,0.32924038,0.32238123,0.36010668,0.32924038,0.28808534,0.25721905,0.21263443,0.14404267,0.06516216,0.041155048,0.034295876,0.05144381,0.07545093,0.07545093,0.06516216,0.082310095,0.116605975,0.14747226,0.14747226,0.18176813,0.22292319,0.29837412,0.40126175,0.51100856,0.64819205,0.72364295,0.805953,0.94656616,1.1900668,1.4027013,1.6084765,1.762808,1.862266,1.9480057,1.8656956,1.7799559,1.7593783,1.8382589,2.0097382,2.0680413,2.0749004,2.085189,2.0886188,1.9891608,1.9651536,2.0063086,2.0165975,1.9582944,1.8245405,1.9308578,1.9548649,2.0097382,2.1229146,2.2498093,2.1091962,2.1091962,2.0577524,1.9685832,2.0234566,1.9239986,1.879414,1.821111,1.7319417,1.6359133,1.6427724,1.6290541,1.6221949,1.6256244,1.6393428,1.6496316,1.6427724,1.6153357,1.611906,1.728512,1.5844694,1.5981878,1.6427724,1.6770682,1.7250825,1.7010754,1.7525192,1.8862731,2.1023371,2.4075704,2.5481834,2.8156912,3.223812,3.5873485,3.5290456,3.4364467,3.3198407,3.5530527,3.7965534,2.9974594,2.5070283,2.5790498,3.1243541,4.245829,6.217842,9.218731,11.880091,14.2190695,16.362562,18.554068,20.683842,22.823904,26.099161,30.711956,35.959225,1.5398848,1.8691251,2.177788,1.7525192,0.91227025,1.0014396,1.097468,0.94999576,0.86082643,0.91912943,1.0185875,1.2415106,1.5810398,1.9308578,2.2258022,2.4658735,2.3424082,2.1503513,1.9308578,1.6770682,1.3238207,1.1763484,1.0117283,0.89855194,0.9294182,1.2243627,1.4404267,1.8279701,2.0886188,2.1640697,2.2223728,2.1057668,1.9480057,1.7147937,1.4335675,1.214074,1.4164196,1.7490896,2.3835633,3.690236,6.23499,5.8405876,5.0277753,4.2389703,3.8377085,4.091498,4.6676683,5.096367,4.3933015,2.942586,2.4761622,4.249259,5.8200097,6.025785,5.3878818,6.121814,5.305572,4.9591837,4.7259717,4.698535,5.4324665,7.932636,10.405369,12.188754,11.976119,7.8126,4.046913,2.4384367,2.095478,2.318401,2.6133456,2.301253,2.74367,3.1483612,3.1552205,2.8396983,2.0714707,1.587899,1.4610043,1.5981878,1.7216529,1.8759843,2.0577524,2.2909644,2.5241764,2.6064866,2.6613598,2.6613598,2.7916842,2.9254382,2.603057,2.651071,2.6545007,2.726522,2.8465576,2.8465576,2.702515,2.2738166,1.8073926,1.5158776,1.5776103,1.879414,1.8725548,1.8862731,2.0028791,2.0749004,1.9102802,1.728512,1.4747226,1.1592005,0.85739684,0.8162418,0.89855194,1.1454822,1.4472859,1.5227368,1.2106444,1.2175035,1.6942163,2.153781,1.4850113,0.8196714,0.65505123,0.83681935,1.1729189,1.4541451,1.8691251,2.0920484,2.0680413,1.9685832,2.1674993,2.1057668,2.2909644,2.6476414,2.9494452,2.7882545,2.16064,1.646202,1.4918705,1.845118,2.7573884,2.1160555,2.0646117,2.8122618,4.5270553,7.3393173,8.045813,7.8091707,8.272165,9.427936,9.616563,10.110424,12.80608,16.338554,20.560377,26.569014,39.975273,52.229187,59.252983,58.402447,48.47036,37.48196,27.611609,21.740154,20.323736,21.37662,25.708187,27.807095,26.34266,22.216867,18.547209,16.657507,14.688923,12.439114,10.028113,7.8846216,6.7974424,6.3310184,6.1972647,6.0154963,5.336438,5.73427,6.958633,8.47451,9.760606,10.319629,11.732618,12.744347,13.677195,14.750656,16.091625,14.784951,15.415996,17.189093,19.582945,22.343761,20.265432,23.125708,25.372087,25.01884,23.660725,23.60928,23.379498,22.408924,21.681852,23.725885,26.174612,24.500973,24.075705,25.889956,26.551867,29.789396,37.379074,41.48429,38.89838,31.017189,39.690617,35.67457,30.24896,29.583622,34.717712,31.548775,34.285587,42.784103,56.992886,76.942795,96.985306,94.049576,78.89766,62.10297,54.03658,48.919636,35.756878,20.968498,10.089847,7.7542973,9.084977,7.250148,8.416207,12.164746,11.523414,5.0620713,8.217292,14.061309,15.861842,7.082098,7.205563,4.420738,2.7059445,2.9631636,3.0248961,2.609916,5.2815647,6.461343,4.9214582,2.7882545,2.1263442,1.8691251,1.7182233,1.5330256,1.313532,4.033195,8.594546,11.118723,10.823778,10.017825,7.016936,5.6210938,5.552502,6.540223,8.337327,7.613684,11.129011,14.13676,13.725209,8.824328,14.832966,21.801888,21.44864,15.566897,16.023033,11.629731,8.196714,5.8405876,6.756287,15.21022,11.125582,14.188204,23.35206,35.365906,44.776695,52.318356,58.697388,62.363617,62.487083,58.964897,44.73211,33.050934,28.506731,29.641924,28.945719,26.534718,26.27064,24.240324,20.241425,17.802988,24.734184,39.15903,42.372555,35.49966,39.4917,38.949825,26.819374,16.03675,12.415107,14.63062,14.308239,13.056439,12.075578,12.1921835,13.834956,18.516342,20.008213,17.881868,14.373401,14.3974085,13.615462,15.117621,15.930434,15.086755,13.6086035,14.126471,17.312557,21.572105,26.099161,30.897154,19.236557,21.987085,39.978703,59.62681,52.95969,27.275509,19.301718,19.390888,19.582945,13.588025,11.231899,18.550638,22.511812,21.208569,23.873358,53.227196,57.874287,43.49746,22.913074,16.081335,15.117621,16.005884,15.988737,14.7026415,14.198492,19.336014,15.951012,13.015285,13.639469,15.076467,14.229359,14.819247,15.590904,15.848124,15.419425,15.930434,13.972139,13.173045,15.4742985,21.12283,28.002583,25.913963,20.220848,14.071597,8.419638,11.331357,11.029553,10.151579,10.412228,12.617453,13.347955,13.954991,14.894698,15.601193,14.493437,12.614022,12.915827,14.229359,14.970149,13.166186,10.106995,8.546532,8.255017,8.625413,8.656279,8.237869,8.4264965,9.582268,11.105004,11.451392,10.113853,7.4936485,5.3158607,4.1463714,3.4055803,4.3933015,4.1943855,3.758828,3.6936657,4.2526884,4.513337,4.331569,4.0606318,4.2183924,5.5113473,5.7274113,6.64997,8.292743,10.323058,12.082437,9.39707,8.968371,9.962952,11.30049,11.646879,9.431366,8.752307,9.115844,9.753747,9.595985,9.139851,8.89635,9.499957,10.000677,7.857185,10.05898,13.042721,14.983868,15.539461,15.834405,13.749216,12.295071,10.628291,9.294182,10.261326,11.108434,12.257345,12.22305,10.436234,7.2432885,8.028665,8.618553,8.433355,7.829748,8.1041155,4.8734436,3.7965534,3.4638834,3.426158,4.197815,4.3349986,4.7808447,5.3158607,5.65539,5.429037,5.435896,4.9351764,4.40359,3.8171308,2.6579304,2.1229146,2.1297739,2.1503513,2.1674993,2.6647894,2.9803114,3.3438478,3.426158,3.2718265,3.3026927,2.2635276,2.136633,2.2360911,2.1469216,1.7353712,2.5824795,2.4418662,2.2292318,2.4212887,3.0489032,2.5001693,3.3232703,4.07435,4.1017866,3.542764,5.103226,8.207003,19.44919,32.82115,29.748241,22.398636,15.127911,7.023795,0.69963586,2.2600982,5.3913116,3.5221863,1.1729189,0.31895164,0.39440256,0.4389872,0.37382504,0.2777966,0.20577525,0.17833854,0.2777966,0.21263443,0.1371835,0.11317638,0.09945804,0.16804978,0.3566771,0.4424168,0.3806842,0.30866286,0.36353627,0.33609957,0.33952916,0.4046913,0.4664239,0.5590228,0.83681935,1.1180456,1.2826657,1.2689474,1.1729189,1.155771,1.138623,1.0837497,0.97400284,0.823101,0.8025235,0.8162418,0.84367853,0.9294182,0.90884066,1.0082988,1.1111864,1.138623,1.039165,0.9877212,0.8711152,0.7613684,0.6790583,0.5727411,0.5727411,0.72364295,0.85396725,0.922559,1.0117283,1.0494537,1.0494537,1.1043272,1.1832076,1.1249046,1.1729189,1.1489118,1.0906088,0.97400284,0.72364295,0.6859175,0.6241849,0.548734,0.48357183,0.45956472,0.38754338,0.39097297,0.36010668,0.28808534,0.2709374,0.29494452,0.33609957,0.4115505,0.5212973,0.65505123,0.52815646,0.41840968,0.37039545,0.39097297,0.4424168,0.39097297,0.4081209,0.39097297,0.29837412,0.16804978,0.08916927,0.041155048,0.024007112,0.030866288,0.030866288,0.044584636,0.041155048,0.048014224,0.07545093,0.08916927,0.09945804,0.116605975,0.14404267,0.17490897,0.19891608,0.25378948,0.37382504,0.5178677,0.6859175,0.91912943,1.1249046,1.3169615,1.4404267,1.546744,1.8039631,1.6667795,1.5673214,1.6256244,1.7765263,1.7456601,1.821111,1.8999915,1.9891608,2.0131679,1.821111,1.7593783,1.845118,1.8931323,1.8245405,1.6599203,1.8519772,1.9445761,2.0268862,2.136633,2.2841053,2.0817597,1.9891608,1.8519772,1.6942163,1.704505,1.611906,1.5570327,1.546744,1.5364552,1.4232788,1.3992717,1.3958421,1.3924125,1.3786942,1.3375391,1.3306799,1.3203912,1.3306799,1.4095604,1.6359133,1.529596,1.4095604,1.3786942,1.4267083,1.4267083,1.4438564,1.611906,1.8142518,2.0165975,2.277246,2.2978237,2.2600982,2.6304936,3.210094,3.1586502,2.7985435,2.6785078,2.6853669,2.6167753,2.1743584,2.020027,2.3801336,3.216953,4.756838,7.4936485,10.851214,13.262215,14.723219,15.999025,18.602083,20.567236,23.156574,26.428402,29.950588,32.773136,0.9911508,0.78537554,1.4918705,1.5913286,0.9294182,0.7339317,1.2209331,1.1043272,0.89169276,0.83681935,0.94656616,1.1283343,1.3203912,1.546744,1.7833855,1.9548649,1.8691251,1.8931323,1.8245405,1.6187652,1.371835,1.2620882,1.08032,0.9328478,0.9294182,1.1763484,1.5776103,1.9891608,2.270387,2.369845,2.318401,2.318401,2.201795,1.8759843,1.4472859,1.1900668,1.471293,2.037175,3.1826572,4.976331,7.2467184,6.1972647,5.3673043,4.804852,4.605936,4.897451,5.288424,5.0483527,4.0777793,2.9391565,2.8534167,4.355576,6.159539,6.7700057,6.327589,6.6225333,6.012067,5.8405876,5.720552,5.994919,7.750868,10.926665,15.388559,17.405157,14.977009,7.874333,4.2835546,2.901431,2.452155,2.0886188,1.4027013,1.2586586,2.037175,2.452155,2.153781,1.7388009,1.6667795,1.5741806,1.3375391,1.0734608,1.1592005,1.8416885,2.4247184,2.6956558,2.7642474,3.083199,3.2649672,3.74168,4.2526884,4.5201964,4.2252517,4.715683,4.461893,3.7519686,3.0043187,2.760818,2.3835633,1.8965619,1.5364552,1.430138,1.6016173,1.6496316,1.8005334,1.8862731,1.8176813,1.587899,1.4541451,1.2998136,1.1214751,1.039165,1.2963841,1.138623,1.1523414,1.1763484,1.0837497,0.77851635,0.8265306,1.4061309,2.0063086,2.1091962,1.2037852,0.8505377,0.8162418,1.0082988,1.2963841,1.5398848,1.6633499,1.7319417,1.7422304,1.7525192,1.862266,2.0440342,2.2086544,2.318401,2.386993,2.4727325,2.5447538,2.3904223,2.5001693,2.9665933,3.4776018,2.7093742,2.7368107,3.3712845,4.3349986,5.2644167,5.6656785,7.1061053,8.790032,9.884071,9.506817,10.703742,15.63206,21.980227,29.569902,40.373104,49.78389,54.317806,53.964558,49.41007,42.039883,31.33271,24.562706,21.829325,21.85333,21.987085,20.841602,20.388897,19.325726,17.384579,15.333686,12.394529,10.906088,9.791472,8.471081,6.8969,5.9434752,5.844017,5.305572,4.3349986,4.2252517,5.422178,6.883182,8.186425,8.745448,7.8434668,7.7714453,8.519095,9.856634,11.293632,12.099585,13.173045,14.321958,15.916716,16.997036,15.289101,15.241087,15.247946,16.321407,18.752985,22.11055,25.077143,29.233803,30.831991,28.520449,23.345201,24.11343,24.562706,24.586712,24.35693,24.308916,31.559063,40.784653,44.941315,42.760098,38.757767,42.921288,34.703995,28.119188,30.42044,42.115334,39.268776,41.14133,45.424885,53.580444,70.81755,112.342995,135.76022,131.34634,105.93652,82.930855,72.38145,50.71331,27.44013,11.231899,9.901219,7.9120584,7.2432885,8.81061,14.232788,25.817934,9.191295,14.308239,21.260014,19.764713,9.170717,6.3618846,5.24041,4.4516044,3.7691166,4.07435,3.9508848,7.4353456,8.841476,6.608815,3.3266997,2.3492675,2.0886188,2.5619018,3.1312134,2.4727325,2.0680413,2.6476414,3.7451096,4.8940215,5.6005163,7.0889573,7.39762,7.438775,7.8983397,9.2153015,8.189855,9.050681,19.054789,29.309254,14.771234,18.005335,20.433481,21.699,21.918493,21.699,14.435134,10.422516,7.795452,7.6171136,13.855534,10.521975,11.4376745,16.383139,24.243753,33.02007,42.015877,53.37467,62.93979,66.18075,58.19667,48.70014,38.26048,33.390465,33.92548,33.033787,39.33394,34.738293,25.509272,18.512913,21.208569,24.175161,30.58506,34.08324,34.58739,38.284485,34.83089,22.182571,12.106443,9.283894,11.321068,11.664027,10.943813,10.127572,11.005547,16.204802,18.742695,17.309128,15.12448,14.363112,16.143068,12.627741,15.062748,20.76958,25.423532,23.053686,19.198832,23.86307,26.767931,24.621008,21.1194,20.78673,27.206917,34.450207,38.274197,36.08955,22.683292,15.350834,13.745787,16.105343,19.239986,15.066177,16.732958,17.024471,20.334024,42.64692,85.1155,78.036835,47.091667,17.525192,14.1299,21.174273,18.293419,12.041282,8.584257,13.687484,17.78927,18.310568,17.350283,15.906426,13.855534,12.902108,13.395968,13.118172,12.123591,12.771784,13.46799,13.310229,12.812939,15.179354,26.335802,34.84461,28.962866,19.750994,13.032433,9.383351,7.6274023,8.752307,10.5597,11.821788,12.298501,12.689473,13.337666,13.783512,13.663476,12.710052,12.199042,13.231348,15.563468,17.21653,14.496866,12.542002,11.540562,11.674315,11.952112,10.206452,8.255017,7.5931067,8.165848,9.668007,11.537132,9.205012,6.6705475,4.5647807,3.2718265,2.9288676,3.758828,4.3795834,4.2389703,3.7176728,4.1189346,5.3158607,5.926327,5.6142344,4.681387,4.0606318,5.1340923,7.6342616,9.709162,10.580277,10.542552,12.593445,12.531713,11.96926,11.674315,11.550851,10.429376,9.513676,8.97866,9.414218,11.856084,8.889491,8.2310095,8.512236,8.848335,8.834618,8.796892,10.628291,13.241637,14.586036,11.657167,10.851214,12.188754,12.926115,12.408247,12.055,13.862392,11.372512,9.709162,10.268185,10.7586155,11.513125,11.338216,9.115844,6.5882373,8.347616,9.139851,7.1129646,5.1855364,4.540774,4.6402316,4.3933015,4.5167665,4.972902,5.501058,5.6005163,5.638242,5.079219,4.417309,3.6970954,2.486451,1.9137098,1.9239986,2.1503513,2.4315774,2.8225505,2.750529,2.942586,2.952875,2.7402403,2.6545007,2.0440342,1.8999915,1.9068506,1.8828435,1.786815,2.6407824,2.3767042,2.369845,2.9871707,3.5873485,2.6579304,2.8568463,3.7553983,4.32471,2.9460156,4.15323,5.3981705,9.270175,13.2690735,9.829198,8.241299,12.703192,9.647429,0.19891608,0.19891608,2.7128036,3.9268777,2.6579304,0.22292319,0.4424168,0.31895164,0.24350071,0.20920484,0.20577525,0.22978236,0.32581082,0.23321195,0.12689474,0.08916927,0.07545093,0.12346515,0.29151493,0.42869842,0.42869842,0.26064864,0.4424168,0.42526886,0.34638834,0.3806842,0.7476501,0.77165717,0.8711152,1.0117283,1.1489118,1.2209331,1.1351935,0.94999576,0.9431366,1.0597426,0.90198153,0.7888051,0.7990939,0.7922347,0.83338976,1.1763484,1.1626302,1.0940384,1.1489118,1.2860953,1.2346514,1.1249046,0.97057325,0.72021335,0.4629943,0.42869842,0.6241849,0.8711152,1.0117283,1.0254467,1.039165,1.0734608,1.1008976,1.1797781,1.2723769,1.2346514,0.980862,0.8162418,0.7099246,0.6379033,0.5658819,0.6241849,0.58645946,0.48357183,0.4115505,0.53501564,0.51100856,0.4938606,0.48700142,0.4664239,0.3806842,0.26064864,0.2194936,0.274367,0.40126175,0.53501564,0.6310441,0.59331864,0.5007198,0.41840968,0.3806842,0.31895164,0.38754338,0.4115505,0.34981793,0.29151493,0.1920569,0.09602845,0.041155048,0.030866288,0.030866288,0.0548734,0.05144381,0.044584636,0.05144381,0.07545093,0.08916927,0.082310095,0.06859175,0.06516216,0.07545093,0.11317638,0.17833854,0.25721905,0.33266997,0.3806842,0.52815646,0.8025235,1.0528834,1.2037852,1.2655178,1.3169615,1.3272504,1.3101025,1.3169615,1.4644338,1.4541451,1.4575747,1.4575747,1.4198492,1.2963841,1.2346514,1.313532,1.3546871,1.3443983,1.4027013,1.5741806,1.7833855,2.0131679,2.1983654,2.1983654,2.0749004,1.9445761,1.7490896,1.5570327,1.5570327,1.4953002,1.4267083,1.4507155,1.5090185,1.371835,1.3992717,1.3478279,1.2929544,1.2517995,1.1900668,1.214074,1.2483698,1.2723769,1.2929544,1.3443983,1.4404267,1.3272504,1.255229,1.2895249,1.3272504,1.5090185,1.7319417,1.8828435,1.9582944,2.0440342,1.99602,1.8554068,1.7696671,1.8759843,2.3046827,2.8054025,2.6167753,2.311542,2.1983654,2.318401,1.9891608,2.510458,3.7142432,5.761707,9.153569,13.440554,16.496315,17.826996,18.21111,19.713268,22.312897,25.382378,29.446438,33.58938,35.444786,0.6859175,0.607037,0.8196714,0.8196714,0.59674823,0.6344737,1.2003556,1.4644338,1.430138,1.2106444,1.0082988,1.1214751,1.2963841,1.5261664,1.7490896,1.8416885,1.7662375,1.8382589,1.879414,1.8039631,1.6290541,1.4507155,1.2517995,1.1249046,1.1111864,1.2003556,1.4747226,1.9137098,2.1126258,2.037175,2.037175,2.07833,2.0131679,1.7765263,1.4232788,1.1180456,1.4953002,2.311542,3.7485392,5.73427,7.956643,7.3839016,6.351596,5.7136927,5.953764,7.191845,5.9434752,4.32471,3.1209247,2.8396983,3.7313912,5.4667625,5.3227196,5.3398676,6.0223556,6.355026,7.3839016,7.39762,7.7577267,9.050681,11.070708,15.388559,19.46291,20.076805,16.578627,10.88894,7.0375133,4.870014,3.9200184,3.57363,3.07634,3.457024,2.719663,1.8245405,1.2723769,1.0940384,1.2346514,1.313532,1.138623,0.8745448,1.039165,1.8176813,1.9720128,1.9685832,2.1880767,2.935727,4.1155047,4.232111,3.8479972,3.5016088,3.724532,4.1155047,3.7965534,3.0729103,2.3081124,1.9068506,1.7250825,1.4027013,1.1214751,1.0151579,1.1866373,1.3443983,1.6736387,1.9685832,2.0577524,1.8073926,1.5844694,1.6599203,1.8348293,1.8999915,1.6393428,1.1008976,0.78537554,0.75450927,0.91227025,0.99801,1.3992717,1.6256244,1.5981878,1.3032433,0.7888051,0.72021335,0.7579388,0.8779744,1.0425946,1.2003556,1.1351935,1.1797781,1.2312219,1.3306799,1.6530612,2.0337453,2.311542,2.5447538,2.8499873,3.4227283,3.7211025,3.2855449,2.9082901,2.860276,2.9048605,3.0043187,3.7553983,4.4550343,4.7945633,4.8734436,4.5819287,5.5902276,6.9689217,8.399059,10.179015,13.9309845,19.685833,27.021719,35.194427,43.14421,50.154285,52.87052,50.973957,45.356293,38.119865,28.225504,22.398636,18.814716,16.03675,13.015285,10.542552,8.97523,8.220721,7.932636,7.5245147,7.257007,6.7700057,6.444195,6.310441,6.0532217,6.2658563,6.2555676,5.6656785,4.7499785,4.386442,5.2609873,6.025785,6.9552035,8.018375,8.8929205,8.244728,9.853205,11.458252,12.360233,13.430264,15.138199,16.952452,18.03277,18.276272,18.303709,17.014183,17.772121,18.516342,19.11995,21.400625,22.786179,25.814505,26.754211,25.10801,23.60242,22.974806,26.164322,28.664492,28.667921,27.076593,31.613937,37.358498,38.551994,37.33106,43.73753,45.575787,37.042973,28.661062,27.128036,35.31446,38.672028,46.405746,51.903378,56.653355,70.26539,141.15497,195.55508,196.58395,150.32568,105.8405,87.94148,64.12643,36.97095,14.078457,8.05953,5.171818,5.5422134,7.3701835,13.440554,31.126936,14.55174,15.21365,18.650097,17.141079,9.709162,14.153908,9.6988735,5.90232,6.1286726,7.517656,6.9552035,10.878652,11.965831,8.659708,5.1683884,3.3541365,2.668219,3.4776018,4.4721823,2.6785078,2.0714707,2.3321195,3.7005248,6.2212715,9.760606,11.008976,11.406808,10.39508,9.0369625,10.034973,14.565458,15.817257,22.77246,29.813404,16.760393,22.065966,22.295748,18.221397,13.265644,13.495427,12.092726,12.267634,15.028452,18.413456,17.490896,15.254805,15.666355,18.838724,24.185452,30.430729,35.756878,39.25506,42.585186,45.273983,44.72182,42.73266,40.088448,37.341347,36.32276,40.139893,49.924503,43.408287,31.2504,22.343761,23.808197,26.579304,31.291555,34.66627,35.448215,34.40219,26.054577,17.415445,11.156448,8.477941,9.102125,9.832627,10.257896,9.72288,9.918367,14.874121,16.407146,14.750656,13.543441,13.869251,14.277372,13.279363,18.139088,26.815945,32.526207,23.76361,14.644339,14.850114,20.515793,28.414133,35.972942,26.620459,21.174273,19.058218,19.507494,21.561817,16.047039,13.543441,16.78783,22.158566,19.682402,18.269413,21.232576,22.885637,33.699127,80.3278,111.89029,86.645096,45.592937,17.021042,16.496315,20.94449,16.153357,10.796341,10.508256,17.885298,21.263443,20.491785,17.031332,13.032433,11.351934,11.105004,12.895248,12.710052,10.521975,10.281903,10.899229,12.027563,16.019604,26.02714,46.011345,48.13426,32.886314,18.835295,13.618892,13.9138365,9.956093,8.014946,7.671987,8.433355,9.6988735,10.988399,11.653738,12.089295,12.205902,11.427385,10.525404,10.628291,11.029553,11.592006,12.7272,14.191633,15.141628,14.740367,13.766364,14.627191,12.449403,9.942374,8.611694,8.838047,9.877212,7.81603,5.360445,3.758828,3.3952916,3.7965534,4.479041,4.99005,4.9214582,4.4550343,4.3521466,4.523626,5.871454,6.166398,5.2747054,5.1683884,5.9812007,7.706283,9.414218,10.991828,13.1421795,15.673215,14.939283,12.024134,8.98209,8.841476,8.556821,8.347616,8.735159,9.791472,11.0981455,10.192734,10.216741,11.211322,12.380811,12.092726,11.540562,12.127021,12.281353,11.06042,8.179566,9.80519,9.887501,8.80718,7.2021337,5.9880595,9.14328,8.272165,8.549961,10.943813,12.233338,10.834066,9.962952,9.304471,8.625413,7.7851634,8.539673,7.425057,6.8591747,6.7802944,4.664239,4.5270553,4.7328305,4.9831905,5.06893,4.90431,5.3227196,4.8940215,4.0709205,3.07634,1.937717,1.6564908,1.7147937,1.9480057,2.2258022,2.4315774,2.2326615,2.311542,2.4452958,2.4487255,2.177788,1.920569,1.7182233,1.8108221,2.085189,2.0646117,2.0406046,2.1812177,2.2155135,2.3218307,3.1346428,2.959734,2.750529,3.4398763,4.3007026,2.9803114,3.9646032,4.3109913,5.4736214,7.250148,7.8126,6.2075534,9.129561,7.174697,0.7442205,0.05144381,1.3546871,3.6353626,3.0900583,0.31552204,0.31895164,0.36353627,0.29151493,0.21263443,0.16462019,0.12003556,0.30523327,0.26064864,0.13375391,0.030866288,0.0274367,0.058302987,0.24007112,0.42526886,0.48014224,0.31895164,0.34638834,0.37725464,0.4355576,0.5727411,0.8711152,1.0220171,1.1214751,1.1866373,1.2449403,1.3169615,1.1660597,0.9774324,0.980862,1.1043272,0.97400284,0.83338976,0.85739684,0.9259886,0.980862,1.0288762,1.0734608,1.1249046,1.1489118,1.1420527,1.1146159,1.0528834,1.0185875,0.9945804,0.96371406,0.9259886,0.86082643,0.85396725,0.939707,1.0631721,1.0734608,1.0906088,1.1592005,1.1729189,1.1317638,1.1146159,0.85739684,0.7133542,0.65162164,0.6379033,0.66191036,0.607037,0.5658819,0.58988905,0.66876954,0.7407909,0.64819205,0.6379033,0.65162164,0.66876954,0.7099246,0.548734,0.35324752,0.25378948,0.29494452,0.44927597,0.48700142,0.5521636,0.52815646,0.432128,0.4046913,0.33609957,0.32581082,0.33952916,0.3841138,0.51100856,0.4698535,0.29837412,0.12689474,0.030866288,0.030866288,0.044584636,0.048014224,0.0548734,0.06516216,0.05144381,0.07545093,0.08573969,0.082310095,0.06859175,0.05144381,0.058302987,0.072021335,0.106317215,0.16462019,0.22292319,0.28122616,0.38754338,0.548734,0.7407909,0.88826317,1.0048691,1.1146159,1.2963841,1.4644338,1.3684053,1.4129901,1.3478279,1.255229,1.2003556,1.2243627,1.1934965,1.2312219,1.3375391,1.4404267,1.4027013,1.4678634,1.5810398,1.7113642,1.8348293,1.9514352,1.7525192,1.5810398,1.4232788,1.3169615,1.3375391,1.4129901,1.4335675,1.4095604,1.371835,1.3855534,1.2620882,1.1694894,1.1660597,1.2037852,1.1420527,1.1454822,1.2277923,1.1866373,1.0288762,0.9534253,1.0220171,0.9877212,0.9774324,1.0425946,1.155771,1.4095604,1.6290541,1.7936742,1.8759843,1.8725548,1.7353712,1.7147937,1.7216529,1.8073926,2.1469216,2.9871707,2.8054025,2.393852,2.177788,2.2223728,2.2052248,2.5550427,3.3952916,5.0277753,7.936065,12.504276,17.031332,20.337454,22.319756,23.948809,29.724234,35.033237,38.699467,40.369675,40.537724,0.4355576,0.45956472,0.53501564,0.5521636,0.5761707,0.8471081,1.471293,1.8519772,2.1126258,2.1674993,1.7559488,1.3752645,1.5055889,1.8519772,2.2120838,2.4830213,2.3458378,2.194936,2.0131679,1.821111,1.6770682,1.4953002,1.2483698,1.1934965,1.371835,1.6256244,1.8348293,2.095478,2.153781,2.0028791,1.8691251,1.8725548,1.786815,1.5810398,1.3101025,1.1180456,1.5913286,2.644212,4.331569,6.444195,8.508806,7.9257765,6.6225333,6.042933,6.444195,6.8866115,4.7019644,3.3815732,3.450165,4.623084,5.809721,5.936616,4.695105,4.338428,5.377593,6.560801,7.431916,7.966932,8.608265,10.031544,13.128461,18.331144,21.527521,22.083115,20.779871,19.826445,17.20281,14.212211,12.0138445,10.840926,9.993818,8.940934,6.0532217,3.4913201,2.1434922,1.6187652,1.5501735,1.4232788,1.1592005,0.89512235,0.9877212,1.7936742,1.7147937,1.5124481,1.7422304,2.74367,3.2786856,3.3609958,3.0969174,2.8122618,3.069481,3.3061223,2.9940298,2.3458378,1.670209,1.3546871,1.2415106,1.0117283,0.83338976,0.8128122,0.9842916,1.1592005,1.4095604,1.704505,1.8691251,1.605047,1.5090185,1.6873571,1.8279701,1.7147937,1.2209331,0.8128122,0.65505123,0.8162418,1.155771,1.3169615,1.2860953,1.2792361,1.2655178,1.1523414,0.7956643,0.91227025,0.84367853,0.7956643,0.86082643,1.039165,1.0837497,1.0494537,0.99801,1.0254467,1.2620882,1.7353712,2.1469216,2.5413244,2.9803114,3.5530527,3.474172,2.9700227,2.4555845,2.1983654,2.3218307,2.74367,3.5461934,4.5784993,5.535354,5.967482,6.5950966,6.8111606,7.56567,9.095266,10.930096,13.927555,19.438902,26.726774,34.72114,42.015877,48.31603,49.554108,45.177956,36.528538,26.85024,19.041069,15.858413,12.830087,8.879202,6.3138704,5.1340923,4.3590055,4.2355404,4.417309,3.9474552,4.629943,5.055212,5.861165,6.6465406,5.970912,6.8454566,6.5333643,6.025785,5.9434752,6.5127864,6.7940125,7.0478024,8.577398,10.909517,11.818358,11.917816,12.583157,13.121602,13.330807,13.505715,15.244516,16.856422,18.413456,19.915615,21.311457,20.443771,20.464348,21.013083,22.333473,25.27263,26.479845,27.01829,25.979126,24.933102,27.913412,29.508171,31.32928,31.353289,29.796255,29.106909,31.881445,33.699127,34.042084,34.896053,40.764076,42.862984,37.39965,29.864847,25.632736,29.960876,35.92493,46.371452,52.596153,55.727367,66.75006,144.14214,202.63031,203.84782,155.69984,112.38758,94.16618,69.15763,41.011005,17.703531,11.55428,6.4133286,6.4373355,8.683716,13.529722,24.665592,13.958421,16.228807,17.71039,13.989287,10.007536,15.271953,9.640571,5.4941993,6.262427,6.3893213,8.282454,11.7257595,12.065289,8.862054,5.9126086,4.7602673,3.9131594,4.8494368,6.135532,3.40901,2.7779658,2.9322972,3.782835,5.295283,7.4696417,10.858074,13.588025,15.261664,17.240536,22.624989,26.383816,24.638157,27.128036,29.984882,15.721229,17.87501,20.138538,19.932762,16.918156,13.018714,13.2690735,13.38911,15.858413,19.11309,17.532051,18.437462,19.332584,19.404606,19.582945,22.52553,22.991955,23.554407,25.828222,29.604198,32.865738,35.098396,38.6686,38.589718,37.018967,43.271107,62.596832,54.44813,38.74748,27.793377,26.246634,25.883097,29.192648,32.16953,32.24155,28.242653,20.882757,14.198492,9.424506,7.1952744,7.5279446,9.170717,9.932085,9.767465,10.216741,14.387119,13.838386,12.127021,11.732618,13.697772,17.655516,22.237446,25.9414,28.153484,26.260351,15.645778,11.4205265,11.869802,18.814716,31.76141,47.88047,30.7634,16.96617,10.64201,11.626302,15.419425,13.207341,15.244516,20.879328,25.584723,20.96164,26.174612,33.270428,41.57003,63.546825,124.823265,118.173294,79.12058,39.275635,16.945591,17.117071,17.237106,12.662037,11.965831,17.916164,27.467566,26.719915,20.598103,14.634049,11.574858,11.38623,13.2690735,15.3817,14.911846,12.144169,10.463672,11.458252,14.54831,24.164873,41.81353,66.084724,51.646156,31.219534,18.584934,16.143068,14.887839,12.30536,9.72631,8.093826,8.14527,10.422516,11.626302,11.019264,10.525404,10.878652,11.612583,8.81747,7.39762,7.466212,8.872343,11.177026,13.341095,15.62863,15.87899,14.009865,12.024134,10.1652975,8.093826,7.0615206,7.3427467,8.213862,7.301592,5.9469047,4.5030484,3.7553983,4.928317,4.8734436,5.1238036,5.3398676,5.038064,3.6147852,3.8720043,4.712253,5.3570156,6.094377,8.285883,8.042382,8.217292,8.868914,10.347065,13.310229,15.861842,14.843254,11.574858,8.179566,7.548522,7.73372,6.914048,6.866034,7.7440085,8.073249,7.0752387,7.579388,9.544542,11.859513,12.332796,12.452832,13.149038,11.914387,9.071259,7.740579,14.572317,13.982429,9.932085,5.7891436,4.32471,5.353586,5.7274113,7.2604365,9.499957,9.702303,8.968371,8.272165,8.848335,9.774324,7.9463544,8.31675,7.455923,7.226141,7.5382333,6.334448,5.0174866,4.3658648,4.040054,3.8617156,3.841138,4.2526884,4.139512,3.6627994,2.8739944,1.728512,1.8656956,1.9171394,1.9239986,1.9925903,2.2978237,2.2841053,2.5447538,2.6990852,2.5996273,2.3252604,2.7333813,2.551613,2.4247184,2.4830213,2.3389788,1.9548649,2.0989075,2.0440342,1.8965619,2.609916,3.3815732,3.199805,3.5976372,4.2835546,3.1449318,4.190956,5.2266912,5.2335505,5.0243454,7.2535777,5.4976287,7.9189177,6.790583,1.7902447,0.01371835,0.42183927,2.170929,2.4761622,1.0837497,0.24350071,0.5041494,0.47328308,0.31895164,0.16119061,0.06516216,0.14061308,0.11317638,0.0548734,0.006859175,0.006859175,0.037725464,0.15090185,0.33266997,0.48700142,0.44584638,0.432128,0.5624523,0.6310441,0.64133286,0.8265306,0.9877212,1.0117283,1.0494537,1.1351935,1.1763484,1.0940384,0.99801,1.0082988,1.0837497,1.0185875,0.881404,0.89855194,0.9431366,0.94999576,0.90884066,0.9774324,1.0631721,1.1283343,1.1626302,1.2106444,1.039165,0.9945804,1.0528834,1.1454822,1.1454822,0.9877212,1.0014396,1.0871792,1.1454822,1.0563129,1.155771,1.2380811,1.2003556,1.0494537,0.89169276,0.6790583,0.6276145,0.6756287,0.7373613,0.7133542,0.61389613,0.5555932,0.5418748,0.5761707,0.6276145,0.71678376,0.7956643,0.7956643,0.7407909,0.7579388,0.65162164,0.52815646,0.38754338,0.274367,0.2709374,0.3018037,0.3841138,0.39097297,0.33609957,0.3566771,0.31895164,0.32924038,0.34638834,0.37382504,0.47328308,0.5007198,0.42183927,0.3018037,0.18519773,0.10288762,0.06516216,0.048014224,0.05144381,0.0548734,0.044584636,0.07888051,0.09945804,0.10288762,0.08573969,0.044584636,0.037725464,0.030866288,0.044584636,0.082310095,0.12689474,0.1371835,0.17490897,0.25378948,0.37039545,0.5178677,0.6824879,0.90198153,1.1180456,1.2312219,1.0940384,1.2655178,1.2895249,1.2209331,1.1317638,1.1146159,1.0837497,1.1454822,1.2449403,1.3203912,1.313532,1.430138,1.5090185,1.5536032,1.5913286,1.6633499,1.5673214,1.4918705,1.4198492,1.3546871,1.3375391,1.3889829,1.4507155,1.4472859,1.3889829,1.3786942,1.2586586,1.2346514,1.2106444,1.155771,1.1008976,1.1180456,1.1523414,1.0837497,0.922559,0.7990939,0.8162418,0.805953,0.82996017,0.90884066,1.0220171,1.255229,1.5158776,1.7971039,1.9891608,1.9137098,1.587899,1.5227368,1.6221949,1.8588364,2.2806756,3.1723683,3.1792276,2.7779658,2.3835633,2.3801336,2.527606,2.6990852,3.1620796,4.197815,6.101236,9.595985,14.520873,19.490345,24.332924,30.070623,43.795834,50.55898,51.46439,48.854473,46.31315,0.2469303,0.28122616,0.36353627,0.45270553,0.6379033,1.1660597,1.6324836,1.8759843,2.335549,2.819121,2.5070283,1.9411465,1.9068506,2.2635276,2.8122618,3.2786856,3.2375305,3.0248961,2.633923,2.1846473,1.9308578,1.5741806,1.2003556,1.1729189,1.5193073,1.920569,2.0920484,2.0920484,1.9857311,1.8313997,1.6770682,1.7216529,1.6736387,1.5570327,1.4369972,1.4095604,2.1400626,3.5599117,5.422178,7.3873315,9.019815,8.179566,6.708273,5.9914894,6.046363,5.545643,3.642222,3.433017,5.0003386,6.9620624,6.468202,5.3673043,4.2835546,4.1326528,5.144381,6.835168,7.0786686,7.9189177,8.964942,10.63858,14.160767,18.825006,20.4472,21.177702,22.758743,26.510712,27.409264,27.60132,26.665043,24.281479,20.241425,16.105343,11.334786,6.9689217,3.8514268,2.644212,2.1846473,1.8519772,1.5810398,1.3615463,1.2312219,1.8245405,1.728512,1.529596,1.6667795,2.4452958,2.5927682,2.5721905,2.3972816,2.218943,2.3389788,2.3629858,2.177788,1.821111,1.4644338,1.4095604,1.0837497,0.8265306,0.6790583,0.67219913,0.82996017,0.9534253,1.0220171,1.155771,1.2929544,1.2209331,1.2072148,1.3478279,1.2929544,0.97400284,0.59331864,0.5521636,0.52472687,0.71678376,1.0940384,1.3684053,1.138623,1.0597426,1.1111864,1.1660597,0.980862,1.1934965,1.1111864,1.0323058,1.0597426,1.0940384,1.1797781,1.0631721,1.0117283,1.1146159,1.2826657,1.5536032,1.9102802,2.2155135,2.510458,3.0351849,2.9700227,2.603057,2.3081124,2.253239,2.4075704,2.6750782,3.3266997,4.976331,7.2707253,8.89635,9.849775,9.4862385,9.784613,11.430815,13.817808,15.837835,19.432043,23.842491,28.616478,33.599667,39.176178,39.423107,34.131256,24.936531,15.309678,10.573419,9.650859,8.076678,5.3227196,4.8014226,4.65395,4.2869844,4.290414,4.496189,3.974892,4.170378,5.3570156,6.4304767,6.8969,6.8626046,7.64798,7.4181976,7.6205435,8.608265,9.661148,10.515115,10.72775,11.965831,13.941273,14.4145565,15.313108,15.837835,16.492886,16.835844,15.453721,16.774113,17.312557,18.015623,19.092514,20.015072,21.109112,20.258574,19.888178,21.596113,26.174612,29.26467,29.806545,27.944279,26.35295,30.221525,32.635956,34.25472,31.740831,27.258362,28.486153,31.222963,31.198957,31.16809,32.409603,34.700565,36.607418,34.16898,29.391565,25.495554,26.915403,32.893173,43.034462,49.163136,51.738758,59.86688,125.03933,173.98297,176.43855,139.81743,109.21521,91.61457,66.02642,38.97726,17.995045,11.595435,7.3084507,7.099246,10.357354,16.2974,23.931662,12.439114,16.21509,16.828985,10.950673,10.31277,16.324837,9.163857,4.187526,5.2335505,4.619654,7.7440085,10.484249,10.398509,7.798882,5.7479887,5.518206,5.0174866,6.4304767,8.021805,4.139512,3.7931237,3.6147852,4.616225,6.917478,9.746887,15.337115,20.978786,25.063425,28.59247,35.16356,34.189556,27.059444,24.082563,24.61072,17.014183,14.754086,15.806969,17.902447,18.87302,16.636929,17.04162,16.108772,16.835844,19.099373,19.661825,23.550978,20.237995,16.602633,15.9578705,18.03963,14.466,14.7026415,19.006773,25.313786,29.237232,32.15581,35.966084,37.48196,38.66174,46.604664,74.055084,64.41451,44.831566,30.746252,25.886526,25.61559,27.206917,27.44013,25.039417,20.673553,17.230247,12.140739,8.210432,6.8454566,8.028665,8.553391,9.177576,10.2236,11.766914,13.646329,11.952112,10.374502,10.1652975,12.682614,19.363451,27.673342,28.952578,25.632736,19.658396,12.47341,11.677745,10.988399,15.899568,27.44356,42.20793,26.205479,13.505715,8.203573,9.997248,14.181344,13.457702,18.36544,24.476965,27.450418,23.03654,32.17296,42.64006,58.19324,86.96405,141.46362,107.10944,65.9784,32.306713,14.441993,14.808959,13.495427,13.214201,17.754974,26.918833,36.514816,29.76196,19.308577,13.070158,12.778643,13.992717,16.115631,17.521763,16.647217,14.339106,13.862392,15.0250225,21.153696,38.06156,62.308746,81.216064,50.233166,27.693918,17.412016,16.2974,14.321958,13.039291,10.425946,9.108984,10.213311,13.365103,13.416546,12.048141,11.238758,11.633161,12.545431,8.899779,6.5470824,6.334448,8.186425,11.101575,12.0309925,14.116182,14.836395,13.296511,10.233889,8.927217,8.224151,7.8949103,7.8194594,8.001227,8.704293,7.3530354,5.597087,4.787704,5.98463,4.746549,4.5270553,5.007198,5.188966,3.4192986,3.7005248,3.7862647,4.479041,6.2144127,9.067829,9.304471,8.97866,9.431366,10.81006,12.05157,14.29452,13.865822,11.513125,8.831187,8.2653055,8.179566,5.9297566,4.647091,4.9180284,4.8082814,5.1512403,5.1409516,6.39961,8.89635,10.971251,12.000127,12.953552,11.681175,9.112414,9.239308,15.971589,14.915276,10.405369,6.3207297,6.0566516,6.1904054,6.0737996,6.8454566,7.750868,6.1492505,7.2295704,7.1712675,8.086967,9.335337,7.5210853,6.927767,6.6533995,7.157549,7.970361,7.6651278,6.5710897,4.928317,3.5770597,2.9940298,3.2683969,3.9131594,3.673088,3.0283258,2.2566686,1.4335675,1.9514352,2.170929,2.1332035,2.1434922,2.760818,2.4315774,2.6956558,2.9665933,2.9734523,2.7299516,3.3266997,3.2443898,3.0557625,2.9494452,2.702515,1.8073926,1.8725548,1.9651536,1.8313997,1.9239986,3.3678548,3.566771,3.9680326,4.5167665,3.6525106,4.791134,6.6739774,6.2727156,4.8288593,7.8537555,6.1046658,6.869464,6.0326443,2.884283,0.106317215,0.034295876,0.8676856,1.8142518,1.9582944,0.2503599,0.4972902,0.51100856,0.3841138,0.20577525,0.058302987,0.0274367,0.006859175,0.0034295875,0.006859175,0.006859175,0.041155048,0.08916927,0.21263443,0.4046913,0.5727411,0.6310441,0.7613684,0.8265306,0.8265306,0.9294182,0.96371406,0.85396725,0.89512235,1.0734608,1.0734608,1.0460242,1.0563129,1.0563129,1.0425946,1.0563129,0.94656616,0.9774324,1.0323058,1.0323058,0.97057325,1.0323058,1.0528834,1.0906088,1.1729189,1.2860953,1.1111864,1.1146159,1.1626302,1.1832076,1.1454822,1.08032,1.1489118,1.214074,1.196926,1.0666018,1.2106444,1.2277923,1.1043272,0.89512235,0.72021335,0.61389613,0.6379033,0.72707254,0.7956643,0.7339317,0.64819205,0.5761707,0.52472687,0.51100856,0.5727411,0.7442205,0.8471081,0.8711152,0.84367853,0.823101,0.7133542,0.6379033,0.53844523,0.39440256,0.23664154,0.21263443,0.2503599,0.2709374,0.26064864,0.2709374,0.24007112,0.26064864,0.28465575,0.29837412,0.33266997,0.42869842,0.51100856,0.48014224,0.3566771,0.274367,0.17147937,0.12689474,0.09602845,0.06516216,0.05144381,0.06859175,0.09259886,0.106317215,0.10288762,0.08916927,0.05144381,0.034295876,0.030866288,0.037725464,0.061732575,0.058302987,0.08573969,0.12003556,0.16804978,0.26407823,0.3806842,0.58988905,0.7922347,0.922559,0.9362774,1.1729189,1.3066728,1.3203912,1.2655178,1.2586586,1.1694894,1.1660597,1.2106444,1.2723769,1.3238207,1.4610043,1.5055889,1.4610043,1.3821237,1.3649758,1.371835,1.3684053,1.3615463,1.3478279,1.3375391,1.3786942,1.4267083,1.4198492,1.3684053,1.3238207,1.2758065,1.2792361,1.214074,1.1008976,1.0940384,1.0666018,1.0597426,1.0425946,0.9877212,0.89169276,0.88826317,0.82996017,0.82996017,0.9259886,1.0768905,1.2895249,1.6153357,1.8862731,1.99602,1.9068506,1.6873571,1.5981878,1.7319417,2.085189,2.5721905,3.093488,3.2512488,3.0969174,2.8225505,2.7539587,2.9665933,3.1072063,3.4192986,4.1017866,5.31929,7.332458,11.2593355,16.918156,24.751333,35.85634,52.081715,57.750824,56.831696,53.2855,51.06313,0.11317638,0.10288762,0.20920484,0.34638834,0.6001778,1.2312219,1.4267083,1.4438564,1.8965619,2.620205,2.6819375,2.4967396,2.3458378,2.633923,3.3026927,3.8479972,3.9131594,3.7691166,3.3609958,2.8294096,2.5070283,1.8897027,1.4129901,1.3855534,1.7422304,2.061182,2.153781,1.903421,1.6530612,1.5433143,1.5227368,1.6427724,1.6907866,1.7353712,1.8519772,2.0989075,3.3747141,5.079219,6.8043017,8.333898,9.609704,8.621983,7.099246,6.0737996,5.597087,4.73969,4.046913,5.2266912,7.366754,8.47451,5.5147767,4.290414,4.012617,4.448175,5.518206,7.3084507,7.5245147,8.134981,9.328478,11.434244,14.932424,17.981327,17.672665,18.152807,21.472647,27.556736,32.94462,39.694046,42.921288,40.4074,32.58451,24.387796,17.569777,11.314209,6.108095,3.7382503,2.7916842,2.4075704,2.2978237,2.201795,1.8965619,2.1572106,2.153781,2.0749004,2.0508933,2.1640697,2.4624438,2.1915064,1.8279701,1.6153357,1.5810398,1.4918705,1.5021594,1.5398848,1.5981878,1.7182233,1.0871792,0.78537554,0.61389613,0.53501564,0.6756287,0.71678376,0.66876954,0.65505123,0.72707254,0.8779744,0.7990939,0.7956643,0.61046654,0.30523327,0.26407823,0.45613512,0.4046913,0.45956472,0.7476501,1.155771,1.1111864,1.0700313,1.1077567,1.2037852,1.2449403,1.4267083,1.4404267,1.471293,1.5124481,1.3546871,1.3443983,1.2758065,1.3855534,1.6427724,1.7490896,1.6770682,1.8245405,1.920569,2.0337453,2.5893385,2.9288676,2.7745364,2.8568463,3.2032347,3.1586502,2.9185789,3.4124396,5.586798,8.930646,11.465111,11.852654,11.7086115,12.185325,13.920695,17.062197,18.173384,18.44775,18.214539,18.159666,19.339443,22.998814,22.748453,18.934752,12.956982,7.2638664,5.7479887,5.967482,6.166398,6.101236,7.0478024,6.7871537,6.23156,6.125243,6.3824625,6.1046658,5.528495,7.0546613,7.5588107,6.9552035,8.210432,8.903209,9.355915,10.436234,12.024134,13.001566,15.374841,16.280252,16.674654,17.027903,17.326277,18.20425,19.521212,21.654415,23.156574,20.735287,21.170843,20.087093,18.313997,16.684942,16.03675,18.70154,17.556059,16.21166,17.439453,23.156574,28.585611,30.50618,28.980015,26.496992,27.947708,28.815393,32.601658,30.375856,24.03455,26.301506,29.981453,30.056904,29.154922,28.832542,29.600769,31.126936,29.67622,27.200058,25.643026,26.963417,30.780548,38.1473,43.425438,46.508636,52.829365,99.132225,137.61563,142.98636,119.43539,100.634384,83.18465,58.460747,34.035225,15.707511,7.514226,6.3378778,6.279575,10.55284,19.263992,29.42929,11.091286,14.205351,15.004445,8.930646,10.6317215,17.892159,9.674867,3.6765177,4.540774,3.8479972,6.0737996,8.2310095,8.279024,6.5196457,5.6039457,5.6313825,5.754848,7.534804,9.043822,4.856296,4.822,4.1120753,5.4907694,9.836057,16.153357,22.875349,29.028028,32.622234,34.24443,37.046402,31.305275,21.44864,15.649208,15.9921665,18.482046,14.3974085,11.80464,12.264205,15.584045,19.792149,20.316875,19.493774,19.325726,20.714708,23.44123,28.496443,18.574646,12.05157,14.733508,19.847023,13.618892,14.3974085,22.175713,31.535057,31.641375,33.561943,34.59082,37.289906,43.524895,54.44813,86.07578,74.35689,49.53353,30.228384,23.417223,25.783638,25.996273,22.847912,17.703531,14.517444,14.647768,10.882081,7.781734,7.366754,9.108984,7.56567,8.611694,11.351934,13.858963,13.166186,10.9541025,9.403929,9.1810055,11.509696,18.163095,25.821363,25.711617,23.153145,20.721567,18.279701,15.285671,10.621432,10.971251,17.103354,23.852781,15.762384,11.516555,10.909517,12.607163,14.174485,15.151917,20.834743,26.215767,28.304386,26.116308,34.67999,46.683544,67.27821,95.59632,124.77868,86.298706,51.491825,25.111439,10.978109,11.955542,14.318527,21.225718,29.419,36.89207,42.89728,28.280378,17.034761,13.54687,16.235666,17.53891,16.983316,17.000465,16.095055,15.268523,17.998474,20.556948,31.562494,53.78965,77.69388,81.428696,44.05648,23.76361,15.388559,13.694343,13.38911,12.233338,9.647429,9.760606,12.912396,15.6526375,14.232788,13.872682,13.88983,13.738928,13.032433,10.593996,8.625413,7.891481,8.875772,11.790922,11.485688,12.164746,12.747777,12.511135,11.084427,11.238758,11.626302,11.159878,9.863494,8.872343,10.323058,8.042382,6.0978065,5.960623,6.5196457,5.055212,4.3452873,4.6573796,5.1683884,3.9611735,4.016047,3.6044965,4.033195,5.518206,7.181556,9.218731,9.592556,10.405369,11.4376745,10.14129,11.814929,12.590015,11.602294,9.760606,9.740028,9.297611,6.2727156,4.0709205,3.542764,2.959734,5.4084597,4.8014226,4.5682106,6.012067,8.309891,9.839486,10.569988,10.7757635,10.882081,11.482259,12.6757555,11.101575,8.683716,7.449064,9.523964,10.340206,8.443645,7.2432885,6.842027,4.033195,5.7891436,6.3481665,7.040943,7.764586,6.9826403,5.885172,5.953764,6.9963584,8.100685,7.6342616,8.100685,6.39961,4.098357,2.6373527,3.3266997,4.0434837,3.2958336,2.1915064,1.4267083,1.2860953,1.7765263,2.1469216,2.2463799,2.3629858,3.2478194,2.3972816,2.4590142,2.860276,3.1483612,2.9803114,3.3712845,3.3884325,3.3369887,3.3061223,3.1792276,1.728512,1.6359133,1.9308578,1.9891608,1.5501735,3.0248961,3.6593697,4.2766957,4.8082814,4.280125,5.2266912,7.281014,6.9723516,5.435896,8.405919,8.152129,6.7974424,5.381023,3.683377,0.23321195,0.048014224,0.25721905,1.4027013,2.3595562,0.32238123,0.31895164,0.3841138,0.37725464,0.25721905,0.06859175,0.01371835,0.0,0.0034295875,0.01371835,0.01371835,0.048014224,0.07888051,0.1371835,0.2777966,0.59331864,0.7613684,0.83338976,0.91227025,1.0151579,1.08032,0.96371406,0.7888051,0.83338976,1.0357354,1.0185875,1.0048691,1.1111864,1.1420527,1.0906088,1.1249046,1.0906088,1.1420527,1.214074,1.2449403,1.1626302,1.1900668,1.1351935,1.1146159,1.1797781,1.3169615,1.2346514,1.3375391,1.3649758,1.2517995,1.155771,1.2655178,1.2758065,1.2620882,1.2449403,1.1626302,1.2037852,1.1146159,0.922559,0.72707254,0.6893471,0.72021335,0.7407909,0.7682276,0.78537554,0.72364295,0.6756287,0.6173257,0.5727411,0.5658819,0.6344737,0.72707254,0.764798,0.83338976,0.922559,0.9328478,0.77165717,0.65848076,0.6173257,0.58645946,0.4115505,0.3018037,0.2503599,0.24007112,0.23664154,0.18519773,0.13032432,0.13032432,0.16119061,0.19548649,0.21263443,0.34638834,0.52472687,0.5521636,0.44927597,0.45270553,0.34295875,0.2709374,0.19891608,0.13032432,0.09602845,0.07888051,0.07888051,0.09259886,0.11317638,0.15433143,0.08573969,0.058302987,0.041155048,0.020577524,0.020577524,0.0274367,0.058302987,0.08573969,0.1097468,0.14061308,0.16119061,0.2503599,0.41840968,0.64476246,0.8745448,1.0940384,1.2723769,1.371835,1.4335675,1.5638919,1.4781522,1.3512574,1.2998136,1.3581166,1.4541451,1.5398848,1.5638919,1.4850113,1.3341095,1.2277923,1.2312219,1.2483698,1.2758065,1.3066728,1.3478279,1.4198492,1.3855534,1.3169615,1.2655178,1.2449403,1.3066728,1.2689474,1.1729189,1.1008976,1.1660597,1.0666018,1.0563129,1.1077567,1.1592005,1.1249046,1.1523414,1.0563129,1.0151579,1.1077567,1.2963841,1.4815818,1.8416885,2.0097382,1.937717,1.8828435,1.978872,1.9239986,1.9994495,2.301253,2.7128036,2.6716487,2.8225505,3.000889,3.0969174,3.0523329,3.4227283,3.806842,4.2423997,4.8494368,5.8062916,6.6533995,8.786603,13.783512,22.762173,36.381065,47.753574,51.38208,51.560417,51.649586,54.05716,0.01371835,0.06516216,0.14061308,0.21263443,0.31552204,0.53501564,0.7305021,0.7682276,0.9568549,1.3649758,1.8142518,2.352697,2.551613,2.935727,3.566771,4.0434837,3.690236,3.2718265,3.059192,3.093488,3.2032347,2.6545007,2.4075704,2.4555845,2.620205,2.5481834,2.3767042,1.9582944,1.6599203,1.5947582,1.6324836,1.646202,1.7388009,1.9239986,2.318401,3.1723683,5.4084597,6.725421,7.5759587,8.546532,10.39165,9.8429165,8.241299,7.140401,6.776865,6.0566516,6.39961,9.047252,9.798331,7.723431,5.171818,4.122364,3.724532,4.389872,6.1492505,8.652849,10.22703,10.024684,10.024684,11.842365,16.739817,18.948471,17.2131,16.822126,19.696121,24.384367,31.781986,43.106483,50.929375,51.848503,46.477768,34.24786,23.461807,15.134769,9.242738,4.715683,3.1037767,2.7745364,2.901431,3.018037,3.0043187,3.2512488,3.1826572,3.0489032,2.8225505,2.2120838,1.845118,1.4267083,1.138623,0.9945804,0.823101,1.0185875,1.1489118,1.3443983,1.4987297,1.2655178,0.8025235,0.65162164,0.5212973,0.4046913,0.5658819,0.5761707,0.66191036,0.8093826,0.91569984,0.7922347,0.53844523,0.37382504,0.35324752,0.48357183,0.70306545,0.5555932,0.5555932,0.6824879,0.88826317,1.0837497,0.8505377,0.84024894,1.1008976,1.488441,1.6496316,1.587899,1.5433143,1.5741806,1.6736387,1.7696671,1.7593783,2.0920484,2.3732746,2.3972816,2.1503513,2.07833,2.1332035,2.4624438,3.0043187,3.4947495,3.6147852,3.4913201,3.6970954,4.1120753,3.8925817,2.9391565,3.1963756,5.055212,7.6685576,8.927217,9.438225,10.940384,12.679185,14.143619,15.059319,12.80265,9.510246,6.776865,5.425607,5.5079174,5.3878818,5.0277753,4.2286816,3.3198407,3.175798,3.6010668,4.4687524,6.121814,7.73029,7.2775846,6.8626046,7.380472,8.303031,8.848335,7.9943686,8.351046,9.3079,9.650859,9.184435,8.759167,11.115293,12.47341,13.234778,14.05102,15.806969,18.787281,21.352612,22.885637,23.502962,24.079134,23.626429,24.308916,27.1006,30.221525,29.158352,28.01287,25.4544,21.328604,17.305698,16.890718,17.024471,16.208231,16.060759,17.724108,21.849901,26.246634,24.799347,22.309467,21.294308,22.004232,22.041958,27.477856,29.26467,26.545008,26.641035,29.960876,29.281818,26.661613,25.135447,28.68507,33.239563,30.194088,25.543568,24.363789,30.821703,30.125496,33.229275,37.375645,42.74638,52.476116,93.27106,132.5364,137.43729,110.30239,88.62397,74.07223,53.70734,33.08866,16.462019,6.7459984,4.7808447,4.32471,7.98065,15.6697855,24.645016,7.0786686,9.431366,11.842365,9.119273,10.741467,14.514014,9.873782,6.39961,6.108095,3.433017,4.9351764,6.619104,7.051232,6.543653,7.140401,6.15268,6.4544835,7.06495,7.15069,6.025785,5.662249,4.7088237,4.3658648,6.728851,14.784951,21.647556,21.575535,20.550089,20.419764,18.907316,13.828096,12.9707,13.886399,13.965281,10.436234,10.864933,11.31078,12.205902,13.96871,16.983316,17.851004,19.339443,19.510923,19.253704,22.292318,25.60187,16.925014,10.484249,13.258785,24.963966,16.578627,17.62122,29.120626,40.39368,29.052036,32.26213,37.790623,44.186806,53.498135,71.25654,105.521545,89.81061,56.10462,28.43471,22.841053,22.868488,23.94538,22.2786,17.87501,14.5414505,14.321958,10.100135,7.366754,7.2158523,6.3618846,6.509357,10.261326,13.735497,15.193072,15.0456,10.333347,8.1212635,8.968371,12.72034,18.492336,20.985645,22.851341,27.6802,32.416462,27.374968,19.829874,11.499407,8.22758,11.266195,17.274832,12.072148,13.509145,18.080786,20.069946,11.550851,15.700651,20.601532,24.92967,28.18092,30.670801,37.15272,50.308617,72.77585,95.65119,98.49775,67.782364,33.68541,14.359683,12.336226,14.496866,25.481834,38.123295,47.249428,50.490387,48.292023,22.412354,13.924125,15.608052,19.871029,18.722118,13.852104,12.524854,12.689473,13.910407,17.364002,26.092302,44.96189,62.706577,68.523155,52.095432,28.571894,18.62609,14.243076,11.873232,12.435684,11.64345,9.914937,10.844356,13.540011,12.648318,11.012405,14.140189,15.659496,13.80066,11.382801,11.701753,11.71547,11.190743,10.484249,10.5597,12.096155,11.760056,12.13731,12.816368,10.374502,14.562028,14.685493,12.579727,10.007536,8.652849,7.699424,6.0154963,5.3261495,5.785714,5.9812007,7.8983397,7.130112,6.252138,5.768566,4.1189346,4.4996185,3.8514268,3.724532,4.6779575,6.3035817,8.683716,9.441654,9.016385,8.186425,8.1041155,9.006097,10.569988,10.511685,9.057541,8.9100685,9.668007,8.988949,7.8777623,6.427047,3.8137012,4.1943855,5.504488,6.756287,6.636252,3.525616,4.8322887,4.773986,8.038953,13.2862215,13.152468,11.2250395,8.958082,7.582818,8.327039,12.404818,11.502836,8.759167,7.349606,7.257007,5.2781353,3.7039545,4.280125,5.422178,6.6533995,8.604835,9.764035,7.7680154,6.5333643,6.81802,6.193835,6.7185616,7.2364297,5.15467,2.0097382,3.450165,2.644212,1.7559488,1.3581166,1.5913286,2.1674993,1.6290541,1.5673214,1.5433143,1.5981878,2.2566686,2.1126258,2.194936,2.3458378,2.49331,2.6407824,3.3609958,3.3369887,3.2272418,3.350707,3.6936657,2.534465,1.9137098,1.7490896,1.9651536,2.503599,3.1380725,3.707384,4.214963,4.523626,4.3624353,4.461893,5.7754254,6.385892,6.169828,6.8043017,11.897239,11.547421,8.244728,3.9680326,0.18176813,0.037725464,0.037725464,0.84367853,1.6907866,0.39783216,0.17833854,0.30523327,0.37725464,0.2503599,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.024007112,0.11317638,0.17833854,0.22635277,0.33609957,0.5555932,0.72021335,0.7613684,0.72707254,0.7613684,0.7133542,0.78537554,0.77851635,0.70306545,0.7613684,0.83681935,1.039165,1.2689474,1.4061309,1.2963841,1.4198492,1.4129901,1.3581166,1.2963841,1.2346514,1.1763484,1.2586586,1.3272504,1.3649758,1.5090185,1.3032433,1.3615463,1.4575747,1.5090185,1.5707511,1.7182233,1.488441,1.3615463,1.4198492,1.3581166,1.0768905,0.9877212,0.90884066,0.8128122,0.823101,0.922559,0.864256,0.8196714,0.8093826,0.6859175,0.6379033,0.6241849,0.59674823,0.548734,0.548734,0.6241849,0.6036074,0.6276145,0.72707254,0.823101,0.7510797,0.61389613,0.58302987,0.66876954,0.71678376,0.607037,0.42526886,0.2709374,0.18519773,0.1371835,0.09945804,0.09259886,0.12346515,0.17833854,0.21263443,0.29837412,0.34638834,0.3841138,0.41498008,0.42869842,0.4629943,0.40126175,0.31552204,0.25378948,0.22978236,0.20577525,0.14404267,0.09945804,0.106317215,0.16804978,0.106317215,0.082310095,0.06516216,0.044584636,0.044584636,0.034295876,0.058302987,0.07545093,0.07888051,0.09259886,0.09259886,0.1097468,0.17147937,0.31552204,0.59674823,0.8162418,0.9328478,1.0666018,1.2689474,1.5261664,1.7936742,1.6873571,1.5090185,1.4438564,1.5398848,1.6153357,1.7250825,1.7902447,1.7525192,1.5570327,1.4335675,1.5227368,1.6016173,1.605047,1.6187652,1.6290541,1.4404267,1.2517995,1.1729189,1.2209331,1.4267083,1.3992717,1.3169615,1.2998136,1.371835,1.313532,1.3066728,1.3169615,1.3203912,1.2963841,1.3821237,1.4027013,1.4232788,1.4541451,1.4815818,1.529596,1.8142518,2.0714707,2.1743584,2.1503513,2.201795,2.1297739,2.0817597,2.1160555,2.2120838,2.0063086,1.9891608,2.1469216,2.428148,2.7470996,3.724532,4.6916757,5.360445,5.7822843,6.3310184,6.8454566,7.870903,10.789482,16.21509,24.003683,29.59391,35.211575,40.095306,45.66839,55.55589,0.05144381,0.061732575,0.061732575,0.116605975,0.23321195,0.37382504,0.4355576,0.5041494,0.607037,0.7922347,1.155771,2.037175,2.4212887,2.719663,3.0454736,3.2375305,2.668219,2.1743584,2.0303159,2.2978237,2.8259802,2.8225505,2.5378947,2.3629858,2.4007113,2.4761622,2.2463799,2.061182,2.0303159,2.1126258,2.1194851,2.1023371,2.177788,2.6476414,3.806842,5.919468,8.203573,8.772884,9.033533,9.791472,11.231899,10.868362,9.89093,9.081548,8.597976,7.9737906,9.321619,11.46854,11.2421875,8.608265,6.660259,5.0277753,4.413879,4.897451,6.5196457,9.273604,11.159878,11.249047,11.4754,13.656617,19.510923,20.858751,18.893597,17.971039,19.03421,19.61038,22.789608,28.650774,34.210136,38.209034,41.120754,37.66716,28.959436,19.761284,12.713481,8.340756,5.919468,4.557922,3.858286,3.6593697,4.057202,4.3487167,4.4550343,4.4584637,4.249259,3.532475,3.3884325,2.5996273,1.5981878,0.77851635,0.48357183,0.58988905,0.72707254,0.89855194,1.1729189,1.6804979,1.3649758,0.99801,0.6893471,0.5418748,0.66191036,0.77165717,0.7339317,0.6756287,0.59331864,0.35324752,0.23321195,0.20577525,0.25721905,0.4081209,0.7133542,0.66533995,0.72707254,0.8676856,0.980862,0.864256,0.77851635,0.97057325,1.3032433,1.6153357,1.7456601,1.762808,1.6221949,1.5707511,1.6153357,1.5364552,1.9651536,2.5413244,2.668219,2.4212887,2.5790498,2.2120838,1.9514352,1.9342873,2.2463799,2.9220085,3.100347,2.7779658,2.5619018,2.6304936,2.74367,2.6613598,2.901431,3.5359046,4.3521466,4.835718,4.773986,5.363875,6.0635104,6.7494283,7.7131424,6.848886,5.627953,3.7485392,1.8862731,1.6873571,1.4404267,1.4198492,1.6324836,2.0817597,2.784825,4.0709205,5.137522,5.720552,5.9297566,6.2418494,6.7357097,8.937505,10.933525,11.399949,9.619993,9.191295,9.14328,8.556821,7.3118806,6.0840883,7.8949103,9.3079,11.276484,14.212211,17.991615,20.131678,20.635828,20.831314,21.328604,22.038528,22.642136,24.747904,27.872257,30.818274,31.648233,31.497332,28.01973,23.297188,19.483486,18.79414,20.12139,18.728977,18.54378,20.70785,23.585274,24.03455,23.081123,23.760181,25.622448,24.737614,23.290329,23.722456,23.585274,22.86163,23.955667,26.671902,27.062874,24.679312,21.997374,24.425522,27.594461,25.571005,22.148275,20.601532,23.671013,24.408375,26.407824,29.960876,35.118977,41.672916,71.805275,110.42586,122.31624,102.791595,77.72474,63.807476,45.140232,28.393555,16.341984,7.8537555,5.8508763,5.336438,5.446185,8.1212635,18.087645,6.4304767,6.6876955,9.56512,10.508256,9.729739,13.248496,10.950673,8.577398,7.3564653,4.0194764,4.846007,5.07236,5.2301207,5.7308407,6.8969,7.3530354,7.0272245,7.1369715,7.5931067,7.0272245,5.3158607,4.0846386,3.5873485,4.7191124,9.0369625,13.231348,14.280802,12.576297,10.069269,10.264755,9.297611,7.5245147,6.9723516,7.3839016,6.2384195,7.06495,8.886061,11.588576,14.987297,18.800999,22.587263,28.92857,29.250952,23.931662,22.292318,20.21056,17.439453,15.484588,18.924463,35.376194,20.066517,16.427725,19.696121,25.317215,28.966295,37.927807,47.897617,57.36328,68.13561,85.32127,105.12372,93.71348,61.94864,30.207806,28.34897,25.365229,23.20802,20.728426,18.279701,17.689812,19.03421,13.21763,8.176137,6.5230756,5.56965,9.191295,13.193623,15.656067,15.258235,11.273054,8.601405,8.776315,11.787492,16.064188,18.468328,16.252815,24.171732,37.622574,44.22453,23.835632,14.033872,8.155559,10.443094,17.398296,17.809847,18.430603,17.161655,15.6252,14.448852,13.272504,17.960749,22.628418,27.001143,30.869717,34.110676,40.1639,51.241467,62.463078,68.862686,65.42967,41.559742,23.725885,15.4742985,16.317978,21.723007,35.383053,43.723812,49.365482,50.600132,41.360825,17.473747,16.304258,21.884197,24.0174,18.269413,11.026124,9.2153015,11.1393,14.644339,17.134218,29.875137,43.82327,48.90249,42.585186,29.916292,20.402617,15.865272,13.251926,11.454823,11.314209,10.762046,11.331357,12.322508,12.394529,9.547972,10.052121,12.343085,13.289652,12.634601,12.9809885,13.7697935,11.763485,9.407358,8.14527,8.423067,9.414218,9.496528,8.927217,8.604835,10.069269,14.033872,12.504276,10.978109,10.957532,9.932085,5.9434752,4.232111,4.338428,5.188966,5.0895076,5.552502,5.456474,5.312431,5.3227196,5.363875,6.6431108,5.0929375,4.0057583,4.7671266,6.852316,8.381912,7.98408,7.2158523,7.8126,11.691463,10.278474,10.72775,11.039842,10.597425,10.168727,10.738038,9.242738,7.0375133,5.144381,4.2423997,5.7925735,7.8366075,8.210432,6.715132,5.137522,6.7459984,7.4524937,10.583707,14.802099,14.092175,10.278474,7.7542973,6.557371,7.3358874,11.355364,10.549411,8.652849,7.1232533,6.0840883,4.3041325,3.7039545,4.372724,5.470192,6.433906,6.9826403,8.172707,7.2775846,6.4990683,6.7940125,7.891481,6.9723516,6.416758,5.7891436,5.038064,4.4859004,3.875434,2.2292318,1.3958421,1.6530612,1.728512,1.5913286,1.5707511,1.670209,1.8999915,2.294394,2.020027,2.2258022,2.5447538,2.7470996,2.7368107,3.0077481,3.292404,3.3129816,3.117495,3.069481,2.4487255,2.4075704,2.428148,2.417859,2.7230926,3.0626216,3.8479972,4.465323,4.804852,5.2438393,5.2918534,5.007198,5.5730796,6.526505,5.754848,14.459141,18.478617,15.501736,8.028665,3.357566,0.69963586,0.020577524,0.4355576,1.3341095,2.3732746,0.5727411,0.25378948,0.37725464,0.34981793,0.041155048,0.006859175,0.0,0.0,0.006859175,0.037725464,0.05144381,0.1371835,0.19891608,0.22978236,0.29837412,0.5761707,0.6310441,0.65505123,0.7099246,0.72707254,0.805953,0.84024894,0.823101,0.78194594,0.77508676,0.91569984,1.097468,1.3649758,1.6016173,1.5398848,1.5947582,1.5055889,1.4164196,1.3889829,1.4061309,1.4335675,1.4747226,1.4781522,1.4404267,1.3992717,1.3409687,1.3546871,1.471293,1.6256244,1.6564908,1.7147937,1.6256244,1.5604624,1.4953002,1.2003556,0.88826317,0.7407909,0.64476246,0.5624523,0.5555932,0.70306545,0.7373613,0.7133542,0.67219913,0.6379033,0.6001778,0.6241849,0.6241849,0.61389613,0.72021335,0.72364295,0.6379033,0.58302987,0.6207553,0.7373613,0.6756287,0.66533995,0.70649505,0.78537554,0.864256,0.7442205,0.52815646,0.3566771,0.26407823,0.18519773,0.14061308,0.106317215,0.09259886,0.10288762,0.12689474,0.22292319,0.32581082,0.38754338,0.39440256,0.37725464,0.36696586,0.33952916,0.34981793,0.39097297,0.42526886,0.33952916,0.29494452,0.2503599,0.20234565,0.15433143,0.13375391,0.12689474,0.10288762,0.06859175,0.06859175,0.06859175,0.058302987,0.058302987,0.06859175,0.07888051,0.07888051,0.082310095,0.106317215,0.16462019,0.29151493,0.4115505,0.5796003,0.77851635,1.0048691,1.2689474,1.4507155,1.4472859,1.4644338,1.5741806,1.7010754,1.6084765,1.6084765,1.6221949,1.5981878,1.5193073,1.5536032,1.6359133,1.6290541,1.529596,1.4815818,1.4164196,1.3409687,1.3066728,1.3341095,1.3924125,1.5193073,1.5501735,1.5364552,1.4815818,1.3615463,1.2723769,1.2655178,1.2483698,1.2106444,1.2243627,1.3684053,1.5364552,1.6873571,1.7902447,1.8348293,1.8725548,1.9445761,2.0749004,2.1846473,2.1023371,2.0646117,2.0886188,2.1023371,2.061182,1.9445761,1.786815,1.8108221,1.937717,2.1743584,2.6476414,3.5290456,4.331569,5.3432975,6.368744,6.7219915,6.824879,7.6376915,9.458802,12.020704,14.507155,17.71382,22.436361,29.501312,41.508297,62.833473,0.034295876,0.034295876,0.030866288,0.08573969,0.20234565,0.34638834,0.42869842,0.5212973,0.5658819,0.6036074,0.7888051,1.5055889,2.0028791,2.2600982,2.3218307,2.3149714,2.0268862,1.762808,1.7147937,1.9685832,2.503599,2.884283,2.8705647,2.836269,2.867135,2.750529,2.3801336,2.301253,2.411,2.6133456,2.819121,2.7162333,3.2135234,4.705394,6.9689217,9.170717,9.414218,9.218731,9.585697,10.72089,12.010415,11.180455,10.39165,9.860064,9.668007,9.770895,11.567999,12.7272,11.612583,8.772884,6.9346256,5.90575,5.751418,6.334448,7.6616983,9.897789,10.593996,11.125582,12.432255,15.450292,21.109112,22.61127,20.189981,17.741257,16.973028,17.391438,18.533491,21.482935,24.679312,27.93742,32.457615,38.274197,36.796043,29.51846,20.104242,14.411126,9.434795,6.773435,5.3878818,4.6402316,4.3007026,4.297273,4.2938433,4.180667,3.8925817,3.4021509,3.8377085,3.8720043,3.2546785,2.1023371,0.89855194,0.6036074,0.5624523,0.66533995,0.9328478,1.5090185,1.5673214,1.2929544,0.9328478,0.67219913,0.65848076,0.69963586,0.5796003,0.48014224,0.42526886,0.28122616,0.18862732,0.20920484,0.24007112,0.274367,0.4046913,0.5212973,0.97057325,1.2517995,1.1626302,0.83681935,0.91912943,0.99801,1.1694894,1.3958421,1.4953002,1.4232788,1.371835,1.4164196,1.5090185,1.4987297,2.020027,2.2155135,1.9823016,1.6667795,2.054323,2.170929,2.0268862,2.0474637,2.417859,3.0900583,2.6990852,2.393852,2.3492675,2.510458,2.603057,2.6647894,3.0557625,3.3712845,3.3850029,3.0626216,2.6304936,2.8019729,3.000889,3.0420442,3.117495,2.644212,2.2806756,1.5433143,0.65848076,0.58645946,0.5624523,0.823101,1.4369972,2.270387,2.9974594,3.333559,3.6936657,4.297273,5.137522,5.9914894,6.3447366,8.203573,9.126132,8.529384,7.671987,6.4990683,5.8405876,5.3707337,5.0655007,5.195825,7.016936,8.899779,12.30193,16.835844,20.27915,19.70298,19.569225,19.61724,20.12139,21.915064,22.079683,24.720467,28.17749,31.133795,32.59137,32.557076,29.034887,24.754763,22.306036,24.134007,25.406384,24.555847,24.43238,25.063425,23.677872,22.196291,21.980227,22.878778,24.538698,26.428402,26.037428,24.963966,24.134007,23.873358,23.897366,24.871368,24.634727,22.844482,20.992504,22.408924,22.724447,21.596113,20.53294,20.059656,19.709839,19.236557,20.145397,22.234016,26.047716,32.893173,53.021423,82.98916,101.989075,99.53006,75.44406,57.404434,40.527435,26.531288,16.064188,8.7283,6.2658563,5.1855364,4.4413157,6.6636887,18.12537,8.7283,6.433906,8.930646,12.212761,10.583707,14.46943,13.680624,10.323058,6.475061,4.1943855,4.389872,4.6916757,4.73969,4.8185706,5.874883,7.8194594,7.7680154,7.380472,7.1712675,6.5196457,4.9351764,3.5839188,3.0111778,4.0537724,7.846896,11.862943,16.602633,16.228807,11.619442,10.343636,9.235879,7.8503256,6.6876955,5.9297566,5.4153185,7.016936,9.942374,14.29452,19.099373,22.333473,28.534168,34.9132,35.650562,31.102928,27.813953,21.513802,17.672665,16.187653,18.30028,26.610168,20.049368,19.353163,21.4555,25.114868,30.9143,38.119865,48.63841,59.03006,70.128204,87.02578,93.37395,81.16119,59.287277,38.555424,31.67567,27.381826,23.585274,21.493225,21.20514,21.69214,20.728426,15.556609,9.619993,6.025785,7.5416627,13.313659,17.686382,17.737827,14.04759,10.686595,10.569988,13.347955,15.522313,16.448301,18.362011,14.654627,21.52066,36.607418,45.538063,21.915064,10.583707,8.97866,17.082775,26.709627,21.486366,17.46003,13.564018,11.451392,11.616013,13.38225,15.947581,18.787281,22.734735,26.980564,29.076042,34.700565,43.686085,47.523792,44.111355,37.7529,26.706198,21.301168,19.250275,20.433481,26.887966,35.89749,42.413708,49.331184,51.78334,37.173298,23.091412,22.518671,24.590141,23.907654,20.512363,14.102464,10.528833,9.764035,11.348505,14.393978,24.987974,32.317,32.34101,26.208908,20.248285,15.758954,13.876111,12.641459,11.533703,11.434244,13.077017,13.697772,12.435684,9.904649,8.207003,12.672326,14.21564,14.448852,15.145059,18.224829,16.307688,11.958971,8.594546,7.31531,6.927767,7.466212,7.1129646,6.166398,5.8680243,8.4093485,13.203912,12.792361,12.144169,12.346515,10.63858,5.9126086,4.105216,4.232111,4.8494368,4.0709205,5.305572,5.689686,6.307011,7.1026754,6.883182,7.610255,5.5559316,4.1360826,4.6848164,6.447624,7.058091,6.0395036,5.761707,7.0958166,9.403929,9.287323,10.14129,10.789482,10.813489,10.556271,9.887501,7.7680154,6.392751,6.3173003,6.464772,7.6925645,7.133542,5.9297566,5.020916,5.164959,6.5024977,7.4696417,10.203023,13.341095,12.003556,7.747438,6.883182,6.893471,6.790583,7.1026754,5.9983487,5.360445,5.0620713,4.976331,5.0003386,4.7499785,4.6848164,4.3692946,3.923448,4.033195,5.6519604,7.4696417,7.390761,6.217842,7.658269,8.937505,7.9086285,6.4819202,5.6313825,5.3878818,5.6005163,4.588788,3.5564823,2.8259802,1.8176813,1.5261664,1.5501735,1.704505,1.8725548,2.0097382,1.7936742,2.1229146,2.527606,2.7333813,2.6716487,2.7573884,3.3987212,3.6113555,3.2718265,3.1346428,3.0283258,3.0248961,2.9803114,2.9460156,3.199805,3.275256,4.245829,4.897451,5.144381,6.029215,5.7136927,4.7431192,5.3741636,6.728851,4.7774153,10.97468,15.347404,13.29994,7.829748,9.534253,1.9514352,0.034295876,0.24007112,1.1180456,3.2889743,1.0185875,0.31895164,0.31552204,0.3806842,0.09945804,0.0274367,0.0034295875,0.0034295875,0.017147938,0.044584636,0.08573969,0.17490897,0.23664154,0.26750782,0.33609957,0.5178677,0.5624523,0.58302987,0.67219913,0.881404,0.84367853,0.8471081,0.84024894,0.83681935,0.90541106,1.0494537,1.1900668,1.3855534,1.5707511,1.5638919,1.6084765,1.5330256,1.3889829,1.2929544,1.4404267,1.4747226,1.5124481,1.488441,1.4198492,1.3992717,1.4129901,1.3992717,1.4987297,1.6599203,1.6324836,1.6324836,1.6084765,1.5090185,1.3032433,0.94999576,0.70649505,0.5796003,0.5144381,0.47328308,0.42526886,0.5521636,0.6036074,0.58645946,0.53501564,0.50757897,0.47671264,0.53844523,0.58645946,0.61389613,0.6893471,0.7442205,0.6962063,0.65505123,0.67219913,0.7339317,0.6962063,0.66876954,0.66191036,0.6859175,0.72707254,0.66876954,0.52815646,0.4115505,0.33609957,0.23664154,0.22292319,0.18176813,0.13032432,0.09602845,0.106317215,0.18862732,0.30866286,0.37725464,0.37725464,0.32924038,0.33609957,0.34981793,0.37039545,0.39783216,0.4081209,0.39097297,0.40126175,0.4081209,0.3841138,0.31895164,0.2469303,0.2194936,0.20577525,0.18519773,0.14061308,0.1097468,0.07888051,0.061732575,0.061732575,0.058302987,0.058302987,0.05144381,0.058302987,0.082310095,0.13032432,0.19891608,0.30523327,0.432128,0.5796003,0.77508676,1.0082988,1.1111864,1.2415106,1.4335675,1.611906,1.5193073,1.4678634,1.4369972,1.4061309,1.371835,1.4404267,1.4815818,1.4575747,1.3855534,1.3306799,1.3478279,1.3752645,1.430138,1.4815818,1.4267083,1.4918705,1.4987297,1.4472859,1.371835,1.3409687,1.3581166,1.4164196,1.4369972,1.430138,1.4610043,1.5981878,1.7765263,1.9548649,2.0989075,2.170929,2.1846473,2.1160555,2.085189,2.1023371,2.0646117,2.0680413,2.1160555,2.1915064,2.2258022,2.1160555,1.937717,1.9308578,2.0337453,2.2635276,2.6887965,3.3678548,3.981751,4.7191124,5.5662203,6.327589,6.691125,7.421627,8.237869,8.97523,9.585697,11.495977,14.438563,19.843594,30.125496,48.71386,0.010288762,0.034295876,0.10288762,0.17833854,0.2503599,0.3566771,0.490431,0.5555932,0.5590228,0.548734,0.61389613,1.0220171,1.4232788,1.6804979,1.7765263,1.7936742,1.8554068,1.8931323,1.937717,2.0406046,2.301253,2.5824795,2.668219,2.836269,3.07634,3.0866287,3.0111778,3.1586502,3.3026927,3.350707,3.333559,3.275256,4.3795834,6.3378778,8.443645,9.585697,8.927217,8.920357,9.688584,10.851214,11.523414,10.782623,10.336777,10.254466,10.683165,11.845795,13.306799,13.097594,11.1393,8.388771,6.848886,7.016936,7.4181976,7.997798,8.855195,10.268185,10.299051,11.592006,14.225929,18.005335,22.487804,24.11343,22.12427,20.145397,19.723558,20.340883,20.382038,21.43835,22.563255,23.797907,26.167753,33.242992,37.708313,35.66771,28.26323,21.671564,15.169065,10.408798,7.5107965,5.994919,4.7774153,4.513337,4.232111,3.8479972,3.4707425,3.3952916,3.7485392,4.2252517,4.245829,3.5221863,2.07833,1.2655178,0.881404,0.83338976,0.9877212,1.1797781,1.3341095,1.3546871,1.1694894,0.85739684,0.6241849,0.5624523,0.41498008,0.32924038,0.33952916,0.34295875,0.26407823,0.33952916,0.36010668,0.28808534,0.25378948,0.39097297,1.0357354,1.4095604,1.2277923,0.70306545,0.72707254,0.7099246,0.83681935,1.0597426,1.1111864,1.0082988,1.039165,1.1351935,1.2620882,1.4198492,1.8519772,1.8519772,1.5536032,1.3066728,1.646202,2.2155135,2.534465,2.750529,2.952875,3.1689389,2.8499873,3.0248961,3.340418,3.4913201,3.2135234,2.860276,2.9803114,3.210094,3.2066643,2.6236343,1.7765263,1.611906,1.5330256,1.2723769,0.90884066,0.65848076,0.58645946,0.5624523,0.5658819,0.6893471,0.823101,1.1900668,1.7902447,2.4007113,2.5893385,2.335549,2.1915064,2.5619018,3.3850029,4.122364,4.6093655,5.5490727,5.6245236,4.9523244,5.096367,4.5442033,4.1943855,4.170378,4.537344,5.295283,7.5759587,10.237319,13.992717,17.778982,18.735836,17.401728,17.250826,17.772121,18.999914,21.517231,23.492674,25.869379,28.475864,30.783978,31.891733,30.657082,28.201498,26.407824,26.613598,29.621347,29.34012,27.872257,27.114319,26.706198,24.027689,22.079683,21.380049,21.503513,22.796469,26.366669,27.402405,26.586163,25.348082,24.43924,23.921373,24.572994,23.677872,21.969936,20.673553,21.493225,19.397747,19.047928,19.61038,19.730417,17.521763,15.141628,15.090185,16.942162,20.755863,27.076593,39.453976,60.44648,84.018036,97.46887,81.44585,56.402996,39.282494,26.548437,16.410576,8.80718,5.888602,4.496189,3.875434,6.3790326,17.484037,10.072699,7.082098,9.990388,14.743796,11.766914,14.232788,14.538021,11.393089,6.48535,4.4447455,5.2815647,5.5490727,5.147811,4.6916757,5.4907694,7.966932,8.327039,7.740579,7.208993,7.579388,5.1340923,3.3952916,2.6064866,3.3712845,6.6431108,11.581717,16.081335,18.279701,17.562918,14.592895,10.127572,8.48137,7.953213,7.5416627,6.9620624,7.8194594,10.302481,14.808959,20.11796,23.413794,30.814844,35.67457,36.689728,33.65454,27.453848,21.167414,17.38115,17.494326,19.421753,17.562918,20.872469,22.892496,25.790497,29.614489,32.292995,36.209583,44.094208,54.098312,66.053856,81.48357,73.64353,60.617958,50.895077,44.670376,33.860317,30.59192,27.584171,25.663603,25.35837,26.922262,25.252052,18.890167,11.4033785,7.455923,12.833516,20.27915,21.476076,17.912735,13.224489,13.152468,12.401388,14.822677,15.484588,15.028452,19.692692,16.832415,23.561266,37.125286,44.591496,22.841053,9.97324,10.518545,18.430603,24.710178,17.391438,11.499407,8.704293,8.971801,11.194174,13.179905,13.440554,15.676644,19.60695,23.499533,24.144297,28.280378,34.103817,34.048943,27.906553,22.851341,20.560377,22.354052,22.964518,22.518671,26.548437,31.775127,37.804344,44.21424,45.699253,32.066643,27.056015,26.558725,25.173172,21.434921,17.820137,14.706071,10.734609,8.580828,9.427936,12.939834,20.001354,22.823904,20.711279,16.088194,14.493437,11.921246,12.055,12.590015,12.994707,14.503725,17.353712,15.868701,11.756626,8.213862,9.921797,14.651197,15.038741,15.371411,17.689812,21.801888,16.427725,11.444533,8.570539,7.6342616,6.56766,6.4579134,5.669108,4.4756117,3.957744,6.018926,11.214751,14.071597,14.870691,13.660047,10.240748,6.5162163,4.856296,4.6573796,4.8768735,4.029765,5.6176643,6.842027,7.8366075,8.467651,8.323608,8.580828,6.759717,5.288424,5.113515,5.6965446,5.5833683,5.113515,5.6142344,6.9071894,7.291303,8.48137,9.146709,9.132992,8.820899,9.132992,7.623973,6.0532217,6.385892,8.279024,9.0644,8.182996,6.159539,4.7774153,4.3658648,3.8274195,5.0414934,6.492209,8.213862,9.407358,8.457363,6.3207297,6.8454566,7.010077,5.658819,3.5050385,4.7602673,5.1169443,4.8322887,4.7842746,6.478491,6.989499,5.2918534,3.1449318,1.762808,1.7971039,5.675967,8.505377,7.610255,4.647091,5.586798,8.923786,8.285883,6.2658563,5.329579,7.8091707,7.857185,6.9346256,5.4496145,3.7313912,2.020027,1.5673214,1.5055889,1.5536032,1.587899,1.646202,1.6187652,1.9308578,2.311542,2.5550427,2.5310357,2.411,3.018037,3.316411,3.1312134,3.1277838,3.3781435,3.1586502,3.0489032,3.292404,3.7965534,3.5702004,3.9680326,4.2869844,4.465323,5.079219,4.962613,4.4447455,5.295283,6.6053853,4.7602673,7.284444,10.4533825,9.115844,5.744559,10.432805,2.836269,0.38754338,0.1097468,1.0940384,4.4859004,1.3889829,0.32924038,0.25378948,0.3841138,0.216064,0.0548734,0.006859175,0.006859175,0.024007112,0.05144381,0.12346515,0.19891608,0.26064864,0.32924038,0.48357183,0.5761707,0.5418748,0.5521636,0.69963586,0.99801,0.88826317,0.90541106,0.922559,0.91912943,0.9602845,1.0528834,1.2449403,1.430138,1.5261664,1.4987297,1.5193073,1.4095604,1.2929544,1.2655178,1.4164196,1.3752645,1.4850113,1.5021594,1.4198492,1.4507155,1.5364552,1.4747226,1.5158776,1.6633499,1.6804979,1.6976458,1.5604624,1.3169615,1.0254467,0.75450927,0.61046654,0.5658819,0.5521636,0.52815646,0.44927597,0.548734,0.6207553,0.607037,0.52472687,0.4629943,0.44584638,0.51100856,0.58988905,0.6310441,0.61046654,0.7133542,0.7099246,0.70649505,0.72707254,0.72364295,0.69963586,0.6344737,0.6173257,0.65162164,0.65162164,0.64133286,0.5693115,0.4972902,0.432128,0.32581082,0.34981793,0.3018037,0.20920484,0.12346515,0.11317638,0.14747226,0.23664154,0.33266997,0.3806842,0.33609957,0.33952916,0.34295875,0.33609957,0.32581082,0.32924038,0.40126175,0.44584638,0.47328308,0.47671264,0.4629943,0.3841138,0.33609957,0.3018037,0.26407823,0.22635277,0.216064,0.15090185,0.09259886,0.06859175,0.05144381,0.041155048,0.034295876,0.034295876,0.044584636,0.058302987,0.08573969,0.13375391,0.1920569,0.26407823,0.37382504,0.58988905,0.7099246,0.85396725,1.0563129,1.2586586,1.2826657,1.3581166,1.4061309,1.4129901,1.3992717,1.3512574,1.2998136,1.2449403,1.1934965,1.1660597,1.2415106,1.3821237,1.4850113,1.4987297,1.4061309,1.4335675,1.4472859,1.4129901,1.3821237,1.4850113,1.5501735,1.6290541,1.6599203,1.646202,1.6393428,1.7593783,1.9445761,2.095478,2.1743584,2.2052248,2.2155135,2.1640697,2.095478,2.061182,2.1057668,2.16064,2.2292318,2.3561265,2.510458,2.5790498,2.369845,2.318401,2.3629858,2.486451,2.702515,3.1586502,3.6216443,4.0263357,4.479041,5.2266912,6.1766872,6.790583,7.1369715,7.3873315,7.8263187,8.913498,10.693454,14.009865,20.220848,31.202387,0.0,0.0548734,0.18862732,0.2777966,0.29837412,0.35324752,0.47671264,0.47671264,0.45956472,0.48014224,0.53844523,0.6962063,0.864256,1.1283343,1.4541451,1.6770682,1.8965619,2.136633,2.2360911,2.1812177,2.0920484,1.9754424,1.9411465,2.253239,2.8568463,3.3850029,3.9337368,4.372724,4.4516044,4.1429415,3.6182148,4.057202,5.8371577,7.3358874,7.8434668,7.5553813,7.9257765,8.995808,10.100135,10.72775,10.532263,10.751757,10.984968,11.283342,12.0309925,13.9309845,14.592895,12.936404,10.323058,7.9943686,7.06838,8.2653055,8.899779,9.23245,9.647429,10.6317215,10.80663,13.022143,17.04505,21.877338,25.77335,27.292658,26.665043,27.693918,30.495892,31.497332,29.988314,28.534168,27.117748,25.646456,23.952238,24.806206,29.991743,33.726562,33.116096,28.17406,21.77102,14.959861,10.14129,7.699424,5.98463,5.288424,4.616225,3.9611735,3.5050385,3.6010668,3.350707,3.4947495,3.899441,4.149801,3.5599117,2.5413244,1.862266,1.5604624,1.471293,1.2346514,1.0288762,1.2792361,1.3649758,1.0734608,0.6001778,0.4698535,0.33952916,0.30866286,0.37382504,0.4629943,0.35324752,0.44584638,0.48700142,0.41840968,0.3841138,0.42869842,0.96714365,1.3341095,1.196926,0.5555932,0.37382504,0.33609957,0.48357183,0.69963586,0.72021335,0.7682276,0.82996017,0.8848336,0.9774324,1.2312219,1.5707511,1.7936742,1.8519772,1.8416885,2.0097382,2.5961976,3.3301294,3.7005248,3.6044965,3.3301294,3.4433057,4.081209,4.5201964,4.4447455,3.9714622,3.5153272,3.4604537,3.5702004,3.57363,3.1655092,1.7250825,1.0700313,0.7442205,0.52472687,0.44584638,0.5212973,0.5658819,0.70306545,0.9259886,1.1317638,1.214074,1.471293,1.8176813,2.0234566,1.6942163,1.7559488,1.6084765,1.3615463,1.2037852,1.3992717,2.2841053,2.644212,2.9563043,3.426158,3.981751,4.9180284,5.1855364,5.3432975,5.638242,6.029215,8.834618,12.360233,16.012743,18.632948,18.492336,17.820137,16.678083,16.561478,17.988186,20.519222,26.431831,28.94229,30.489033,31.905453,32.39588,29.26124,27.896265,28.907993,31.559063,33.729992,31.613937,28.294096,25.920822,24.974257,24.281479,22.587263,20.749004,20.53294,22.261452,24.792488,26.77136,26.822803,25.317215,23.588703,23.948809,25.619019,24.096281,21.524092,19.795578,20.574095,18.228258,18.821575,19.6241,18.95533,16.160215,13.073587,12.154458,14.441993,19.05136,23.170294,30.372427,45.095646,69.051315,91.751755,90.49652,59.969765,39.91011,26.370098,16.321407,7.6514096,5.0414934,3.8514268,3.4638834,5.4770513,13.680624,12.006986,10.110424,12.850664,17.494326,13.725209,14.212211,14.651197,12.915827,9.338767,6.711703,8.285883,7.740579,6.4407654,5.6793966,6.6876955,8.7145815,9.040393,8.30646,7.7371492,9.112414,6.23499,3.9714622,2.668219,2.7230926,4.5853586,10.041832,11.55771,15.824117,21.644127,19.919044,13.056439,9.304471,8.824328,9.949233,9.191295,8.841476,9.873782,12.874671,17.322845,21.554956,30.118637,34.854897,35.90435,32.176388,21.349182,17.610931,16.400288,20.409475,24.751333,16.969599,21.496655,22.957659,26.208908,31.555634,34.74515,37.58828,40.781223,47.592384,58.11779,69.301674,50.853924,40.79151,41.439705,45.39402,35.530525,34.35761,33.620247,31.891733,30.43759,33.212124,31.716825,21.884197,13.05301,11.129011,18.578075,24.871368,21.345753,15.717799,12.9707,15.364552,12.542002,14.212211,14.476289,14.061309,20.313446,20.217419,29.209797,39.107586,40.48285,22.69701,11.1393,11.249047,13.7697935,13.176475,7.6685576,5.446185,6.416758,9.191295,12.199042,13.666906,12.751206,14.901558,18.38259,21.218857,21.174273,23.01596,25.536709,24.497543,20.474638,18.852442,19.53493,23.324625,24.415234,22.607841,23.307476,26.19176,31.360147,35.22872,34.937206,28.342112,26.130028,25.546997,22.841053,17.367432,11.571428,11.780633,9.132992,8.279024,10.672876,14.565458,17.590355,18.169954,15.206791,10.655728,9.517105,8.152129,10.388221,12.665466,14.613472,19.068506,20.793589,17.19938,11.763485,8.868914,13.807519,14.894698,14.212211,15.518884,19.11652,21.843042,14.5414505,10.762046,9.290752,8.700864,7.366754,6.680836,5.579939,3.9714622,2.7402403,3.7382503,8.399059,14.363112,16.94902,14.688923,9.3079,7.0306544,5.686256,5.1580997,5.1752477,5.31929,6.111525,7.5416627,8.30646,8.457363,9.39021,9.671436,8.694004,7.377043,6.210983,5.267846,4.695105,5.363875,6.3173003,6.8763227,6.615674,8.028665,8.1212635,7.2295704,6.2555676,6.667118,5.206114,5.23698,6.866034,9.146709,10.062409,6.8454566,5.312431,4.9660425,4.6573796,2.5756202,3.6387923,5.288424,5.6965446,5.0174866,5.411889,6.3961806,7.0958166,6.3447366,4.3487167,2.668219,7.689135,8.344186,6.6122446,5.2747054,7.9086285,8.7317295,5.3913116,2.2360911,1.1797781,1.6976458,7.394191,8.604835,6.0326443,2.5893385,3.4192986,6.5059276,6.310441,5.2781353,6.142391,11.924676,9.770895,7.6514096,5.7719955,4.149801,2.6407824,2.0989075,1.6942163,1.4541451,1.3684053,1.3786942,1.5673214,1.6942163,1.9685832,2.318401,2.3595562,2.054323,2.3424082,2.6407824,2.7711067,2.9734523,3.1792276,2.7642474,2.7470996,3.3712845,4.1326528,3.6593697,3.0900583,2.935727,3.1277838,3.0317552,3.57363,3.9646032,4.928317,6.046363,5.785714,5.65539,7.2467184,6.210983,3.4844608,5.295283,3.1243541,1.0323058,0.0034295875,0.9877212,4.887162,1.5398848,0.33952916,0.20577525,0.36696586,0.37382504,0.10288762,0.01371835,0.006859175,0.0274367,0.06859175,0.17147937,0.22635277,0.28122616,0.3841138,0.59331864,0.6276145,0.5041494,0.5590228,0.8196714,1.0048691,0.88826317,0.9294182,1.0048691,1.0357354,0.9842916,0.99801,1.2449403,1.4575747,1.4987297,1.3992717,1.3581166,1.196926,1.1866373,1.3443983,1.4198492,1.3375391,1.5055889,1.5673214,1.4815818,1.5330256,1.6599203,1.5810398,1.587899,1.7182233,1.7799559,1.821111,1.4987297,1.1214751,0.85739684,0.7613684,0.6824879,0.6756287,0.6756287,0.64819205,0.5796003,0.6173257,0.7339317,0.7476501,0.6344737,0.53158605,0.5178677,0.5727411,0.67219913,0.7407909,0.65162164,0.6962063,0.69963586,0.71678376,0.7373613,0.6893471,0.66533995,0.58988905,0.61389613,0.72364295,0.7442205,0.69963586,0.64819205,0.6001778,0.5453044,0.45613512,0.4664239,0.39783216,0.28808534,0.17490897,0.13032432,0.106317215,0.14747226,0.2503599,0.35324752,0.34638834,0.33266997,0.30523327,0.2709374,0.25721905,0.28808534,0.39440256,0.4424168,0.45270553,0.45613512,0.4972902,0.48357183,0.45613512,0.39097297,0.32238123,0.33609957,0.36010668,0.25721905,0.16462019,0.12003556,0.082310095,0.05144381,0.037725464,0.034295876,0.030866288,0.030866288,0.0274367,0.05144381,0.08573969,0.12346515,0.17147937,0.274367,0.32924038,0.42526886,0.59331864,0.8025235,0.9911508,1.2826657,1.5021594,1.587899,1.5844694,1.3821237,1.2346514,1.1351935,1.0734608,1.039165,1.0940384,1.2723769,1.3684053,1.3546871,1.3581166,1.4061309,1.488441,1.5398848,1.5741806,1.7113642,1.7010754,1.7422304,1.7319417,1.6599203,1.6290541,1.7525192,1.9342873,2.0234566,1.99602,1.9651536,1.978872,2.0406046,2.0714707,2.0920484,2.2155135,2.2463799,2.3801336,2.5996273,2.867135,3.1243541,2.9048605,2.7951138,2.726522,2.6750782,2.6476414,2.9391565,3.292404,3.549623,3.7382503,4.0709205,5.3432975,5.8645945,6.2658563,6.8385973,7.5416627,8.032094,9.489669,11.80464,15.282242,20.642687,0.0,0.024007112,0.058302987,0.07545093,0.12346515,0.30523327,0.32924038,0.29151493,0.28465575,0.35324752,0.48700142,0.5007198,0.5590228,0.7613684,1.0906088,1.4198492,1.5398848,1.762808,1.879414,1.8005334,1.5570327,1.4575747,1.4815818,1.937717,2.8122618,3.7382503,4.530485,4.9488945,4.846007,4.3761535,3.998899,5.7925735,8.375052,9.033533,7.750868,7.2021337,8.899779,10.80663,11.862943,11.924676,11.763485,13.251926,14.256795,14.191633,13.783512,15.090185,15.371411,12.668896,9.932085,8.495089,8.056101,9.2153015,9.4862385,9.451943,9.877212,11.718901,11.413667,14.222499,19.94648,27.374968,34.271866,36.103268,36.724022,41.40541,49.475227,54.334953,49.279743,42.96587,36.610847,30.410152,23.513252,20.255144,19.514353,23.461807,29.700228,31.2504,25.0257,18.423744,13.083877,9.671436,7.888051,5.7754254,4.5819287,3.8720043,3.309552,2.6236343,2.5378947,2.352697,2.7128036,3.6182148,4.4241676,4.166949,3.6387923,2.976882,2.4315774,2.335549,1.4438564,1.4507155,1.5090185,1.2243627,0.6241849,0.4046913,0.34981793,0.47328308,0.67219913,0.7339317,0.37725464,0.2709374,0.3018037,0.4081209,0.5796003,0.65162164,1.1111864,1.4095604,1.313532,0.8848336,0.7510797,0.5418748,0.34638834,0.25721905,0.36696586,0.7442205,0.91227025,0.96714365,0.9842916,1.0220171,1.4610043,2.0028791,2.5756202,3.0866287,3.4021509,3.549623,3.9508848,4.2766957,4.465323,4.746549,3.7931237,3.683377,3.549623,3.3609958,3.9200184,5.2644167,6.7700057,6.824879,5.579939,4.9591837,2.7368107,1.3752645,0.7888051,0.7373613,0.823101,1.0082988,1.1523414,1.3375391,1.546744,1.6942163,1.670209,1.6256244,1.6564908,1.7559488,1.8142518,2.0234566,1.845118,1.6633499,1.646202,1.7559488,1.9754424,2.4247184,3.4227283,4.73969,5.56965,6.5333643,5.9983487,5.579939,6.090947,7.507367,10.206452,14.387119,20.025362,26.733635,33.75057,30.235243,24.751333,19.984205,18.04306,20.4472,28.417562,33.778008,37.204166,39.15903,39.91697,35.863197,33.1744,32.852016,34.57367,36.696587,35.14641,30.876575,26.10945,22.645567,21.849901,20.179693,19.157675,19.912186,21.897917,22.889067,25.804216,26.77136,25.77678,24.511261,26.366669,27.673342,24.027689,19.630959,17.329706,18.584934,19.696121,21.915064,22.127699,19.442331,15.182784,14.400838,12.521424,12.679185,15.306249,18.1288,21.77788,31.294985,50.836777,75.72872,92.499405,64.911804,40.033573,22.77932,12.88839,4.928317,4.5270553,3.782835,3.758828,5.295283,9.019815,21.503513,20.049368,17.676094,18.732407,18.890167,21.70929,19.823015,17.370861,15.902997,14.387119,13.227919,11.399949,9.002667,7.5450926,9.949233,11.485688,10.9198065,9.331907,7.490219,5.830299,8.282454,6.012067,3.7965534,3.5976372,4.5613513,8.553391,13.1593275,16.300829,18.86959,24.703318,23.69159,15.525743,10.511685,10.669447,9.764035,11.729189,12.644889,13.498857,15.4742985,19.94305,32.687397,41.347107,42.372555,34.98522,21.177702,16.064188,14.685493,22.02824,31.192099,23.389786,15.494876,14.88441,18.351723,26.582733,44.159367,49.674145,47.65069,44.660088,44.179947,46.57037,31.483612,30.639935,37.464813,43.199085,36.90922,35.726013,35.99695,36.41879,37.15615,39.84152,32.50563,20.076805,13.944703,15.96816,18.492336,15.234227,13.138749,12.288212,12.010415,10.847785,11.729189,20.560377,22.78275,16.88043,14.404267,19.006773,27.635616,29.912863,23.160004,12.404818,11.465111,11.561139,11.396519,10.158438,7.5210853,6.7665763,8.371623,10.703742,13.032433,15.532601,14.71636,13.073587,13.104454,14.726648,15.289101,15.618341,17.580065,17.70696,15.741806,14.616901,19.099373,21.143406,21.935642,22.926792,25.831654,20.731855,22.422644,27.731644,33.040646,34.285587,26.058006,19.716698,14.565458,11.327928,12.147599,11.585147,10.062409,10.206452,13.258785,19.058218,14.555169,11.626302,10.532263,10.093276,7.675417,5.672538,9.431366,11.828648,13.035862,20.508932,19.03078,17.545769,14.829536,12.854094,16.7844,15.443433,15.234227,17.573206,20.745575,19.929333,14.373401,11.897239,10.851214,10.076128,8.879202,8.525954,6.6053853,4.256118,2.5790498,2.6407824,6.2658563,11.201033,15.155347,15.54632,9.489669,7.085528,5.761707,5.144381,5.4667625,7.5519514,7.56567,6.0669403,5.9400454,7.7680154,9.8429165,9.928656,9.839486,9.0644,7.5862474,5.888602,4.972902,5.586798,5.9983487,5.3844523,3.8445675,5.8234396,7.4696417,8.018375,7.2775846,5.6313825,4.616225,6.0840883,7.0615206,6.8283086,6.914048,4.5442033,2.6167753,2.061182,2.867135,4.0880685,3.9303071,3.7176728,3.4776018,3.6765177,5.2026844,6.0703697,6.029215,5.363875,4.681387,4.914599,9.56512,9.6645775,7.0889573,5.137522,8.529384,6.4407654,3.3198407,1.488441,1.978872,4.5167665,5.6519604,4.0777793,2.0028791,1.5021594,4.5167665,4.5167665,2.942586,4.7671266,10.545981,16.417435,9.544542,5.3844523,4.3041325,5.0449233,4.715683,3.7622573,2.6545007,2.0028791,1.7833855,1.3443983,1.5981878,1.4335675,1.6221949,2.1400626,2.1503513,2.0406046,2.4075704,2.7985435,3.0454736,3.2649672,2.6785078,2.3767042,2.651071,3.2889743,3.5702004,3.1689389,2.7093742,2.6613598,2.9220085,2.8225505,3.3850029,3.5702004,3.9611735,5.0277753,7.140401,4.773986,4.3281393,3.6147852,2.095478,0.90198153,3.2821152,1.5501735,0.0,0.19891608,0.9911508,1.2963841,0.6241849,0.17147937,0.3018037,0.53501564,0.20577525,0.048014224,0.006859175,0.034295876,0.106317215,0.26407823,0.31552204,0.34638834,0.37382504,0.33609957,0.22635277,0.29837412,0.6173257,0.9911508,0.9911508,0.7099246,0.65848076,0.84367853,1.1283343,1.2517995,1.2277923,1.2380811,1.2895249,1.3238207,1.2517995,1.1523414,1.1008976,1.1763484,1.3581166,1.5398848,1.6633499,1.6942163,1.6324836,1.5673214,1.6770682,1.6770682,1.7250825,1.845118,1.9239986,1.6942163,1.6084765,1.3203912,1.0837497,1.0185875,1.1283343,0.97057325,0.77508676,0.6824879,0.70306545,0.70306545,0.5555932,0.6756287,0.764798,0.7133542,0.5796003,0.5555932,0.6241849,0.805953,1.0082988,1.0082988,0.7888051,0.7613684,0.77165717,0.7510797,0.70306545,0.6790583,0.5796003,0.5796003,0.70649505,0.85396725,0.67219913,0.6173257,0.6241849,0.6276145,0.5796003,0.4698535,0.36010668,0.31209245,0.29151493,0.16804978,0.14404267,0.14747226,0.14747226,0.15090185,0.19891608,0.23664154,0.26407823,0.274367,0.28808534,0.33609957,0.3841138,0.42526886,0.44927597,0.44927597,0.4115505,0.4972902,0.53844523,0.53158605,0.50757897,0.5178677,0.44584638,0.36353627,0.3018037,0.25378948,0.16804978,0.106317215,0.072021335,0.048014224,0.030866288,0.030866288,0.017147938,0.024007112,0.024007112,0.024007112,0.061732575,0.09602845,0.13375391,0.19548649,0.32581082,0.59674823,0.90198153,1.2037852,1.4747226,1.646202,1.6324836,1.4507155,1.3306799,1.2758065,1.2243627,1.0528834,1.0768905,1.0185875,1.0254467,1.1249046,1.2346514,1.4198492,1.611906,1.6907866,1.6633499,1.6633499,1.5638919,1.5776103,1.5158776,1.4232788,1.5570327,1.6907866,1.704505,1.7010754,1.7216529,1.7696671,1.7456601,1.8039631,1.9308578,2.1057668,2.287535,2.201795,2.4830213,2.9185789,3.309552,3.4776018,3.309552,3.018037,2.8054025,2.7093742,2.6236343,2.8568463,3.1072063,3.2958336,3.5221863,4.057202,4.6093655,5.3227196,5.8337283,6.1732574,6.759717,7.016936,7.939495,9.918367,13.560589,19.713268,0.01371835,0.12346515,0.12003556,0.12346515,0.18519773,0.28122616,0.30523327,0.34638834,0.4046913,0.44584638,0.41498008,0.48700142,0.5521636,0.7682276,1.039165,1.0288762,1.1420527,1.3546871,1.4164196,1.313532,1.2758065,1.4610043,1.8108221,2.4041407,3.3129816,4.5922174,6.293293,7.2604365,7.1541195,6.228131,5.3398676,7.058091,9.290752,9.640571,8.553391,9.314759,11.382801,12.614022,13.509145,14.507155,15.999025,18.327715,18.135658,16.530611,14.88441,14.822677,13.725209,12.377381,11.341646,10.738038,10.240748,9.283894,8.320179,9.23245,11.907528,14.256795,14.109323,16.39,22.316326,31.569353,42.303963,46.6321,52.7059,62.53853,71.7504,69.56918,57.6205,46.079937,36.7446,30.111778,25.382378,20.96164,17.971039,17.497755,19.339443,22.021381,18.588364,14.54831,11.4376745,9.427936,7.31531,5.7582774,4.4241676,3.3369887,2.5207467,2.0131679,1.646202,1.6016173,1.7319417,1.9445761,2.2052248,2.49331,3.0386145,3.1209247,2.6990852,2.4075704,1.546744,1.2586586,1.1489118,0.99801,0.7613684,0.47328308,0.4081209,0.5521636,0.764798,0.7579388,0.432128,0.31895164,0.34981793,0.45613512,0.5796003,0.61389613,0.7099246,0.8128122,0.85739684,0.7613684,0.7442205,0.59674823,0.4389872,0.39097297,0.548734,0.45956472,0.41498008,0.48357183,0.6962063,1.0357354,1.6016173,2.0714707,2.6476414,3.292404,3.707384,3.6216443,3.7313912,4.040054,4.389872,4.4756117,4.0434837,3.9371665,4.2869844,4.8425775,4.996909,6.697984,9.139851,11.207891,11.80121,9.8429165,6.252138,3.4878905,1.9102802,1.3752645,1.2277923,1.4575747,1.8588364,2.4247184,3.0557625,3.57363,3.4913201,3.117495,2.6647894,2.270387,1.9994495,2.1674993,2.1572106,2.2463799,2.5001693,2.767677,3.40901,4.650521,5.4016004,5.422178,5.3261495,6.835168,7.4044795,8.673427,11.204462,14.466,19.53493,26.397535,35.304173,43.89872,47.21513,37.07041,26.983994,21.143406,20.594673,23.252604,28.51016,29.885426,30.7634,31.634514,30.067194,28.396984,28.698788,31.977474,37.276188,41.666058,40.544582,33.16754,25.735624,21.386908,20.2037,19.761284,19.809298,20.834743,22.432932,23.304047,26.737064,27.916842,28.047167,27.851679,27.539587,26.843382,25.34122,22.878778,19.994495,17.912735,20.604961,21.699,21.702429,20.296299,16.328266,14.239647,14.2362175,16.228807,18.53692,17.919594,18.845583,21.976797,33.25328,52.20861,71.969894,50.20916,30.722244,16.681513,8.508806,3.8925817,3.4398763,3.0660512,3.192946,3.9131594,4.99005,10.710602,14.805529,14.956431,13.077017,15.313108,19.11995,16.835844,13.649758,13.13532,17.257685,13.245067,11.72233,10.477389,8.985519,8.4093485,10.419086,10.9198065,10.388221,8.573969,4.523626,8.1487,9.81205,10.285333,9.595985,7.016936,6.341307,9.3593445,12.404818,15.556609,22.642136,19.812727,17.7927,17.775553,18.989626,18.70154,16.05733,14.637479,15.6252,20.320305,30.146074,46.5738,52.397236,43.696373,26.483274,16.698662,15.745236,16.400288,19.572655,23.334913,22.916504,24.703318,24.655304,28.331821,35.695145,41.09675,46.409176,43.49403,36.319332,31.394444,37.770046,34.117535,34.16212,36.92294,40.08159,39.975273,39.32708,36.429077,35.918068,43.264244,64.76433,40.839527,27.786518,21.747015,18.735836,14.671775,10.203023,9.019815,10.13786,12.0138445,12.531713,22.436361,34.631973,33.284145,18.897026,8.327039,10.9369545,15.37827,17.511473,16.047039,12.538571,14.246507,15.141628,14.2533655,12.504276,12.710052,12.120162,9.798331,8.848335,10.515115,14.177915,14.658057,12.566009,12.298501,14.531162,16.204802,14.922135,15.21365,16.170506,17.960749,21.808746,25.51613,23.736176,21.050808,20.61182,24.11343,21.421204,22.412354,26.380386,29.662502,25.643026,20.327166,14.990726,11.046701,9.884071,12.878101,12.902108,11.334786,11.218181,12.785502,13.46799,11.345076,10.734609,11.050131,10.813489,7.6274023,6.756287,8.255017,9.417647,12.21619,23.280039,22.076254,16.45516,12.068718,11.674315,15.138199,15.786391,19.078794,21.129688,19.816156,14.788382,11.7257595,10.542552,10.549411,10.827208,10.233889,7.3427467,5.07236,3.5770597,2.8156912,2.5550427,4.2938433,7.7542973,10.943813,12.079007,9.589127,7.438775,6.324159,5.7274113,5.675967,6.7459984,5.6176643,4.07435,3.9508848,5.545643,7.6205435,7.675417,7.250148,8.083538,9.623423,9.050681,11.063849,10.367643,9.80519,9.89093,8.800322,6.8043017,6.307011,6.800872,7.0615206,5.178677,4.1360826,6.118384,7.133542,6.2041235,5.360445,5.579939,4.5990767,4.15323,4.48933,4.383013,3.7142432,3.1415021,3.1860867,4.1017866,5.861165,5.079219,5.284994,7.5588107,9.592556,5.693115,8.635701,7.6788464,5.3570156,3.683377,4.1463714,3.1826572,1.821111,1.255229,1.7593783,2.6853669,2.3664153,1.7388009,2.4555845,4.588788,6.6293926,4.4516044,2.6990852,5.627953,11.197603,11.084427,6.1149545,4.091498,4.9248877,6.540223,4.8597255,4.835718,4.619654,3.2889743,1.4610043,1.2929544,1.5021594,1.5604624,1.6256244,1.7490896,1.8588364,2.1503513,2.3801336,2.503599,2.609916,2.9494452,3.0660512,3.0866287,3.117495,3.0729103,2.6785078,2.5790498,2.5550427,2.5961976,2.627064,2.5310357,2.7882545,2.8396983,3.3712845,4.7774153,7.1541195,5.2644167,5.501058,6.1046658,5.178677,0.6927767,2.2635276,1.3409687,0.2777966,0.041155048,0.20920484,0.7305021,0.41840968,0.12346515,0.16804978,0.34981793,0.16804978,0.048014224,0.010288762,0.05144381,0.15433143,0.3841138,0.47671264,0.4629943,0.4081209,0.4081209,0.5727411,0.7133542,1.0220171,1.2998136,0.96714365,1.1077567,0.939707,0.82996017,0.9568549,1.3238207,1.3684053,1.2723769,1.2037852,1.2003556,1.1660597,1.3032433,1.2346514,1.1729189,1.2346514,1.4678634,1.6290541,1.6839274,1.6359133,1.6153357,1.862266,1.7250825,1.5913286,1.5913286,1.6393428,1.4369972,1.4198492,1.2826657,1.196926,1.1694894,1.0425946,0.9842916,0.91569984,0.8162418,0.7133542,0.66533995,0.6173257,0.7305021,0.85739684,0.89169276,0.7888051,0.84024894,0.86082643,0.8745448,0.8848336,0.8848336,0.7922347,0.7956643,0.8128122,0.7956643,0.72707254,0.7510797,0.7305021,0.7133542,0.7510797,0.9294182,0.8711152,0.71678376,0.6001778,0.5624523,0.5418748,0.4629943,0.4046913,0.432128,0.4629943,0.25378948,0.18862732,0.16804978,0.16462019,0.16462019,0.17490897,0.2194936,0.28808534,0.30866286,0.29837412,0.34638834,0.44584638,0.5178677,0.59674823,0.66876954,0.6790583,0.64819205,0.64476246,0.66876954,0.6962063,0.6790583,0.5555932,0.47671264,0.41840968,0.36696586,0.3018037,0.2709374,0.216064,0.15090185,0.09945804,0.07888051,0.048014224,0.0274367,0.017147938,0.017147938,0.024007112,0.041155048,0.06516216,0.09259886,0.1371835,0.24007112,0.41840968,0.58988905,0.8196714,1.0734608,1.2175035,1.3066728,1.3443983,1.371835,1.371835,1.2483698,1.2346514,1.1660597,1.1420527,1.1797781,1.2106444,1.3272504,1.4198492,1.4953002,1.5570327,1.6256244,1.5981878,1.6564908,1.6633499,1.6187652,1.6530612,1.7113642,1.6976458,1.6976458,1.7079345,1.6599203,1.6564908,1.6804979,1.786815,1.9137098,1.9239986,2.0817597,2.3149714,2.6304936,2.9974594,3.3438478,3.5633414,3.5118976,3.3747141,3.2409601,3.07634,3.0043187,3.2821152,3.6147852,3.8891523,4.180667,4.770556,5.411889,5.892031,6.1629686,6.358455,6.3001523,6.3035817,7.507367,10.628291,15.978448,0.06859175,0.13032432,0.15090185,0.14061308,0.1371835,0.20234565,0.36353627,0.44584638,0.47671264,0.4664239,0.37725464,0.41840968,0.5212973,0.6859175,0.8471081,0.8676856,0.97057325,1.155771,1.2003556,1.1592005,1.3615463,1.5673214,1.8176813,2.386993,3.4467354,5.099797,6.8591747,8.1487,8.323608,7.56567,6.8763227,7.658269,8.89635,9.129561,8.673427,9.650859,11.252477,12.994707,14.874121,16.839275,18.770132,20.803877,20.86904,19.020493,16.396858,15.2033615,14.267084,14.730078,15.357693,15.05246,12.857523,10.995257,10.096705,11.4376745,14.493437,16.979887,18.094503,22.43979,32.306713,45.63066,55.991444,60.17211,68.30023,78.547844,83.836266,71.82242,56.070324,41.98501,31.751122,25.821363,22.899355,18.900457,15.46744,13.334236,12.679185,13.1421795,11.616013,10.295622,8.947794,7.5039372,6.0532217,5.2609873,4.314421,3.3541365,2.5619018,2.1640697,2.0406046,1.7559488,1.4027013,1.1283343,1.1523414,1.3306799,1.8725548,2.3149714,2.469303,2.4247184,1.8142518,1.3752645,1.0734608,0.8471081,0.6207553,0.42526886,0.4355576,0.66191036,0.91569984,0.78194594,0.44927597,0.26750782,0.2709374,0.39440256,0.48700142,0.58645946,0.66533995,0.7133542,0.72707254,0.7133542,0.7407909,0.66533995,0.6001778,0.61389613,0.7339317,0.53844523,0.3806842,0.4046913,0.6241849,0.90198153,1.2860953,1.7662375,2.2669573,2.6853669,2.9048605,2.9117198,3.0386145,3.350707,3.6765177,3.5942078,4.2355404,5.137522,6.1629686,6.848886,6.39961,6.7871537,8.213862,9.860064,10.696883,9.469091,6.6225333,4.0023284,2.3492675,1.7593783,1.6770682,2.0440342,2.627064,3.4810312,4.431027,5.079219,5.178677,5.079219,4.7362604,4.245829,3.8479972,3.7725463,3.391862,3.2581081,3.5599117,4.1189346,5.267846,6.307011,6.869464,7.010077,7.2158523,8.275595,8.340756,9.966381,13.509145,17.130789,19.45262,23.184011,28.280378,32.886314,33.352737,24.963966,19.253704,17.29884,18.766703,21.904776,26.051146,27.220636,27.60132,27.954567,27.594461,27.76594,30.653652,35.41392,40.729782,44.831566,40.366245,31.284697,24.37065,22.079683,22.52896,21.681852,21.253153,21.808746,23.259462,24.871368,27.409264,27.213776,25.8488,24.590141,24.418663,22.378057,21.87048,21.424633,20.148827,17.737827,19.895037,18.965618,18.015623,17.816708,16.835844,14.177915,14.695783,16.732958,18.03277,15.745236,17.034761,18.21111,25.125158,37.58142,49.331184,31.689388,18.169954,9.901219,5.9640527,3.3747141,3.0146074,3.3472774,3.8102717,4.3795834,5.5559316,6.012067,10.30934,11.008976,8.186425,9.458802,11.334786,9.407358,7.4181976,7.8777623,12.05157,10.947243,11.348505,12.332796,12.017275,7.5416627,9.256456,8.872343,10.813489,13.022143,6.989499,10.47396,12.754636,13.927555,13.72178,11.492548,9.31133,11.523414,14.030442,17.343424,26.555296,20.817596,20.855322,23.794477,27.128036,28.705647,22.690151,20.152256,21.318316,26.472986,35.948936,50.9671,50.45609,38.267338,23.434372,20.165974,24.212887,25.670462,25.975695,25.495554,23.557837,34.67999,45.349434,49.38949,45.418026,36.83034,37.09099,35.383053,32.5022,32.23812,41.364254,41.38826,39.2482,38.085567,39.67347,44.392582,47.307728,44.046192,43.367134,49.314037,61.20442,44.612072,35.719154,28.774239,20.755863,11.372512,8.035523,7.864044,9.417647,12.346515,17.405157,29.652214,35.67114,30.962317,18.605513,9.294182,9.253027,10.340206,11.859513,12.932974,12.517994,14.3974085,15.22051,13.917266,11.832077,12.71691,11.163307,9.921797,10.4533825,12.020704,11.670886,13.419975,12.795791,12.651748,14.229359,17.158226,16.95931,17.995045,20.598103,24.288338,27.752222,33.18126,28.139765,21.880768,19.11309,20.001354,19.87789,26.140316,32.74227,33.58595,22.53239,17.339994,13.046151,10.182446,9.270175,10.81006,11.660598,11.478829,12.041282,13.083877,12.288212,11.547421,11.489118,11.135871,10.39165,10.05898,9.47938,8.450503,8.405919,12.085866,23.52354,22.53582,15.199932,10.556271,11.362224,14.119612,14.695783,17.04848,17.720678,15.5085945,11.434244,11.067279,11.012405,11.482259,11.7257595,10.024684,6.495639,5.1855364,4.1600895,3.1517909,3.549623,3.4776018,4.945465,6.6396813,7.7885933,8.131552,6.461343,5.871454,5.7308407,5.627953,5.3570156,3.940596,2.9254382,2.8019729,3.5804894,4.7842746,4.3590055,4.722542,6.0052075,7.5690994,8.038953,10.398509,10.415657,9.760606,9.153569,8.375052,6.159539,5.470192,6.543653,7.8537555,6.118384,4.3795834,4.8905916,5.7102633,5.895461,5.48734,5.5833683,4.2526884,4.2115335,5.501058,5.470192,3.083199,2.5447538,2.9322972,3.9165888,5.7719955,4.290414,4.1017866,7.0546613,10.203023,5.8062916,5.672538,4.7534084,3.5702004,2.644212,2.5207467,2.7813954,2.4967396,2.5721905,3.192946,3.8205605,3.9851806,3.9508848,4.3933015,5.254128,5.7377,3.2718265,2.335549,4.3487167,7.4456344,6.464772,4.887162,5.1683884,6.1732574,6.358455,3.782835,4.479041,5.586798,5.6210938,4.125794,1.646202,1.5433143,1.6804979,1.7353712,1.6907866,1.8416885,2.510458,2.5790498,2.3595562,2.2566686,2.767677,3.1483612,3.3609958,3.275256,2.9288676,2.5310357,2.5138876,2.5721905,2.7299516,2.976882,3.2821152,3.2512488,3.234101,3.6113555,5.4667625,10.590566,9.9698105,9.496528,10.028113,10.401938,7.4524937,3.6353626,1.2106444,0.14404267,0.006859175,0.006859175,0.2503599,0.20920484,0.2194936,0.33952916,0.34295875,0.14404267,0.044584636,0.0274367,0.09259886,0.22292319,0.4389872,0.5144381,0.4698535,0.42183927,0.6001778,0.6927767,0.8505377,1.1660597,1.4061309,0.99801,1.2860953,1.3752645,1.3546871,1.3375391,1.471293,1.488441,1.3821237,1.5124481,1.8039631,1.7593783,1.704505,1.4678634,1.2929544,1.3066728,1.5227368,1.5776103,1.5810398,1.5707511,1.6016173,1.7422304,1.6667795,1.5227368,1.4129901,1.3649758,1.3101025,1.3101025,1.2243627,1.1454822,1.0768905,0.922559,1.0014396,1.0871792,1.0185875,0.8265306,0.7305021,0.66876954,0.7133542,0.8265306,0.9328478,0.8848336,0.9945804,0.980862,0.9362774,0.9294182,1.0117283,0.97057325,0.89512235,0.83681935,0.8265306,0.8779744,0.8848336,0.84024894,0.8025235,0.8265306,0.97400284,0.90541106,0.86082643,0.7922347,0.6962063,0.6241849,0.5521636,0.53501564,0.5624523,0.5521636,0.34638834,0.23664154,0.1920569,0.16804978,0.15776102,0.15090185,0.20577525,0.25721905,0.28808534,0.30866286,0.34981793,0.4389872,0.52815646,0.6379033,0.7613684,0.85739684,0.7510797,0.7099246,0.70649505,0.70306545,0.6344737,0.5796003,0.5727411,0.5418748,0.47671264,0.40126175,0.37382504,0.31552204,0.25721905,0.22635277,0.23664154,0.19548649,0.116605975,0.058302987,0.037725464,0.01371835,0.020577524,0.024007112,0.030866288,0.048014224,0.07888051,0.16119061,0.2469303,0.39440256,0.6036074,0.84024894,0.9911508,1.1351935,1.2517995,1.3169615,1.3238207,1.2620882,1.2723769,1.2929544,1.2929544,1.2586586,1.2415106,1.2998136,1.3649758,1.430138,1.5433143,1.5913286,1.6153357,1.6633499,1.7216529,1.704505,1.704505,1.6839274,1.6290541,1.5227368,1.3306799,1.3752645,1.4575747,1.5536032,1.6324836,1.6839274,1.8759843,2.153781,2.428148,2.7162333,3.1277838,3.3781435,3.4673128,3.450165,3.350707,3.1517909,3.0489032,3.1483612,3.4433057,3.8857226,4.3590055,4.8254294,5.3878818,5.909179,6.169828,5.871454,5.8474464,6.094377,7.14726,9.3936405,13.059869,0.09602845,0.09259886,0.12346515,0.12003556,0.08916927,0.14747226,0.34295875,0.39097297,0.38754338,0.37725464,0.35324752,0.37725464,0.4664239,0.5727411,0.6824879,0.84367853,0.97400284,1.1832076,1.2072148,1.1454822,1.4644338,1.6804979,1.9171394,2.4658735,3.4707425,4.9214582,6.193835,7.3564653,7.699424,7.3290286,7.143831,7.699424,8.464222,8.848335,8.930646,9.455373,10.6488695,13.37882,16.561478,19.45262,21.647556,24.254042,24.562706,22.041958,18.163095,16.383139,15.803539,17.233677,18.578075,18.427174,16.050468,15.529172,14.802099,15.278812,17.12736,19.305147,22.590693,30.952026,46.72127,64.826065,72.82043,70.978745,72.94389,76.27746,75.337746,61.26958,46.018204,33.26014,24.696459,20.27572,18.20768,15.285671,12.71691,11.050131,9.952662,8.196714,7.4765005,7.267296,6.636252,5.5319247,4.7842746,4.15666,3.5564823,3.0111778,2.5001693,1.9514352,1.9754424,1.605047,1.1043272,0.72021335,0.6790583,0.7133542,0.9842916,1.4095604,1.8245405,1.9857311,1.8245405,1.6324836,1.3924125,1.0563129,0.5761707,0.42526886,0.42869842,0.65162164,0.9362774,0.90884066,0.50757897,0.32581082,0.34638834,0.47671264,0.5418748,0.5418748,0.6207553,0.66533995,0.65505123,0.65162164,0.64133286,0.59674823,0.59331864,0.65848076,0.7682276,0.7133542,0.59331864,0.5796003,0.6927767,0.8196714,1.0048691,1.3615463,1.6736387,1.8828435,2.0680413,2.4830213,3.0214665,3.415869,3.6044965,3.7485392,5.0414934,6.4579134,7.5519514,7.98408,7.5416627,6.7631464,6.7665763,6.9860697,6.931196,6.1801167,4.6093655,3.1037767,2.1983654,1.9582944,1.9925903,2.5413244,3.192946,4.0709205,5.07236,5.8337283,6.2487082,6.783724,7.023795,6.8214493,6.327589,5.8371577,5.528495,5.5730796,5.888602,6.159539,6.5779486,7.5931067,8.1487,8.186425,8.628842,9.054111,8.371623,9.325048,12.21962,14.925565,14.092175,14.29795,15.738377,17.638369,18.241976,15.206791,15.004445,16.901007,19.949911,22.998814,24.391226,25.426962,25.876238,25.958548,26.34952,28.283808,33.832882,38.219322,40.48628,43.511177,36.706875,28.35583,22.837624,21.332033,21.839613,21.177702,21.150267,21.554956,22.498095,24.408375,25.824793,24.974257,22.463799,20.052797,20.652975,18.945042,19.078794,19.819586,19.805868,17.55263,18.687822,16.616352,14.678635,14.452282,15.738377,14.143619,14.006435,14.784951,15.597764,15.223939,15.837835,16.921585,20.2037,25.029129,28.359259,19.006773,11.115293,6.807731,5.3878818,3.3369887,2.7882545,3.1963756,3.923448,4.7534084,5.9126086,4.5442033,7.143831,7.613684,5.1752477,4.372724,6.217842,5.0174866,4.0846386,4.8494368,6.8557453,8.309891,10.333347,13.042721,14.023583,8.357904,8.251588,9.712592,15.169065,19.562366,10.371073,13.059869,15.042171,16.928444,17.765263,15.031882,13.282792,15.501736,17.720678,20.104242,26.953129,24.374079,25.152594,28.294096,32.66682,37.015537,32.41989,30.766829,32.43018,35.681427,36.65886,47.420906,45.39059,36.230164,27.402405,28.167202,32.5948,33.884323,34.09353,33.92205,32.704548,44.24511,61.43763,66.73634,56.19722,39.48484,38.119865,38.219322,38.363365,40.040432,47.626682,47.520363,42.468582,39.56715,42.88699,53.46384,59.46562,55.20607,53.189472,57.061478,61.615967,55.007153,44.40973,32.317,20.388897,9.445084,9.568549,11.132441,12.816368,15.573756,22.652426,30.845709,28.92857,22.570116,16.46545,14.318527,12.826657,10.100135,9.510246,11.022695,11.201033,13.443983,14.105893,12.771784,10.446524,9.571979,7.486789,7.6342616,10.021255,13.197053,14.280802,16.914726,14.96329,13.207341,14.064738,17.576635,18.362011,20.35803,24.500973,29.569902,32.220974,35.02638,27.93399,20.714708,17.569777,17.12736,19.233126,32.118088,41.796383,39.659748,22.456938,14.5243025,10.672876,9.22216,9.047252,9.582268,10.302481,11.314209,12.233338,12.325937,10.525404,11.122152,11.790922,11.194174,10.203023,11.897239,12.517994,9.743458,8.577398,11.962401,20.776442,19.915615,14.232788,11.0981455,12.22305,13.663476,12.812939,13.183334,12.895248,11.47197,9.853205,11.218181,12.761495,13.296511,12.0138445,8.491658,5.720552,5.446185,4.839148,3.923448,5.562791,4.2389703,3.549623,3.5187566,4.15323,5.4633327,4.866585,4.911169,5.1752477,5.1855364,4.4275975,3.1552205,2.7573884,2.6956558,2.719663,2.867135,2.2360911,3.1895163,4.2081037,4.756838,5.2506986,7.4113383,8.073249,7.6274023,6.7871537,6.550512,5.5319247,5.178677,6.166398,7.517656,6.6053853,5.6485305,5.360445,5.3878818,5.7411294,6.800872,5.1100855,3.474172,3.940596,5.8817425,5.98463,2.7402403,2.085189,2.644212,3.7965534,5.662249,4.4275975,3.7794054,5.267846,7.1712675,4.506478,3.9131594,4.057202,3.3644254,2.0920484,2.301253,3.2272418,3.625074,4.461893,5.994919,7.7680154,7.8434668,7.1541195,5.8543057,4.417309,3.625074,2.6407824,2.8225505,4.040054,5.2575574,4.557922,5.1409516,5.813151,6.101236,5.597087,3.9508848,5.425607,5.909179,5.6999745,4.6093655,1.9720128,1.6084765,1.6427724,1.7079345,1.704505,1.8142518,2.4007113,2.5207467,2.2498093,1.9891608,2.4624438,2.9117198,3.3198407,3.4295874,3.2443898,3.0248961,3.2032347,3.2203827,3.4878905,4.016047,4.40359,4.4241676,4.7259717,5.15467,6.7459984,11.736049,14.363112,15.8138275,20.913624,27.85854,28.228935,8.803751,1.5810398,0.0034295875,0.017147938,0.0548734,0.058302987,0.09259886,0.22978236,0.39783216,0.39783216,0.16462019,0.0548734,0.048014224,0.14404267,0.37039545,0.4664239,0.490431,0.5144381,0.58988905,0.7476501,0.72364295,0.85739684,1.1317638,1.4095604,1.4267083,1.7216529,1.6633499,1.5364552,1.488441,1.488441,1.6187652,1.5913286,1.8485477,2.294394,2.3081124,2.054323,1.7079345,1.4610043,1.3992717,1.5090185,1.5055889,1.4815818,1.4781522,1.5124481,1.5707511,1.5501735,1.488441,1.3752645,1.2620882,1.2620882,1.3375391,1.2723769,1.1592005,1.0528834,0.9774324,1.0528834,1.1866373,1.1660597,0.9911508,0.88826317,0.77851635,0.72707254,0.78537554,0.89855194,0.90884066,1.0014396,0.9911508,0.97400284,1.0151579,1.1454822,1.0871792,0.94999576,0.88826317,0.9294182,0.97057325,0.9911508,1.0151579,1.0048691,0.97057325,0.980862,0.85739684,0.922559,0.922559,0.8162418,0.764798,0.7305021,0.6824879,0.6344737,0.5727411,0.45613512,0.34638834,0.2709374,0.20920484,0.15776102,0.1371835,0.16804978,0.19891608,0.23664154,0.2777966,0.31895164,0.4115505,0.5418748,0.6927767,0.84367853,0.96714365,0.8676856,0.83338976,0.7956643,0.72021335,0.6173257,0.6173257,0.65162164,0.65505123,0.61046654,0.5658819,0.5007198,0.4664239,0.42869842,0.3841138,0.36696586,0.33609957,0.26750782,0.19548649,0.12346515,0.041155048,0.030866288,0.01371835,0.006859175,0.010288762,0.017147938,0.041155048,0.07545093,0.14061308,0.25721905,0.4664239,0.6344737,0.8505377,1.0528834,1.196926,1.2826657,1.2758065,1.3889829,1.4781522,1.4918705,1.4850113,1.3752645,1.3169615,1.3101025,1.3752645,1.5501735,1.6359133,1.6084765,1.6290541,1.704505,1.6804979,1.6873571,1.6530612,1.5364552,1.3478279,1.1729189,1.3238207,1.4472859,1.5055889,1.5090185,1.5501735,1.6427724,1.8519772,2.054323,2.2463799,2.5721905,2.8328393,3.0557625,3.1860867,3.2272418,3.2375305,3.2032347,3.1517909,3.2992632,3.6936657,4.2286816,4.7191124,5.219832,5.658819,5.857735,5.5113473,5.627953,6.159539,7.14726,8.64256,10.714031,0.06859175,0.0548734,0.07888051,0.08916927,0.08573969,0.1371835,0.2469303,0.23664154,0.22635277,0.26064864,0.30866286,0.34638834,0.45613512,0.53501564,0.61046654,0.84367853,1.0151579,1.2929544,1.3341095,1.2277923,1.4644338,1.7216529,2.095478,2.6476414,3.3678548,4.1635194,5.3913116,6.632822,6.773435,6.036074,5.970912,7.1987042,8.320179,9.098696,9.482809,9.568549,10.803201,14.435134,18.674105,22.374628,25.035988,29.75167,29.978024,25.93797,20.234566,17.840714,17.566347,18.897026,20.11796,20.553518,20.546658,21.551527,20.800447,19.764713,19.552078,20.886189,26.291218,37.83864,56.330975,75.26916,80.85938,72.1208,64.20874,57.493603,51.03569,42.57147,31.418451,23.129137,17.929884,15.13134,13.121602,11.533703,10.419086,10.017825,9.592556,7.4524937,6.420188,5.7754254,5.1683884,4.530485,4.0777793,3.1620796,2.5619018,2.3252604,2.1572106,1.4541451,1.2826657,1.0460242,0.75450927,0.50757897,0.47328308,0.53158605,0.66533995,0.89855194,1.1592005,1.2860953,1.4472859,1.6736387,1.7182233,1.4644338,0.9328478,0.6344737,0.5178677,0.6036074,0.8162418,0.980862,0.548734,0.4389872,0.53844523,0.69963586,0.7339317,0.48014224,0.4424168,0.48357183,0.52815646,0.5727411,0.4972902,0.44927597,0.45270553,0.5144381,0.6241849,0.7407909,0.75450927,0.7305021,0.72364295,0.764798,0.83338976,0.9259886,1.0460242,1.2826657,1.8279701,2.8396983,3.9303071,4.671098,5.038064,5.422178,6.5813785,7.8983397,8.868914,9.304471,9.328478,7.939495,6.5779486,5.1752477,3.7862647,2.5824795,1.8691251,1.605047,1.6873571,1.9411465,2.1469216,2.7059445,3.2786856,3.998899,4.835718,5.6039457,6.0635104,6.9654922,7.8023114,8.186425,7.8434668,7.2295704,7.689135,8.529384,9.050681,8.567109,7.010077,7.7920227,8.330468,8.093826,8.591117,8.824328,7.8366075,7.7611566,8.872343,9.592556,8.22758,7.500508,8.285883,10.528833,13.234778,15.405707,17.851004,21.002794,24.329493,26.34266,24.703318,25.090862,25.53328,25.238335,24.600431,27.371538,34.64569,37.783764,36.09984,36.854347,30.653652,24.669024,20.162544,17.878439,18.04649,19.089085,19.991066,20.433481,20.875898,22.563255,22.343761,21.822466,19.847023,17.586924,18.519772,18.005335,18.355152,19.524641,20.124819,17.412016,17.641798,16.012743,13.869251,12.610593,13.718349,14.109323,13.008426,12.1921835,12.895248,15.7966795,15.79325,17.058767,17.171944,15.786391,14.637479,14.5414505,10.377932,6.944915,5.501058,3.765687,2.7128036,2.4212887,3.0351849,4.0709205,4.413879,4.3178506,5.2815647,5.5147767,4.256118,1.786815,5.6073756,5.744559,5.254128,5.363875,5.4667625,7.034084,9.235879,12.017275,13.543441,10.203023,8.186425,12.538571,19.843594,23.756752,15.028452,15.426285,16.839275,19.967058,22.542679,19.339443,16.660936,19.665255,22.103691,22.223726,22.796469,28.043737,29.199507,31.065203,36.05868,44.238247,47.228848,46.834446,47.32488,46.69726,36.67944,42.98645,44.53662,41.3231,37.385933,40.798374,40.870396,39.200184,39.107586,42.019306,47.47578,55.326103,69.63777,75.588104,68.303665,52.829365,53.223766,54.050297,52.585865,50.0514,51.587856,48.607544,41.690063,40.07816,48.06567,64.99411,71.42116,65.628586,61.10496,64.3082,74.65183,70.65293,52.06114,32.052925,17.55263,9.208443,12.240198,15.46744,17.988186,20.45406,25.056566,25.464687,19.301718,14.081886,13.612033,17.974468,16.87014,11.592006,9.074688,10.100135,9.321619,12.13731,12.377381,11.149589,8.934075,5.610805,3.8788633,4.0674906,6.924337,12.181894,18.554068,21.400625,17.62465,14.466,14.863832,17.466888,17.357141,19.401176,24.600431,31.25726,34.978363,31.360147,23.753323,17.902447,16.033321,16.846134,20.70442,36.555973,46.680115,41.950714,21.85333,11.650309,7.888051,7.6925645,8.855195,9.825768,9.640571,10.957532,11.773774,10.854645,7.7268605,9.571979,11.032983,11.022695,10.429376,12.113303,14.634049,11.602294,9.908078,12.30536,17.405157,16.204802,13.941273,13.347955,14.335675,14.009865,11.592006,10.906088,10.422516,9.846346,10.124143,11.482259,14.081886,14.280802,11.170166,6.574519,5.717122,6.2384195,5.9812007,5.336438,7.226141,5.346727,3.2786856,2.095478,2.1400626,3.0283258,3.5187566,3.8685746,4.249259,4.496189,4.125794,3.4604537,3.7965534,3.7794054,3.0557625,2.2978237,2.352697,3.5702004,3.923448,3.1449318,2.7299516,4.90431,5.2815647,4.887162,4.5784993,5.038064,5.2472687,5.086078,5.254128,5.802862,6.142391,7.5279446,7.5416627,6.375603,5.5319247,7.798882,4.3761535,2.877424,3.782835,5.686256,5.305572,2.585909,1.7079345,2.3046827,3.8102717,5.453044,4.866585,3.899441,3.2649672,3.07634,2.8534167,4.482471,5.4187484,4.15323,1.8554068,2.3561265,3.3952916,3.9440255,5.3501563,8.069819,11.667457,10.556271,8.48137,5.720552,3.2203827,2.5927682,4.0023284,5.3570156,6.341307,6.39961,4.722542,5.521636,4.8117113,4.530485,4.98662,4.856296,6.948344,5.7068334,3.7348208,2.4727325,2.201795,1.7353712,1.5501735,1.587899,1.7250825,1.7696671,1.8176813,2.07833,2.0474637,1.8348293,2.1743584,2.5241764,3.0523329,3.5118976,3.7313912,3.6319332,4.201245,4.280125,4.5270553,4.972902,5.0003386,5.3878818,6.427047,7.490219,8.587687,10.38479,16.585485,22.69701,35.465363,49.907356,49.320896,14.853543,2.5001693,0.010288762,0.058302987,0.26064864,0.14061308,0.07888051,0.116605975,0.24007112,0.37039545,0.20577525,0.08573969,0.06516216,0.20577525,0.5624523,0.4629943,0.47671264,0.6276145,0.7922347,0.70306545,0.7133542,0.84024894,1.0220171,1.3169615,1.8759843,2.061182,1.6187652,1.313532,1.3786942,1.5227368,1.7902447,1.8142518,1.9823016,2.311542,2.4212887,2.1674993,1.8554068,1.5810398,1.4061309,1.3546871,1.3684053,1.3546871,1.3306799,1.3341095,1.4198492,1.4164196,1.4575747,1.4267083,1.3272504,1.2620882,1.4267083,1.3992717,1.2963841,1.2037852,1.1797781,1.1420527,1.214074,1.2209331,1.1283343,1.0425946,0.922559,0.8128122,0.77508676,0.8128122,0.8471081,0.881404,0.91569984,0.96371406,1.0460242,1.1832076,1.0906088,0.99801,1.0185875,1.097468,0.9911508,1.0528834,1.1866373,1.2312219,1.155771,1.039165,0.9259886,0.96371406,0.9431366,0.8471081,0.8711152,0.86082643,0.75450927,0.64133286,0.5693115,0.5453044,0.48014224,0.39440256,0.3018037,0.2194936,0.17490897,0.1371835,0.14061308,0.16462019,0.19891608,0.24007112,0.34638834,0.5144381,0.7099246,0.8779744,0.9431366,0.9259886,0.94656616,0.90541106,0.7990939,0.70649505,0.67219913,0.6756287,0.6927767,0.70649505,0.7339317,0.6379033,0.66191036,0.65162164,0.5590228,0.4698535,0.4629943,0.4389872,0.37039545,0.25378948,0.12346515,0.1097468,0.06859175,0.030866288,0.010288762,0.0034295875,0.0,0.006859175,0.017147938,0.05144381,0.15090185,0.31209245,0.5418748,0.77851635,0.96714365,1.0563129,1.2312219,1.4610043,1.6359133,1.7456601,1.8691251,1.7662375,1.5330256,1.3958421,1.4541451,1.6667795,1.7902447,1.7490896,1.6873571,1.6633499,1.6256244,1.6153357,1.6016173,1.4918705,1.3341095,1.3101025,1.5261664,1.6256244,1.6221949,1.5604624,1.546744,1.5158776,1.5364552,1.5981878,1.7010754,1.8279701,2.1126258,2.4418662,2.6922262,2.8911421,3.216953,3.3541365,3.3198407,3.3369887,3.5153272,3.8479972,4.437886,4.9008803,5.188966,5.302142,5.271276,5.4736214,5.9228973,6.691125,7.7440085,8.934075,0.044584636,0.06859175,0.10288762,0.09602845,0.07545093,0.1371835,0.2469303,0.274367,0.29151493,0.29494452,0.19891608,0.2469303,0.607037,0.7305021,0.59674823,0.7339317,0.8676856,1.1832076,1.4267083,1.5021594,1.4644338,1.6221949,1.9274281,2.3492675,2.843128,3.357566,6.6636887,9.716022,9.1810055,5.809721,4.4550343,6.0669403,7.8537555,9.122703,9.798331,10.422516,12.05843,16.081335,20.817596,25.084003,28.198069,35.863197,36.52511,31.020618,22.892496,18.403166,19.233126,20.234566,21.60983,23.832203,27.663052,25.210897,24.826784,23.708738,21.764162,21.606401,27.3441,36.32276,45.89474,53.919975,58.7797,55.45643,47.781013,38.89838,30.9143,24.85765,18.814716,15.46401,13.101024,10.950673,9.156999,9.266746,9.266746,8.886061,8.244728,7.8434668,5.5593615,4.852866,4.863155,4.8940215,4.3933015,3.8205605,2.8534167,2.2429502,2.1160555,1.9685832,1.3443983,1.097468,0.823101,0.51100856,0.53501564,0.53501564,0.65162164,0.90884066,1.1626302,1.1146159,0.85739684,0.94999576,1.1694894,1.4575747,1.9239986,1.2037852,0.96714365,0.864256,0.72364295,0.5658819,0.37039545,0.3018037,0.48357183,0.78537554,0.8093826,0.4046913,0.22292319,0.23664154,0.37725464,0.548734,0.5007198,0.4972902,0.47328308,0.41498008,0.36696586,0.42869842,0.45956472,0.45956472,0.44927597,0.47328308,0.4115505,0.34981793,0.48357183,1.0597426,2.3664153,3.9508848,5.1100855,6.7871537,8.4264965,7.949784,8.412778,10.268185,12.586586,14.29795,14.174485,11.72233,8.453933,5.4187484,3.1312134,1.5570327,0.97057325,0.9534253,1.1763484,1.5638919,2.2566686,2.2566686,2.5961976,3.2855449,4.040054,4.273266,3.8342788,3.8137012,4.4859004,5.5730796,6.2555676,6.708273,8.165848,9.942374,11.080997,10.360784,6.883182,5.305572,5.288424,6.3207297,7.7371492,8.711152,7.857185,7.431916,7.346176,5.171818,7.284444,8.772884,10.343636,12.380811,14.970149,19.473198,21.578964,23.27661,24.86451,24.963966,25.989414,27.755651,28.328392,27.152044,25.039417,25.564144,31.106358,33.8123,31.126936,25.817934,22.316326,17.686382,13.6086035,12.593445,17.974468,21.85676,21.095392,20.45063,21.733295,23.835632,19.696121,18.71526,18.636377,18.557497,18.934752,17.826996,17.007324,18.900457,21.404055,17.912735,16.94902,17.010754,16.345413,14.658057,13.107883,14.095605,13.245067,11.976119,11.4754,12.696333,18.492336,19.613811,19.661825,19.164536,15.563468,13.37882,8.841476,5.055212,3.6319332,4.6676683,3.1552205,2.054323,1.8588364,2.3492675,2.5927682,4.2183924,4.1120753,4.417309,4.7259717,2.0920484,5.336438,8.282454,8.735159,7.298162,7.3701835,8.529384,9.112414,9.637141,10.251037,10.72775,10.371073,10.6145735,13.039291,17.984756,24.548986,18.814716,18.28656,22.20315,27.896265,30.777119,20.460918,24.905664,27.906553,24.61415,21.513802,29.292107,29.587051,31.967184,40.623463,54.38297,70.309975,67.48056,60.8546,55.28152,45.517487,50.2023,52.70247,50.895077,49.818188,61.660553,57.874287,46.584087,38.521126,40.359386,54.70192,72.96447,78.91138,81.18176,81.8231,76.291176,73.47205,72.04534,67.37082,59.472477,53.03857,42.64006,36.08612,38.42167,50.9671,71.30455,74.638115,70.39914,64.140144,64.887794,85.112076,77.61842,54.54073,30.046616,13.701202,10.4533825,10.086417,12.6757555,17.549198,21.928782,20.965069,14.898128,11.358793,10.686595,11.845795,12.421966,12.956982,11.115293,11.187314,12.521424,9.506817,10.432805,8.872343,7.3393173,6.1629686,3.4638834,2.3149714,2.568761,5.425607,9.595985,11.293632,13.454271,16.684942,18.36887,18.04306,17.394867,13.7697935,14.867262,20.845032,29.401854,35.798035,29.85113,23.310905,17.86815,15.453721,18.248835,23.585274,33.393894,38.692604,33.74371,16.067617,10.854645,7.922347,7.3839016,8.399059,9.156999,8.862054,9.815479,11.091286,11.180455,7.9943686,9.949233,10.124143,9.80862,10.062409,11.732618,14.675205,13.214201,12.562579,14.743796,18.602083,15.87899,14.685493,15.806969,17.549198,15.731518,13.313659,12.994707,12.30536,11.273054,12.421966,11.626302,12.079007,11.372512,8.906639,5.888602,8.158989,9.825768,9.472521,7.4456344,5.861165,3.9303071,2.7539587,2.136633,2.1983654,3.357566,3.4192986,3.07634,3.340418,4.016047,3.724532,4.6402316,6.368744,6.1492505,3.9337368,2.3972816,4.5201964,6.790583,6.210983,3.316411,2.1812177,4.012617,3.6010668,2.7299516,2.486451,3.2821152,4.3178506,4.2835546,4.0777793,4.3624353,5.56965,8.879202,8.477941,6.495639,4.9934793,5.9812007,3.2718265,1.7971039,2.9220085,5.038064,3.5873485,1.6942163,1.1489118,1.9411465,3.415869,4.256118,3.6113555,2.3218307,1.7902447,2.4384367,3.707384,6.3824625,5.336438,3.0969174,1.5124481,1.7696671,3.0523329,2.668219,3.0900583,5.528495,9.932085,8.042382,5.7651367,3.707384,3.0351849,5.4633327,8.601405,11.351934,11.451392,8.433355,3.6456516,4.0366244,2.5413244,3.0420442,4.90431,2.976882,4.8425775,4.8425775,3.450165,1.99602,2.6545007,2.1194851,1.7559488,1.7010754,1.8691251,1.9514352,1.4541451,1.4815818,1.6187652,1.821111,2.4555845,2.3458378,2.620205,3.0797696,3.450165,3.3884325,4.3761535,4.852866,4.729401,4.2423997,3.9371665,4.6676683,6.591667,9.112414,11.286773,11.825217,17.429163,27.10403,41.535732,51.176304,36.271317,14.527733,3.666229,0.044584636,0.18519773,0.7476501,0.2469303,0.07545093,0.05144381,0.06516216,0.07545093,0.18519773,0.11317638,0.08916927,0.25721905,0.67219913,0.37725464,0.5693115,0.7099246,0.59331864,0.33609957,0.6276145,0.8471081,0.96371406,1.0460242,1.2655178,1.1077567,1.196926,1.4267083,1.7319417,2.061182,2.037175,1.8382589,1.8073926,1.9685832,2.0303159,1.9925903,1.8005334,1.5501735,1.3066728,1.097468,1.0631721,1.0425946,1.0254467,1.039165,1.1763484,1.3101025,1.3992717,1.4267083,1.3958421,1.2963841,1.3443983,1.4232788,1.471293,1.4369972,1.2655178,1.2655178,1.2655178,1.2312219,1.1420527,1.0082988,0.9945804,0.90884066,0.78194594,0.66533995,0.64133286,0.7133542,0.77851635,0.8505377,0.96371406,1.1592005,1.1351935,1.2106444,1.2723769,1.2483698,1.1146159,1.1249046,1.0940384,1.1523414,1.2929544,1.3443983,1.4164196,1.2586586,1.0220171,0.83681935,0.823101,0.66533995,0.6241849,0.6207553,0.59674823,0.53501564,0.4972902,0.4698535,0.44584638,0.4046913,0.31895164,0.18519773,0.106317215,0.082310095,0.09602845,0.106317215,0.14404267,0.23664154,0.42869842,0.6379033,0.6241849,0.7339317,0.8093826,0.85739684,0.8745448,0.84024894,0.66876954,0.5521636,0.52815646,0.58645946,0.67219913,0.6824879,0.7888051,0.823101,0.7613684,0.70306545,0.66533995,0.5555932,0.42183927,0.31895164,0.31895164,0.34638834,0.24007112,0.12346515,0.05144381,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.01371835,0.041155048,0.15433143,0.29151493,0.4081209,0.5178677,0.9568549,1.3341095,1.6496316,1.9411465,2.2566686,2.294394,1.9925903,1.7250825,1.6667795,1.8005334,2.0817597,2.1160555,2.0097382,1.845118,1.6633499,1.4198492,1.5124481,1.5981878,1.5776103,1.6016173,1.6153357,1.6256244,1.5947582,1.5844694,1.7559488,1.6942163,1.5947582,1.529596,1.4987297,1.4507155,1.4987297,1.7765263,2.0337453,2.2155135,2.4727325,3.059192,3.2306714,3.3644254,3.566771,3.6765177,3.9954693,4.4687524,4.839148,4.99005,4.928317,5.0620713,5.3707337,5.871454,6.6636887,7.9189177,0.06859175,0.09602845,0.08573969,0.06516216,0.06516216,0.1371835,0.22635277,0.29494452,0.31209245,0.2777966,0.19891608,0.51100856,0.52815646,0.5007198,0.607037,0.91569984,1.313532,1.2277923,1.1592005,1.2895249,1.4781522,1.6564908,2.1846473,2.7230926,3.0523329,3.07634,6.3447366,8.1487,6.9517736,3.9954693,3.2821152,5.1100855,7.023795,8.546532,9.716022,11.080997,12.2093315,16.071047,21.592682,26.548437,27.549875,37.259037,38.781776,32.42332,22.803328,18.87645,20.889618,23.039968,25.348082,27.879116,30.715385,30.42044,30.142645,28.976585,26.733635,23.948809,28.19464,35.66428,39.954693,39.91011,39.615166,40.0713,35.698574,29.525318,24.295198,22.43979,18.12537,15.018164,12.065289,9.352485,8.1041155,8.340756,8.330468,7.438775,5.8200097,4.400161,3.57363,2.9220085,2.7985435,3.0420442,2.9906003,2.867135,2.4727325,2.1126258,1.9823016,2.1743584,1.8073926,1.6084765,1.5433143,1.3786942,0.6790583,0.4664239,0.4938606,0.77165717,1.0734608,0.96714365,0.66191036,0.64476246,0.72364295,0.8848336,1.2998136,1.313532,1.2586586,1.1214751,0.91569984,0.69963586,0.42526886,0.26407823,0.26750782,0.39440256,0.5144381,0.28808534,0.22978236,0.23321195,0.23321195,0.2194936,0.29837412,0.4355576,0.52472687,0.52815646,0.48700142,0.45270553,0.36696586,0.41498008,0.4972902,0.22978236,0.14747226,0.22292319,0.48357183,0.85739684,1.155771,1.8931323,2.6990852,3.590778,4.588788,5.703404,7.750868,11.201033,14.599753,16.606062,15.995596,12.555719,8.621983,5.1100855,2.5584722,1.1420527,0.6927767,0.5624523,0.72364295,1.138623,1.7593783,2.0508933,2.6236343,3.083199,3.223812,3.0283258,2.5481834,2.469303,3.2683969,4.7191124,5.90232,7.191845,7.281014,7.2158523,7.1232533,6.1972647,4.184097,3.9337368,4.9214582,6.992929,10.360784,9.139851,8.81404,8.357904,7.425057,6.3447366,7.205563,10.038403,12.788932,14.726648,16.444872,17.87501,20.244854,22.186,23.396646,24.645016,26.35638,28.108898,29.302395,29.549326,28.678211,31.34986,34.607967,35.3419,32.85888,28.904564,24.94339,19.915615,16.256245,15.920145,20.36832,23.077694,19.630959,16.386568,16.722668,21.04052,18.053349,16.462019,17.000465,18.900457,19.87446,18.831865,16.808409,17.487467,19.895037,18.427174,16.280252,17.20967,18.550638,18.663815,16.928444,16.060759,14.064738,12.737488,12.634601,13.073587,14.095605,14.256795,14.171056,13.773223,12.343085,11.914387,11.022695,8.7317295,5.73427,4.3521466,2.9254382,1.7079345,1.3992717,1.9685832,2.644212,3.1140654,2.9906003,4.8734436,7.606825,6.276145,4.1326528,8.110974,10.696883,10.840926,13.96185,13.810948,14.009865,14.328816,15.055889,16.976458,16.640358,15.371411,16.11906,21.260014,32.58451,26.593021,19.637817,18.30028,22.690151,26.418112,21.04395,22.103691,24.206028,24.058556,20.440342,26.274069,29.67279,33.194977,42.16678,64.67173,86.25413,92.50969,88.06495,73.96591,47.63011,50.2366,55.219788,58.649376,62.552246,74.8919,71.33199,58.87573,50.243458,51.474678,61.890335,84.97832,92.02955,96.20336,101.45749,102.548096,100.27428,96.378265,89.23101,77.33034,59.27699,46.827587,39.56715,40.410828,50.143997,67.43598,65.72804,57.20552,52.092003,55.247223,66.17046,57.462738,37.848927,23.725885,18.636377,13.258785,19.689262,20.94792,18.825006,16.29054,17.473747,21.407484,15.817257,11.067279,9.904649,7.500508,6.7700057,6.7048435,9.349055,13.437123,14.376831,16.640358,12.80608,8.803751,6.48535,3.6113555,3.858286,3.5153272,3.9063,5.610805,8.460793,12.504276,17.63494,21.551527,21.829325,15.930434,14.112752,17.909306,28.376408,41.631763,48.857903,39.632313,29.079472,19.562366,13.560589,13.660047,19.562366,24.754763,26.35981,22.53239,12.442543,7.298162,4.5956473,4.496189,6.2555676,8.203573,8.340756,8.22758,7.6857057,7.5210853,9.5205345,11.629731,10.844356,9.650859,9.873782,12.648318,13.581166,12.500846,12.655178,14.531162,15.87899,11.849225,12.13731,14.891269,17.288551,15.536031,12.854094,12.80608,13.639469,14.04759,13.166186,11.777204,11.588576,10.285333,8.47451,9.6988735,10.151579,8.632272,7.2295704,6.3618846,4.7842746,3.4227283,2.8328393,3.275256,4.588788,6.1766872,3.7862647,2.620205,2.3046827,2.9288676,5.0174866,6.831738,6.2658563,4.547633,3.426158,5.178677,6.0806584,6.1801167,4.619654,2.5996273,3.3781435,4.770556,4.3658648,2.935727,2.0028791,3.8308492,5.9812007,5.295283,4.4447455,4.434457,4.616225,8.073249,7.2775846,5.2335505,4.0366244,4.8597255,3.9646032,4.2698364,4.7431192,4.331569,1.961724,1.6324836,3.841138,4.9591837,3.9474552,2.3767042,2.7642474,1.8245405,1.3615463,1.9137098,2.74367,3.981751,3.7348208,2.620205,1.6633499,2.3321195,4.7259717,4.4447455,3.0489032,2.4144297,4.722542,3.309552,2.5138876,2.8980014,3.7862647,3.2786856,7.870903,11.907528,10.683165,5.717122,4.770556,2.3972816,1.6599203,2.8054025,4.5613513,4.1463714,3.2512488,3.5942078,5.627953,7.6959944,6.012067,2.9460156,1.7971039,1.5398848,1.9857311,3.758828,2.0474637,1.6290541,1.5844694,1.7936742,2.9563043,3.1895163,2.8911421,2.884283,3.3198407,3.6696587,4.3624353,4.437886,3.8720043,3.275256,3.8891523,4.338428,5.1340923,6.1904054,7.0203657,6.7494283,8.182996,13.344524,17.809847,19.267422,17.53548,13.224489,6.4819202,1.728512,0.29837412,0.42869842,0.4664239,0.29151493,0.116605975,0.041155048,0.06516216,0.12346515,0.082310095,0.116605975,0.26407823,0.41498008,0.47328308,0.6379033,0.607037,0.39097297,0.31209245,0.4972902,0.5521636,0.66191036,0.8505377,0.97400284,1.039165,1.1900668,1.3169615,1.3752645,1.3992717,1.4644338,1.786815,2.095478,2.1400626,1.6770682,1.4815818,1.4267083,1.3615463,1.2963841,1.3924125,1.3066728,1.2037852,1.1592005,1.1797781,1.1866373,1.2826657,1.2963841,1.2998136,1.3101025,1.2620882,1.3478279,1.3615463,1.3409687,1.3238207,1.3409687,1.4095604,1.3889829,1.2929544,1.1592005,1.0563129,1.2380811,1.1729189,0.9568549,0.75450927,0.7990939,0.71678376,0.7133542,0.84024894,1.097468,1.4404267,1.3375391,1.2483698,1.1146159,0.9945804,1.0666018,1.2449403,1.2723769,1.2895249,1.2963841,1.1592005,1.155771,1.0460242,0.8676856,0.6756287,0.5555932,0.58302987,0.6036074,0.5727411,0.50757897,0.48357183,0.50757897,0.5693115,0.5727411,0.490431,0.3566771,0.24350071,0.16119061,0.116605975,0.09945804,0.082310095,0.09945804,0.16462019,0.30523327,0.48357183,0.58988905,0.5624523,0.64476246,0.7373613,0.764798,0.66876954,0.61389613,0.6241849,0.6379033,0.6379033,0.6344737,0.6276145,0.6893471,0.7373613,0.7407909,0.7373613,0.77851635,0.7339317,0.65162164,0.5727411,0.5041494,0.42183927,0.33266997,0.26750782,0.21263443,0.1371835,0.08573969,0.058302987,0.034295876,0.01371835,0.01371835,0.010288762,0.061732575,0.14747226,0.2469303,0.34638834,0.5418748,0.7099246,0.90198153,1.1626302,1.5364552,1.7422304,1.8897027,1.879414,1.7456601,1.6530612,1.786815,1.7422304,1.6359133,1.5673214,1.5913286,1.4438564,1.4541451,1.5055889,1.5398848,1.5536032,1.5741806,1.7353712,1.8519772,1.862266,1.8279701,1.6187652,1.4129901,1.3203912,1.3684053,1.4850113,1.4953002,1.5673214,1.6804979,1.821111,1.9720128,2.136633,2.3389788,2.620205,2.9734523,3.3472774,3.7142432,4.170378,4.5167665,4.7019644,4.804852,4.619654,4.6916757,5.0174866,5.535354,6.1492505,0.058302987,0.07545093,0.08916927,0.09945804,0.1097468,0.14747226,0.24007112,0.34638834,0.37039545,0.30866286,0.23664154,0.48014224,0.432128,0.47328308,0.6790583,0.8162418,1.0528834,0.9945804,0.939707,1.0528834,1.371835,1.5536032,2.0303159,2.6853669,3.1449318,2.7779658,3.7005248,4.1017866,3.4638834,2.3561265,2.4590142,4.07435,6.046363,7.9463544,9.496528,10.587136,11.718901,15.656067,21.45893,26.791937,27.909983,37.190445,37.807774,31.291555,22.419212,19.198832,21.249723,24.319204,27.529299,30.389574,32.786858,33.383606,34.968075,34.58739,31.120077,25.258911,27.721355,33.908333,36.57998,34.5188,32.51249,33.616817,29.741383,24.326063,20.083664,18.969048,15.206791,12.586586,10.566559,8.985519,8.080108,7.970361,7.31531,6.0086374,4.2869844,2.726522,2.2600982,2.037175,2.7299516,4.105216,5.0003386,5.9983487,5.778855,5.144381,4.5956473,4.3041325,3.7382503,3.6216443,3.474172,2.959734,1.8965619,1.2346514,0.83338976,0.67219913,0.66533995,0.6756287,0.52472687,0.50757897,0.5624523,0.7099246,1.0528834,1.1660597,1.1900668,1.1317638,1.0220171,0.91569984,0.70306545,0.48014224,0.4046913,0.4938606,0.6241849,0.37725464,0.23321195,0.16804978,0.16119061,0.20920484,0.22635277,0.30866286,0.36696586,0.3806842,0.4081209,0.34638834,0.30866286,0.36353627,0.41840968,0.23321195,0.17490897,0.20234565,0.30523327,0.42869842,0.4698535,0.75450927,1.0151579,1.3101025,1.7490896,2.4795918,4.064061,6.8111606,9.740028,11.897239,12.356804,9.314759,6.245279,3.8171308,2.1572106,0.84367853,0.61389613,0.6379033,0.90541106,1.3581166,1.8965619,2.417859,2.9906003,3.1895163,2.9254382,2.4144297,2.1983654,2.5001693,3.0523329,3.8274195,5.0449233,6.5539417,6.4304767,5.720552,4.928317,4.040054,3.5942078,4.3007026,5.754848,7.7542973,10.2921915,9.424506,9.043822,8.498518,7.4524937,5.878313,7.3427467,10.590566,14.812388,18.763273,20.76958,22.220297,24.703318,26.452408,27.652763,30.444448,31.751122,30.790836,30.18723,30.67766,31.106358,31.380726,32.961765,35.791176,38.24333,37.111565,30.735962,23.129137,18.45804,17.775553,19.044498,21.013083,18.732407,16.307688,15.786391,17.165085,16.2974,15.217079,15.4914465,17.326277,19.562366,20.800447,19.963629,19.342873,19.178253,17.648657,16.61292,16.12249,17.106783,18.900457,19.263992,17.765263,15.765814,14.589465,14.688923,15.649208,15.031882,13.622321,13.88983,15.29253,14.2533655,14.016724,14.987297,13.841815,10.062409,5.919468,3.9303071,2.4041407,1.5055889,1.3203912,1.8691251,2.4247184,2.5447538,4.7328305,9.379922,14.757515,11.228469,12.754636,13.107883,11.996697,15.05246,21.28402,21.60983,21.139977,22.384918,25.269201,23.845922,20.436913,17.833855,17.864721,21.390337,22.967947,19.689262,15.9921665,15.933864,23.18744,24.051697,23.52354,23.489244,24.127148,23.917942,29.950588,34.848038,38.356506,45.81586,68.15962,105.6896,113.09408,103.07282,81.80595,48.95393,48.47722,55.19578,61.77373,65.56686,68.63634,68.63976,64.291046,60.196117,61.485645,73.81501,93.17846,98.77212,106.01884,112.10293,96.00787,87.53679,85.67452,80.93484,70.11449,56.28639,46.714413,40.040432,39.546574,44.95846,52.441822,48.35718,44.944744,44.931026,46.879032,45.2294,36.130703,27.457277,21.253153,17.449741,13.834956,19.833303,19.901896,15.704081,12.281353,18.02934,20.934202,13.954991,7.7028537,5.6999745,4.40359,4.5853586,4.945465,7.363324,11.444533,14.514014,15.817257,13.605173,10.021255,6.4819202,3.673088,4.6916757,5.7239814,5.6313825,5.0449233,6.385892,11.965831,19.095943,23.039968,21.726437,15.755525,17.141079,24.717037,41.213352,59.153526,60.837452,45.695824,33.044075,22.731306,15.066177,10.847785,14.2533655,17.806417,19.654966,18.022482,11.214751,8.220721,6.667118,5.501058,5.171818,7.654839,9.613133,9.798331,7.613684,5.65539,9.729739,11.732618,10.7586155,10.278474,11.266195,12.2093315,12.394529,12.116733,13.13189,14.887839,14.510585,11.619442,11.797781,13.419975,14.733508,13.848674,11.622872,12.418536,13.704632,14.040731,13.094165,12.099585,12.4974165,12.229909,11.091286,10.714031,10.64201,8.577398,6.6396813,5.5730796,4.746549,4.482471,4.32471,4.6882463,5.6176643,6.7802944,4.0194764,2.8156912,2.3492675,2.7162333,4.945465,6.7528577,5.24041,3.4776018,3.3266997,5.4633327,5.6519604,4.5819287,3.5393343,3.4295874,4.7774153,4.8768735,3.6525106,2.3458378,2.1194851,4.057202,5.219832,4.7362604,4.523626,4.8322887,4.2698364,5.130663,4.547633,3.3438478,2.5001693,3.1483612,2.702515,3.4947495,4.4756117,4.448175,2.061182,3.1963756,8.508806,9.242738,4.712253,2.2841053,3.3678548,2.0474637,1.138623,1.4918705,1.9994495,2.270387,3.642222,3.474172,2.277246,3.724532,4.064061,3.1415021,1.9651536,1.4781522,2.5481834,1.6942163,2.0337453,2.750529,3.1209247,2.5207467,5.8508763,8.587687,7.1369715,3.083199,3.1826572,1.862266,1.7010754,3.350707,5.5593615,5.209543,3.40901,3.6799474,5.669108,7.706283,6.7974424,4.1155047,3.100347,3.0900583,3.7211025,4.9523244,3.3712845,2.4761622,2.218943,2.5207467,3.2649672,3.3129816,3.059192,3.0317552,3.3198407,3.5839188,3.5016088,3.3541365,2.819121,2.1880767,2.3561265,2.6545007,3.0523329,3.7108135,4.372724,4.3521466,3.8788633,5.844017,6.9346256,6.632822,7.226141,8.556821,6.7494283,3.5839188,0.8196714,0.18519773,0.4972902,0.42526886,0.20577525,0.034295876,0.07888051,0.08573969,0.0548734,0.11317638,0.2469303,0.32238123,0.5007198,0.61389613,0.5418748,0.35324752,0.29494452,0.4389872,0.52472687,0.6276145,0.7682276,0.91912943,1.1934965,1.2620882,1.2209331,1.2209331,1.4747226,1.587899,1.7456601,1.7422304,1.546744,1.2929544,1.2517995,1.2620882,1.2620882,1.255229,1.3101025,1.3512574,1.4850113,1.5604624,1.488441,1.2449403,1.2929544,1.1900668,1.2415106,1.4129901,1.3341095,1.313532,1.3272504,1.3375391,1.3478279,1.3855534,1.3169615,1.2312219,1.1832076,1.1900668,1.2312219,1.3409687,1.4027013,1.2860953,1.0563129,0.9842916,0.9431366,0.85396725,0.90884066,1.1111864,1.2998136,1.2517995,1.255229,1.2175035,1.1694894,1.255229,1.3924125,1.4129901,1.3684053,1.2758065,1.1146159,0.94999576,0.83338976,0.72364295,0.6036074,0.48014224,0.47328308,0.53158605,0.5658819,0.53844523,0.490431,0.53501564,0.5796003,0.58988905,0.5453044,0.44927597,0.39783216,0.3018037,0.216064,0.15776102,0.11317638,0.08916927,0.1097468,0.17490897,0.2777966,0.39783216,0.47328308,0.53501564,0.6001778,0.66191036,0.66191036,0.6241849,0.65505123,0.71678376,0.77851635,0.7990939,0.7956643,0.864256,0.9534253,0.9945804,0.91227025,0.91569984,0.8848336,0.83338976,0.77508676,0.7339317,0.66533995,0.59674823,0.4938606,0.37725464,0.30523327,0.22292319,0.17833854,0.13375391,0.07888051,0.041155048,0.017147938,0.024007112,0.061732575,0.12003556,0.20577525,0.31552204,0.42183927,0.5453044,0.7099246,0.94656616,1.0734608,1.3169615,1.488441,1.5536032,1.6359133,1.5707511,1.471293,1.3889829,1.3752645,1.4610043,1.4129901,1.3546871,1.3889829,1.4987297,1.5398848,1.4918705,1.6016173,1.7730967,1.8759843,1.7559488,1.5913286,1.4541451,1.3409687,1.2826657,1.3306799,1.4987297,1.4781522,1.5261664,1.704505,1.8656956,1.903421,1.9582944,2.1194851,2.4212887,2.8156912,3.1586502,3.7108135,4.046913,4.0846386,4.108646,3.957744,4.0023284,4.2938433,4.73969,5.1100855,0.044584636,0.06859175,0.10288762,0.12689474,0.14061308,0.15776102,0.24007112,0.34981793,0.37725464,0.32924038,0.31552204,0.45956472,0.39097297,0.4629943,0.6893471,0.75450927,0.72364295,0.8676856,0.9602845,1.0082988,1.2415106,1.2792361,1.430138,1.8554068,2.2978237,2.0680413,1.5501735,1.2655178,1.1763484,1.3478279,1.9274281,3.1106358,4.7191124,6.7357097,8.652849,9.493098,11.194174,15.265094,20.62211,25.543568,27.649334,36.689728,35.564823,29.161781,22.374628,20.100813,21.294308,24.061985,27.158903,29.820263,31.792276,35.019516,38.56914,38.167877,33.136673,26.383816,27.553307,32.35816,34.457066,32.50906,30.18037,30.783978,26.706198,21.434921,17.46003,16.276823,13.21763,11.396519,10.600855,10.22703,9.270175,8.320179,6.619104,4.8117113,3.292404,2.218943,2.3149714,2.9117198,4.232111,6.1561093,8.2310095,9.678296,9.482809,8.64942,7.7611566,6.9963584,6.0395036,5.5113473,5.0106273,4.2389703,2.9906003,2.2738166,1.4061309,0.8265306,0.6310441,0.5521636,0.45613512,0.39440256,0.42869842,0.58988905,0.8711152,0.97057325,1.0185875,0.9911508,0.9328478,0.9568549,0.939707,0.77165717,0.61046654,0.5418748,0.5521636,0.35324752,0.1920569,0.11317638,0.12346515,0.22292319,0.20234565,0.21263443,0.2469303,0.3018037,0.39097297,0.39440256,0.38754338,0.4629943,0.5555932,0.45270553,0.29837412,0.2469303,0.25378948,0.28465575,0.33609957,0.37039545,0.29494452,0.29151493,0.40126175,0.51100856,1.08032,2.301253,3.858286,5.3398676,6.2418494,4.5647807,3.117495,2.1434922,1.5193073,0.75450927,0.7305021,0.9431366,1.3478279,1.879414,2.4590142,2.9906003,3.391862,3.3369887,2.9494452,2.7813954,2.9322972,3.4673128,3.7176728,3.806842,4.65395,6.001778,5.8337283,5.0620713,4.273266,3.7485392,4.506478,5.6039457,6.9689217,8.477941,9.928656,10.412228,10.415657,9.650859,8.158989,6.2864337,7.9086285,10.645439,14.606613,18.756414,20.934202,22.985096,24.963966,26.428402,28.10204,31.878016,32.138664,31.26412,30.986322,31.747692,32.711407,30.002031,29.878567,34.155262,40.938984,44.632652,37.41337,26.843382,19.555508,17.103354,15.944152,18.11165,17.480608,16.170506,15.268523,14.850114,15.038741,14.754086,14.88098,16.026463,18.506054,22.168854,24.013971,22.837624,19.672113,17.751545,18.468328,17.182234,17.264544,19.54522,22.28546,21.11597,19.582945,17.679523,16.101913,16.245956,15.107333,13.88983,15.402277,18.410025,17.63151,15.429714,15.066177,14.747226,12.761495,7.500508,4.73969,3.2821152,2.2395205,1.4541451,1.488441,2.0131679,2.6956558,4.6848164,9.678296,19.929333,19.871029,16.763824,14.424845,14.284232,15.388559,24.902235,26.229485,24.672453,24.082563,26.874247,27.889406,24.645016,20.207129,15.913286,11.369082,18.067066,20.12139,17.700102,15.145059,20.985645,24.76848,25.996273,26.390675,26.843382,27.42641,32.18325,38.675457,43.775253,50.154285,66.31107,103.16199,109.44157,97.24938,75.21428,48.508083,45.702682,52.901386,58.237823,57.791977,55.6039,58.855152,61.75658,62.408203,64.352776,76.59984,87.88661,88.346176,90.86006,90.70916,65.59429,56.756245,57.61021,57.318695,51.663307,43.048183,36.295322,32.800575,33.10581,35.355618,35.31446,32.82458,33.8466,36.518246,36.81319,28.534168,21.990515,20.587814,21.356041,21.472647,18.259123,17.977898,16.108772,13.797231,13.896688,20.958208,16.856422,9.678296,4.8322887,3.7931237,4.1292233,5.2266912,6.1629686,7.0032177,8.498518,12.065289,14.023583,14.033872,11.454823,7.2604365,4.033195,5.1100855,6.8111606,8.011517,8.584257,9.407358,14.411126,19.905325,21.568676,19.010202,15.7795315,18.04649,26.833092,43.3054,59.222115,56.920864,40.770935,28.76052,19.737276,13.210771,9.321619,11.705182,14.5585985,16.770683,16.427725,10.782623,8.165848,8.412778,6.927767,4.2081037,5.8337283,8.838047,9.770895,7.888051,5.7377,9.156999,10.521975,10.1652975,10.768905,11.958971,10.299051,10.185875,11.074138,13.077017,14.994157,14.308239,12.905538,12.336226,12.147599,12.089295,12.103014,11.701753,13.413116,14.575747,14.009865,12.0138445,11.478829,12.600305,13.166186,12.1921835,9.945804,9.22902,8.471081,7.442205,6.3824625,6.001778,5.4324665,5.4084597,5.3878818,5.5250654,6.6465406,5.2918534,4.139512,3.4673128,3.433017,4.091498,5.23698,3.6765177,2.3801336,2.9460156,5.610805,4.32128,3.0557625,2.976882,3.998899,4.7808447,4.5270553,2.884283,1.9582944,2.3732746,3.2546785,3.3609958,3.5393343,4.4756117,5.3673043,3.9097297,2.9700227,2.6819375,2.218943,1.6736387,2.0646117,2.1297739,3.0557625,4.547633,5.1512403,2.2841053,3.9063,8.639131,8.64942,3.9371665,2.3321195,3.5393343,2.07833,0.96714365,1.1489118,1.4610043,1.8588364,3.4124396,3.6010668,2.6990852,3.7622573,2.860276,1.8759843,1.3169615,1.3238207,1.6873571,1.7559488,2.2292318,2.2429502,1.8279701,1.9102802,3.940596,4.839148,3.8925817,2.318401,3.275256,2.836269,2.2841053,3.3301294,5.31929,5.223262,3.6456516,3.673088,4.6882463,5.8062916,5.857735,5.195825,4.8768735,4.7602673,4.763697,4.880303,3.957744,3.018037,2.6167753,2.8054025,3.117495,2.9220085,2.7333813,2.668219,2.726522,2.784825,2.3595562,2.177788,1.9137098,1.5261664,1.2517995,1.313532,1.6427724,2.1880767,2.7779658,3.117495,2.3767042,2.5721905,2.877424,3.1449318,3.899441,4.9523244,5.003768,3.7485392,1.7216529,0.32581082,0.35324752,0.36353627,0.26407823,0.12346515,0.14747226,0.082310095,0.06859175,0.16119061,0.31552204,0.3841138,0.432128,0.48357183,0.432128,0.32238123,0.33266997,0.5007198,0.6241849,0.7099246,0.78194594,0.90541106,1.196926,1.2723769,1.255229,1.2929544,1.5913286,1.5981878,1.5673214,1.3924125,1.138623,1.0323058,1.1214751,1.1214751,1.1146159,1.1660597,1.2963841,1.3443983,1.5055889,1.6290541,1.5741806,1.2037852,1.2106444,1.1077567,1.1317638,1.2723769,1.255229,1.2449403,1.2415106,1.3066728,1.4232788,1.471293,1.2998136,1.1180456,1.0837497,1.2175035,1.3924125,1.4953002,1.6187652,1.5055889,1.2106444,1.1249046,1.1043272,0.9945804,0.9602845,1.0185875,1.0494537,1.1043272,1.2243627,1.2998136,1.3101025,1.2963841,1.3684053,1.3752645,1.3375391,1.255229,1.0837497,0.8676856,0.71678376,0.6276145,0.5658819,0.490431,0.4389872,0.5007198,0.61046654,0.67219913,0.5693115,0.5453044,0.5555932,0.5761707,0.5658819,0.490431,0.44927597,0.34981793,0.26750782,0.22635277,0.20577525,0.12689474,0.1097468,0.1097468,0.13032432,0.19548649,0.30866286,0.3806842,0.45956472,0.5521636,0.6241849,0.6001778,0.64133286,0.7407909,0.8505377,0.90884066,0.9294182,0.9842916,1.0563129,1.1043272,1.0460242,1.0357354,1.0323058,1.0117283,0.96714365,0.90884066,0.89855194,0.90198153,0.8265306,0.6790583,0.5727411,0.4698535,0.3806842,0.29494452,0.216064,0.15776102,0.08916927,0.044584636,0.030866288,0.05144381,0.09945804,0.17833854,0.26750782,0.37382504,0.50757897,0.66533995,0.6962063,0.8711152,1.0494537,1.2003556,1.4027013,1.3512574,1.3341095,1.3032433,1.2655178,1.2792361,1.2449403,1.1729189,1.1900668,1.2860953,1.3272504,1.2895249,1.3478279,1.5330256,1.7147937,1.6084765,1.4850113,1.4815818,1.4232788,1.3101025,1.3066728,1.4164196,1.3581166,1.3958421,1.5741806,1.7250825,1.7490896,1.704505,1.8313997,2.153781,2.4761622,2.8225505,3.3541365,3.5942078,3.4604537,3.2718265,3.2615378,3.3952916,3.7005248,4.098357,4.4104495,0.05144381,0.082310095,0.12003556,0.14404267,0.16462019,0.2194936,0.26750782,0.30523327,0.31552204,0.32581082,0.40126175,0.5144381,0.4046913,0.4115505,0.6036074,0.764798,0.61389613,0.8711152,1.0597426,1.0494537,1.0906088,0.9294182,0.7373613,0.7133542,0.8779744,1.0837497,0.8093826,0.6310441,0.64819205,0.939707,1.5501735,2.3252604,3.3541365,5.1340923,7.274155,8.48137,10.840926,14.808959,19.171394,23.070835,26.003132,34.861755,32.59137,26.949697,22.748453,21.815605,21.925352,23.125708,24.86451,26.881107,29.192648,35.98666,39.742058,37.972393,32.056355,27.244642,27.961426,31.452747,33.06808,31.514479,28.870268,28.880556,24.981115,20.20027,16.667795,15.594335,14.153908,13.423406,13.248496,12.953552,11.317638,8.913498,6.186976,4.1155047,3.1826572,3.357566,4.4687524,5.504488,6.3893213,7.7097125,10.707172,12.154458,12.377381,11.821788,10.744898,9.205012,7.970361,6.557371,5.3981705,4.417309,3.0283258,2.668219,1.7525192,1.1592005,1.0254467,0.72021335,0.48700142,0.31552204,0.29151493,0.42183927,0.6310441,0.8093826,0.8745448,0.8128122,0.72021335,0.8025235,0.96371406,0.90198153,0.6824879,0.41498008,0.25721905,0.1920569,0.12689474,0.09602845,0.11317638,0.17833854,0.2469303,0.26064864,0.31552204,0.41498008,0.47671264,0.5624523,0.5453044,0.6379033,0.78537554,0.66533995,0.39097297,0.36010668,0.4355576,0.5144381,0.53501564,0.42526886,0.33266997,0.3018037,0.31895164,0.28122616,0.20234565,0.20577525,0.37039545,0.66876954,0.9568549,0.7613684,0.7613684,0.7888051,0.7682276,0.7339317,0.8471081,1.1592005,1.611906,2.2052248,2.9906003,3.6868064,4.057202,3.7485392,3.1723683,3.5050385,3.9063,4.605936,4.866585,4.7259717,5.0277753,6.200694,6.0737996,5.535354,5.1855364,5.329579,7.0786686,8.196714,9.136421,10.124143,11.153018,12.830087,13.536582,12.548861,10.278474,8.272165,8.7145815,10.419086,12.686044,14.990726,16.993607,18.903887,19.86074,21.225718,23.729315,27.453848,26.562155,28.496443,30.406723,31.192099,31.500761,28.400414,27.392115,31.356718,40.304512,51.35464,45.613514,31.442457,19.898466,14.980438,13.63604,16.245956,16.11906,14.932424,14.126471,14.874121,14.400838,14.493437,15.326826,16.496315,17.014183,22.093403,26.980564,26.202047,20.982216,19.274282,21.500084,20.323736,20.04251,22.432932,26.737064,25.413242,23.914513,20.872469,17.12736,15.738377,15.086755,14.96672,16.780972,19.356592,18.962189,15.141628,12.171606,11.838936,12.319078,8.182996,5.504488,4.256118,3.4021509,2.6545007,2.4624438,2.2258022,3.316411,5.1855364,9.47938,20.04251,25.673891,18.358582,15.049029,18.506054,17.29884,24.02083,26.569014,24.267761,20.20027,21.20514,25.996273,25.900244,23.201159,18.770132,12.085866,17.648657,22.323185,23.067406,20.824455,20.502073,23.478956,27.639046,30.152933,30.355278,29.7551,30.42044,37.71517,44.684093,50.171436,58.807137,76.942795,83.65107,76.77474,60.635105,46.028492,44.035904,51.841644,52.589294,44.766407,42.22851,47.48264,51.683884,54.34524,57.05462,63.450798,66.36252,60.971207,54.430984,46.875603,31.397873,28.17406,29.823692,32.526207,32.457615,25.790497,19.898466,21.561817,23.643576,23.314335,22.065966,23.262892,24.473536,26.126596,25.996273,19.20569,16.969599,16.249386,21.678423,28.911423,24.627867,17.106783,13.570878,14.764374,18.972477,22.04539,11.297061,5.6519604,4.2081037,5.288424,6.4407654,7.3084507,8.381912,7.473071,6.2041235,10.0041065,14.092175,14.592895,11.976119,7.829748,4.839148,4.870014,5.7239814,8.961512,13.80409,17.144508,19.106232,19.274282,17.364002,14.819247,14.812388,16.273392,23.43094,33.534508,41.37797,39.303074,27.556736,18.36544,11.770344,8.282454,8.899779,11.832077,13.690913,15.230798,15.172495,10.179015,7.4936485,9.918367,9.3593445,4.98662,3.223812,5.693115,7.0923867,7.157549,6.8145905,8.152129,8.515666,9.246168,10.796341,11.523414,7.6857057,7.39762,9.582268,12.600305,14.88098,14.918706,13.978998,12.46998,10.957532,10.13786,10.827208,12.668896,15.066177,15.937293,14.424845,10.926665,11.080997,12.713481,13.166186,11.578287,8.872343,7.5245147,8.666568,9.373062,8.7317295,7.8263187,5.7411294,5.4976287,5.06893,4.5853586,6.3001523,7.0306544,5.720552,4.9694724,4.9591837,3.4604537,3.316411,2.0817597,1.3615463,2.3561265,5.8543057,3.1346428,2.3767042,2.8739944,3.8034124,4.245829,4.4584637,2.860276,2.2326615,2.7882545,2.1743584,2.1229146,2.7299516,4.180667,5.2335505,3.2032347,2.3218307,2.2360911,2.1469216,1.903421,1.9925903,2.9494452,3.7759757,5.1238036,5.662249,2.0749004,2.952875,4.48933,4.1635194,2.3767042,2.452155,2.8739944,1.7422304,0.88826317,0.91912943,1.2072148,2.2498093,2.6922262,2.8396983,2.7745364,2.3458378,1.9857311,1.7593783,1.529596,1.3306799,1.3615463,2.5721905,2.5893385,1.6976458,0.7956643,1.4027013,3.6970954,3.6765177,3.3541365,3.7794054,5.055212,3.9783216,3.0317552,3.0077481,3.7211025,4.029765,3.415869,3.532475,3.882293,4.1463714,4.187526,5.446185,5.9469047,5.411889,4.2835546,3.7279615,3.5770597,3.2135234,2.8637056,2.6579304,2.6407824,2.3664153,2.0886188,1.8416885,1.6907866,1.7079345,1.5330256,1.3546871,1.313532,1.3203912,1.08032,0.91569984,1.1489118,1.4575747,1.7353712,2.1091962,1.9548649,1.6427724,1.6221949,2.2806756,3.9508848,3.6113555,2.6785078,2.270387,2.1332035,0.6173257,0.15090185,0.15433143,0.26407823,0.29151493,0.22978236,0.10288762,0.116605975,0.25721905,0.4355576,0.4629943,0.31895164,0.31552204,0.30523327,0.29494452,0.44584638,0.6310441,0.7510797,0.83681935,0.8848336,0.864256,0.980862,1.1454822,1.2860953,1.3821237,1.4507155,1.2929544,1.2929544,1.2586586,1.1180456,0.9294182,1.0151579,0.97400284,0.94656616,1.0494537,1.3786942,1.3066728,1.2826657,1.3581166,1.4027013,1.1214751,1.1214751,1.097468,1.0117283,0.9259886,1.0014396,1.1351935,1.1180456,1.214074,1.4267083,1.4987297,1.3443983,1.138623,1.1077567,1.2895249,1.5227368,1.6873571,1.762808,1.5570327,1.214074,1.2003556,1.1283343,1.0700313,0.99801,0.9259886,0.9259886,1.0220171,1.1592005,1.255229,1.255229,1.1317638,1.1694894,1.1626302,1.1797781,1.1763484,0.9911508,0.89512235,0.7133542,0.5761707,0.52815646,0.5144381,0.48357183,0.5178677,0.66533995,0.8162418,0.7133542,0.58302987,0.5521636,0.5727411,0.5761707,0.4938606,0.4115505,0.31552204,0.26750782,0.2777966,0.31209245,0.18519773,0.14747226,0.116605975,0.082310095,0.07545093,0.09259886,0.18862732,0.3018037,0.40126175,0.48700142,0.5007198,0.5693115,0.66533995,0.7613684,0.83338976,0.89855194,0.91227025,0.91912943,0.94999576,1.0117283,1.0666018,1.1146159,1.1283343,1.0940384,0.99801,1.0082988,1.0906088,1.1043272,1.0117283,0.88826317,0.7888051,0.66191036,0.53501564,0.42526886,0.36353627,0.24350071,0.14747226,0.08573969,0.05144381,0.044584636,0.07888051,0.14404267,0.2503599,0.40126175,0.58302987,0.65505123,0.7133542,0.7510797,0.8025235,0.9568549,1.0837497,1.2346514,1.2826657,1.2037852,1.0940384,1.0494537,1.0117283,1.0014396,1.0082988,1.0185875,1.0666018,1.1351935,1.2929544,1.4610043,1.4267083,1.3203912,1.4267083,1.4850113,1.4369972,1.4267083,1.2826657,1.2209331,1.255229,1.3581166,1.4815818,1.4918705,1.4678634,1.6873571,2.1023371,2.3389788,2.7470996,3.1037767,3.1895163,2.9871707,2.6887965,2.7230926,2.9151495,3.210094,3.542764,3.841138,0.07545093,0.08916927,0.16462019,0.20920484,0.24350071,0.42869842,0.42869842,0.29151493,0.24007112,0.32581082,0.4115505,0.4972902,0.41840968,0.4046913,0.51100856,0.59674823,0.65505123,0.69963586,0.7305021,0.7613684,0.8093826,0.7339317,0.69963586,0.6001778,0.47328308,0.47328308,0.47328308,0.5007198,0.5178677,0.6344737,1.097468,1.7936742,2.7745364,4.166949,6.025785,8.347616,10.4705305,13.694343,17.075916,20.183123,23.087982,28.897703,27.988863,24.967398,23.050257,24.061985,23.976246,23.225166,22.913074,24.542128,29.998602,36.67601,36.799473,32.879456,28.208357,26.83995,27.889406,30.770258,32.694256,32.042637,28.379837,27.84482,24.53184,21.19485,18.999914,17.545769,18.842154,19.394318,18.680964,16.568336,13.320518,8.621983,5.48734,4.2423997,5.003768,7.689135,9.482809,8.999237,7.81603,7.716572,10.679735,13.474849,15.309678,15.762384,14.280802,10.192734,9.14328,6.958633,4.729401,2.9185789,1.3443983,1.1592005,1.2243627,1.2963841,1.2586586,1.097468,0.67219913,0.42869842,0.32924038,0.33952916,0.4115505,0.66876954,0.7613684,0.71678376,0.6310441,0.65505123,0.6790583,0.58645946,0.48700142,0.40126175,0.24350071,0.17147937,0.12346515,0.106317215,0.13032432,0.22978236,0.45956472,0.58302987,0.6379033,0.6241849,0.48700142,0.52472687,0.5624523,0.5624523,0.5178677,0.45613512,0.39783216,0.58302987,0.764798,0.7888051,0.59674823,0.44927597,0.47671264,0.52472687,0.52472687,0.48700142,0.48700142,0.38754338,0.26064864,0.16119061,0.1371835,0.23664154,0.4424168,0.5761707,0.5624523,0.42869842,0.5624523,0.8779744,1.1900668,1.6599203,2.8088322,4.722542,5.744559,5.127233,3.5290456,2.9906003,3.2478194,4.8117113,5.8062916,5.7994323,5.7994323,7.2638664,8.097256,8.114404,7.932636,8.958082,12.22648,13.584596,14.208781,14.754086,15.364552,17.29541,17.758404,16.849564,14.54831,10.72775,9.177576,10.134431,11.893809,13.759505,16.067617,16.969599,17.058767,18.739265,22.04539,24.658733,23.180582,24.94682,25.85566,24.6896,23.101702,24.590141,25.85223,30.276398,41.395123,62.864338,58.8723,38.212463,20.841602,14.623761,15.319967,16.698662,16.03675,14.5585985,13.910407,16.143068,14.020154,13.516005,16.365992,19.52807,15.182784,20.406046,27.361248,27.515581,21.897917,21.1194,24.487255,21.997374,22.20315,27.066305,31.93632,27.371538,24.315775,21.723007,19.802439,20.03565,22.683292,20.488356,17.61436,15.913286,14.922135,15.398848,13.786942,11.55428,9.547972,8.011517,7.963502,6.025785,4.5201964,4.4413157,5.4770513,3.9028704,4.2046742,6.444195,11.132441,19.226267,26.623888,19.428614,17.333136,22.727877,20.6907,23.400076,25.735624,24.02083,18.993055,15.806969,16.722668,21.181131,24.69303,25.039417,22.292318,23.098272,27.409264,28.990303,26.445549,23.225166,25.457829,27.865398,28.616478,28.911423,32.9892,27.717926,31.50762,35.22872,37.276188,43.5489,49.008804,59.709118,62.644844,54.561306,41.97815,46.944195,58.7797,55.96401,38.65145,28.640486,36.453087,35.962654,36.92637,39.584297,34.655983,32.810863,27.892836,23.911083,22.85477,24.658733,20.752434,19.932762,20.018501,19.589804,17.991615,12.205902,18.4649,19.003344,12.826657,15.731518,17.610931,17.734396,18.430603,19.301718,17.226818,16.54433,15.247946,18.804428,24.823355,23.039968,15.704081,13.697772,16.283682,19.178253,14.527733,5.127233,3.2889743,5.096367,7.8091707,9.873782,9.225591,7.332458,5.40503,5.8165803,12.116733,15.608052,13.512574,8.862054,5.086078,6.012067,3.1792276,2.7573884,6.9071894,15.179354,24.504402,22.004232,16.763824,12.120162,10.127572,11.567999,15.54632,21.318316,25.721907,27.474424,27.206917,18.71183,12.603734,8.824328,7.654839,9.705732,10.412228,10.563129,11.873232,12.912396,9.078118,12.363663,17.082775,17.412016,11.694893,2.4418662,3.3678548,4.4241676,5.7136927,6.831738,6.883182,6.4544835,8.076678,10.635151,11.396519,6.012067,5.8543057,9.0369625,12.843805,15.433144,15.824117,13.663476,10.9541025,8.858624,8.241299,9.644,11.571428,14.352823,15.055889,13.454271,12.037852,14.369971,16.657507,16.438013,13.413116,9.445084,9.153569,11.05699,12.178465,11.204462,8.484799,6.029215,5.2506986,4.122364,3.1380725,5.3090014,6.9209075,5.346727,5.470192,6.999788,4.4859004,2.201795,1.1008976,1.2106444,2.386993,4.3041325,3.059192,3.0214665,3.1072063,3.6593697,6.4544835,5.953764,3.7691166,3.0729103,3.8857226,3.0660512,3.642222,3.426158,3.2135234,3.0214665,2.1057668,1.7525192,1.9274281,2.318401,2.6167753,2.5173173,3.9337368,3.7005248,4.1155047,4.6402316,1.8931323,1.196926,3.0729103,3.9165888,3.3301294,4.1360826,2.452155,1.6187652,1.1111864,0.89169276,1.4027013,1.8313997,2.4418662,2.935727,2.836269,1.4815818,1.3821237,1.879414,1.9823016,1.6427724,1.7388009,3.74168,4.1772375,2.767677,1.0117283,2.1983654,6.835168,7.658269,7.2295704,6.3721733,4.149801,2.1846473,3.5873485,4.2423997,3.1140654,2.2600982,3.2958336,4.6093655,4.5030484,3.223812,2.9288676,3.8102717,4.7431192,4.3590055,2.9563043,2.5173173,3.2375305,3.9851806,4.040054,3.309552,2.335549,2.1400626,1.879414,1.5124481,1.2586586,1.587899,1.6359133,1.2003556,0.9842916,1.08032,0.94656616,0.94656616,0.75450927,0.6790583,0.8025235,0.9602845,1.3169615,1.313532,1.1592005,1.1454822,1.6324836,2.5241764,2.0886188,1.1283343,0.33609957,0.274367,0.10288762,0.024007112,0.17833854,0.40126175,0.22978236,0.09602845,0.16119061,0.30866286,0.40126175,0.30523327,0.26750782,0.26750782,0.31209245,0.42183927,0.64133286,0.6893471,0.85739684,1.0357354,1.0837497,0.84024894,0.7888051,0.86082643,0.9568549,1.0460242,1.1454822,1.0940384,1.1660597,1.1111864,0.939707,0.91569984,0.96371406,0.94999576,0.9294182,0.9774324,1.1592005,1.1351935,1.2586586,1.3375391,1.3169615,1.2655178,1.3272504,1.2517995,1.0871792,0.90198153,0.7922347,0.9774324,1.0666018,1.1283343,1.1797781,1.2037852,1.1214751,1.1797781,1.3203912,1.5090185,1.7559488,1.704505,1.6667795,1.5673214,1.4061309,1.2346514,1.1763484,1.1763484,1.1283343,1.0460242,1.0837497,1.0357354,1.0666018,1.1283343,1.1454822,1.0220171,1.0117283,0.9328478,0.89855194,0.89512235,0.8093826,0.9568549,0.75450927,0.5418748,0.4664239,0.5041494,0.490431,0.5144381,0.6379033,0.8128122,0.8848336,0.7613684,0.64133286,0.59331864,0.6036074,0.5796003,0.50757897,0.4046913,0.33266997,0.31209245,0.33609957,0.20234565,0.15776102,0.13375391,0.09945804,0.07545093,0.06516216,0.06859175,0.09945804,0.17147937,0.30523327,0.31895164,0.3841138,0.45270553,0.5041494,0.5658819,0.69963586,0.7133542,0.70306545,0.70649505,0.7339317,0.90198153,1.0014396,1.0323058,1.0220171,1.0220171,0.97400284,0.9602845,0.980862,1.0220171,1.0837497,1.0220171,0.980862,0.8745448,0.71678376,0.59674823,0.48357183,0.3841138,0.26407823,0.13032432,0.044584636,0.020577524,0.034295876,0.07545093,0.15433143,0.29151493,0.64476246,0.5693115,0.4629943,0.5041494,0.6241849,0.78537554,0.9431366,1.0700313,1.1180456,1.0082988,1.1283343,1.1043272,1.0666018,1.0666018,1.0666018,1.1043272,1.1489118,1.1763484,1.1797781,1.2037852,1.2655178,1.3924125,1.5124481,1.546744,1.3889829,1.255229,1.2483698,1.2175035,1.2003556,1.4198492,1.3821237,1.4198492,1.6084765,1.8862731,2.0440342,2.5207467,2.7128036,2.726522,2.6750782,2.702515,2.5310357,2.534465,2.7642474,3.1346428,3.4021509,0.06516216,0.048014224,0.10288762,0.15776102,0.18176813,0.15776102,0.14747226,0.16462019,0.26407823,0.40126175,0.38754338,0.5624523,0.5693115,0.53844523,0.53501564,0.5693115,0.5727411,0.5658819,0.6276145,0.7682276,0.90541106,0.91227025,0.7407909,0.52472687,0.37039545,0.34981793,0.52815646,0.5555932,0.5007198,0.4698535,0.6241849,1.4369972,2.428148,3.5873485,5.0449233,7.1026754,9.89093,12.236768,14.160767,16.256245,19.716698,23.11542,22.974806,21.812176,21.61326,23.808197,23.485815,22.412354,21.94936,23.732746,29.655643,33.07151,33.17097,30.75997,27.1932,24.35007,22.61813,24.898806,27.76594,29.069183,27.906553,27.786518,26.462696,25.581293,25.979126,27.690489,28.544456,27.368109,23.955667,19.219408,15.199932,11.760056,10.494537,9.088407,7.905199,9.983529,11.526843,11.533703,11.513125,12.288212,14.027013,13.461131,14.417986,15.309678,14.30138,9.314759,6.917478,4.8117113,3.199805,2.1023371,1.3684053,1.3409687,1.471293,1.605047,1.611906,1.4027013,1.0151579,0.7510797,0.64133286,0.64819205,0.6927767,0.84024894,0.90541106,0.78194594,0.52815646,0.37382504,0.33266997,0.30866286,0.28465575,0.26407823,0.28122616,0.34295875,0.39783216,0.4629943,0.53158605,0.5693115,0.490431,0.39440256,0.30866286,0.29151493,0.4389872,0.5727411,0.52472687,0.4698535,0.490431,0.5693115,0.6036074,0.66191036,0.65505123,0.58988905,0.5693115,0.4629943,0.34638834,0.26750782,0.23664154,0.2194936,0.18176813,0.12003556,0.07545093,0.058302987,0.06516216,0.12346515,0.22635277,0.31895164,0.4081209,0.53844523,0.72021335,0.89512235,1.5261664,2.5653315,3.4776018,4.7499785,5.192395,4.6402316,3.5770597,3.1380725,3.6970954,4.4721823,5.3330083,6.40304,8.093826,11.05356,13.262215,13.395968,12.627741,14.620332,14.7369375,15.6526375,16.609491,17.267973,17.686382,20.100813,21.479506,21.139977,18.766703,14.387119,12.624311,12.466551,14.123041,16.732958,18.37573,21.016512,20.382038,18.578075,17.604073,19.349733,20.985645,23.499533,24.94682,24.813065,24.0174,22.978235,25.663603,29.830551,36.73774,51.14887,50.027393,33.194977,19.250275,14.928994,15.086755,15.042171,14.997586,15.337115,16.599203,19.476627,16.139639,15.29939,17.089634,18.355152,12.63117,18.451181,25.10115,25.269201,19.977346,18.591793,18.893597,18.180243,19.678972,23.835632,28.27352,25.886526,23.406935,22.179142,21.839613,20.303158,19.260563,15.896138,11.423956,7.4765005,6.0875177,7.31531,8.23444,7.9909387,6.608815,4.9831905,4.787704,4.122364,3.9646032,5.7651367,11.4205265,10.405369,8.940934,10.38479,13.728639,13.612033,19.233126,21.098822,20.594673,20.052797,22.727877,23.876787,26.02714,27.234354,26.150604,21.997374,17.754974,18.639809,21.558388,25.080574,29.43272,33.41104,30.749681,25.927681,21.94593,20.306587,21.973368,25.989414,30.50618,33.280716,31.68253,28.870268,30.207806,32.128376,35.25273,44.37886,53.885677,59.335293,54.95914,44.13536,39.351086,46.985348,56.608772,56.680794,45.654667,31.974045,30.029469,26.719915,31.322422,38.442245,28.01287,24.60729,20.189981,17.339994,17.099922,18.993055,14.863832,14.3974085,14.147048,12.97413,12.05843,9.592556,11.029553,13.828096,16.276823,17.501184,14.586036,12.127021,12.72034,16.13621,19.315437,23.513252,25.317215,23.60585,19.78529,17.816708,15.29596,17.449741,18.79757,16.510035,10.425946,4.249259,3.216953,3.7211025,4.290414,5.6005163,6.711703,8.501947,10.172156,11.80464,14.373401,14.232788,11.135871,7.2021337,4.249259,3.789694,3.9646032,6.8111606,13.4645605,20.745575,21.184563,13.567448,9.499957,9.22902,11.252477,12.312219,15.745236,17.38115,17.326277,16.019604,14.267084,11.170166,8.30646,6.6465406,6.526505,7.630832,7.9875093,10.765475,12.864383,12.644889,9.932085,24.789059,34.25472,28.558174,12.758065,6.7391396,4.698535,4.184097,5.2918534,6.8797526,6.5779486,7.349606,10.64201,13.732068,13.869251,8.268735,7.6925645,9.757176,11.80464,13.039291,14.5414505,13.347955,9.921797,7.449064,6.756287,6.276145,8.995808,10.837497,11.015835,11.008976,14.555169,19.325726,20.766151,18.79071,14.095605,8.128122,9.729739,11.1393,11.149589,9.201583,5.394741,4.7088237,3.6936657,2.8019729,2.5378947,3.4295874,4.8082814,4.149801,4.2081037,5.007198,3.8514268,1.9308578,1.7525192,3.059192,4.372724,3.0077481,1.6667795,1.5158776,2.0474637,2.9940298,4.355576,3.875434,3.3129816,3.7211025,4.557922,3.7005248,2.9460156,3.940596,4.15666,2.8980014,1.2998136,1.3478279,1.8725548,2.5653315,3.1620796,3.4467354,3.806842,3.74168,3.6216443,3.309552,2.1846473,1.1763484,2.435007,3.9680326,4.1292233,1.5844694,1.1900668,0.8745448,0.91912943,1.2586586,1.488441,1.6907866,1.7319417,1.9548649,2.1297739,1.4678634,1.0494537,1.9411465,2.534465,2.428148,2.4487255,3.199805,3.2443898,2.218943,1.2072148,2.7230926,5.826869,4.448175,3.4021509,3.8445675,3.2821152,3.9440255,5.3330083,4.9694724,2.8877127,1.6221949,4.341858,4.9523244,4.122364,2.884283,2.6476414,2.901431,2.8225505,2.5481834,2.5721905,3.7622573,4.033195,3.8137012,3.2649672,2.719663,2.6407824,2.7470996,2.270387,1.5981878,1.0940384,1.1111864,1.1900668,0.96371406,0.70649505,0.5521636,0.50757897,0.5761707,0.6790583,0.805953,0.91569984,0.94999576,0.8848336,1.0014396,1.0357354,1.0117283,1.2655178,1.5433143,1.9480057,1.6873571,0.7922347,0.116605975,0.034295876,0.0034295875,0.0548734,0.12689474,0.082310095,0.06516216,0.15433143,0.23664154,0.25378948,0.19548649,0.15776102,0.19548649,0.25721905,0.36353627,0.59331864,0.6001778,0.64133286,0.66191036,0.70649505,0.89855194,0.78194594,0.6756287,0.72707254,0.9259886,1.0700313,1.1214751,1.0837497,0.91912943,0.72364295,0.72021335,0.9534253,1.2209331,1.4129901,1.4541451,1.2929544,1.3855534,1.3924125,1.4335675,1.529596,1.6084765,1.4918705,1.2620882,1.1043272,1.0563129,1.0254467,1.0117283,1.2037852,1.3615463,1.3821237,1.2895249,1.3409687,1.2998136,1.1934965,1.1214751,1.2175035,1.4438564,1.587899,1.5844694,1.4232788,1.1763484,1.2895249,1.5501735,1.5741806,1.3786942,1.3752645,1.1900668,1.196926,1.2689474,1.3066728,1.255229,1.155771,1.0117283,0.8711152,0.7476501,0.61389613,0.7407909,0.77508676,0.7339317,0.6344737,0.5041494,0.4046913,0.4938606,0.6344737,0.7682276,0.90884066,0.8162418,0.7442205,0.70306545,0.6790583,0.65162164,0.5590228,0.4629943,0.36010668,0.29494452,0.36010668,0.34295875,0.30866286,0.25721905,0.1920569,0.08916927,0.08573969,0.07888051,0.082310095,0.10288762,0.15776102,0.17147937,0.22292319,0.30866286,0.42869842,0.5761707,0.66191036,0.6207553,0.61046654,0.66876954,0.7339317,0.85396725,0.99801,1.0631721,1.0425946,1.0220171,0.96371406,0.94999576,0.939707,0.94999576,1.0597426,1.0940384,1.0906088,1.0014396,0.89512235,0.94999576,0.7510797,0.53501564,0.36696586,0.26407823,0.16804978,0.09602845,0.05144381,0.030866288,0.037725464,0.09602845,0.19548649,0.26750782,0.33952916,0.42526886,0.52815646,0.6173257,0.71678376,0.805953,0.8711152,0.89855194,1.0288762,1.0288762,1.0768905,1.1763484,1.1763484,1.3203912,1.4164196,1.3821237,1.2723769,1.2655178,1.2895249,1.3889829,1.3855534,1.2860953,1.3032433,1.3341095,1.3101025,1.3238207,1.3958421,1.4815818,1.3752645,1.4472859,1.6496316,1.8965619,2.0440342,2.1880767,2.3424082,2.4144297,2.4144297,2.469303,2.4727325,2.5207467,2.5756202,2.6373527,2.719663,0.05144381,0.048014224,0.082310095,0.116605975,0.1371835,0.1371835,0.20577525,0.18519773,0.2503599,0.38754338,0.3806842,0.67219913,0.6756287,0.59674823,0.5521636,0.59331864,0.50757897,0.53844523,0.59331864,0.65505123,0.7922347,0.8848336,0.77851635,0.6001778,0.45613512,0.42869842,0.71678376,0.7888051,0.6379033,0.40126175,0.36696586,1.0460242,2.0165975,3.100347,4.434457,6.468202,9.335337,11.115293,12.288212,14.057879,18.351723,19.312008,20.21399,20.320305,20.087093,21.170843,22.316326,22.501524,23.163433,25.804216,31.970613,32.042637,30.626217,28.198069,25.282919,22.453508,20.36832,22.381487,25.60187,28.043737,28.626766,29.42243,29.888855,31.703106,35.482513,40.774364,40.287365,37.09099,31.233253,24.511261,20.478067,18.12194,15.415996,13.025573,12.531713,16.434584,17.86815,16.678083,14.970149,13.63604,12.325937,10.4533825,10.690024,11.417097,11.005547,7.822889,5.7891436,4.547633,3.875434,3.3541365,2.3629858,2.3389788,2.5001693,2.5653315,2.4041407,2.037175,1.7182233,1.4815818,1.3512574,1.3272504,1.3958421,1.5330256,1.4267083,1.138623,0.764798,0.45956472,0.30523327,0.2194936,0.17833854,0.1920569,0.31895164,0.5761707,0.66876954,0.6927767,0.6859175,0.6276145,0.6173257,0.6344737,0.6310441,0.6241849,0.72021335,0.8196714,0.6379033,0.47328308,0.4424168,0.45613512,0.47328308,0.47328308,0.42869842,0.3806842,0.41840968,0.3806842,0.28465575,0.20577525,0.16119061,0.13375391,0.07888051,0.044584636,0.034295876,0.05144381,0.09259886,0.12689474,0.18862732,0.29494452,0.50757897,0.922559,1.196926,1.3684053,1.9171394,2.8534167,3.7279615,4.2835546,4.40702,4.338428,4.201245,4.0057583,4.9214582,6.327589,8.687145,11.063849,11.146159,12.80265,14.229359,14.531162,14.445422,16.355703,16.016174,17.768692,20.20027,21.904776,21.486366,21.681852,21.956219,21.260014,19.281141,16.410576,16.540901,16.640358,17.508043,18.910746,19.582945,20.148827,20.049368,19.95334,20.244854,21.02337,21.44864,25.51956,29.00402,29.453297,26.205479,22.820475,23.132568,24.552416,28.074602,38.277626,41.703785,30.729103,20.03908,15.587475,14.610043,13.457702,14.369971,16.156786,17.96761,19.294859,18.108221,16.774113,16.492886,16.13278,12.202472,14.057879,16.856422,17.648657,16.503176,16.503176,16.29054,16.695232,18.152807,21.705858,29.00745,33.65111,28.822252,22.580404,18.187103,14.099034,10.655728,8.289313,5.675967,2.9665933,1.8073926,2.767677,3.724532,4.2766957,4.15323,3.199805,3.0660512,2.9940298,3.9646032,7.2432885,14.38369,11.996697,12.730629,13.951562,13.745787,10.906088,12.288212,18.835295,22.038528,19.754423,16.19794,18.231688,20.244854,23.537258,26.654755,25.392666,22.865059,20.049368,19.222837,21.160555,25.10458,29.919722,28.311245,24.819925,21.94593,20.135109,21.390337,22.9508,23.849352,24.566135,27.045727,26.658184,27.831102,27.85511,28.856548,37.794052,45.373444,46.124523,41.53916,36.13756,37.48882,36.6863,43.994747,46.127953,39.91354,32.286137,29.724234,29.220085,33.6614,39.687187,37.67745,30.00546,21.973368,16.019604,13.498857,14.675205,13.96871,16.925014,15.902997,11.89038,14.493437,11.736049,10.611144,12.744347,17.079346,19.884748,17.998474,14.942713,12.857523,13.7697935,19.579515,22.70044,24.398085,22.453508,18.231688,16.691803,16.6335,14.651197,12.106443,10.278474,10.350495,8.457363,5.2026844,3.2203827,3.2375305,4.07435,5.9983487,9.033533,11.187314,11.705182,11.094715,10.014396,9.6645775,8.261876,5.857735,4.341858,5.936616,10.871792,16.482597,19.003344,13.591455,7.781734,6.4407654,8.639131,12.0309925,12.864383,14.510585,13.687484,12.085866,10.432805,8.467651,7.48336,7.023795,8.035523,10.175586,11.835506,9.400499,10.22703,11.910957,13.38225,14.908417,34.892624,47.787872,37.965534,13.920695,8.261876,6.8900414,5.442755,5.586798,6.701414,5.878313,7.010077,10.456812,13.317088,13.440554,9.431366,8.39563,9.115844,10.096705,11.122152,13.2690735,12.154458,9.716022,7.6616983,6.601956,6.046363,8.992378,9.431366,9.325048,10.950673,16.931873,18.718689,17.195951,14.7197895,12.421966,10.213311,11.235329,11.362224,9.781183,6.924337,4.4859004,4.1600895,3.5359046,3.0111778,3.6216443,7.051232,4.2698364,3.7965534,4.1463714,4.1189346,2.8054025,2.5481834,2.7539587,3.8377085,4.4927597,1.7147937,1.1454822,1.3546871,1.7113642,1.9754424,2.311542,1.8931323,1.7696671,2.1880767,2.7470996,2.3767042,3.0420442,3.3129816,2.976882,2.194936,1.5021594,1.4267083,1.4061309,1.8073926,2.7402403,4.0263357,4.0709205,3.2478194,3.3301294,4.098357,3.3198407,1.7936742,1.6496316,2.1332035,2.270387,0.8711152,0.88826317,0.7442205,0.96371406,1.4369972,1.4267083,1.5364552,1.3581166,1.5330256,1.9685832,1.8313997,0.97057325,1.6359133,2.153781,1.9480057,1.5536032,1.9651536,2.061182,1.7113642,1.4644338,2.551613,4.8254294,3.5393343,2.4315774,2.6990852,2.983741,3.4467354,4.5990767,4.1120753,2.1640697,1.4198492,3.7279615,4.0194764,3.3369887,2.6476414,2.8088322,2.8465576,2.8877127,2.836269,2.9082901,3.6353626,3.6696587,3.199805,2.6853669,2.428148,2.5893385,3.6044965,3.117495,2.1640697,1.3581166,0.90884066,1.0323058,0.9294182,0.6962063,0.44584638,0.33266997,0.39783216,0.45270553,0.53158605,0.6276145,0.71678376,0.6927767,0.7373613,0.89169276,1.1420527,1.3958421,1.3409687,1.879414,1.7936742,0.90884066,0.09602845,0.020577524,0.0,0.01371835,0.030866288,0.017147938,0.05144381,0.14061308,0.19891608,0.1920569,0.15776102,0.17490897,0.20577525,0.24350071,0.31209245,0.48014224,0.48014224,0.41840968,0.40126175,0.48357183,0.65162164,0.53844523,0.51100856,0.67219913,0.88826317,0.7956643,0.8128122,0.7888051,0.7579388,0.8128122,1.0837497,1.1523414,1.2963841,1.4678634,1.5741806,1.4815818,1.5844694,1.6016173,1.5741806,1.5604624,1.6496316,1.5193073,1.371835,1.3101025,1.3341095,1.3684053,1.2175035,1.2517995,1.3443983,1.4095604,1.3752645,1.4267083,1.3992717,1.2826657,1.1832076,1.3306799,1.3101025,1.3341095,1.3684053,1.3375391,1.1420527,1.3581166,1.5604624,1.6359133,1.6290541,1.7319417,1.3306799,1.2312219,1.2037852,1.1592005,1.138623,1.0666018,0.980862,0.9259886,0.8745448,0.7305021,0.7476501,0.7682276,0.77165717,0.72707254,0.58645946,0.52815646,0.5418748,0.6001778,0.70649505,0.88826317,0.91227025,0.86082643,0.8025235,0.764798,0.72707254,0.607037,0.52472687,0.4664239,0.42183927,0.3841138,0.34638834,0.30523327,0.2709374,0.22978236,0.1371835,0.12346515,0.1097468,0.09945804,0.09945804,0.11317638,0.116605975,0.1371835,0.1920569,0.29494452,0.4424168,0.4938606,0.51100856,0.5624523,0.65505123,0.7133542,0.8093826,0.85739684,0.8505377,0.8162418,0.8196714,0.8471081,0.90541106,0.96371406,1.0082988,1.0425946,1.0323058,1.0563129,1.0425946,1.0014396,1.0460242,0.8711152,0.7682276,0.64476246,0.4972902,0.40126175,0.29151493,0.16804978,0.07545093,0.034295876,0.0274367,0.041155048,0.09259886,0.14747226,0.20920484,0.29151493,0.36010668,0.45613512,0.5624523,0.66191036,0.7510797,0.8779744,0.9362774,1.0151579,1.1111864,1.1317638,1.214074,1.2929544,1.3238207,1.3066728,1.3101025,1.2620882,1.3306799,1.3581166,1.3409687,1.4369972,1.371835,1.2449403,1.2243627,1.313532,1.3409687,1.3786942,1.5364552,1.646202,1.7147937,1.9342873,1.9754424,2.1057668,2.2120838,2.2566686,2.2738166,2.3149714,2.4212887,2.5824795,2.7711067,2.9322972,0.12003556,0.072021335,0.082310095,0.106317215,0.13032432,0.17490897,0.23664154,0.23321195,0.28465575,0.3806842,0.36353627,0.58988905,0.6241849,0.6241849,0.64476246,0.6173257,0.4972902,0.53158605,0.5453044,0.52815646,0.6241849,0.82996017,1.1077567,1.2346514,1.0906088,0.66191036,0.6790583,0.69963586,0.5727411,0.34638834,0.26407823,0.6962063,1.6084765,2.7162333,4.046913,5.9434752,8.519095,10.007536,11.4205265,13.742357,17.926455,16.729528,17.576635,18.094503,17.71039,17.672665,20.015072,22.36434,24.621008,27.501862,32.533066,30.965746,28.959436,27.062874,25.296637,23.149715,21.993944,23.643576,26.428402,28.945719,30.074053,30.941738,33.712845,38.77149,46.045643,55.02087,54.046867,49.169994,41.443134,33.1744,27.94085,25.423532,21.064526,18.45804,19.514353,24.44953,23.969387,20.471207,16.400288,13.203912,11.331357,9.818909,9.280463,9.211872,8.913498,7.466212,6.6705475,6.6122446,6.7665763,6.526505,5.1992545,5.267846,5.178677,4.6608095,3.789694,2.9906003,2.5378947,2.2120838,1.9994495,1.8897027,1.8828435,1.937717,1.7388009,1.4198492,1.0528834,0.66876954,0.4081209,0.28465575,0.20577525,0.18519773,0.34638834,0.66191036,0.75450927,0.7373613,0.66876954,0.5693115,0.65848076,0.77165717,0.83681935,0.85739684,0.90884066,0.90541106,0.70649505,0.5212973,0.432128,0.37725464,0.34295875,0.29494452,0.25378948,0.22978236,0.26064864,0.26407823,0.26064864,0.2503599,0.2194936,0.15776102,0.106317215,0.082310095,0.06516216,0.06859175,0.13375391,0.22292319,0.274367,0.39097297,0.65505123,1.1592005,1.4781522,1.845118,2.3561265,3.100347,4.1429415,5.2026844,6.0326443,6.2967224,5.9983487,5.4907694,6.135532,7.490219,10.155008,12.9707,13.029003,14.517444,15.638919,16.331696,16.80155,17.521763,18.132229,19.805868,22.035099,23.389786,21.517231,20.584383,20.148827,19.936192,19.442331,17.902447,18.921034,20.471207,22.017952,23.132568,23.496103,21.489796,20.982216,22.141417,24.175161,25.313786,24.487255,28.698788,33.218983,34.275295,29.01774,24.645016,22.2786,20.419764,20.546658,27.09374,33.561943,26.702768,18.509483,14.483148,13.594885,12.123591,12.840376,14.514014,16.163645,17.082775,16.359133,14.959861,14.061309,13.101024,9.767465,9.194724,9.877212,11.269625,12.617453,12.9707,12.500846,13.454271,14.96329,19.442331,32.601658,48.027943,39.121304,23.821915,12.3533745,7.1952744,3.9337368,3.474172,3.6559403,3.0969174,1.1832076,1.2758065,1.587899,2.435007,3.426158,3.450165,3.8377085,3.1415021,3.4604537,6.4544835,13.327377,12.346515,16.194511,18.993055,17.439453,10.840926,8.309891,16.060759,23.952238,24.710178,13.927555,15.367981,16.39,19.20912,22.957659,23.69159,22.882208,22.474087,22.508383,22.957659,23.729315,26.047716,24.727325,22.961088,21.729866,19.79901,20.968498,21.78474,19.569225,17.233677,23.266321,25.457829,25.968836,25.917393,26.565584,29.326403,33.390465,30.396433,27.954567,28.290667,28.249512,21.181131,25.255482,28.503302,27.450418,27.10403,26.69248,27.882545,29.971165,33.472775,40.08159,31.308704,20.159115,12.833516,11.132441,12.490558,13.766364,16.750105,15.223939,11.955542,18.70497,15.532601,14.256795,15.501736,18.04306,18.811287,22.11055,19.020493,14.493437,12.662037,16.859852,17.597214,18.019053,17.425734,16.530611,17.473747,15.522313,9.911508,7.654839,10.340206,14.1299,14.87755,9.14328,4.8117113,4.3178506,4.6402316,4.99005,6.8145905,8.416207,9.290752,10.127572,11.080997,11.461681,10.264755,7.905199,6.228131,8.272165,13.330807,16.53404,14.994157,7.7920227,6.3961806,7.3393173,9.935514,12.55229,12.607163,12.017275,10.360784,8.937505,7.8606143,6.046363,5.717122,6.8866115,9.743458,13.05301,14.177915,11.379372,11.303921,13.176475,16.431154,20.70099,41.624905,52.891098,40.290794,14.04759,8.793462,8.460793,6.90033,6.1732574,6.451054,6.029215,7.284444,10.117283,11.856084,11.303921,8.721441,8.073249,8.639131,9.023245,9.314759,11.070708,10.515115,9.650859,8.337327,7.0923867,7.1129646,9.136421,8.467651,8.011517,10.017825,16.071047,14.496866,12.271064,11.214751,11.502836,11.646879,11.201033,9.72631,7.5416627,5.641671,5.7239814,5.4016004,4.4516044,4.0846386,5.1683884,8.261876,3.8617156,3.9303071,4.2595477,3.309552,2.201795,2.668219,2.9871707,3.350707,3.1552205,1.0117283,0.85396725,1.762808,2.7642474,3.069481,2.061182,1.0906088,0.70649505,0.77165717,1.0460242,1.1694894,2.5413244,2.74367,2.5378947,2.287535,1.9651536,1.2998136,0.84367853,1.0357354,1.9857311,3.4810312,3.7485392,2.860276,3.3815732,4.8082814,3.5770597,1.9102802,1.0494537,0.8162418,0.90541106,0.8848336,0.91569984,0.85739684,0.94999576,1.2312219,1.5433143,1.7971039,1.4815818,1.4198492,1.7525192,1.9274281,0.8162418,1.0048691,1.3992717,1.4095604,0.94999576,1.0425946,1.1729189,1.6290541,2.1640697,1.99602,4.016047,3.4535947,2.4898806,2.1880767,2.4830213,2.4830213,3.175798,2.8568463,1.5810398,1.2003556,2.527606,3.0660512,2.9151495,2.6064866,3.1243541,3.57363,3.9783216,3.6970954,3.0146074,3.1517909,2.9974594,2.609916,2.386993,2.3904223,2.3629858,3.4776018,2.8980014,2.0920484,1.5707511,0.89169276,0.91227025,0.83338976,0.6962063,0.53501564,0.4115505,0.39783216,0.31895164,0.29151493,0.34638834,0.44927597,0.53501564,0.5418748,0.72021335,1.0700313,1.3341095,1.255229,1.4369972,1.2346514,0.59674823,0.06859175,0.01371835,0.0,0.006859175,0.01371835,0.006859175,0.041155048,0.11317638,0.16119061,0.16119061,0.15090185,0.20234565,0.22978236,0.2469303,0.2709374,0.33952916,0.4355576,0.37725464,0.3566771,0.42526886,0.48357183,0.48014224,0.59331864,0.75450927,0.823101,0.607037,0.6036074,0.6276145,0.72364295,0.9259886,1.2895249,1.3169615,1.4164196,1.5776103,1.7216529,1.7079345,1.7250825,1.7422304,1.6290541,1.4438564,1.4404267,1.4027013,1.4027013,1.488441,1.587899,1.4781522,1.313532,1.255229,1.255229,1.2826657,1.2963841,1.2826657,1.3512574,1.3169615,1.2346514,1.4267083,1.2312219,1.1214751,1.1283343,1.1934965,1.1660597,1.4644338,1.5330256,1.611906,1.7730967,1.9239986,1.5398848,1.4129901,1.2895249,1.1077567,1.0151579,0.9945804,0.9431366,0.939707,0.9534253,0.84367853,0.89512235,0.7990939,0.7305021,0.77165717,0.922559,0.78194594,0.6344737,0.5796003,0.64133286,0.77851635,0.89512235,0.94656616,0.91569984,0.84367853,0.8162418,0.7579388,0.72364295,0.6756287,0.59331864,0.48700142,0.3841138,0.32581082,0.30523327,0.28808534,0.20577525,0.17147937,0.14747226,0.13032432,0.11317638,0.11317638,0.106317215,0.10288762,0.12003556,0.17833854,0.2777966,0.34295875,0.42526886,0.5212973,0.61389613,0.6824879,0.72364295,0.71678376,0.6927767,0.6859175,0.70649505,0.78194594,0.8779744,0.9842916,1.0666018,1.0666018,1.0357354,1.0460242,1.0494537,1.039165,1.0528834,0.9259886,0.91912943,0.8676856,0.7407909,0.64476246,0.51100856,0.33952916,0.19891608,0.11317638,0.044584636,0.030866288,0.020577524,0.0274367,0.0548734,0.1097468,0.15776102,0.23664154,0.33609957,0.4424168,0.5624523,0.6790583,0.7682276,0.8505377,0.9328478,1.0117283,1.0357354,1.0631721,1.1214751,1.196926,1.2312219,1.2826657,1.3203912,1.3443983,1.371835,1.4438564,1.3443983,1.1797781,1.1214751,1.1832076,1.2312219,1.3032433,1.4815818,1.5364552,1.5193073,1.762808,1.8039631,1.9480057,2.1126258,2.2326615,2.2498093,2.3046827,2.3732746,2.5447538,2.7951138,2.9940298,0.216064,0.10288762,0.09602845,0.12003556,0.1371835,0.17147937,0.16462019,0.2469303,0.32924038,0.36696586,0.33952916,0.34638834,0.44927597,0.64133286,0.7888051,0.64476246,0.5144381,0.5418748,0.5418748,0.48357183,0.48357183,0.7579388,1.5124481,2.0165975,1.8416885,0.84367853,0.42183927,0.32924038,0.33952916,0.32924038,0.28465575,0.44927597,1.255229,2.3629858,3.6593697,5.2609873,7.421627,8.968371,11.183885,14.270514,17.339994,14.5414505,14.459141,14.87755,14.812388,14.534592,16.846134,21.019941,24.699888,27.254932,29.789396,28.784527,27.868828,27.584171,27.470995,26.044287,25.814505,27.17262,29.563044,31.991192,33.00635,34.144974,39.700905,48.449783,59.37645,71.68867,71.50004,64.81235,55.336395,46.05593,39.23791,35.811752,30.084341,27.302946,29.079472,33.34588,29.710516,24.260902,19.03764,15.529172,14.644339,12.788932,10.861504,9.575408,9.009526,8.635701,9.455373,10.467101,10.981539,10.655728,9.499957,9.458802,8.868914,7.73372,6.245279,4.7774153,3.6353626,2.952875,2.5550427,2.318401,2.16064,2.0303159,1.8485477,1.6187652,1.3306799,0.9294182,0.6036074,0.490431,0.37725464,0.2709374,0.39783216,0.6207553,0.6962063,0.6790583,0.607037,0.52472687,0.5727411,0.6310441,0.6824879,0.75450927,0.88826317,0.78537554,0.6927767,0.6001778,0.5144381,0.42869842,0.32581082,0.22978236,0.17833854,0.17147937,0.19891608,0.1920569,0.24350071,0.29151493,0.29151493,0.20577525,0.17490897,0.16119061,0.14747226,0.16804978,0.29151493,0.45270553,0.53501564,0.67219913,0.94656616,1.3581166,1.7250825,2.510458,3.2855449,4.166949,5.802862,7.9292064,9.441654,9.321619,7.932636,7.040943,7.6274023,8.433355,10.052121,12.418536,14.815818,17.566347,18.986197,19.8676,20.231136,19.312008,20.272291,20.930773,21.589252,21.60983,19.397747,19.188541,19.404606,21.047379,23.153145,22.78275,22.985096,25.217756,27.649334,29.223515,29.659073,26.373528,24.638157,24.583282,25.996273,28.304386,28.25637,30.633076,34.56338,36.933228,32.385593,27.230925,23.410364,19.613811,17.141079,19.895037,25.18346,20.04251,14.270514,12.020704,11.780633,10.6317215,10.175586,10.467101,11.516555,13.313659,11.177026,10.120712,10.089847,9.523964,5.336438,5.3844523,6.6293926,7.98408,8.64599,8.069819,7.208993,8.275595,10.131001,16.232237,34.64226,60.41904,48.250866,24.895376,7.3290286,2.7299516,1.4918705,2.633923,5.0414934,6.3790326,3.07634,2.4727325,2.5961976,4.2081037,6.355026,6.375603,6.711703,4.461893,2.9151495,4.7019644,11.794352,15.018164,19.363451,25.26577,28.074602,18.03963,10.247607,15.021593,25.68761,31.246971,16.396858,16.115631,16.307688,17.463459,19.089085,19.720127,18.327715,23.743034,28.777668,30.139215,28.43471,26.315224,22.055677,19.967058,20.234566,18.921034,19.823015,22.978235,21.109112,16.770683,22.343761,27.498432,25.34122,26.404394,29.803116,23.252604,24.94682,19.456049,18.183672,20.78673,15.179354,9.040393,10.371073,14.195063,16.986746,16.695232,18.28656,19.805868,19.696121,20.364891,28.198069,24.044838,13.773223,8.22758,10.065839,13.773223,13.341095,12.452832,11.0981455,11.996697,20.598103,17.778982,17.607502,18.362011,18.241976,15.385129,23.427511,20.96164,15.8138275,12.651748,12.994707,12.439114,11.592006,12.164746,14.781522,18.969048,13.666906,8.862054,10.762046,17.168514,17.487467,19.394318,13.114742,7.7714453,6.252138,5.1855364,3.1277838,2.877424,4.1326528,7.2878733,13.433694,17.230247,15.237658,11.71547,9.091836,7.963502,9.760606,13.450842,14.54831,11.550851,5.953764,7.936065,10.106995,11.742908,12.178465,10.792912,8.748878,7.5039372,7.010077,6.6876955,5.439326,5.209543,6.8969,10.031544,12.9638405,12.878101,12.840376,14.455711,17.394867,21.143406,25.0257,44.6498,50.257175,36.305614,13.646329,9.510246,9.2153015,7.9943686,6.8385973,6.4098988,7.0306544,8.495089,10.436234,10.48082,8.587687,7.0478024,7.4456344,8.862054,9.112414,8.23444,8.484799,8.7283,8.958082,8.364764,7.5382333,8.47451,8.927217,7.490219,6.327589,7.226141,11.609154,9.043822,9.030104,10.237319,11.375941,11.214751,9.280463,6.6396813,5.171818,5.6485305,7.740579,8.083538,6.5333643,6.1046658,6.910619,6.159539,3.2786856,4.0503426,4.1017866,2.5378947,1.9514352,1.8313997,2.2326615,2.1332035,1.4095604,0.84367853,0.548734,1.8519772,3.6936657,4.7328305,3.3198407,1.3581166,0.53844523,0.33609957,0.44927597,0.7990939,1.3752645,2.386993,3.093488,3.0489032,2.1091962,0.8848336,0.490431,0.7956643,1.5604624,2.4555845,2.651071,2.4727325,3.309552,4.3624353,2.6545007,1.4369972,0.83338976,0.7476501,0.9294182,0.9534253,0.89512235,0.89855194,0.7613684,0.7373613,1.5364552,2.194936,1.9308578,1.4781522,1.313532,1.6530612,0.6001778,0.37382504,0.7613684,1.2586586,1.0631721,0.7373613,0.72707254,1.7353712,2.8534167,1.5741806,3.1826572,3.3884325,2.7539587,1.9857311,1.9445761,2.16064,2.4007113,2.1503513,1.5055889,1.1523414,2.2498093,3.340418,3.415869,2.9048605,3.707384,4.5099077,4.722542,3.9783216,2.9220085,3.210094,2.8294096,2.5413244,2.5653315,2.6785078,2.2292318,2.4761622,1.7936742,1.4095604,1.4815818,1.1043272,0.805953,0.7510797,0.70306545,0.58645946,0.5007198,0.42183927,0.30866286,0.24007112,0.23664154,0.2503599,0.34295875,0.40126175,0.52472687,0.7339317,0.9877212,0.9842916,0.6927767,0.34981793,0.10288762,0.01371835,0.0034295875,0.0,0.0034295875,0.01371835,0.017147938,0.037725464,0.09259886,0.13375391,0.14404267,0.15776102,0.1920569,0.2194936,0.22978236,0.23321195,0.2503599,0.4664239,0.48357183,0.44927597,0.44584638,0.47671264,0.6241849,0.78537554,0.82996017,0.7407909,0.6207553,0.64476246,0.72364295,0.83338976,0.9877212,1.2483698,1.5055889,1.7559488,1.9411465,2.0097382,1.8999915,1.8245405,1.7936742,1.611906,1.3272504,1.2106444,1.2620882,1.3238207,1.4987297,1.6530612,1.4129901,1.2723769,1.2209331,1.1489118,1.0666018,1.0940384,1.0631721,1.2175035,1.2449403,1.1729189,1.3958421,1.2517995,1.1008976,1.039165,1.097468,1.2312219,1.5913286,1.6221949,1.6942163,1.879414,1.9342873,1.728512,1.6667795,1.5055889,1.2243627,1.0357354,1.0460242,1.0048691,0.9774324,0.96714365,0.91227025,1.0768905,0.88826317,0.69963586,0.7510797,1.1763484,0.922559,0.7133542,0.6036074,0.6001778,0.6379033,0.78194594,0.96371406,0.9945804,0.90541106,0.9328478,1.0048691,1.0254467,0.90541106,0.70649505,0.6310441,0.53844523,0.45613512,0.4081209,0.37039545,0.26750782,0.22292319,0.19548649,0.16804978,0.1371835,0.12689474,0.1097468,0.09259886,0.09259886,0.11317638,0.15433143,0.26407823,0.36696586,0.45270553,0.52472687,0.6241849,0.6207553,0.64476246,0.67219913,0.6893471,0.6790583,0.7305021,0.82996017,0.9362774,1.0151579,1.0288762,1.0597426,1.0288762,0.9842916,0.9602845,0.980862,0.90884066,0.90541106,0.91569984,0.89512235,0.82996017,0.70649505,0.52815646,0.36353627,0.23321195,0.12689474,0.07888051,0.030866288,0.01371835,0.024007112,0.041155048,0.058302987,0.09602845,0.15090185,0.22978236,0.34638834,0.45613512,0.5727411,0.65505123,0.72021335,0.83681935,0.8711152,0.8711152,0.922559,1.0220171,1.0837497,1.3066728,1.313532,1.2792361,1.2758065,1.2689474,1.2826657,1.1763484,1.0871792,1.0768905,1.1214751,1.0734608,1.2003556,1.2998136,1.3684053,1.5947582,1.6633499,1.8142518,2.0303159,2.2360911,2.3321195,2.4487255,2.4247184,2.428148,2.5173173,2.6304936,0.16804978,0.13032432,0.13032432,0.12003556,0.09602845,0.12346515,0.19548649,0.21263443,0.21263443,0.24007112,0.34981793,0.24007112,0.36010668,0.6276145,0.8505377,0.71678376,0.45956472,0.66191036,0.7613684,0.59331864,0.39783216,0.50757897,1.2483698,1.7010754,1.4541451,0.6241849,0.31895164,0.2709374,0.36353627,0.4664239,0.4424168,0.39440256,0.9842916,1.8828435,2.976882,4.3933015,6.310441,8.419638,10.854645,13.395968,15.470869,11.821788,11.780633,12.548861,12.80265,12.679185,13.790371,17.648657,22.103691,25.173172,25.039417,26.02714,26.93598,28.324963,29.473875,28.34897,27.642475,29.525318,33.431618,37.67059,39.426537,44.433735,52.48641,64.8775,80.341515,95.07503,96.038734,85.825424,73.496056,64.140144,58.86544,55.85083,46.951054,40.99386,41.035015,44.354855,39.41282,34.690277,31.17152,28.25637,23.725885,16.45173,11.640019,9.126132,8.745448,10.343636,13.018714,14.575747,14.733508,13.992717,13.625751,12.442543,11.413667,10.984968,10.55284,8.453933,5.5730796,4.1017866,3.4124396,3.07634,2.867135,2.5619018,2.3492675,2.1194851,1.7936742,1.3443983,0.9877212,0.85396725,0.6790583,0.4698535,0.5178677,0.7133542,0.75450927,0.7305021,0.6824879,0.61046654,0.4629943,0.39097297,0.4389872,0.607037,0.84024894,0.71678376,0.7133542,0.7510797,0.7339317,0.5658819,0.33266997,0.1920569,0.14404267,0.18519773,0.31895164,0.2469303,0.1920569,0.1920569,0.216064,0.16804978,0.16804978,0.20577525,0.31552204,0.52472687,0.85396725,0.9259886,1.1111864,1.3924125,1.7490896,2.1503513,2.760818,4.187526,5.579939,7.1712675,10.285333,11.430815,10.738038,8.958082,7.346176,7.675417,10.751757,12.984418,14.730078,16.828985,20.61525,22.70044,22.628418,22.450079,22.374628,20.752434,18.71183,19.603521,20.759293,21.592682,23.61957,23.705309,25.464687,29.628206,34.868614,37.811203,37.211025,35.58883,34.43649,34.018078,33.369884,30.317553,29.00745,26.881107,24.703318,26.534718,29.124056,28.818823,31.771698,37.08413,36.802902,27.5876,23.132568,20.53294,18.71183,18.416885,16.050468,12.730629,11.22161,11.132441,8.9100685,7.9943686,7.226141,6.6533995,6.550512,7.414768,6.708273,5.7719955,5.693115,5.6793966,3.0660512,3.690236,4.770556,4.8905916,4.0880685,3.8445675,3.9440255,4.8837323,6.3618846,11.694893,27.831102,56.262383,45.572357,22.895926,5.586798,1.2072148,1.0597426,2.3492675,5.90232,9.14328,6.1046658,6.1149545,6.9792104,11.05699,15.542891,12.466551,9.853205,6.279575,4.307562,6.9963584,17.899017,23.475527,21.647556,30.461596,45.932465,42.05017,21.482935,16.780972,23.643576,29.141205,11.736049,13.200482,15.690363,18.440891,20.649546,21.45207,19.414894,22.422644,27.92027,32.32729,31.020618,26.332373,19.805868,17.785841,20.018501,19.654966,18.945042,24.470106,24.404943,19.696121,24.079134,32.85545,25.804216,25.985985,32.92061,22.566685,24.11686,17.593784,14.589465,16.304258,13.519434,12.260776,15.004445,19.78872,19.939621,4.0606318,8.06296,14.79524,15.704081,11.375941,11.537132,16.979887,13.937843,10.233889,11.345076,20.399187,15.175924,11.965831,11.588576,14.054449,18.571217,15.175924,14.904987,14.105893,13.039291,15.885849,20.70785,21.133118,17.549198,12.932974,12.847235,12.22648,10.422516,11.900668,16.808409,20.995934,18.70154,18.163095,20.62897,21.843042,12.055,16.657507,13.358243,9.431366,6.8214493,2.1229146,1.3992717,1.4129901,2.9082901,7.380472,17.058767,19.929333,16.050468,11.4033785,8.827758,8.011517,8.803751,11.355364,11.784062,9.321619,6.3310184,7.699424,10.80663,11.71547,9.55826,6.5299344,5.4941993,5.195825,5.6313825,6.5127864,7.2947326,6.584808,6.931196,8.659708,11.084427,12.511135,14.904987,18.259123,21.860191,24.92624,26.610168,44.313698,46.05593,32.900032,14.88098,10.984968,10.254466,8.899779,7.5931067,6.9689217,7.630832,9.424506,10.429376,8.971801,6.375603,6.9723516,7.840037,9.338767,10.106995,9.4862385,7.507367,6.9689217,6.800872,6.691125,7.2432885,9.962952,9.791472,7.2707253,4.7191124,3.882293,5.919468,5.164959,7.226141,8.683716,9.006097,10.542552,7.2707253,4.9248877,4.6882463,6.2487082,7.8126,10.511685,10.288762,9.901219,9.551401,6.866034,3.350707,3.532475,3.8137012,2.74367,1.0220171,0.5212973,1.1660597,1.4267083,0.939707,0.48700142,0.39097297,0.61389613,0.7956643,1.4164196,3.782835,1.3924125,0.5007198,0.29837412,0.36010668,0.64133286,0.7888051,1.3546871,2.294394,2.8396983,1.5090185,0.71678376,0.6276145,1.1900668,2.1400626,3.0043187,1.3821237,1.2072148,2.0406046,2.7882545,1.6770682,1.3478279,1.0460242,0.94999576,0.9877212,0.85396725,0.72021335,0.58645946,0.432128,0.34295875,0.48700142,1.7696671,2.1812177,1.6564908,0.90884066,1.4335675,0.70306545,0.37382504,0.6824879,1.2072148,0.85396725,0.64819205,0.47671264,1.1660597,2.2566686,2.0131679,1.6976458,3.210094,3.4055803,2.1743584,2.4555845,2.9082901,3.1415021,2.726522,2.0063086,2.1057668,4.852866,6.077229,5.219832,3.7211025,5.051782,4.57507,3.340418,2.9117198,3.625074,4.5784993,3.9440255,3.5564823,3.525616,3.474172,2.5481834,2.061182,1.7010754,1.2895249,1.08032,1.7388009,0.922559,1.0837497,0.9602845,0.35324752,0.12346515,0.17147937,0.22978236,0.25378948,0.22635277,0.15090185,0.17833854,0.25721905,0.32924038,0.4629943,0.85396725,0.58645946,0.23664154,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.07888051,0.12689474,0.15090185,0.15776102,0.18176813,0.15776102,0.12346515,0.13032432,0.20234565,0.33609957,0.44584638,0.4629943,0.42183927,0.36696586,0.36696586,0.5727411,0.58988905,0.6310441,0.7407909,0.77851635,0.8162418,0.9602845,1.0357354,1.1008976,1.4815818,2.0920484,2.435007,2.4830213,2.2806756,1.937717,1.8999915,1.8656956,1.6942163,1.4438564,1.3581166,1.3203912,1.2586586,1.2517995,1.3649758,1.6324836,1.3272504,1.1214751,0.96371406,0.8848336,1.0082988,1.1523414,1.2723769,1.2483698,1.2346514,1.6633499,1.529596,1.3684053,1.2312219,1.1832076,1.2826657,1.611906,1.7936742,1.9720128,2.1057668,1.9823016,1.6290541,1.5673214,1.471293,1.2655178,1.1454822,1.2037852,1.2860953,1.2963841,1.2312219,1.1454822,1.1934965,0.9945804,0.78194594,0.6379033,0.5041494,0.5658819,0.6790583,0.70649505,0.6379033,0.6241849,0.7613684,0.85739684,0.91912943,0.97057325,1.0666018,1.2277923,1.2380811,0.9877212,0.64476246,0.65505123,0.77851635,0.6893471,0.548734,0.42869842,0.30523327,0.28122616,0.26407823,0.24007112,0.20234565,0.15090185,0.10288762,0.072021335,0.06859175,0.082310095,0.106317215,0.20577525,0.29151493,0.34295875,0.3806842,0.5041494,0.5761707,0.64133286,0.6344737,0.5590228,0.47328308,0.48357183,0.6241849,0.7407909,0.7613684,0.6859175,0.7956643,0.77851635,0.69963586,0.6379033,0.6859175,0.72364295,0.7339317,0.77508676,0.85396725,0.91569984,0.89169276,0.7305021,0.52815646,0.36010668,0.274367,0.17833854,0.08916927,0.041155048,0.0274367,0.01371835,0.01371835,0.034295876,0.058302987,0.09259886,0.15090185,0.26407823,0.51100856,0.607037,0.5418748,0.5796003,0.65162164,0.7442205,0.8779744,1.0220171,1.0837497,1.1797781,1.1317638,1.1317638,1.196926,1.1592005,1.2826657,1.1934965,1.039165,0.89169276,0.7339317,0.6344737,0.7579388,0.96371406,1.2037852,1.5090185,1.5947582,1.6804979,1.821111,2.0268862,2.2566686,2.503599,2.5173173,2.4144297,2.311542,2.3492675,0.12003556,0.11317638,0.08916927,0.09259886,0.1097468,0.08573969,0.1097468,0.16119061,0.2194936,0.25721905,0.22978236,0.29494452,0.3841138,0.4389872,0.4664239,0.5453044,0.6310441,0.70649505,0.66876954,0.5453044,0.50757897,0.50757897,0.5727411,0.5555932,0.42183927,0.2469303,0.32238123,0.33266997,0.34981793,0.37039545,0.30866286,0.29837412,0.7305021,1.471293,2.49331,3.8685746,6.56766,9.136421,10.755186,11.183885,10.748327,10.244178,11.214751,11.756626,11.252477,10.347065,10.707172,13.125031,16.660936,20.131678,22.086544,22.43979,24.206028,26.8571,29.00402,28.400414,29.556185,32.440468,36.16157,40.006138,43.446014,51.28262,62.562534,84.13807,113.52963,138.9463,136.61761,122.02472,109.12261,101.625534,92.98298,78.95596,66.57515,62.754593,67.00385,71.41773,68.39626,61.180412,52.84651,43.250526,29.0246,21.729866,17.754974,15.371411,13.701202,12.713481,14.116182,13.649758,13.035862,12.758065,12.05157,11.122152,9.884071,9.112414,8.680285,7.5862474,5.994919,4.976331,4.506478,4.40702,4.3452873,4.0709205,3.5050385,2.9220085,2.417859,1.9171394,1.3684053,1.1043272,0.94999576,0.82996017,0.7510797,0.89855194,0.7990939,0.6276145,0.5178677,0.5624523,0.6310441,0.5796003,0.5521636,0.6241849,0.8265306,0.9774324,0.97057325,0.7956643,0.548734,0.4046913,0.33952916,0.2709374,0.274367,0.3566771,0.4424168,0.37039545,0.2777966,0.2469303,0.2777966,0.2777966,0.29837412,0.33952916,0.58645946,1.0906088,1.7833855,1.8176813,1.8519772,2.020027,2.386993,2.9460156,4.698535,6.23156,6.931196,7.4010496,9.47938,11.8869505,11.897239,11.355364,10.772334,9.335337,15.251375,19.397747,21.318316,21.939072,23.557837,24.500973,23.760181,23.160004,23.60585,25.097721,23.478956,23.406935,24.305487,25.540138,26.414682,26.69591,29.737953,35.25273,41.73122,46.440044,51.89652,53.63875,50.8745,43.86442,33.93234,30.540476,31.67567,32.022057,30.070623,28.132906,27.93742,24.243753,25.238335,30.561054,31.288126,23.917942,20.604961,18.917604,18.475187,20.94449,17.54234,13.567448,12.308789,12.229909,6.9826403,6.4098988,6.9620624,6.368744,4.5201964,3.474172,4.033195,3.8479972,3.6799474,3.566771,2.7985435,3.666229,3.4433057,3.8891523,5.9983487,10.021255,11.015835,11.266195,11.204462,12.2093315,16.588915,26.740494,20.642687,10.834066,4.4859004,3.4021509,2.8156912,4.7945633,7.2707253,8.587687,7.531374,9.078118,10.600855,12.037852,12.80608,11.818358,16.149927,13.046151,11.015835,13.687484,19.816156,34.981792,26.274069,25.653315,39.00127,46.093655,28.541027,15.433144,12.826657,19.243416,25.660173,30.132355,21.688711,14.949572,16.13621,23.053686,19.637817,27.536158,34.141544,33.6614,27.10403,25.011982,22.751883,22.504953,23.931662,24.168303,19.154245,17.761833,16.400288,16.516893,24.579853,23.153145,17.401728,15.405707,16.527182,11.399949,14.562028,15.536031,13.2690735,10.618003,14.335675,17.494326,13.540011,10.017825,8.848335,6.355026,16.479168,16.146498,12.600305,10.175586,10.264755,18.825006,14.476289,9.499957,11.101575,21.390337,20.687271,17.55263,13.862392,12.075578,15.223939,15.316538,18.54035,19.630959,16.942162,12.442543,12.850664,10.117283,10.796341,14.123041,12.006986,14.54831,10.501397,7.473071,7.73372,8.241299,10.028113,7.9120584,9.595985,13.419975,8.354475,10.408798,9.527394,7.3050213,4.6882463,1.961724,1.9445761,3.532475,5.802862,8.618553,12.603734,14.856973,12.823228,10.021255,7.891481,5.813151,6.7048435,8.951223,10.028113,9.012956,6.5882373,6.7357097,7.06838,6.6705475,5.5147767,4.479041,3.549623,3.508468,5.394741,8.268735,9.1981535,8.999237,9.80519,11.334786,14.068168,19.288,18.54378,19.517782,22.20315,25.584723,27.659622,44.179947,45.092216,31.524769,13.656617,10.731179,9.568549,8.529384,7.805741,7.689135,8.594546,9.606275,9.482809,8.56368,7.641121,7.9257765,7.805741,8.1212635,8.419638,8.519095,8.484799,5.192395,4.57507,5.754848,7.699424,9.218731,14.311668,10.285333,4.863155,2.4590142,4.173808,4.99005,6.495639,6.742569,6.029215,6.893471,6.591667,4.7602673,3.9303071,4.482471,4.6402316,9.544542,10.456812,9.551401,8.008087,6.036074,2.4727325,4.7808447,6.725421,5.5422134,1.9239986,0.90884066,0.8128122,0.8471081,0.65162164,0.31895164,1.529596,2.0577524,1.488441,0.88826317,2.8088322,1.99602,0.864256,0.28122616,0.39440256,0.6173257,0.7133542,1.6564908,2.435007,2.2806756,0.65505123,0.7613684,1.2792361,1.7422304,1.9102802,1.7593783,0.7510797,1.6804979,2.620205,2.469303,0.9568549,0.980862,1.6976458,1.7490896,1.0288762,0.67219913,0.5453044,0.37725464,0.30523327,0.34295875,0.39097297,1.4369972,1.5261664,1.0357354,0.64476246,1.3375391,0.53501564,0.2194936,0.32581082,0.6241849,0.70649505,1.0666018,0.5761707,0.42183927,1.5638919,4.7362604,1.4027013,1.7936742,3.1723683,3.7519686,2.726522,4.280125,5.425607,5.48734,4.6093655,3.7279615,4.7774153,4.437886,3.474172,3.2066643,5.5147767,5.223262,3.99204,3.6765177,4.5201964,5.1512403,3.6765177,3.0351849,3.2135234,3.415869,2.0474637,1.4507155,1.313532,1.2517995,1.0323058,0.5796003,0.5418748,1.1797781,1.0666018,0.216064,0.061732575,0.14747226,0.2469303,0.26407823,0.20577525,0.15090185,0.12003556,0.1920569,0.30866286,0.4115505,0.4389872,0.2503599,0.08573969,0.006859175,0.0034295875,0.0,0.0,0.006859175,0.017147938,0.034295876,0.06859175,0.09602845,0.12689474,0.15433143,0.1920569,0.24350071,0.2194936,0.16462019,0.17147937,0.2709374,0.432128,0.5727411,0.6276145,0.64819205,0.65505123,0.64819205,0.64133286,0.6893471,0.78537554,0.86082643,0.7888051,0.8676856,1.196926,1.4267083,1.5158776,1.7353712,1.7113642,1.8897027,2.1743584,2.4315774,2.5001693,2.3664153,2.3321195,2.1469216,1.8005334,1.529596,1.3752645,1.2449403,1.1694894,1.2483698,1.646202,1.7113642,1.4164196,1.1317638,0.9877212,0.8848336,0.922559,1.097468,1.1351935,1.1283343,1.5158776,1.6839274,1.546744,1.4541451,1.488441,1.488441,1.6530612,1.6839274,1.6324836,1.5501735,1.5090185,1.4575747,1.3478279,1.2586586,1.2517995,1.3649758,1.4164196,1.3101025,1.2620882,1.3581166,1.546744,1.7216529,1.3443983,1.0220171,0.91227025,0.7099246,0.5178677,0.45270553,0.44927597,0.48014224,0.5658819,0.58988905,0.6927767,0.7613684,0.8162418,0.9842916,1.2689474,1.3409687,1.1832076,0.9602845,1.0220171,0.9294182,0.7442205,0.6276145,0.5727411,0.39097297,0.32581082,0.274367,0.2194936,0.16804978,0.12689474,0.1097468,0.09259886,0.08573969,0.08573969,0.082310095,0.10288762,0.19891608,0.274367,0.31895164,0.42869842,0.52472687,0.61389613,0.64133286,0.61046654,0.58302987,0.5178677,0.5555932,0.5693115,0.4972902,0.3566771,0.3806842,0.4424168,0.48014224,0.4972902,0.5761707,0.6241849,0.72364295,0.823101,0.91569984,1.0254467,0.9328478,0.8128122,0.6790583,0.5418748,0.39783216,0.26064864,0.17490897,0.11317638,0.058302987,0.0274367,0.0274367,0.024007112,0.024007112,0.034295876,0.0548734,0.09602845,0.17147937,0.25721905,0.3566771,0.53158605,0.5178677,0.6001778,0.64819205,0.6859175,0.91227025,1.1763484,1.2209331,1.2312219,1.2860953,1.3684053,1.1489118,1.0117283,0.91227025,0.84367853,0.82996017,0.6824879,0.66191036,0.71678376,0.8162418,0.9259886,1.097468,1.3375391,1.5055889,1.5981878,1.7319417,2.0165975,2.2258022,2.335549,2.3252604,2.1674993,0.041155048,0.10288762,0.09945804,0.106317215,0.1371835,0.15776102,0.11317638,0.14404267,0.1920569,0.20577525,0.15090185,0.22635277,0.24350071,0.2194936,0.22635277,0.4115505,0.58302987,0.5590228,0.52472687,0.5658819,0.69963586,0.53501564,0.4046913,0.2469303,0.11317638,0.15090185,0.33952916,0.32238123,0.26064864,0.2194936,0.17490897,0.22635277,0.59331864,1.1866373,2.037175,3.309552,6.1801167,8.508806,10.134431,10.621432,9.266746,8.80718,9.318189,9.438225,8.886061,8.436785,8.954653,10.618003,13.13189,15.951012,18.30028,20.440342,23.232025,26.239773,28.324963,27.642475,30.10149,33.623676,37.461384,41.350536,45.527775,52.572147,63.910362,88.85032,126.45232,165.56334,176.23279,164.50702,149.38597,136.74109,119.30506,97.37971,86.401596,89.162415,98.250824,96.04559,82.57418,70.183075,59.078075,47.904476,33.73685,27.724785,24.216316,21.380049,18.20082,14.476289,13.234778,12.267634,11.211322,10.021255,8.958082,8.2310095,7.48336,6.948344,6.543653,5.8680243,5.0449233,4.513337,4.2869844,4.3281393,4.530485,4.431027,3.9543142,3.3541365,2.760818,2.16064,1.6942163,1.3924125,1.1523414,0.9294182,0.7442205,0.805953,0.7442205,0.64133286,0.5693115,0.5693115,0.5212973,0.5727411,0.6756287,0.7956643,0.9259886,0.96714365,0.8676856,0.72021335,0.5761707,0.4115505,0.32238123,0.25721905,0.28808534,0.39097297,0.47328308,0.4938606,0.41840968,0.34981793,0.33609957,0.37039545,0.44584638,0.66533995,1.2003556,1.961724,2.6167753,2.9494452,2.9734523,3.2478194,3.8342788,4.32471,6.9037595,8.069819,8.06296,8.220721,10.960961,12.079007,12.46312,14.466,17.926455,20.169403,21.891056,23.18744,24.799347,26.949697,29.374416,28.420992,26.733635,25.879667,25.317215,22.402065,21.832754,23.256033,24.535269,25.485264,27.865398,29.549326,32.27242,36.466805,42.026165,48.30574,55.737656,62.78203,63.12156,53.745064,34.933777,28.071173,27.299517,28.667921,30.327843,32.51592,32.203827,27.337242,23.928232,23.28347,21.997374,21.27716,23.02625,22.275171,19.558937,20.927343,18.084215,13.776653,12.442543,13.114742,9.431366,10.134431,12.788932,13.666906,10.63858,3.1655092,3.0386145,3.6456516,3.724532,2.9700227,2.037175,5.336438,9.31133,11.88352,13.063298,14.953001,14.29795,12.229909,11.80121,14.63062,20.920483,20.186552,14.112752,9.8429165,9.39707,9.6817255,10.707172,15.073037,15.450292,11.8115,11.441104,11.729189,12.020704,12.895248,13.629181,12.205902,13.138749,11.653738,11.814929,15.035312,20.083664,25.543568,17.425734,16.37285,25.684181,31.312134,21.729866,15.443433,18.104792,31.226395,52.194893,50.973957,32.464474,15.398848,10.082987,18.389448,14.411126,22.059107,27.707638,26.414682,21.928782,26.215767,25.313786,24.346642,23.983105,20.409475,20.382038,20.28601,18.022482,18.855871,35.39677,29.079472,17.947031,11.526843,11.163307,10.014396,11.14273,13.821238,13.80409,11.317638,11.063849,17.168514,13.46799,9.023245,8.31675,11.266195,23.612709,19.387459,13.073587,11.043272,11.540562,15.885849,10.816919,9.355915,15.014734,21.764162,19.54179,16.7844,13.419975,11.660598,15.9921665,12.583157,14.733508,16.033321,13.443983,7.3050213,13.495427,10.906088,14.496866,21.356041,10.707172,12.758065,10.240748,7.7680154,7.5210853,9.280463,8.683716,4.791134,10.837497,20.135109,6.1046658,5.4976287,4.9077396,4.3761535,3.9886103,3.8720043,5.8165803,6.81802,7.9292064,9.0644,8.992378,10.628291,11.516555,10.734609,8.735159,7.3598948,8.752307,8.282454,6.989499,5.669108,4.8940215,4.437886,3.940596,3.782835,4.0091877,4.341858,3.357566,3.6182148,6.327589,10.4533825,12.713481,11.043272,11.183885,14.486577,21.52066,32.08379,25.344652,21.503513,21.928782,25.166313,26.942839,43.57977,47.921627,35.894062,16.012743,9.403929,8.22758,7.1849856,6.8591747,7.2432885,7.716572,9.129561,9.966381,9.277034,7.7748747,7.8537555,8.556821,8.378482,8.045813,7.7783046,7.301592,5.2164025,5.2472687,6.910619,9.122703,10.196163,13.251926,9.414218,5.0312047,3.782835,6.6876955,6.5985265,6.684266,6.6876955,6.416758,5.744559,7.2432885,10.755186,9.119273,3.4638834,3.1963756,6.776865,7.9257765,7.6342616,6.725421,5.8474464,2.527606,2.983741,5.919468,7.5107965,1.3924125,0.7133542,0.64133286,0.7682276,0.77165717,0.3841138,1.3958421,1.8519772,1.4747226,0.9568549,1.9514352,1.7182233,0.7956643,0.26064864,0.33609957,0.39097297,0.39440256,1.2860953,1.6496316,1.1111864,0.34981793,0.8505377,1.3409687,1.5227368,1.3443983,0.9911508,0.66533995,1.4472859,2.4418662,2.7230926,1.3443983,1.2517995,1.2620882,1.0940384,0.7613684,0.5796003,0.39097297,0.25721905,0.23321195,0.28808534,0.31209245,1.8862731,1.9308578,1.2415106,0.59331864,0.75450927,0.29494452,0.13032432,0.19548649,0.58302987,1.5330256,1.0494537,0.47671264,0.216064,0.90884066,3.4227283,1.1111864,0.8848336,2.218943,3.5873485,2.4452958,3.0969174,4.636802,5.1821065,4.3521466,3.2649672,4.1017866,3.3952916,2.4658735,2.3218307,3.6353626,3.9268777,3.1449318,2.6613598,2.901431,3.3644254,2.2498093,1.7662375,1.8005334,1.9239986,1.3924125,1.2175035,1.1008976,1.0014396,0.82996017,0.4629943,0.548734,0.70649505,0.58302987,0.22292319,0.082310095,0.39097297,0.45270553,0.32924038,0.15776102,0.16119061,0.12689474,0.24007112,0.33609957,0.31895164,0.16119061,0.072021335,0.020577524,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.05144381,0.09602845,0.09602845,0.1097468,0.13375391,0.16119061,0.18519773,0.19891608,0.24007112,0.31895164,0.4115505,0.45613512,0.5453044,0.6379033,0.64133286,0.5658819,0.5144381,0.7476501,0.7579388,0.7956643,0.91569984,0.9945804,1.196926,1.4678634,1.6427724,1.6839274,1.6907866,1.704505,1.8691251,2.0920484,2.2738166,2.318401,2.270387,2.2395205,2.1160555,1.8759843,1.5810398,1.4129901,1.3512574,1.3443983,1.4164196,1.6667795,1.7971039,1.6907866,1.471293,1.2380811,1.0563129,1.1043272,1.2003556,1.2758065,1.3786942,1.7010754,1.8931323,1.7971039,1.6873571,1.670209,1.704505,1.8279701,1.6084765,1.3855534,1.2998136,1.2963841,1.3272504,1.3066728,1.2792361,1.2723769,1.2826657,1.2998136,1.2449403,1.2003556,1.2620882,1.5570327,1.7353712,1.5433143,1.2929544,1.0940384,0.881404,0.6344737,0.45270553,0.36696586,0.3806842,0.4664239,0.52472687,0.58988905,0.6756287,0.7888051,0.9431366,1.0254467,1.0871792,1.1351935,1.1934965,1.3238207,1.1489118,1.0014396,0.90198153,0.8128122,0.6310441,0.5007198,0.42526886,0.3566771,0.274367,0.18519773,0.14404267,0.12346515,0.10288762,0.082310095,0.07545093,0.06859175,0.106317215,0.16119061,0.22978236,0.34638834,0.5178677,0.6276145,0.66191036,0.64133286,0.6379033,0.5521636,0.52472687,0.5178677,0.4972902,0.40126175,0.34295875,0.37382504,0.42869842,0.47671264,0.5041494,0.6756287,0.89169276,1.0357354,1.1043272,1.1797781,1.1660597,1.0631721,0.922559,0.7682276,0.6001778,0.4629943,0.33266997,0.216064,0.13375391,0.10288762,0.08916927,0.0548734,0.0274367,0.017147938,0.020577524,0.030866288,0.05144381,0.09259886,0.16804978,0.2709374,0.30866286,0.5178677,0.6173257,0.58302987,0.66876954,0.83338976,0.9431366,1.039165,1.1454822,1.255229,1.1763484,1.1592005,1.097468,0.97057325,0.85396725,0.7099246,0.66876954,0.6756287,0.70306545,0.7510797,0.89512235,1.1283343,1.3169615,1.4438564,1.5741806,1.7216529,1.8519772,2.0063086,2.153781,2.194936,0.041155048,0.1097468,0.12003556,0.116605975,0.12689474,0.15776102,0.11317638,0.14061308,0.17147937,0.17147937,0.15090185,0.16804978,0.1371835,0.14061308,0.19548649,0.26407823,0.40126175,0.4046913,0.42183927,0.53501564,0.7305021,0.51100856,0.40126175,0.274367,0.15090185,0.20234565,0.4355576,0.39097297,0.25721905,0.15090185,0.13032432,0.18176813,0.4664239,0.91569984,1.5810398,2.644212,5.586798,7.7542973,9.410788,10.30591,9.668007,7.9292064,7.6514096,7.507367,7.140401,7.1884155,8.018375,9.019815,10.6145735,12.737488,14.826107,17.86815,21.45893,24.706749,26.68562,26.428402,28.914852,32.954906,37.35507,41.748367,46.604664,52.09886,62.250443,84.851425,123.78067,178.97302,212.2503,204.49258,182.8073,159.2426,130.7736,102.92878,95.654625,104.29033,115.23071,105.946815,88.651405,74.39118,60.782578,47.009354,33.82259,27.913412,24.308916,21.308027,17.936743,13.972139,11.458252,10.13786,8.920357,7.507367,6.375603,5.919468,5.6999745,5.501058,5.171818,4.6127954,3.998899,3.6456516,3.5153272,3.5942078,3.8788633,3.9646032,3.7931237,3.4535947,3.0043187,2.4487255,2.0749004,1.6770682,1.3272504,1.0563129,0.8711152,0.8162418,0.7305021,0.6893471,0.6859175,0.6173257,0.52472687,0.6310441,0.823101,0.980862,0.96714365,0.8779744,0.77851635,0.7476501,0.7407909,0.5693115,0.38754338,0.31552204,0.36353627,0.47328308,0.53501564,0.5693115,0.53158605,0.50757897,0.53844523,0.607037,0.72364295,1.0734608,1.7971039,2.7128036,3.3129816,3.9200184,4.2115335,4.715683,5.3570156,5.429037,7.5279446,8.364764,8.2481575,8.450503,11.218181,12.229909,14.033872,17.528622,21.959648,24.919382,23.68473,23.160004,24.151155,26.428402,28.733084,26.737064,26.208908,26.651323,26.147175,21.36633,22.28546,24.672453,26.304935,27.813953,32.68054,33.397324,33.18469,34.350746,38.23647,45.198532,57.747395,69.55889,69.77839,56.11834,34.872044,28.51702,27.690489,29.038317,30.708527,32.371876,32.488483,30.002031,26.215767,21.599543,15.7966795,18.680964,24.696459,25.780209,21.973368,21.424633,19.843594,14.904987,12.932974,14.260224,13.231348,14.003006,15.673215,16.335125,13.564018,4.4413157,3.0077481,3.7691166,4.0709205,4.1189346,6.9654922,10.686595,14.054449,16.177364,18.015623,22.36777,24.394655,20.20027,15.8138275,16.369421,26.088871,22.36777,16.067617,12.929544,13.347955,12.370522,15.570327,21.897917,21.743584,16.242527,17.264544,15.028452,12.085866,11.526843,12.586586,10.655728,8.64942,9.448513,10.912948,12.435684,14.946142,12.761495,9.301042,10.909517,16.719238,18.608942,17.645227,20.172834,26.75764,38.41481,56.61563,50.737316,33.867176,16.647217,7.5279446,12.758065,10.213311,14.243076,17.833855,18.694681,19.250275,27.306376,25.317215,21.664703,19.178253,15.138199,19.713268,24.4461,22.227156,19.308577,35.307602,32.797146,19.675543,9.832627,8.014946,9.794902,9.026674,10.861504,13.567448,14.843254,11.8115,15.896138,13.4645605,9.815479,9.153569,14.586036,22.035099,16.53747,10.666017,9.966381,12.946692,11.914387,7.922347,10.741467,18.845583,19.435472,15.319967,13.516005,11.664027,11.070708,16.681513,11.108434,13.972139,15.391989,11.375941,3.8102717,23.506393,17.106783,14.7197895,19.668684,8.515666,9.126132,8.303031,7.4113383,7.8366075,10.984968,8.152129,6.3173003,18.410025,31.116648,4.852866,3.117495,2.7059445,3.2889743,4.482471,5.844017,7.8777623,8.656279,9.253027,9.270175,6.842027,6.8283086,9.156999,10.6317215,10.501397,10.425946,11.177026,7.623973,4.540774,3.6970954,3.858286,2.8808534,2.1640697,2.2978237,3.2203827,4.214963,4.372724,6.1458206,9.56512,13.728639,16.798119,13.440554,12.860953,18.386019,29.374416,41.2305,29.045176,21.993944,20.807306,23.36235,24.703318,37.51626,43.720383,34.861755,16.448301,7.9429245,6.4819202,5.878313,6.121814,6.7357097,6.790583,8.357904,9.829198,9.407358,7.5588107,7.010077,8.621983,9.15014,8.320179,6.8557453,6.464772,6.543653,7.9086285,9.825768,11.207891,10.618003,10.669447,7.4936485,5.1409516,5.5490727,8.546532,7.2192817,6.135532,6.2864337,6.9723516,5.802862,6.2418494,10.72775,9.253027,2.6064866,2.3835633,4.1429415,5.0586414,5.295283,5.1066556,4.8288593,3.690236,2.5447538,3.799983,5.4153185,0.89855194,0.6241849,0.71678376,0.8128122,0.72021335,0.44584638,0.8711152,1.0837497,1.1008976,1.0906088,1.3821237,1.5638919,0.88826317,0.42183927,0.42183927,0.35324752,0.30523327,0.75450927,0.7613684,0.28808534,0.19891608,0.65848076,0.9945804,1.0014396,0.7682276,0.7099246,0.8128122,1.255229,2.170929,2.9185789,2.07833,1.5638919,1.0666018,0.7682276,0.6379033,0.45613512,0.29494452,0.19891608,0.19548649,0.25378948,0.29837412,2.2806756,2.301253,1.4438564,0.5796003,0.37039545,0.1920569,0.1097468,0.14061308,0.4698535,1.4575747,0.7922347,0.35324752,0.18176813,0.61046654,2.2909644,1.1454822,0.5658819,1.4438564,3.0523329,3.0660512,2.318401,3.1620796,3.724532,3.350707,2.6133456,3.2718265,2.5893385,1.8485477,1.6393428,1.8897027,2.1846473,1.8348293,1.4610043,1.3786942,1.5810398,1.1592005,0.99801,0.9259886,0.8676856,0.8471081,0.9842916,0.9362774,0.89512235,0.8848336,0.7339317,0.5727411,0.33609957,0.2503599,0.28465575,0.12346515,0.5624523,0.7613684,0.5693115,0.18176813,0.15090185,0.15090185,0.26064864,0.2777966,0.16462019,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.041155048,0.061732575,0.09602845,0.08573969,0.1097468,0.15090185,0.18176813,0.16119061,0.22635277,0.31209245,0.41498008,0.4972902,0.47671264,0.45270553,0.4972902,0.5007198,0.4389872,0.4046913,0.71678376,0.82996017,0.8779744,0.9328478,1.0323058,1.2106444,1.4129901,1.6084765,1.7593783,1.7936742,1.8382589,1.9239986,1.9857311,2.0063086,1.9891608,1.9857311,1.9994495,1.9445761,1.7902447,1.5673214,1.4472859,1.430138,1.4815818,1.5741806,1.6839274,1.7319417,1.7525192,1.6324836,1.4061309,1.2689474,1.3512574,1.3615463,1.4644338,1.6633499,1.7971039,2.0063086,2.0097382,1.8931323,1.8073926,1.9754424,2.095478,1.6633499,1.2929544,1.1934965,1.1489118,1.1523414,1.196926,1.2346514,1.2346514,1.1900668,1.1111864,1.1729189,1.2106444,1.2655178,1.5673214,1.7353712,1.6770682,1.4747226,1.2243627,1.0151579,0.8848336,0.5796003,0.3566771,0.3018037,0.34638834,0.45270553,0.5590228,0.67219913,0.7888051,0.89512235,0.8779744,0.9362774,1.0288762,1.1351935,1.2620882,1.155771,1.1934965,1.2243627,1.1489118,0.9568549,0.8196714,0.71678376,0.61389613,0.47671264,0.3018037,0.20234565,0.17147937,0.14404267,0.10288762,0.09602845,0.072021335,0.06516216,0.08916927,0.15433143,0.25721905,0.48014224,0.59331864,0.61389613,0.58988905,0.6207553,0.59331864,0.5453044,0.52472687,0.53501564,0.52472687,0.45270553,0.432128,0.44927597,0.47671264,0.5041494,0.6962063,0.94999576,1.1454822,1.2620882,1.3889829,1.4164196,1.2826657,1.1283343,1.0185875,0.9362774,0.7339317,0.5590228,0.4046913,0.28465575,0.23321195,0.15776102,0.106317215,0.06859175,0.041155048,0.0274367,0.024007112,0.0274367,0.034295876,0.048014224,0.07545093,0.13375391,0.33266997,0.44927597,0.44584638,0.48014224,0.58988905,0.7339317,0.8471081,0.939707,1.0768905,1.1797781,1.2826657,1.2483698,1.0871792,0.96371406,0.8196714,0.7579388,0.7305021,0.71678376,0.72021335,0.77165717,0.89169276,1.0460242,1.2277923,1.4472859,1.5776103,1.6324836,1.7696671,1.99602,2.170929,0.08573969,0.106317215,0.1097468,0.10288762,0.08573969,0.072021335,0.10288762,0.14061308,0.16119061,0.16804978,0.19891608,0.15776102,0.12003556,0.16804978,0.2469303,0.12346515,0.2469303,0.33952916,0.40126175,0.4698535,0.6207553,0.48700142,0.45956472,0.4046913,0.31895164,0.29151493,0.53844523,0.51100856,0.39097297,0.28465575,0.19891608,0.17147937,0.32581082,0.6344737,1.1454822,1.9480057,4.880303,7.157549,8.632272,9.489669,10.254466,7.750868,6.8900414,6.6533995,6.584808,6.8043017,7.4936485,7.64798,8.522525,10.285333,12.034423,14.421415,18.331144,21.767591,23.852781,24.85079,26.514141,30.543905,35.41392,40.451984,45.836437,50.46981,59.225548,75.92078,109.27695,172.91637,65535.0,221.48276,194.41989,160.97455,124.610634,93.95012,90.74689,102.03023,111.49932,99.5232,86.08951,72.79985,57.34613,40.764076,27.416122,21.37662,17.676094,15.05246,12.744347,10.494537,8.872343,7.4044795,6.4133286,5.7891436,4.976331,4.887162,5.003768,5.0312047,4.7945633,4.2389703,3.4844608,3.0111778,2.7916842,2.7779658,2.8980014,3.093488,3.2512488,3.2821152,3.1277838,2.7573884,2.3732746,1.845118,1.4507155,1.2860953,1.2449403,1.0563129,0.82996017,0.7442205,0.77508676,0.6893471,0.7373613,0.823101,0.97057325,1.0906088,0.9568549,0.88826317,0.864256,0.881404,0.8779744,0.7339317,0.53158605,0.4629943,0.5007198,0.5796003,0.6173257,0.6173257,0.65505123,0.77508676,0.97057325,1.1866373,1.3924125,1.7799559,2.503599,3.4192986,4.105216,4.8734436,5.576509,6.125243,6.4579134,6.526505,7.5553813,7.9429245,8.035523,8.453933,10.110424,12.411677,15.614912,18.574646,20.399187,20.460918,19.692692,19.517782,19.912186,20.742146,21.78131,20.886189,22.769032,24.891945,25.4544,23.406935,25.60873,28.225504,31.01033,34.457066,39.820942,36.778896,32.9309,31.2504,33.109238,38.277626,55.37755,67.5663,64.55512,48.250866,32.74913,30.828562,32.00491,32.85888,31.627655,28.18435,27.721355,28.300955,27.741934,23.976246,15.038741,16.695232,23.454948,26.287788,23.657295,21.52066,21.146837,16.163645,13.570878,14.678635,15.086755,15.854982,14.79524,13.653188,12.006986,7.2604365,3.9954693,3.6765177,3.8617156,5.535354,13.107883,14.928994,14.562028,15.522313,20.059656,29.161781,39.505417,36.590267,25.859089,17.29884,25.430391,23.118849,18.252264,15.7966795,15.536031,12.05157,17.343424,24.61072,25.135447,20.591244,23.019392,18.025911,11.231899,8.056101,8.4264965,6.8111606,5.7891436,8.378482,9.866923,8.930646,7.658269,6.1629686,7.507367,11.0981455,15.049029,16.170506,20.755863,26.160892,29.67965,31.34643,33.942627,28.990303,24.212887,16.96617,9.551401,9.201583,9.136421,9.301042,11.019264,15.0456,21.568676,26.534718,22.504953,17.525192,14.932424,13.334236,16.835844,25.52985,25.005123,17.590355,22.343761,27.625326,18.718689,8.656279,4.705394,8.368194,7.531374,7.606825,11.609154,17.405157,17.730967,15.227368,12.099585,8.745448,7.781734,14.0750265,14.3974085,9.554831,6.842027,8.916927,13.7938,10.017825,7.284444,12.061859,19.630959,14.088745,10.388221,9.81205,9.427936,9.784613,14.932424,11.149589,17.034761,18.694681,12.175035,3.4638834,33.82602,21.328604,8.766026,10.264755,11.279913,8.669997,6.691125,5.641671,6.3138704,9.9801,6.7185616,9.582268,23.70188,33.74028,3.9200184,3.789694,4.012617,4.506478,5.192395,5.970912,6.7391396,8.501947,10.652299,11.22161,6.8728933,3.9508848,5.6793966,9.431366,12.624311,12.7272,11.118723,6.166398,3.590778,4.2526884,4.139512,2.6990852,1.8348293,1.7319417,2.3801336,3.5359046,6.3824625,10.22703,13.718349,16.352274,18.451181,14.767803,14.46943,21.311457,32.948048,40.938984,27.453848,20.779871,19.651537,21.548098,22.679861,28.249512,31.850578,26.088871,13.560589,6.8454566,4.8117113,4.928317,5.7377,6.3001523,6.193835,7.31531,8.580828,8.697433,7.613684,6.495639,8.340756,9.695444,8.498518,5.9983487,6.7459984,8.100685,10.2921915,12.264205,12.737488,10.203023,9.547972,6.8557453,5.456474,6.4373355,8.652849,6.5882373,5.0106273,5.2815647,6.6293926,6.15268,3.940596,4.448175,3.8925817,2.170929,2.860276,3.2135234,3.4021509,3.4604537,3.3850029,3.1483612,4.7671266,4.3349986,2.6407824,0.91912943,0.84367853,0.77508676,0.90198153,0.77851635,0.44927597,0.45613512,0.45613512,0.4389872,0.65162164,1.0048691,1.097468,1.7353712,1.2243627,0.72707254,0.64133286,0.5658819,0.47671264,0.3806842,0.2469303,0.1097468,0.06859175,0.25721905,0.48700142,0.48357183,0.37725464,0.70306545,0.9911508,1.3375391,1.9582944,2.585909,2.4315774,1.6324836,1.3101025,1.0906088,0.7682276,0.31895164,0.2709374,0.1920569,0.18519773,0.26407823,0.33266997,1.9994495,1.9548649,1.2003556,0.48357183,0.30866286,0.22635277,0.14404267,0.1371835,0.23664154,0.40126175,0.45270553,0.274367,0.16462019,0.6036074,2.2326615,1.2415106,0.6036074,1.1008976,2.585909,4.0057583,2.4967396,2.037175,2.1469216,2.4075704,2.4487255,2.6956558,1.9857311,1.4198492,1.3169615,1.2003556,0.9842916,0.88826317,0.939707,1.0357354,0.9534253,0.86082643,0.9945804,1.0117283,0.823101,0.5693115,0.6824879,0.7339317,0.8779744,1.0288762,0.8779744,0.5144381,0.30866286,0.32581082,0.4081209,0.18519773,0.5041494,0.89512235,0.77851635,0.26064864,0.11317638,0.14061308,0.18862732,0.13375391,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.041155048,0.05144381,0.06516216,0.08573969,0.09602845,0.13032432,0.18176813,0.22292319,0.18176813,0.3018037,0.34295875,0.38754338,0.44584638,0.4664239,0.34295875,0.30866286,0.34638834,0.4081209,0.4355576,0.59674823,0.89169276,1.0288762,0.96371406,0.90884066,0.9911508,1.2037852,1.4541451,1.6873571,1.8725548,1.8416885,1.8588364,1.8485477,1.8039631,1.7971039,1.7765263,1.8108221,1.7662375,1.6256244,1.5055889,1.4610043,1.4232788,1.4815818,1.605047,1.646202,1.6016173,1.6187652,1.5638919,1.4438564,1.3786942,1.4987297,1.4610043,1.5638919,1.7833855,1.7353712,2.0406046,2.136633,2.0440342,1.937717,2.1743584,2.301253,1.7902447,1.2929544,1.08032,1.0631721,1.0666018,1.0906088,1.1351935,1.1832076,1.1866373,1.039165,1.1420527,1.2758065,1.3958421,1.6290541,1.8039631,1.728512,1.5330256,1.3169615,1.1592005,1.1660597,0.7407909,0.39097297,0.29151493,0.2777966,0.3566771,0.5418748,0.6824879,0.7373613,0.7922347,0.8711152,0.939707,0.91569984,0.85396725,0.9294182,0.9534253,1.155771,1.3443983,1.3889829,1.2209331,1.1454822,1.0117283,0.88826317,0.7510797,0.48014224,0.3018037,0.24007112,0.20234565,0.15776102,0.13375391,0.09602845,0.07545093,0.07888051,0.106317215,0.16119061,0.37039545,0.4972902,0.5178677,0.4972902,0.5624523,0.607037,0.5796003,0.5418748,0.53158605,0.5693115,0.5727411,0.5658819,0.5418748,0.53158605,0.59674823,0.65848076,0.83681935,1.0666018,1.2963841,1.5021594,1.5090185,1.3546871,1.2277923,1.196926,1.2072148,0.9602845,0.83338976,0.72707254,0.59674823,0.45270553,0.26407823,0.17833854,0.13032432,0.08916927,0.0548734,0.044584636,0.041155048,0.030866288,0.024007112,0.0274367,0.037725464,0.08573969,0.14747226,0.22635277,0.3566771,0.5212973,0.66533995,0.7373613,0.78537554,0.9534253,1.1043272,1.255229,1.2380811,1.0940384,1.0700313,0.939707,0.85739684,0.8162418,0.7888051,0.7339317,0.6962063,0.6893471,0.75450927,0.90541106,1.1523414,1.3924125,1.488441,1.6153357,1.7971039,1.9239986,0.0,0.0,0.037725464,0.06859175,0.072021335,0.061732575,0.15776102,0.15433143,0.13032432,0.1371835,0.19891608,0.15090185,0.09259886,0.0548734,0.048014224,0.061732575,0.34295875,0.39440256,0.4355576,0.5453044,0.65505123,0.6310441,0.71678376,0.69963586,0.53844523,0.36696586,0.42869842,0.45956472,0.607037,0.7099246,0.31895164,0.18519773,0.216064,0.4046913,0.7888051,1.4335675,3.789694,6.101236,7.4936485,8.080108,8.971801,8.131552,6.8214493,6.3618846,6.914048,7.4765005,7.0615206,6.252138,6.5642304,8.090397,9.506817,11.677745,15.316538,18.20425,20.100813,22.751883,24.27805,26.726774,30.742823,35.890633,40.6509,45.116222,52.424675,63.7526,85.80485,130.80104,176.54144,183.26001,165.7794,135.87683,102.29774,75.3206,75.27602,86.110085,93.703186,85.87687,67.0793,50.672153,36.624565,24.7822,14.832966,12.792361,10.316199,8.258447,6.5779486,4.3178506,4.5510626,4.6436615,4.530485,4.2698364,4.07435,4.355576,4.8288593,5.0346346,4.8117113,4.2869844,3.4947495,2.9391565,2.5481834,2.287535,2.1674993,2.3492675,2.6887965,2.9220085,2.9151495,2.6716487,2.2292318,1.7010754,1.4198492,1.4781522,1.7079345,1.4027013,1.0528834,0.84367853,0.7990939,0.7613684,0.9568549,1.0357354,1.0700313,1.0906088,1.0528834,1.1489118,1.0734608,0.922559,0.7613684,0.6241849,0.6241849,0.5796003,0.5178677,0.4938606,0.5796003,0.72707254,0.96371406,1.2449403,1.6393428,2.335549,2.8705647,3.3369887,3.9200184,4.6779575,5.5079174,6.5230756,7.380472,7.2192817,6.9071894,9.016385,10.837497,9.791472,9.239308,10.110424,10.878652,12.562579,13.653188,14.435134,15.114192,15.824117,15.004445,13.869251,14.167625,16.067617,18.142517,21.486366,22.892496,23.36578,23.345201,22.673002,24.84736,29.539038,36.56283,42.862984,42.496017,35.636845,32.317,30.766829,29.648783,28.060884,34.49479,37.451096,36.291893,32.176388,28.060884,27.302946,26.702768,27.368109,28.67478,28.2598,25.19718,22.46037,21.431492,20.995934,17.576635,17.466888,20.70785,22.343761,20.484926,16.2974,16.479168,14.448852,12.644889,11.900668,11.399949,16.575195,17.566347,16.417435,14.7197895,13.594885,6.8454566,3.6936657,3.1243541,4.0503426,5.295283,6.492209,12.932974,20.128248,24.902235,25.389236,45.421455,51.821068,39.498558,19.764713,20.340883,16.348843,14.078457,16.856422,21.352612,17.593784,25.063425,33.212124,32.32729,24.837072,25.313786,17.86815,9.496528,4.835718,4.064061,2.9288676,2.942586,4.976331,7.5519514,9.208443,8.498518,7.181556,9.067829,12.30193,15.841265,19.456049,23.386356,23.142857,21.390337,17.778982,8.944365,9.870353,14.30481,16.03675,13.251926,8.529384,8.882631,9.410788,11.015835,16.417435,30.149504,23.046827,18.523201,19.733847,23.074265,18.20425,14.040731,21.688711,25.368658,20.522652,13.810948,18.056778,15.110763,9.156999,5.3158607,9.613133,10.113853,7.56567,8.676856,15.0078745,22.978235,13.629181,7.840037,5.5147767,6.276145,9.462232,13.416546,10.329918,10.981539,15.854982,15.138199,12.672326,6.910619,9.205012,15.676644,7.2192817,5.8988905,5.9640527,6.958633,8.488229,10.209882,9.074688,14.997586,15.820687,9.873782,5.967482,25.447538,15.169065,5.188966,10.525404,31.140654,19.154245,10.7757635,6.3138704,6.5367937,12.665466,7.438775,11.279913,15.412566,13.649758,2.3801336,7.349606,7.7748747,6.3001523,4.4104495,2.4555845,4.7774153,7.864044,13.906977,18.344864,9.887501,3.391862,3.9474552,9.465661,14.836395,11.931535,6.6225333,4.040054,4.0846386,5.2164025,4.4721823,3.0797696,2.393852,1.8691251,1.7559488,3.0969174,9.517105,13.522863,14.870691,14.143619,12.7272,11.444533,13.474849,19.562366,26.93941,29.34355,22.456938,19.637817,20.327166,22.789608,24.11,25.293207,21.873909,16.03675,10.031544,6.1492505,3.940596,3.9474552,4.647091,5.096367,4.914599,5.6828265,7.3118806,8.351046,8.423067,8.241299,9.849775,9.5205345,7.7714453,6.135532,7.1712675,8.244728,8.762596,10.072699,11.567999,10.666017,11.787492,9.314759,6.584808,6.135532,9.688584,6.941485,5.2575574,5.3673043,6.468202,6.2247014,4.0537724,3.6456516,3.1655092,3.2512488,7.034084,5.192395,3.6593697,2.8156912,2.6236343,2.6236343,3.199805,5.675967,4.5784993,0.58988905,0.5658819,0.7476501,0.8196714,0.66876954,0.44584638,0.5796003,0.274367,0.19891608,0.34981793,0.64819205,0.91569984,1.611906,1.3546871,0.9328478,0.7339317,0.7476501,0.5041494,0.29494452,0.20920484,0.20577525,0.106317215,0.12003556,0.12346515,0.12689474,0.21263443,0.5178677,1.0940384,1.3821237,1.4267083,1.4198492,1.7250825,1.4815818,1.0700313,0.9259886,0.90541106,0.31895164,0.31895164,0.23664154,0.21263443,0.2709374,0.31895164,0.6379033,0.6241849,0.4424168,0.23664154,0.1371835,0.17490897,0.1920569,0.31552204,0.40126175,0.061732575,0.17147937,0.18862732,0.25721905,0.45270553,0.7922347,0.5727411,0.4355576,0.8093826,1.6873571,2.6407824,1.786815,0.9294182,0.5761707,0.9945804,2.2292318,2.7402403,1.862266,1.1592005,1.0768905,0.9294182,0.78537554,0.939707,1.214074,1.4267083,1.4027013,0.7579388,0.99801,1.2415106,1.08032,0.5796003,0.5178677,0.47671264,0.48357183,0.52472687,0.548734,0.53844523,0.4698535,0.5727411,0.69963586,0.31895164,0.2469303,0.39440256,0.42869842,0.2709374,0.07545093,0.07545093,0.048014224,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.041155048,0.044584636,0.061732575,0.12346515,0.17147937,0.15433143,0.13032432,0.12346515,0.12346515,0.28122616,0.3018037,0.25378948,0.22292319,0.31895164,0.23664154,0.2777966,0.33952916,0.37382504,0.4115505,0.6790583,0.8848336,1.0254467,1.08032,1.0082988,1.3238207,1.5501735,1.488441,1.2277923,1.1283343,1.4095604,1.7456601,1.8862731,1.8108221,1.7250825,1.8108221,1.6667795,1.5124481,1.430138,1.3581166,1.3821237,1.3615463,1.4335675,1.546744,1.4507155,1.4267083,1.5193073,1.5501735,1.4644338,1.3443983,1.5501735,1.4747226,1.4918705,1.6770682,1.786815,2.1743584,2.201795,2.1194851,2.0646117,2.0303159,2.1743584,1.762808,1.1729189,0.82996017,1.2209331,1.4404267,1.3855534,1.3169615,1.2963841,1.1763484,1.2243627,1.2003556,1.255229,1.3855534,1.4335675,1.5673214,1.6016173,1.4987297,1.3546871,1.4027013,1.2929544,0.85396725,0.5418748,0.47328308,0.4115505,0.32581082,0.432128,0.53844523,0.5727411,0.61046654,0.70649505,0.7510797,0.7133542,0.67219913,0.7922347,0.8162418,0.823101,0.939707,1.1351935,1.2209331,1.1832076,1.0460242,1.039165,1.0768905,0.7476501,0.5041494,0.34295875,0.2503599,0.20920484,0.18176813,0.13375391,0.11317638,0.09945804,0.08916927,0.07545093,0.18519773,0.4046913,0.5212973,0.51100856,0.548734,0.53844523,0.52472687,0.52472687,0.53501564,0.53501564,0.6927767,0.7956643,0.8265306,0.8025235,0.77851635,0.70649505,0.6962063,0.8848336,1.1729189,1.2209331,1.2586586,1.2586586,1.2072148,1.1111864,0.9774324,0.96371406,1.1077567,1.2346514,1.196926,0.85396725,0.5007198,0.29151493,0.17833854,0.116605975,0.09259886,0.09259886,0.082310095,0.06516216,0.041155048,0.01371835,0.01371835,0.024007112,0.041155048,0.08916927,0.19891608,0.33266997,0.4389872,0.5796003,0.7442205,0.85396725,1.039165,1.2037852,1.1592005,0.94999576,0.84024894,0.8162418,0.8265306,0.88826317,0.939707,0.85396725,0.8162418,0.7888051,0.764798,0.72707254,0.64133286,0.8128122,1.039165,1.1729189,1.2312219,1.3889829,0.0,0.037725464,0.0274367,0.034295876,0.0548734,0.01371835,0.030866288,0.082310095,0.13032432,0.16462019,0.18519773,0.058302987,0.034295876,0.041155048,0.048014224,0.061732575,0.17490897,0.1920569,0.34981793,0.6036074,0.64476246,0.7476501,0.7305021,0.6790583,0.6379033,0.6241849,0.5555932,0.59674823,0.6927767,0.7099246,0.41840968,0.42183927,0.30866286,0.31209245,0.5521636,1.0425946,2.6956558,4.756838,6.0669403,6.5882373,7.4113383,7.366754,6.375603,5.5662203,5.254128,4.9248877,4.5990767,4.479041,5.0003386,6.186976,7.6514096,9.568549,11.657167,13.38225,15.1862135,18.478617,19.905325,21.599543,24.322634,28.09518,32.19011,37.039543,44.155937,53.895966,71.0199,104.67787,127.95791,128.54437,111.33127,85.259544,63.296467,55.624477,63.001522,73.91104,77.72474,64.67516,46.7247,32.039207,21.098822,13.732068,9.095266,6.800872,4.8905916,3.625074,3.0317552,2.901431,3.5530527,3.789694,3.7142432,3.549623,3.6456516,3.7622573,3.957744,4.1600895,4.2423997,4.029765,3.6970954,3.1826572,2.5721905,2.0234566,1.762808,1.762808,1.8862731,2.0680413,2.2326615,2.2909644,2.1743584,1.9068506,1.7250825,1.6427724,1.4644338,1.2655178,1.1180456,0.9568549,0.7888051,0.7133542,1.0357354,1.2037852,1.3306799,1.4267083,1.371835,0.939707,0.7682276,0.72707254,0.6962063,0.5521636,0.5521636,0.47671264,0.42183927,0.4664239,0.6790583,0.83338976,1.0597426,1.3684053,1.821111,2.5173173,3.210094,3.625074,3.9474552,4.804852,7.267296,8.172707,8.879202,8.457363,7.8777623,10.017825,11.592006,11.657167,11.550851,11.746337,11.832077,14.688923,15.724659,15.573756,15.343974,16.616352,14.791811,14.500296,15.995596,18.571217,20.560377,22.275171,20.927343,20.392326,22.20658,25.567575,28.715937,33.702557,39.40596,44.601784,47.976498,46.282284,38.966972,30.4273,24.096281,22.470657,23.94195,24.120289,23.290329,22.570116,23.873358,21.486366,19.929333,20.330595,21.925352,22.04539,24.68617,23.053686,19.658396,16.324837,14.184773,14.514014,15.265094,15.693792,15.031882,12.476839,12.826657,13.176475,12.734058,11.763485,11.605724,13.402828,11.118723,9.571979,10.528833,12.703192,8.453933,5.120374,3.4398763,3.4433057,4.465323,5.768566,14.222499,20.227707,22.062536,25.879667,38.42167,43.672367,34.961216,18.941612,15.580616,16.431154,15.848124,15.885849,16.12592,13.673765,16.743246,18.437462,18.36544,18.272842,22.017952,13.975569,8.107545,5.6176643,5.219832,3.1380725,3.0900583,3.542764,4.5784993,6.4133286,9.427936,9.349055,9.647429,11.180455,14.109323,17.916164,20.02193,21.136547,20.62211,18.341434,14.678635,15.155347,16.153357,17.03819,15.748666,8.796892,8.584257,7.4936485,8.189855,12.079007,19.301718,12.919256,9.325048,13.865822,20.749004,13.029003,8.906639,13.845244,17.734396,18.766703,23.427511,26.726774,24.562706,16.599203,7.658269,7.6959944,14.640909,13.821238,11.866373,13.190193,19.987637,13.735497,10.343636,9.592556,10.991828,13.80409,17.899017,15.755525,12.048141,9.818909,10.47396,10.048691,6.0223556,9.674867,16.647217,6.9380555,6.5470824,6.5196457,8.06296,11.012405,13.845244,15.062748,23.389786,24.336353,17.95046,18.818146,18.389448,13.430264,17.305698,28.637054,31.277838,19.816156,13.728639,9.071259,6.0497923,9.002667,8.162418,13.5503,16.448301,12.476839,1.611906,15.055889,18.149376,12.7272,4.8082814,4.5922174,6.0326443,14.812388,23.70188,23.708738,4.091498,3.3850029,11.598865,14.627191,10.271614,8.244728,6.7357097,6.0840883,5.960623,6.036074,5.98463,5.099797,3.5359046,2.486451,2.9906003,5.953764,10.988399,15.107333,15.913286,13.848674,12.188754,12.830087,15.0078745,18.6158,21.85676,21.211998,20.255144,21.253153,22.172283,22.035099,20.910194,18.560926,14.291091,10.350495,7.5931067,5.4907694,3.7313912,3.175798,3.5187566,4.232111,4.547633,4.73969,6.15268,8.98209,12.349944,14.29452,12.253916,9.06097,7.006647,6.893471,8.038953,9.033533,10.000677,11.327928,12.932974,14.2533655,11.149589,8.282454,6.0052075,5.164959,7.1266828,5.103226,4.65395,5.0449233,5.0895076,3.1243541,2.1743584,2.527606,3.6010668,5.377593,8.388771,6.3310184,4.3487167,3.1517909,2.6819375,2.136633,2.318401,3.175798,2.5481834,0.69963586,0.34638834,0.42183927,0.31895164,0.22978236,0.26407823,0.45613512,0.2194936,0.41840968,1.5364552,2.6853669,1.587899,1.1214751,1.0563129,1.0494537,1.0220171,1.1489118,0.8265306,0.4629943,0.28465575,0.2709374,0.14404267,0.116605975,0.09602845,0.08573969,0.15090185,0.39783216,0.980862,1.5433143,1.7079345,1.5913286,1.8108221,1.1077567,0.72364295,0.66191036,0.6756287,0.2469303,0.29494452,0.25378948,0.25378948,0.29837412,0.26064864,0.42869842,0.4389872,0.3806842,0.3018037,0.23664154,0.17490897,0.21263443,0.33266997,0.39097297,0.09602845,0.16804978,0.32238123,0.5555932,0.7956643,0.90198153,0.8093826,0.6824879,0.6756287,0.8471081,1.1626302,1.4404267,1.3752645,1.3032433,1.4815818,2.0817597,2.2429502,1.9137098,1.5570327,1.3306799,1.0768905,0.72707254,0.64133286,0.7922347,0.9945804,0.90198153,0.4629943,0.490431,0.53501564,0.4424168,0.36010668,0.5624523,0.4972902,0.36696586,0.34638834,0.58645946,0.6824879,0.64133286,0.77851635,0.864256,0.12346515,0.18862732,0.20234565,0.16804978,0.11317638,0.06516216,0.044584636,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.058302987,0.09259886,0.09259886,0.08573969,0.14747226,0.32238123,0.32238123,0.2469303,0.15433143,0.08573969,0.1371835,0.20577525,0.24350071,0.2503599,0.2709374,0.19548649,0.24007112,0.3018037,0.35324752,0.44927597,0.58988905,0.7407909,0.8471081,0.9328478,1.1043272,0.91569984,0.9774324,1.097468,1.1454822,1.0563129,1.3375391,1.5844694,1.6256244,1.5227368,1.5638919,1.5330256,1.3546871,1.2209331,1.2175035,1.3101025,1.471293,1.6873571,1.7696671,1.646202,1.3512574,1.2895249,1.4095604,1.5364552,1.587899,1.5638919,1.5364552,1.4369972,1.4815818,1.6530612,1.7250825,2.0165975,2.0989075,2.1297739,2.153781,2.07833,1.9308578,2.551613,2.2155135,1.039165,0.9877212,1.1214751,1.2620882,1.3101025,1.2895249,1.3821237,1.5673214,1.4369972,1.3958421,1.4815818,1.3855534,1.2380811,1.1626302,1.2209331,1.3443983,1.3546871,1.255229,0.84024894,0.5590228,0.5624523,0.71678376,0.6036074,0.51100856,0.4698535,0.4664239,0.4629943,0.69963586,0.90541106,0.96714365,0.8848336,0.7922347,0.8093826,1.0254467,1.2758065,1.4267083,1.3684053,1.5364552,1.5227368,1.4095604,1.2277923,0.9568549,0.8265306,0.6893471,0.5521636,0.4664239,0.5007198,0.35324752,0.28465575,0.26064864,0.22635277,0.1371835,0.14061308,0.23664154,0.30523327,0.35324752,0.52472687,0.58988905,0.64133286,0.6756287,0.6824879,0.64476246,0.99801,1.2826657,1.313532,1.1283343,0.99801,0.85739684,0.7339317,0.7888051,1.0117283,1.2449403,1.4575747,1.3992717,1.3992717,1.471293,1.3169615,1.1592005,1.1043272,1.1454822,1.2243627,1.2312219,1.0734608,0.7682276,0.5178677,0.3806842,0.28808534,0.18862732,0.16462019,0.15090185,0.11317638,0.041155048,0.010288762,0.0034295875,0.01371835,0.030866288,0.06516216,0.17833854,0.31895164,0.4629943,0.5624523,0.52472687,0.64133286,0.8676856,1.08032,1.2003556,1.2175035,1.0357354,0.91569984,0.90884066,0.96714365,0.939707,0.9534253,0.84024894,0.7407909,0.7099246,0.7510797,0.7442205,0.7510797,0.8162418,0.96371406,1.1797781,0.0,0.020577524,0.010288762,0.010288762,0.0274367,0.037725464,0.006859175,0.024007112,0.06859175,0.09602845,0.072021335,0.01371835,0.08916927,0.09945804,0.030866288,0.041155048,0.072021335,0.12346515,0.32924038,0.5555932,0.40126175,0.66191036,0.6790583,0.71678376,0.7888051,0.65848076,0.53158605,0.5041494,0.6001778,0.7442205,0.7613684,0.65162164,0.42183927,0.32238123,0.48014224,0.8711152,2.1434922,3.99204,5.086078,5.2506986,5.4633327,6.420188,5.844017,5.0243454,4.5030484,4.0846386,3.2889743,3.083199,3.6079261,4.664239,5.693115,6.9792104,8.429926,9.863494,11.790922,15.450292,15.981877,16.815268,18.842154,22.333473,26.908543,30.5199,37.142433,47.63011,64.966675,94.28279,113.673676,107.56901,86.55936,61.050087,41.285374,37.694595,45.754128,58.892876,66.93526,56.132057,36.96752,23.19773,14.441993,9.496528,6.351596,4.149801,2.7230926,2.3081124,2.8156912,3.8479972,4.9351764,5.288424,5.0826488,4.5784993,4.125794,3.7382503,3.5702004,3.542764,3.5393343,3.3815732,3.309552,3.0626216,2.6819375,2.253239,1.8999915,1.646202,1.5021594,1.5536032,1.7696671,1.978872,2.0886188,2.0268862,1.9137098,1.7388009,1.3855534,1.1351935,1.0014396,0.85739684,0.72021335,0.7305021,1.0185875,1.155771,1.2003556,1.1763484,1.0940384,0.6036074,0.47671264,0.48700142,0.48014224,0.37725464,0.4081209,0.45956472,0.5453044,0.6824879,0.8745448,1.1454822,1.4438564,1.6770682,1.862266,2.1332035,2.5138876,2.603057,2.9048605,3.7519686,5.3158607,6.5333643,8.536243,11.063849,13.978998,17.29884,15.429714,13.965281,13.37882,13.591455,13.982429,15.234227,16.54433,17.556059,18.241976,18.910746,17.189093,17.250826,18.482046,19.939621,20.35803,20.478067,19.061647,20.36832,24.957108,29.713945,29.5116,31.212675,32.24498,32.67025,35.18414,34.607967,28.544456,23.845922,22.117409,19.737276,18.303709,18.482046,17.388008,15.436573,16.317978,15.0250225,15.9578705,17.62808,18.416885,16.592344,18.95876,19.709839,18.166525,15.062748,12.538571,12.744347,13.516005,14.726648,15.477728,14.119612,12.744347,12.099585,11.276484,10.659158,11.931535,11.008976,9.050681,9.534253,12.459691,14.359683,9.657719,6.3378778,3.8925817,3.0729103,5.895461,6.728851,10.275044,14.572317,17.439453,16.479168,23.02625,28.520449,28.160343,23.03654,20.12139,18.79071,15.920145,15.340545,16.746675,15.697222,16.03675,15.237658,13.598314,13.701202,20.399187,14.637479,9.839486,6.560801,4.773986,3.8308492,5.518206,6.8866115,6.2487082,4.887162,7.051232,9.325048,12.260776,13.004995,11.828648,12.113303,13.437123,15.268523,16.506605,17.364002,19.380598,17.051908,14.352823,11.873232,10.271614,10.257896,10.834066,9.599416,11.029553,14.167625,12.63117,8.114404,8.093826,12.397959,16.7844,12.932974,11.756626,13.656617,14.935853,15.762384,20.155685,19.023922,20.409475,17.693241,11.008976,7.2364297,12.452832,13.498857,12.583157,12.744347,17.86815,13.780083,10.4533825,9.112414,11.434244,19.552078,18.506054,13.231348,11.173596,13.594885,15.570327,11.194174,8.268735,10.998687,16.609491,15.361122,8.128122,6.800872,8.224151,11.664027,18.773561,16.331696,21.592682,25.337791,24.387796,21.592682,16.897577,13.426835,15.659496,22.326614,26.394106,22.714157,17.638369,12.000127,8.344186,10.916377,8.498518,10.532263,15.9613,18.440891,6.324159,9.534253,14.273943,18.46147,18.804428,10.786053,7.9257765,22.220297,36.545685,34.779446,1.8073926,2.843128,19.939621,21.260014,6.3173003,5.960623,8.937505,8.882631,7.6033955,6.4373355,6.2898636,4.2286816,2.884283,3.5461934,6.9723516,13.38911,13.653188,12.524854,11.917816,12.360233,12.9981365,14.356253,16.702091,18.53692,18.982767,17.799559,18.272842,19.147387,18.694681,16.664366,14.270514,11.825217,9.1981535,6.992929,5.435896,4.355576,3.0283258,2.5619018,3.350707,4.65395,4.6127954,4.249259,5.4016004,9.458802,15.597764,20.76958,14.688923,8.64256,5.4736214,5.761707,7.8331776,8.532814,9.983529,11.194174,12.05157,13.341095,9.97324,7.130112,5.171818,4.530485,5.689686,4.1155047,3.9337368,5.038064,5.56965,1.9102802,2.3767042,2.9117198,4.307562,6.444195,8.289313,4.8425775,3.093488,2.6064866,2.6785078,2.3252604,1.4507155,1.4267083,1.4164196,1.0700313,0.53844523,0.39440256,0.216064,0.13032432,0.17147937,0.25378948,0.14404267,0.25378948,1.546744,3.1106358,2.1743584,0.97057325,0.6927767,0.6790583,0.66191036,0.7476501,0.5521636,0.31895164,0.23664154,0.26750782,0.16119061,0.17490897,0.106317215,0.072021335,0.15776102,0.4115505,0.9328478,1.9308578,2.1880767,1.821111,2.2806756,1.1317638,0.6344737,0.4629943,0.3566771,0.09259886,0.15090185,0.20577525,0.22292319,0.22635277,0.29151493,0.3566771,0.34638834,0.32581082,0.32924038,0.33266997,0.24007112,0.2469303,0.47328308,0.91227025,1.4438564,0.53158605,0.33266997,0.5041494,0.7510797,0.8196714,0.65848076,0.607037,0.8162418,1.2037852,1.4335675,1.7388009,1.7971039,1.8279701,1.8519772,1.6599203,1.5810398,1.7833855,1.6942163,1.2998136,1.1489118,0.78537554,0.5693115,0.64819205,0.86082643,0.7510797,0.5144381,0.32581082,0.20920484,0.18176813,0.24007112,0.4424168,0.41840968,0.31552204,0.29151493,0.5041494,0.47328308,0.45613512,0.6962063,0.9911508,0.6790583,0.47671264,0.216064,0.06516216,0.048014224,0.05144381,0.034295876,0.020577524,0.010288762,0.0034295875,0.010288762,0.0034295875,0.0,0.010288762,0.0274367,0.041155048,0.0548734,0.12346515,0.18176813,0.19548649,0.15090185,0.22978236,0.2469303,0.26064864,0.28122616,0.26750782,0.21263443,0.22635277,0.25721905,0.274367,0.29494452,0.18519773,0.18519773,0.20920484,0.24007112,0.31895164,0.45270553,0.6344737,0.7990939,0.90541106,0.90884066,0.89169276,1.1866373,1.4438564,1.4850113,1.3032433,1.4438564,1.4644338,1.4472859,1.4575747,1.5536032,1.4335675,1.1214751,0.9259886,0.9602845,1.1317638,1.3786942,1.605047,1.6976458,1.6153357,1.3924125,1.3341095,1.4335675,1.4781522,1.4369972,1.4541451,1.5364552,1.4404267,1.4644338,1.6153357,1.6187652,1.7696671,1.8519772,1.8519772,1.7765263,1.6221949,1.7182233,2.3561265,2.177788,1.2209331,0.9294182,1.0048691,1.0288762,1.0906088,1.1729189,1.1489118,1.2895249,1.4918705,1.6153357,1.611906,1.529596,1.3684053,1.1934965,1.2380811,1.5021594,1.7730967,1.4541451,1.1660597,0.980862,0.8779744,0.7476501,0.6173257,0.50757897,0.4972902,0.58645946,0.7305021,0.8745448,0.9774324,1.0288762,1.0014396,0.8471081,0.8162418,0.94656616,1.0837497,1.1454822,1.1214751,1.214074,1.2415106,1.2483698,1.2175035,1.0700313,0.97400284,0.89512235,0.7922347,0.71678376,0.8162418,0.61046654,0.490431,0.42869842,0.37725464,0.25378948,0.17147937,0.26064864,0.37039545,0.45270553,0.5658819,0.6927767,0.77165717,0.8265306,0.83681935,0.7339317,0.9774324,1.2380811,1.3169615,1.2037852,1.0906088,0.97400284,0.922559,0.99801,1.138623,1.1694894,1.3821237,1.313532,1.2860953,1.3443983,1.2586586,1.2449403,1.3958421,1.430138,1.3032433,1.2175035,1.2243627,1.1489118,1.0117283,0.86082643,0.7579388,0.607037,0.50757897,0.39440256,0.25721905,0.12689474,0.048014224,0.017147938,0.006859175,0.010288762,0.020577524,0.072021335,0.15090185,0.26064864,0.36696586,0.38754338,0.4629943,0.6790583,0.9568549,1.2209331,1.3855534,1.4953002,1.3786942,1.1900668,0.99801,0.7956643,0.84367853,0.8265306,0.8265306,0.8745448,0.97057325,0.91569984,0.8676856,0.89169276,0.9842916,1.0837497,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.006859175,0.01371835,0.030866288,0.030866288,0.0,0.0,0.08916927,0.09945804,0.020577524,0.024007112,0.024007112,0.07888051,0.22292319,0.34638834,0.18862732,0.4664239,0.548734,0.6379033,0.7373613,0.65162164,0.5761707,0.6241849,0.72707254,0.7922347,0.70649505,0.6173257,0.4424168,0.3566771,0.4664239,0.77508676,1.8279701,3.2512488,4.149801,4.32128,4.2526884,5.456474,5.209543,4.40359,3.6765177,3.415869,2.4144297,1.9994495,2.2600982,3.0420442,3.9543142,5.0620713,5.919468,6.9654922,8.742019,11.873232,12.319078,13.543441,15.570327,18.389448,21.969936,26.239773,32.231262,43.212803,62.219574,92.06042,117.62799,104.74989,78.225464,52.733337,32.800575,26.033998,31.106358,43.607204,53.78279,46.518925,29.813404,18.996485,12.572867,8.906639,6.2212715,4.122364,3.1209247,3.4227283,4.6882463,6.0395036,6.773435,6.691125,6.0806584,5.254128,4.554492,4.0194764,3.666229,3.3472774,3.0146074,2.7470996,3.1826572,3.0043187,2.651071,2.3286898,2.0303159,1.6427724,1.3924125,1.3375391,1.4472859,1.587899,1.8862731,1.8759843,1.7216529,1.4987297,1.1832076,1.0151579,0.89855194,0.7990939,0.75450927,0.8505377,0.9842916,0.980862,0.8848336,0.77508676,0.77508676,0.5453044,0.4355576,0.36353627,0.3018037,0.28122616,0.33952916,0.48700142,0.67219913,0.86082643,1.0151579,1.2415106,1.4644338,1.5810398,1.6221949,1.7593783,1.9068506,1.9308578,2.294394,3.0557625,3.8685746,6.2898636,10.220171,15.011304,19.288,20.937632,16.335125,13.461131,12.956982,13.992717,14.270514,14.356253,15.851553,17.20281,17.641798,17.20281,17.748116,18.54035,19.061647,19.1954,19.222837,19.483486,19.558937,22.223726,26.545008,27.85854,26.490133,26.534718,25.495554,23.773901,24.669024,24.367218,22.755312,23.091412,23.983105,19.394318,16.492886,17.353712,16.300829,13.004995,12.459691,12.816368,14.3974085,16.46888,17.727537,16.304258,16.21166,16.952452,16.650646,14.774663,12.130451,13.111313,14.352823,15.563468,16.273392,15.858413,13.3033695,12.21962,11.266195,10.655728,12.171606,9.465661,8.172707,10.446524,14.424845,14.205351,10.034973,8.117833,6.2075534,4.5784993,6.0052075,7.058091,7.740579,10.244178,12.795791,9.685155,12.524854,16.510035,19.576086,20.53294,19.075365,16.331696,12.449403,12.202472,14.994157,14.832966,12.500846,11.821788,10.88894,10.597425,14.637479,12.329367,10.425946,7.579388,4.523626,4.057202,7.9292064,11.780633,11.355364,7.589677,6.6053853,8.934075,12.521424,13.166186,10.662587,8.820899,8.64599,9.712592,12.061859,15.29253,18.581505,16.420864,11.667457,7.6616983,6.7974424,10.532263,10.686595,12.744347,15.854982,16.438013,8.176137,7.5759587,11.941824,14.723219,14.486577,14.915276,13.828096,13.413116,12.843805,12.425395,13.6086035,11.97269,17.031332,18.28656,13.169616,7.06495,10.449953,11.777204,12.415107,14.191633,19.349733,17.947031,14.644339,12.493987,14.452282,23.36578,17.892159,11.183885,11.351934,17.051908,17.480608,11.338216,10.175586,11.482259,13.872682,17.072487,10.779194,10.573419,13.557159,17.20967,19.384027,15.9613,18.722118,26.274069,31.137224,19.744135,22.096832,19.565796,16.033321,14.832966,18.746124,19.308577,15.920145,11.2250395,8.940934,13.869251,10.257896,7.689135,11.4376745,17.63494,13.265644,6.468202,9.3079,16.931873,21.146837,10.412228,7.9875093,20.639257,32.41989,30.070623,3.0043187,9.671436,21.20514,18.053349,3.649081,4.420738,8.237869,8.337327,7.6925645,7.3255987,6.3138704,3.0283258,2.1160555,3.99204,8.279024,13.821238,11.489118,10.545981,10.947243,12.061859,12.686044,14.263655,16.527182,17.36057,16.640358,16.252815,16.815268,16.62321,15.011304,12.21962,9.417647,7.7440085,6.824879,5.686256,4.184097,3.000889,2.1469216,1.879414,2.668219,3.9886103,4.3109913,4.184097,4.8940215,8.501947,14.863832,21.62012,15.13134,8.224151,4.65395,4.9591837,6.468202,6.5299344,8.237869,9.39707,9.55826,10.024684,8.179566,6.193835,5.0586414,5.0483527,5.7068334,3.8137012,3.4638834,4.5956473,5.2644167,1.6736387,3.1586502,3.8925817,4.931747,7.2192817,11.585147,5.40503,3.000889,3.5050385,4.8185706,3.5942078,1.5433143,0.8196714,0.9431366,1.3512574,1.3684053,0.5727411,0.22292319,0.15776102,0.20577525,0.18519773,0.15090185,0.12346515,1.0048691,2.2429502,1.8108221,0.70306545,0.37382504,0.3018037,0.25721905,0.3018037,0.29151493,0.19548649,0.16804978,0.2194936,0.216064,0.20234565,0.15090185,0.15433143,0.41840968,1.2792361,1.2655178,1.6907866,2.3904223,2.976882,2.8054025,1.2998136,0.58645946,0.32581082,0.2194936,0.006859175,0.041155048,0.13032432,0.15433143,0.15433143,0.31895164,0.4389872,0.32581082,0.25378948,0.31552204,0.42526886,0.274367,0.23321195,0.39440256,0.7990939,1.4438564,0.77851635,0.38754338,0.36696586,0.6276145,0.89512235,0.59331864,0.58988905,0.9877212,1.5810398,1.8313997,1.961724,2.095478,2.2841053,2.352697,1.9171394,1.3238207,1.3581166,1.2826657,1.0288762,1.1866373,0.9774324,0.6824879,0.5761707,0.6344737,0.52472687,0.45956472,0.29837412,0.2469303,0.31209245,0.29494452,0.30866286,0.28122616,0.24350071,0.2503599,0.39440256,0.42869842,0.36010668,0.4664239,0.7133542,0.7613684,0.5624523,0.26407823,0.09602845,0.09602845,0.106317215,0.05144381,0.037725464,0.0274367,0.006859175,0.01371835,0.006859175,0.006859175,0.017147938,0.037725464,0.06516216,0.082310095,0.16119061,0.22635277,0.23664154,0.17147937,0.17490897,0.18176813,0.22978236,0.29494452,0.32238123,0.34638834,0.30866286,0.26064864,0.23664154,0.26064864,0.15433143,0.12689474,0.15090185,0.20577525,0.26407823,0.36353627,0.5212973,0.6790583,0.7990939,0.8676856,1.097468,1.4781522,1.6564908,1.5398848,1.2895249,1.3478279,1.313532,1.2895249,1.3203912,1.371835,1.1763484,0.8745448,0.7373613,0.823101,0.97400284,1.2346514,1.4438564,1.5707511,1.5707511,1.4095604,1.3032433,1.3512574,1.3306799,1.2415106,1.3169615,1.546744,1.5707511,1.6187652,1.7216529,1.7147937,1.6599203,1.6427724,1.6359133,1.5673214,1.313532,1.4232788,1.879414,1.8279701,1.2483698,0.9431366,0.9774324,0.8676856,0.864256,0.9842916,1.0151579,1.0528834,1.371835,1.587899,1.6084765,1.6324836,1.6324836,1.4027013,1.3238207,1.5158776,1.8348293,1.3752645,1.1180456,0.9602845,0.8093826,0.5761707,0.48014224,0.42526886,0.45270553,0.58302987,0.7956643,0.8676856,0.8505377,0.8505377,0.89169276,0.9328478,0.97057325,0.96714365,0.89855194,0.8162418,0.8745448,0.9328478,0.91227025,0.9945804,1.1420527,1.0906088,1.0220171,1.0082988,0.9602845,0.89855194,0.97057325,0.91912943,0.823101,0.7133542,0.58988905,0.4115505,0.29494452,0.37725464,0.5212973,0.6207553,0.6001778,0.6756287,0.72364295,0.78194594,0.83681935,0.8093826,0.96714365,1.138623,1.2003556,1.1454822,1.0837497,1.0323058,1.0871792,1.196926,1.2689474,1.2003556,1.3786942,1.2998136,1.2243627,1.2243627,1.196926,1.2758065,1.5055889,1.5741806,1.4232788,1.2586586,1.2963841,1.3203912,1.2723769,1.1763484,1.1523414,1.0700313,1.0185875,0.89512235,0.6824879,0.45270553,0.20577525,0.08916927,0.034295876,0.010288762,0.010288762,0.020577524,0.044584636,0.09945804,0.18519773,0.26064864,0.31209245,0.47328308,0.7099246,0.96714365,1.1763484,1.5158776,1.5261664,1.3992717,1.2106444,0.91912943,0.881404,0.89169276,0.9431366,1.0117283,1.0734608,1.0323058,1.0117283,1.0082988,1.0014396,0.980862,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.041155048,0.024007112,0.010288762,0.0034295875,0.017147938,0.0274367,0.024007112,0.01371835,0.01371835,0.020577524,0.048014224,0.082310095,0.09602845,0.2469303,0.3566771,0.42869842,0.50757897,0.65162164,0.6962063,0.8779744,0.94999576,0.77165717,0.3018037,0.37039545,0.4081209,0.4424168,0.5144381,0.69963586,1.5398848,2.4075704,3.1552205,3.642222,3.7176728,4.482471,4.461893,3.642222,2.5721905,2.393852,1.6393428,1.2037852,1.1008976,1.4507155,2.4555845,3.8788633,4.139512,4.588788,5.885172,8.001227,9.5033865,11.914387,14.116182,15.71437,17.010754,24.079134,29.76196,40.256496,60.720844,95.29452,133.6476,115.71085,81.84711,53.44326,32.900032,22.419212,23.835632,32.039207,38.870945,33.14353,22.254593,15.920145,12.103014,9.523964,7.6376915,5.7651367,5.113515,5.6793966,6.893471,7.630832,7.349606,6.526505,5.610805,4.931747,4.705394,4.506478,4.166949,3.5839188,2.9117198,2.5447538,3.3438478,3.059192,2.5310357,2.1674993,1.9445761,1.5913286,1.4095604,1.3032433,1.2277923,1.1763484,1.5810398,1.5090185,1.2620882,1.0288762,0.864256,0.90884066,0.85396725,0.8162418,0.8505377,0.9568549,0.922559,0.77508676,0.59331864,0.48014224,0.58645946,0.64819205,0.5041494,0.32238123,0.22292319,0.29837412,0.4081209,0.58302987,0.7510797,0.8711152,0.9602845,1.0220171,1.097468,1.1694894,1.2826657,1.5330256,1.704505,2.1023371,2.568761,3.234101,4.5030484,8.279024,13.145609,17.329706,19.188541,17.20624,12.771784,10.371073,10.834066,12.867812,13.011855,13.238208,14.387119,14.421415,13.272504,12.833516,16.62321,17.88873,17.442883,16.859852,18.471758,19.658396,21.462358,24.466677,26.35295,21.911634,22.076254,22.645567,23.019392,23.324625,24.391226,24.518122,26.236343,27.738503,26.802225,20.800447,18.015623,18.53692,17.473747,14.637479,14.555169,15.728088,15.45715,16.170506,18.193962,19.747564,18.145947,16.863281,16.088194,15.326826,13.392539,15.230798,16.077906,15.933864,15.512024,16.273392,13.941273,13.516005,12.902108,11.893809,12.154458,9.016385,7.4970784,9.513676,12.96727,11.753197,10.652299,10.275044,9.451943,7.8023114,5.7308407,6.464772,7.64798,8.669997,9.084977,8.601405,9.736599,10.6488695,11.146159,11.211322,10.984968,10.6488695,9.386781,9.80519,11.766914,12.38424,7.8091707,7.56567,9.469091,10.772334,8.155559,7.534804,8.81404,8.1487,5.4599032,4.4413157,9.06097,14.003006,14.973578,12.144169,10.131001,10.539123,11.30049,11.4754,10.875222,10.069269,8.354475,7.73372,9.424506,12.343085,13.121602,13.71492,9.352485,6.492209,7.1952744,9.139851,8.134981,15.268523,20.978786,19.274282,7.7440085,8.848335,16.654078,18.70497,14.79867,16.993607,13.173045,11.698323,11.231899,10.796341,9.788043,12.22305,18.296848,19.36688,14.037301,8.141841,10.569988,11.108434,12.092726,15.175924,21.321745,24.507832,22.426073,19.459478,19.03764,23.643576,17.46003,11.934964,12.027563,15.501736,12.936404,8.98209,11.362224,12.236768,10.333347,10.9541025,13.224489,16.12249,20.731855,23.410364,15.776102,15.590904,18.430603,27.625326,34.114105,16.479168,26.43526,25.056566,19.226267,13.862392,11.897239,12.507706,11.38623,8.604835,8.176137,18.056778,14.164196,8.357904,6.8214493,11.026124,17.724108,10.799771,10.676306,12.253916,11.406808,4.976331,13.306799,18.053349,18.080786,13.399398,5.195825,20.382038,16.077906,7.250148,2.3595562,3.3541365,4.7671266,4.962613,6.4236174,8.203573,5.9469047,2.5961976,2.054323,3.649081,5.970912,6.8728933,7.099246,12.754636,15.512024,13.334236,10.4705305,12.284782,14.4145565,14.850114,14.003006,14.7197895,15.453721,14.887839,13.173045,10.655728,7.8777623,6.9071894,6.869464,6.077229,4.15666,2.037175,1.5193073,1.2998136,1.4747226,2.1297739,3.3198407,3.99204,4.6265135,6.667118,10.690024,16.410576,13.790371,8.021805,4.8254294,5.1340923,5.0826488,4.3109913,5.672538,6.5230756,6.2830043,6.4407654,6.81802,6.1458206,5.9160385,6.351596,6.4064693,3.7382503,3.3747141,3.8720043,3.789694,1.7113642,3.7759757,4.972902,5.4084597,7.5382333,16.173935,8.652849,4.6402316,5.528495,8.368194,5.871454,2.3972816,1.0563129,0.94656616,1.4335675,2.1469216,0.7339317,0.2503599,0.22635277,0.3018037,0.23321195,0.19548649,0.13375391,0.4081209,0.82996017,0.6893471,0.29494452,0.1920569,0.14404267,0.08573969,0.12689474,0.24350071,0.18862732,0.12689474,0.14404267,0.24350071,0.17490897,0.22978236,0.30523327,0.7888051,2.5481834,1.6736387,0.8848336,2.1812177,4.4516044,3.474172,1.7662375,0.65505123,0.23321195,0.22635277,0.01371835,0.01371835,0.058302987,0.082310095,0.11317638,0.29151493,0.5624523,0.33952916,0.20234565,0.33266997,0.50757897,0.25378948,0.19891608,0.19891608,0.17147937,0.09602845,0.6859175,0.45613512,0.274367,0.5418748,1.2003556,0.8505377,0.7373613,1.0323058,1.5536032,1.7765263,1.8965619,2.2600982,2.5927682,2.7128036,2.5070283,1.4575747,0.84367853,0.5761707,0.64133286,1.0940384,1.0597426,0.7339317,0.42869842,0.2777966,0.20920484,0.23664154,0.30866286,0.4664239,0.58645946,0.37039545,0.20234565,0.14061308,0.13375391,0.17490897,0.31895164,0.59331864,0.52815646,0.3566771,0.2503599,0.31895164,0.45270553,0.32924038,0.20577525,0.17490897,0.17490897,0.06859175,0.06516216,0.058302987,0.020577524,0.01371835,0.017147938,0.017147938,0.024007112,0.048014224,0.08916927,0.14061308,0.20577525,0.2194936,0.18176813,0.18176813,0.20920484,0.21263443,0.20920484,0.21263443,0.20920484,0.3841138,0.33609957,0.23321195,0.16804978,0.16804978,0.11317638,0.09602845,0.16462019,0.28808534,0.3566771,0.42526886,0.52815646,0.6276145,0.7682276,1.0768905,1.3786942,1.5741806,1.5193073,1.2449403,0.9877212,1.0357354,1.0871792,1.0768905,1.0048691,0.96371406,0.7476501,0.6310441,0.67219913,0.8162418,0.89169276,1.1008976,1.3066728,1.4404267,1.4575747,1.3341095,1.1660597,1.1660597,1.1523414,1.1214751,1.2586586,1.5810398,1.8348293,1.9480057,1.9514352,1.9548649,1.7388009,1.611906,1.670209,1.7216529,1.2998136,1.0494537,1.4335675,1.6187652,1.4267083,1.2929544,0.9774324,0.77851635,0.70649505,0.7956643,1.0700313,1.0460242,1.1592005,1.3238207,1.471293,1.5604624,1.6736387,1.4815818,1.3341095,1.3546871,1.4438564,1.039165,0.70649505,0.4972902,0.4081209,0.36696586,0.32581082,0.31895164,0.34295875,0.4115505,0.5624523,0.6379033,0.59331864,0.5555932,0.6310441,0.89855194,1.0425946,1.0014396,0.823101,0.65505123,0.7407909,0.8505377,0.7888051,0.85396725,1.0323058,1.0151579,0.9911508,1.0528834,1.0700313,1.0185875,0.9774324,1.1832076,1.1763484,1.0323058,0.8196714,0.61389613,0.5178677,0.52472687,0.6207553,0.70649505,0.59674823,0.5453044,0.5418748,0.59331864,0.70306545,0.864256,1.0631721,1.1626302,1.1351935,1.039165,1.0151579,1.0254467,1.1351935,1.2277923,1.2689474,1.313532,1.4610043,1.3752645,1.2758065,1.2415106,1.2072148,1.2586586,1.3306799,1.4095604,1.4541451,1.4095604,1.4095604,1.3581166,1.3101025,1.2929544,1.3101025,1.3203912,1.371835,1.3203912,1.1317638,0.864256,0.47328308,0.26407823,0.14404267,0.06859175,0.024007112,0.020577524,0.024007112,0.034295876,0.058302987,0.11317638,0.15090185,0.2469303,0.39783216,0.5590228,0.6859175,1.0014396,1.1660597,1.2998136,1.3821237,1.2655178,1.1111864,1.0563129,1.0528834,1.0597426,1.0460242,1.0666018,1.0666018,1.0323058,0.97400284,0.922559,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.12003556,0.044584636,0.010288762,0.010288762,0.01371835,0.01371835,0.0,0.0,0.010288762,0.020577524,0.037725464,0.061732575,0.072021335,0.14061308,0.24350071,0.3841138,0.5796003,0.70306545,0.66876954,0.6207553,0.5453044,0.29151493,0.29151493,0.51100856,0.6927767,0.7339317,0.6859175,1.1866373,1.7696671,2.318401,2.668219,2.5927682,3.3369887,3.6147852,2.9460156,1.7833855,1.5261664,1.0254467,0.6893471,0.5555932,0.6379033,0.9294182,2.369845,2.8499873,3.192946,4.0949273,6.135532,8.906639,10.981539,12.432255,13.409687,14.1299,23.101702,29.59391,39.74892,61.811455,106.10801,165.47073,147.33508,101.697556,60.01092,35.170418,25.883097,25.93797,29.573332,30.982893,24.3535,16.249386,12.089295,10.347065,9.6645775,8.834618,7.857185,7.4765005,7.39762,7.140401,6.042933,5.127233,4.2835546,4.0229063,4.413879,5.096367,5.267846,4.8905916,4.1326528,3.3747141,3.2032347,2.9974594,2.8705647,2.644212,2.2600982,1.786815,1.529596,1.4095604,1.2758065,1.1008976,0.9911508,1.2620882,1.2277923,1.0323058,0.8162418,0.71678376,0.7888051,0.7442205,0.72707254,0.7613684,0.7613684,0.72707254,0.65162164,0.5178677,0.36696586,0.30523327,0.26750782,0.16804978,0.13032432,0.20234565,0.33609957,0.5796003,0.84367853,0.89169276,0.7305021,0.59674823,0.70649505,0.9534253,1.2209331,1.3478279,1.1283343,1.4095604,2.4418662,3.117495,3.7725463,6.1629686,9.458802,11.8869505,12.106443,10.381361,8.577398,7.6959944,8.40249,9.877212,11.718901,13.917266,14.112752,13.876111,12.199042,10.768905,13.992717,18.54378,17.899017,15.597764,14.956431,19.058218,18.351723,20.61868,25.159454,28.211786,22.9508,21.873909,21.013083,22.11055,25.430391,29.737953,29.189219,26.545008,24.871368,24.52498,23.132568,22.974806,20.817596,18.067066,16.849564,20.03565,20.584383,19.95334,18.152807,16.904436,19.637817,19.980776,19.095943,18.739265,18.886738,17.71382,17.37429,16.417435,15.172495,14.918706,17.899017,16.482597,14.939283,13.588025,12.55915,11.763485,10.079557,8.258447,7.0135064,7.3084507,10.360784,14.033872,11.657167,10.010965,10.772334,10.528833,6.6705475,5.394741,5.658819,6.475061,6.927767,6.989499,6.776865,6.2692857,6.1492505,7.798882,12.034423,16.506605,17.820137,17.058767,19.805868,15.789821,13.056439,14.977009,18.396307,13.612033,8.752307,7.1712675,7.3118806,7.747438,7.1849856,8.711152,8.354475,8.47451,10.816919,16.479168,17.051908,14.706071,12.185325,11.341646,13.121602,12.987847,11.7086115,9.846346,8.471081,9.156999,8.985519,7.130112,5.425607,5.2472687,7.4936485,8.076678,16.839275,26.689049,29.669361,16.935303,8.100685,16.702091,20.680412,16.311117,18.20425,14.664916,13.38568,13.780083,14.033872,11.094715,16.050468,17.545769,17.069057,15.587475,13.5503,9.764035,11.228469,11.465111,10.494537,14.815818,25.814505,26.328943,21.013083,16.321407,20.508932,17.370861,11.698323,9.078118,9.702303,8.347616,5.90575,14.568888,17.182234,11.502836,10.209882,12.771784,16.242527,17.003895,15.0078745,13.762935,15.412566,18.879879,22.87192,23.1943,12.758065,13.660047,11.900668,11.050131,11.55428,10.710602,16.657507,16.239098,11.753197,11.22161,28.396984,19.87446,13.745787,12.504276,14.428274,13.5503,16.722668,20.052797,19.229696,13.985858,8.100685,40.524006,39.91354,27.069735,13.9138365,3.4638834,20.11453,13.684054,4.6573796,1.937717,2.8534167,3.7691166,3.9063,5.48734,7.1678376,4.0434837,2.5653315,2.6545007,3.234101,3.5873485,3.357566,11.718901,21.554956,22.573545,14.534592,7.2467184,9.630281,12.274493,12.493987,11.080997,12.315649,13.008426,13.018714,12.157887,10.319629,7.4627824,7.840037,8.484799,7.7440085,5.360445,2.4418662,1.7079345,1.3889829,1.2175035,1.2346514,1.7696671,2.5893385,4.7602673,6.341307,7.4627824,10.329918,13.114742,8.519095,5.0620713,5.353586,6.0737996,4.6436615,4.588788,4.033195,3.2683969,4.746549,8.090397,7.9909387,7.2604365,6.8557453,5.90575,3.1586502,3.5599117,3.940596,3.0420442,1.5398848,4.2389703,6.094377,5.970912,6.2864337,13.001566,11.180455,6.0395036,5.720552,9.668007,8.604835,2.6613598,1.155771,1.2895249,1.4644338,1.2826657,0.548734,0.39440256,0.37039545,0.26750782,0.12346515,0.08573969,0.11317638,0.106317215,0.06859175,0.09259886,0.16462019,0.20234565,0.17833854,0.116605975,0.09259886,0.17833854,0.18176813,0.12003556,0.048014224,0.061732575,0.15776102,0.34638834,0.41498008,0.8025235,2.609916,1.2175035,0.5144381,1.762808,4.1600895,4.804852,3.0969174,1.196926,0.15090185,0.048014224,0.0,0.0,0.017147938,0.030866288,0.061732575,0.18176813,0.5007198,0.34295875,0.29837412,0.4938606,0.5796003,0.2503599,0.2777966,0.42526886,0.4355576,0.044584636,0.26407823,0.31209245,0.22635277,0.39440256,1.5398848,1.4061309,0.8779744,0.8848336,1.4575747,1.7388009,1.8485477,2.335549,2.469303,2.1297739,1.8005334,1.371835,0.7613684,0.36010668,0.33952916,0.65505123,0.53501564,0.29151493,0.116605975,0.08916927,0.19891608,0.18519773,0.3566771,0.5144381,0.48014224,0.07545093,0.06516216,0.05144381,0.041155048,0.08573969,0.30523327,0.51100856,0.84024894,0.764798,0.40126175,0.48700142,0.7339317,0.5555932,0.29151493,0.12346515,0.07545093,0.041155048,0.07545093,0.082310095,0.041155048,0.01371835,0.0274367,0.030866288,0.041155048,0.06516216,0.07545093,0.15090185,0.24007112,0.22292319,0.12003556,0.106317215,0.15433143,0.21263443,0.25721905,0.25721905,0.18176813,0.18176813,0.16462019,0.15776102,0.16804978,0.16804978,0.13032432,0.11317638,0.216064,0.4046913,0.5041494,0.7476501,0.94656616,1.1489118,1.3101025,1.2963841,1.5776103,1.6393428,1.4747226,1.1729189,0.91569984,0.85396725,0.7922347,0.70649505,0.61046654,0.548734,0.4389872,0.5041494,0.66876954,0.82996017,0.85396725,0.9774324,1.0357354,1.0460242,1.0666018,1.1763484,1.1146159,1.097468,1.1043272,1.1214751,1.1592005,1.6599203,2.16064,2.294394,2.0920484,1.9685832,1.8588364,1.8416885,1.9754424,1.9823016,1.2517995,0.7373613,0.9568549,1.704505,2.503599,2.6236343,1.0014396,0.5693115,0.58645946,0.70649505,0.9602845,0.9842916,1.0014396,1.1592005,1.3649758,1.2655178,1.1077567,1.1043272,1.196926,1.2860953,1.2346514,1.0288762,0.6927767,0.45613512,0.37725464,0.36696586,0.30523327,0.30866286,0.33266997,0.36696586,0.42869842,0.4629943,0.45613512,0.4664239,0.4938606,0.45613512,0.45613512,0.5041494,0.53501564,0.53501564,0.53501564,0.58302987,0.6790583,0.77508676,0.84367853,0.8711152,0.84367853,1.0220171,1.155771,1.1489118,1.039165,1.196926,1.2346514,1.1214751,0.9294182,0.8711152,0.83338976,0.6859175,0.6001778,0.59674823,0.53501564,0.48357183,0.5178677,0.5555932,0.6310441,0.89855194,1.1214751,1.2037852,1.1180456,0.9568549,0.9294182,0.980862,1.0460242,1.0906088,1.1283343,1.2517995,1.313532,1.2620882,1.2037852,1.1489118,1.039165,1.1351935,1.1420527,1.1180456,1.1420527,1.313532,1.4575747,1.5330256,1.5570327,1.4918705,1.2346514,1.0906088,1.0082988,0.9328478,0.8745448,0.89855194,0.75450927,0.59674823,0.42183927,0.24350071,0.12346515,0.061732575,0.0274367,0.0274367,0.05144381,0.07545093,0.11317638,0.16804978,0.22292319,0.26064864,0.26064864,0.41840968,0.59674823,0.7476501,0.9259886,1.2655178,1.2175035,1.2037852,1.1626302,1.0940384,1.0837497,1.2312219,1.1763484,1.1008976,1.0940384,1.1283343,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.010288762,0.0034295875,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0548734,0.24350071,0.09945804,0.11317638,0.15776102,0.18862732,0.23664154,0.29151493,0.38754338,0.5007198,0.5624523,0.45956472,0.39097297,0.45613512,0.4938606,0.48014224,0.52815646,1.1351935,1.5193073,1.7593783,1.8828435,1.8485477,2.8568463,2.784825,2.0680413,1.2792361,1.1111864,0.6893471,0.45270553,0.3566771,0.38754338,0.5658819,2.3081124,3.4707425,3.6559403,3.4055803,4.2046742,7.0546613,9.163857,11.543991,13.690913,13.591455,19.967058,26.949697,38.74062,64.75404,119.644585,177.38855,161.53357,111.053474,59.51706,35.08468,31.401302,31.336142,29.789396,24.339783,15.271953,11.101575,8.848335,7.805741,7.466212,7.517656,7.174697,6.461343,5.672538,4.8837323,3.9303071,3.806842,4.245829,4.7534084,5.099797,5.3158607,4.880303,4.616225,4.273266,3.7451096,3.0454736,2.4487255,2.2258022,2.0920484,1.8931323,1.6016173,1.5021594,1.5158776,1.4610043,1.3478279,1.3958421,1.214074,0.97400284,0.7682276,0.64819205,0.6207553,0.6824879,0.6790583,0.66876954,0.66191036,0.6036074,0.4698535,0.42526886,0.39097297,0.32581082,0.20920484,0.1920569,0.20577525,0.22978236,0.31209245,0.5555932,0.88826317,0.9362774,0.84367853,0.7682276,0.88826317,1.1832076,1.4267083,1.4747226,1.3443983,1.2037852,2.1263442,4.3521466,6.9346256,9.4862385,12.181894,11.688034,10.882081,10.484249,10.628291,10.882081,10.014396,8.954653,8.930646,10.768905,14.928994,16.80498,15.532601,13.258785,11.996697,13.639469,15.038741,15.367981,16.760393,19.28457,20.927343,19.630959,20.896477,21.602972,20.12139,16.283682,17.182234,18.087645,20.049368,22.786179,24.672453,21.548098,19.473198,18.660385,18.87645,19.44576,19.737276,18.015623,16.180794,15.0078745,14.150477,18.02934,22.055677,24.041409,22.745024,17.844143,16.39,16.341984,15.834405,14.860402,15.29939,17.662374,18.115082,16.516893,14.640909,16.153357,15.165636,12.243628,11.540562,12.874671,11.739478,8.618553,9.582268,9.97324,9.2153015,10.813489,11.314209,9.489669,8.961512,9.73317,8.210432,6.228131,6.540223,7.1095347,6.8728933,5.7308407,7.8126,9.136421,10.779194,12.8197975,14.339106,14.805529,14.918706,13.63261,11.567999,11.005547,11.80464,10.089847,8.618553,8.423067,8.81404,8.056101,7.0615206,6.893471,8.515666,12.778643,14.479718,15.391989,15.505165,14.428274,11.4033785,14.239647,15.8138275,15.271953,13.512574,13.197053,14.819247,16.163645,14.267084,10.1652975,8.886061,8.961512,7.9257765,7.0786686,7.407909,9.616563,14.517444,22.909645,33.188118,38.65831,27.51901,14.953001,19.414894,25.135447,25.924252,25.149164,18.221397,14.778092,16.935303,21.02337,17.573206,18.694681,15.752095,12.706621,11.681175,12.9638405,10.556271,11.204462,11.996697,11.331357,8.934075,15.54632,20.855322,17.813278,11.070708,16.955881,14.315098,8.525954,5.9160385,7.1987042,7.455923,4.9934793,12.298501,15.090185,10.707172,8.097256,10.367643,12.21962,12.459691,11.482259,11.273054,10.882081,10.998687,13.663476,16.156786,11.022695,7.805741,6.495639,8.522525,11.828648,10.858074,14.352823,16.486027,15.611482,16.088194,28.26323,19.565796,12.761495,18.530062,30.231813,23.924803,20.652975,22.659285,24.710178,23.400076,17.147938,37.022396,32.9892,19.61038,9.383351,12.740917,41.765514,24.329493,5.90575,2.9940298,3.0969174,4.5990767,4.033195,4.4721823,5.6142344,3.7862647,3.8034124,5.079219,5.07236,4.5442033,7.5553813,21.825895,30.478745,26.253492,12.850664,4.928317,8.052671,10.113853,9.942374,8.388771,8.323608,9.527394,10.278474,9.846346,8.131552,5.65539,5.312431,6.1492505,6.210983,4.866585,2.819121,2.5378947,2.0440342,1.587899,1.3238207,1.2929544,2.3767042,4.7088237,5.8543057,6.4064693,9.9869585,11.7257595,8.532814,5.9743414,5.9743414,6.7802944,6.8866115,5.8371577,4.1155047,2.603057,2.585909,5.353586,6.680836,6.8214493,6.018926,4.5030484,2.428148,3.7485392,4.945465,4.3109913,1.9308578,3.0283258,4.372724,4.6608095,4.2389703,5.103226,6.427047,5.288424,5.4941993,7.5450926,8.64256,4.698535,3.1037767,3.1277838,3.2992632,1.3786942,0.6379033,0.64133286,0.58302987,0.2709374,0.13375391,0.106317215,0.06516216,0.106317215,0.20234565,0.18862732,0.2709374,0.26750782,0.18519773,0.08573969,0.07888051,0.08573969,0.14404267,0.12689474,0.05144381,0.072021335,0.15090185,0.432128,0.6310441,0.8025235,1.3409687,1.4815818,0.88826317,0.66533995,1.2312219,2.3149714,1.7113642,0.9294182,0.33266997,0.06516216,0.037725464,0.0274367,0.0274367,0.030866288,0.06516216,0.20920484,0.41840968,0.23321195,0.18519773,0.39097297,0.5555932,0.16804978,0.17147937,0.22978236,0.17833854,0.020577524,0.5727411,0.548734,0.3018037,0.19891608,0.61389613,0.84024894,1.0048691,1.6976458,2.5070283,1.99602,1.9994495,2.294394,2.1091962,1.4232788,0.9945804,1.1832076,1.0048691,0.6756287,0.4389872,0.5693115,0.39097297,0.1920569,0.14747226,0.31895164,0.6756287,0.2503599,0.14404267,0.16804978,0.17490897,0.07545093,0.044584636,0.0274367,0.020577524,0.048014224,0.15776102,0.36696586,0.7373613,0.7956643,0.5041494,0.25721905,0.33609957,0.23321195,0.14061308,0.14061308,0.20920484,0.13375391,0.082310095,0.05144381,0.048014224,0.05144381,0.034295876,0.030866288,0.041155048,0.07545093,0.12346515,0.17833854,0.25721905,0.28808534,0.25378948,0.1920569,0.20234565,0.22978236,0.2709374,0.28465575,0.18176813,0.17490897,0.15090185,0.15090185,0.16804978,0.16804978,0.14061308,0.16804978,0.25378948,0.38754338,0.5658819,0.8196714,1.0185875,1.2003556,1.4061309,1.6873571,1.7353712,1.5398848,1.2998136,1.0631721,0.72021335,0.66876954,0.66191036,0.6310441,0.5761707,0.5727411,0.5624523,0.5624523,0.61046654,0.71678376,0.8676856,0.939707,0.91227025,0.8711152,0.881404,0.9911508,1.0666018,1.0425946,1.0323058,1.1214751,1.3443983,1.7353712,2.1297739,2.2635276,2.1503513,2.0646117,1.7696671,1.6770682,1.7730967,1.7593783,1.0563129,0.6001778,0.50757897,0.77851635,1.5536032,3.100347,2.6785078,1.3581166,0.58988905,0.6790583,0.7888051,0.8162418,0.8162418,1.0185875,1.3032433,1.2037852,1.0460242,1.08032,1.1317638,1.1111864,1.0048691,0.9431366,0.7613684,0.58988905,0.490431,0.4389872,0.4081209,0.4389872,0.4972902,0.53158605,0.47671264,0.3841138,0.34638834,0.33609957,0.32238123,0.22635277,0.17833854,0.19548649,0.23664154,0.26407823,0.26407823,0.432128,0.6344737,0.77165717,0.83681935,0.91912943,1.0597426,1.08032,1.097468,1.1832076,1.3546871,1.2415106,1.2483698,1.2723769,1.2243627,1.0151579,0.84367853,0.7339317,0.66876954,0.6276145,0.607037,0.5693115,0.5453044,0.5693115,0.65505123,0.8162418,0.89855194,0.99801,0.96714365,0.83681935,0.8196714,0.8711152,0.91569984,0.90884066,0.90884066,1.08032,0.9945804,0.922559,0.91227025,0.9534253,1.0014396,1.3443983,1.5193073,1.4507155,1.255229,1.2380811,1.3272504,1.3855534,1.3512574,1.2346514,1.1146159,1.0563129,1.0254467,0.97400284,0.90884066,0.8745448,0.8471081,0.8093826,0.7888051,0.72364295,0.4629943,0.29494452,0.1920569,0.12346515,0.082310095,0.08916927,0.12346515,0.18862732,0.2469303,0.2709374,0.22292319,0.216064,0.29151493,0.42526886,0.6207553,0.91227025,1.0768905,1.1111864,1.1420527,1.1660597,1.0460242,1.0460242,1.0494537,1.0940384,1.1592005,1.1660597,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.030866288,0.116605975,0.041155048,0.0548734,0.12003556,0.18862732,0.17147937,0.3018037,0.4424168,0.48357183,0.4115505,0.31895164,0.32238123,0.34295875,0.34981793,0.36353627,0.4424168,0.8711152,1.196926,1.3821237,1.4232788,1.371835,1.8862731,1.7971039,1.371835,0.91912943,0.7510797,0.4938606,0.33609957,0.26407823,0.28122616,0.42869842,1.9239986,3.5564823,4.064061,3.542764,3.4398763,5.65539,8.2481575,11.766914,14.891269,14.445422,19.301718,27.326952,39.718052,62.9295,108.69734,155.81645,145.08527,101.31687,53.4364,34.470783,33.476204,31.620796,25.468117,16.074476,9.009526,7.6616983,6.701414,6.018926,5.675967,5.9228973,5.785714,5.470192,4.9934793,4.396731,3.7519686,4.108646,4.7088237,5.24041,5.5490727,5.645101,4.9214582,4.5922174,4.540774,4.4550343,3.8377085,2.8568463,2.0131679,1.4953002,1.2929544,1.1729189,1.3512574,1.4164196,1.5981878,1.8073926,1.6599203,1.2072148,0.94999576,0.8676856,0.84024894,0.66876954,0.65505123,0.7579388,0.7510797,0.61389613,0.5555932,0.4046913,0.32924038,0.28122616,0.23321195,0.16462019,0.21263443,0.26750782,0.34638834,0.48700142,0.7476501,0.84367853,0.7579388,0.6962063,0.84024894,1.2998136,1.8897027,1.786815,2.061182,2.836269,3.2992632,5.07236,6.4304767,8.172707,10.353925,12.257345,10.487679,8.985519,8.323608,8.330468,8.090397,7.73029,9.301042,10.1652975,10.6488695,14.04759,16.87014,15.45715,12.878101,11.533703,13.166186,17.233677,20.04251,20.498644,18.903887,16.969599,17.95389,22.769032,24.936531,22.60441,18.554068,22.151705,21.37319,18.972477,16.482597,14.205351,12.061859,9.952662,9.218731,10.244178,12.46312,12.157887,13.488567,14.493437,14.112752,12.195613,12.775213,15.21365,17.892159,18.739265,15.217079,14.490007,15.899568,16.684942,16.513464,17.487467,14.887839,13.694343,11.962401,9.935514,10.048691,11.273054,9.105555,8.196714,9.72288,11.38623,7.31531,8.169277,9.259886,9.445084,11.118723,9.72631,8.388771,8.258447,8.371623,5.6348124,4.420738,5.271276,5.662249,5.288424,6.0737996,10.329918,11.64345,10.991828,9.839486,10.127572,11.173596,12.991278,14.174485,14.198492,13.443983,16.105343,14.836395,11.897239,9.325048,8.913498,7.6514096,7.2878733,7.414768,8.501947,11.9040985,11.547421,12.668896,14.863832,16.616352,15.275383,13.738928,13.070158,12.199042,11.080997,10.669447,11.413667,12.80265,13.7938,13.773223,12.535142,13.629181,12.840376,12.566009,13.817808,16.19794,25.77678,36.586838,48.418915,53.762215,37.81806,28.640486,24.974257,24.27119,24.000254,21.657845,16.798119,17.676094,22.515242,26.335802,20.971928,21.349182,22.2786,19.600092,13.673765,9.383351,8.625413,7.6171136,8.9100685,11.362224,10.134431,11.712041,16.283682,14.953001,10.041832,15.069608,15.87899,9.942374,7.006647,9.129561,10.676306,5.6313825,7.864044,9.650859,8.1212635,5.2609873,7.7440085,8.381912,9.3764925,10.861504,10.926665,6.550512,5.2026844,8.330468,11.952112,6.6705475,3.7931237,15.031882,17.484037,9.211872,9.22902,11.986408,18.348293,19.86417,19.658396,32.467903,24.61415,16.53747,20.495214,32.85545,34.107246,27.395544,23.917942,24.144297,24.308916,16.414005,20.598103,22.991955,17.63494,12.312219,28.534168,49.71873,24.837072,4.5647807,5.2575574,8.954653,7.723431,6.036074,5.5559316,5.90232,4.6676683,5.751418,6.23499,6.3961806,7.6857057,12.706621,22.734735,26.311794,20.272291,8.934075,4.1120753,6.39961,7.332458,6.8111606,5.535354,4.99005,5.9469047,6.509357,6.8145905,6.4133286,4.297273,3.9783216,5.209543,5.2609873,3.7039545,2.428148,3.093488,2.4144297,1.7147937,1.4232788,1.0460242,1.6667795,3.5461934,5.3158607,7.0032177,10.021255,9.822338,6.81802,4.73969,4.822,5.7754254,7.6788464,5.871454,3.542764,2.2326615,1.8348293,4.914599,6.3138704,6.4819202,5.6039457,3.590778,2.0165975,3.2581081,4.8768735,4.911169,1.8656956,2.2806756,4.214963,4.9831905,3.8720043,2.1297739,3.1860867,4.7842746,5.504488,5.0895076,4.431027,2.6236343,2.386993,3.1963756,3.6559403,1.5124481,0.71678376,0.5007198,0.39783216,0.23664154,0.1371835,0.11317638,0.048014224,0.05144381,0.12003556,0.14061308,0.2194936,0.24007112,0.18862732,0.09945804,0.048014224,0.037725464,0.06859175,0.072021335,0.05144381,0.06859175,0.13375391,0.25378948,0.5212973,0.7407909,0.42869842,1.1214751,1.471293,1.3615463,1.1592005,1.7113642,1.3615463,0.96714365,0.48700142,0.06516216,0.0274367,0.024007112,0.020577524,0.037725464,0.23321195,0.9362774,0.39440256,0.16462019,0.28465575,0.5212973,0.36696586,0.10288762,0.17490897,0.2469303,0.17833854,0.041155048,0.7133542,0.805953,0.71678376,0.7476501,1.0940384,0.8128122,1.2449403,2.153781,2.6716487,1.3272504,1.6633499,1.8382589,1.5638919,1.0185875,0.84024894,0.9259886,0.805953,0.5590228,0.36353627,0.53158605,0.44584638,0.28122616,0.25378948,0.4046913,0.6001778,0.28808534,0.1097468,0.106317215,0.2469303,0.4424168,0.28122616,0.106317215,0.020577524,0.058302987,0.18519773,0.38754338,0.45270553,0.45270553,0.37725464,0.13375391,0.17833854,0.2469303,0.216064,0.12689474,0.18862732,0.16804978,0.08916927,0.037725464,0.041155048,0.05144381,0.041155048,0.034295876,0.041155048,0.06859175,0.09945804,0.17147937,0.2194936,0.2709374,0.30866286,0.28808534,0.24350071,0.24007112,0.25721905,0.26407823,0.22978236,0.28122616,0.28465575,0.20920484,0.1097468,0.10288762,0.1371835,0.30866286,0.48014224,0.6207553,0.8093826,1.0425946,1.1454822,1.1797781,1.2380811,1.4369972,1.4541451,1.3684053,1.255229,1.1077567,0.83681935,0.66876954,0.6207553,0.607037,0.6207553,0.69963586,0.78537554,0.64476246,0.5727411,0.64133286,0.72364295,0.7099246,0.67219913,0.6344737,0.6276145,0.6790583,0.85739684,0.8779744,0.8471081,0.90541106,1.2243627,1.4953002,1.920569,2.1057668,1.9925903,1.8519772,1.9068506,2.0028791,1.937717,1.6016173,0.980862,0.607037,0.53501564,0.58302987,0.805953,1.5158776,1.6084765,1.7353712,1.430138,0.8676856,0.8676856,0.84024894,0.82996017,0.99801,1.2415106,1.1797781,1.1043272,1.0768905,1.0666018,1.0254467,0.90884066,1.0151579,0.85739684,0.66876954,0.5418748,0.42869842,0.42183927,0.5418748,0.59331864,0.52815646,0.45270553,0.48357183,0.4629943,0.432128,0.3841138,0.26750782,0.19891608,0.15433143,0.14747226,0.16462019,0.17147937,0.26407823,0.4424168,0.64133286,0.805953,0.90198153,1.1523414,1.1729189,1.1317638,1.1420527,1.2620882,1.0906088,1.1283343,1.2312219,1.2723769,1.1523414,1.1454822,1.039165,0.881404,0.7133542,0.607037,0.5178677,0.5796003,0.66876954,0.7305021,0.78537554,0.89169276,0.91569984,0.84367853,0.77508676,0.939707,1.0323058,1.0288762,0.9328478,0.8676856,1.0734608,0.89512235,0.8196714,0.881404,0.9945804,0.96371406,1.0666018,1.1934965,1.2243627,1.1249046,0.94656616,0.9328478,1.0357354,1.1317638,1.1660597,1.138623,1.3958421,1.488441,1.3752645,1.1934965,1.255229,1.1283343,0.97400284,0.84367853,0.75450927,0.6962063,0.5796003,0.45270553,0.31552204,0.19548649,0.1371835,0.15090185,0.22292319,0.31895164,0.39097297,0.34981793,0.274367,0.2469303,0.2777966,0.37039545,0.5041494,0.66533995,0.8128122,0.94656616,1.0460242,1.0460242,1.1043272,1.214074,1.3512574,1.488441,1.5673214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.01371835,0.07545093,0.14747226,0.13375391,0.29151493,0.39097297,0.36353627,0.25378948,0.20920484,0.26064864,0.26064864,0.2503599,0.26064864,0.3018037,0.6036074,0.91912943,1.0666018,1.0151579,0.88826317,1.1111864,1.1077567,0.90884066,0.6344737,0.50757897,0.37725464,0.26407823,0.19891608,0.21263443,0.32924038,1.3238207,3.018037,4.0674906,4.0709205,3.5599117,4.7774153,7.6651278,11.770344,15.193072,14.586036,17.806417,27.217207,39.978703,57.798836,86.936615,122.10703,116.907776,85.29727,48.185703,33.383606,32.75942,28.17749,19.52807,10.052121,6.310441,5.936616,5.435896,4.928317,4.57507,4.5613513,4.4241676,4.506478,4.479041,4.32471,4.3178506,4.7945633,5.099797,5.381023,5.576509,5.4016004,4.6608095,4.297273,4.3007026,4.40359,4.064061,3.2478194,2.0749004,1.2037852,0.864256,0.8711152,1.1317638,1.3512574,1.6599203,1.903421,1.6599203,1.2312219,1.1146159,1.0871792,0.96714365,0.6310441,0.70649505,0.7990939,0.72021335,0.53158605,0.5624523,0.4355576,0.34295875,0.26750782,0.21263443,0.18176813,0.31209245,0.51100856,0.77165717,1.0871792,1.4610043,1.5398848,1.7147937,1.8348293,1.9274281,2.1846473,2.5447538,2.7642474,3.3541365,4.431027,5.693115,7.8126,8.48137,8.855195,9.287323,9.349055,7.6445503,6.9380555,7.459353,8.543102,8.625413,8.484799,10.233889,10.906088,10.782623,13.38225,16.808409,16.37285,15.021593,14.373401,14.733508,19.356592,21.181131,20.066517,17.367432,15.920145,18.231688,22.851341,24.19574,22.347193,23.022821,24.319204,21.304598,18.900457,18.36544,17.267973,10.847785,9.674867,8.916927,7.2638664,6.944915,6.9860697,9.253027,11.612583,13.395968,15.422854,11.794352,11.321068,12.109874,13.2690735,14.911846,18.732407,22.511812,26.370098,29.662502,31.000042,17.895588,11.629731,9.585697,9.81205,11.032983,12.905538,12.164746,10.604284,10.192734,13.083877,9.55826,9.194724,10.007536,10.2236,8.292743,7.915488,7.805741,7.548522,7.116394,6.852316,6.8866115,6.1286726,5.861165,6.848886,9.349055,13.320518,15.097044,13.025573,9.105555,8.97866,7.98065,9.088407,11.156448,13.049581,13.642899,18.12537,19.356592,17.95046,14.956431,11.8869505,9.496528,9.637141,9.647429,9.160428,10.117283,10.024684,9.928656,11.499407,14.177915,15.162207,12.421966,10.590566,9.815479,10.113853,11.358793,11.005547,11.653738,13.7938,16.835844,19.109661,23.331484,24.380938,24.84736,25.293207,24.230036,34.556522,45.009907,55.226646,60.84088,53.480988,45.81586,31.061773,20.61525,18.276272,20.234566,21.736725,33.445335,47.033363,51.313488,32.24498,22.847912,24.422092,23.893936,16.575195,6.135532,6.111525,4.8185706,5.9126086,9.108984,10.196163,10.707172,13.88297,12.507706,8.615124,13.450842,15.165636,9.80519,8.772884,12.881531,12.339656,5.5730796,5.7068334,7.6274023,8.22758,6.3893213,7.6925645,7.006647,6.680836,7.3221693,7.795452,3.3609958,2.8396983,7.373613,11.506266,3.1689389,4.7602673,18.03963,18.21111,5.662249,5.926327,9.084977,21.20514,23.969387,18.886738,27.306376,24.600431,19.102802,19.816156,26.754211,30.955456,27.573883,23.60242,21.1194,19.36688,14.754086,12.336226,15.9921665,14.579176,11.828648,26.35295,36.075832,19.027351,6.992929,9.880642,15.71094,10.652299,6.8043017,5.7479887,6.56766,5.844017,5.754848,5.761707,6.8969,9.770895,14.582606,18.269413,18.02934,12.9809885,5.9983487,3.7211025,4.722542,4.7602673,4.290414,3.6936657,3.275256,3.5976372,4.1120753,4.8322887,5.0174866,3.1792276,3.1860867,4.341858,4.190956,2.6990852,2.2326615,2.8019729,2.3629858,1.7456601,1.313532,0.9842916,1.4438564,2.6133456,4.256118,6.4407654,9.534253,8.086967,5.1066556,3.4433057,3.865145,5.020916,6.944915,5.6073756,3.350707,1.8588364,2.1572106,5.096367,6.3207297,5.802862,4.1326528,2.5173173,1.587899,3.0317552,4.605936,4.6402316,2.0474637,2.2600982,4.4927597,4.9214582,3.0386145,1.6599203,3.0283258,5.4736214,6.0086374,4.1943855,2.1297739,2.054323,2.0714707,2.4658735,2.6819375,1.2929544,0.71678376,0.39783216,0.24350071,0.17490897,0.12346515,0.09602845,0.05144381,0.048014224,0.07888051,0.072021335,0.13032432,0.18862732,0.22292319,0.1920569,0.048014224,0.020577524,0.0274367,0.034295876,0.034295876,0.061732575,0.12689474,0.09945804,0.31552204,0.5796003,0.17833854,0.6344737,2.7162333,3.5702004,2.6236343,1.5536032,1.1146159,0.7613684,0.39783216,0.08573969,0.05144381,0.030866288,0.020577524,0.07545093,0.33952916,1.0220171,0.32238123,0.14747226,0.31895164,0.4972902,0.15090185,0.07888051,0.66191036,0.7579388,0.2503599,0.041155048,0.53844523,0.7339317,0.77851635,0.9328478,1.5638919,1.0871792,1.1900668,1.7147937,2.0063086,0.89512235,1.1214751,1.3101025,1.1660597,0.83681935,0.9294182,0.7579388,0.6241849,0.42869842,0.26750782,0.40126175,0.41498008,0.28122616,0.25378948,0.37382504,0.4972902,0.47671264,0.35324752,0.26750782,0.31895164,0.5761707,0.35324752,0.14061308,0.05144381,0.13032432,0.37382504,0.6344737,0.59674823,0.6310441,0.6962063,0.36696586,0.23321195,0.3018037,0.26750782,0.116605975,0.1097468,0.13375391,0.08573969,0.058302987,0.06516216,0.041155048,0.041155048,0.034295876,0.034295876,0.044584636,0.058302987,0.11317638,0.16804978,0.22978236,0.29151493,0.30523327,0.28122616,0.26750782,0.2777966,0.29494452,0.2709374,0.29151493,0.28465575,0.1920569,0.061732575,0.0548734,0.18176813,0.3806842,0.59674823,0.78537554,0.9294182,1.1008976,1.1489118,1.0837497,0.9877212,1.0288762,1.1763484,1.138623,1.0666018,1.0082988,0.8848336,0.77165717,0.6893471,0.6859175,0.7510797,0.78537554,0.89855194,0.69963586,0.5453044,0.5453044,0.5590228,0.5007198,0.4664239,0.45956472,0.47671264,0.4972902,0.66876954,0.72707254,0.6824879,0.65848076,0.8745448,1.0837497,1.4953002,1.8245405,1.9342873,1.8416885,2.2360911,2.417859,2.201795,1.6530612,1.0666018,0.6276145,0.6310441,0.6790583,0.61046654,0.490431,0.6310441,1.4472859,1.5433143,0.89512235,0.84367853,0.8162418,0.8779744,1.08032,1.3169615,1.3272504,1.2312219,1.1454822,1.1043272,1.0837497,1.0185875,1.1214751,0.97400284,0.8265306,0.7339317,0.58988905,0.52472687,0.6001778,0.59331864,0.48014224,0.42869842,0.65505123,0.7099246,0.6790583,0.58302987,0.40126175,0.33952916,0.23664154,0.16804978,0.15090185,0.16462019,0.16119061,0.25378948,0.42183927,0.6310441,0.8128122,1.0700313,1.1694894,1.2072148,1.2312219,1.2483698,1.0357354,1.0563129,1.1694894,1.2723769,1.3169615,1.3581166,1.2586586,1.0563129,0.8265306,0.6790583,0.6207553,0.69963586,0.764798,0.7682276,0.77165717,0.84024894,0.8162418,0.77851635,0.8093826,0.9842916,1.0151579,0.9602845,0.8505377,0.7956643,0.9774324,0.82996017,0.78537554,0.84367853,0.90884066,0.7922347,0.77851635,0.90541106,1.0048691,0.97057325,0.7613684,0.78194594,0.88826317,1.0117283,1.1180456,1.2243627,1.5810398,1.7388009,1.7456601,1.6804979,1.6393428,1.3341095,1.1729189,0.9945804,0.8128122,0.823101,0.75450927,0.64819205,0.548734,0.45613512,0.34638834,0.31209245,0.30523327,0.34981793,0.41498008,0.42869842,0.4046913,0.3566771,0.30523327,0.2777966,0.29494452,0.34638834,0.48357183,0.6379033,0.764798,0.881404,1.0837497,1.1900668,1.2998136,1.4644338,1.6736387,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.05144381,0.13375391,0.15776102,0.15090185,0.15433143,0.20920484,0.22978236,0.20577525,0.17147937,0.14061308,0.12003556,0.4424168,0.72364295,0.77851635,0.6276145,0.50757897,0.7510797,0.78194594,0.6344737,0.42526886,0.35324752,0.2777966,0.18519773,0.12689474,0.14061308,0.2194936,0.7407909,2.177788,3.6970954,4.5167665,3.923448,4.280125,7.034084,10.933525,13.978998,13.413116,15.011304,24.741043,37.211025,50.181725,64.5517,91.0967,89.87577,69.86755,44.433735,31.291555,29.542467,22.36091,13.72178,7.181556,5.861165,5.0620713,4.506478,4.1772375,3.9440255,3.5599117,3.450165,3.6627994,3.8960114,4.245829,5.209543,5.4633327,5.2815647,5.1752477,5.0895076,4.40359,3.8342788,3.542764,3.4433057,3.415869,3.3026927,2.959734,1.9925903,1.1214751,0.7133542,0.77508676,0.96714365,1.3992717,1.6667795,1.6359133,1.4335675,1.2037852,1.2346514,1.1626302,0.8745448,0.4972902,0.77165717,0.7510797,0.5693115,0.41498008,0.5418748,0.4629943,0.40126175,0.33952916,0.29837412,0.32238123,0.6927767,1.2449403,1.821111,2.3835633,2.9906003,3.4021509,4.15666,4.8117113,5.271276,5.7891436,5.051782,5.0449233,5.3878818,6.2692857,8.460793,10.268185,11.026124,10.55284,9.122703,7.425057,6.334448,6.708273,8.838047,11.790922,13.38911,12.648318,10.964391,10.432805,11.808069,14.479718,17.261114,17.247395,17.226818,17.521763,15.999025,18.019053,16.835844,16.029892,16.79469,17.936743,18.416885,18.907316,16.96274,15.827546,24.45296,21.699,19.661825,24.10314,32.210686,32.608517,16.427725,16.242527,15.755525,9.9869585,5.271276,6.358455,7.0203657,9.493098,14.96329,23.571554,14.349394,11.640019,10.336777,10.172156,15.717799,23.955667,29.473875,36.01753,43.14764,46.244556,25.896814,15.834405,14.5243025,18.28656,21.273731,21.006224,20.330595,18.084215,15.440002,15.920145,13.673765,12.233338,12.123591,10.978109,3.5461934,7.4010496,9.39021,8.333898,6.835168,11.283342,12.30536,8.97866,8.412778,11.461681,12.710052,14.225929,16.798119,16.016174,12.881531,13.828096,12.233338,10.333347,10.086417,11.657167,13.419975,16.023033,18.924463,19.853882,17.806417,13.063298,10.854645,11.118723,10.690024,9.136421,8.786603,11.163307,10.326488,9.506817,9.647429,9.3936405,9.719451,9.938945,10.22703,11.369082,14.784951,15.824117,16.441442,17.333136,20.128248,27.381826,38.57943,45.116222,46.083366,41.021297,29.919722,35.66428,42.91786,49.266026,55.257515,64.400795,53.889107,31.696247,16.37971,14.96672,22.919933,33.76429,56.577904,79.72419,86.09637,53.158607,25.495554,20.515793,20.687271,16.177364,4.835718,5.0140567,4.413879,5.363875,7.922347,9.853205,11.526843,13.656617,10.738038,6.40304,13.423406,11.976119,7.016936,9.22902,16.167076,12.267634,5.1100855,6.138962,9.225591,10.9369545,10.542552,8.934075,7.267296,4.4721823,1.8931323,3.2683969,4.0091877,4.2698364,8.021805,11.797781,4.698535,9.825768,12.590015,9.496528,3.5221863,4.1189346,8.014946,22.830763,25.663603,15.889278,15.155347,20.800447,19.78186,18.632948,19.363451,19.442331,21.249723,23.681301,20.165974,13.649758,16.61292,14.946142,13.426835,13.495427,14.188204,12.151029,13.876111,12.4802685,12.151029,14.359683,17.87501,10.4705305,5.5250654,5.212973,7.6788464,7.0443726,4.15323,4.314421,6.4579134,9.517105,12.411677,12.055,10.834066,8.110974,4.7328305,3.0386145,3.1312134,2.8911421,2.860276,3.1072063,3.2546785,2.9803114,3.6936657,4.307562,4.0366244,2.3835633,2.633923,3.3266997,3.1620796,2.3664153,2.6716487,2.1469216,2.2978237,2.0474637,1.3341095,1.1180456,1.7525192,2.3835633,2.983741,4.2698364,7.682276,6.375603,3.998899,3.0043187,3.8960114,5.2301207,5.4907694,5.254128,3.4947495,1.5261664,3.000889,5.144381,6.2075534,4.8734436,2.1572106,1.4164196,1.1900668,3.0557625,4.297273,3.8857226,2.469303,2.5584722,4.290414,3.858286,1.6016173,1.9925903,5.3707337,6.914048,6.5710897,4.8322887,2.7573884,3.6285036,2.750529,1.7696671,1.2963841,0.90541106,0.6756287,0.4389872,0.23664154,0.116605975,0.116605975,0.07888051,0.06859175,0.09602845,0.12003556,0.041155048,0.07888051,0.15433143,0.25721905,0.29151493,0.06859175,0.024007112,0.0274367,0.020577524,0.01371835,0.06516216,0.13375391,0.072021335,0.16119061,0.37039545,0.3806842,0.34638834,3.3781435,4.8837323,3.5153272,1.1729189,0.67219913,0.31552204,0.1371835,0.106317215,0.09602845,0.058302987,0.034295876,0.16119061,0.36353627,0.37382504,0.23321195,0.24007112,0.30523327,0.29151493,0.017147938,0.1371835,1.2380811,1.3101025,0.28465575,0.0274367,0.2503599,0.39440256,0.40126175,0.548734,1.430138,1.3546871,0.89512235,0.8093826,1.1043272,1.039165,0.764798,0.9328478,0.96714365,0.823101,1.0014396,0.70306545,0.58988905,0.44927597,0.26750782,0.23664154,0.25378948,0.15090185,0.13032432,0.26064864,0.48014224,0.66191036,0.66533995,0.4938606,0.29494452,0.33609957,0.18519773,0.10288762,0.09602845,0.2194936,0.5693115,0.88826317,1.0220171,1.1489118,1.1626302,0.66876954,0.41498008,0.31895164,0.23321195,0.116605975,0.05144381,0.09259886,0.09602845,0.116605975,0.12346515,0.030866288,0.030866288,0.030866288,0.024007112,0.017147938,0.030866288,0.041155048,0.116605975,0.1920569,0.22978236,0.24007112,0.28808534,0.2777966,0.29494452,0.33266997,0.26750782,0.17833854,0.13375391,0.08573969,0.041155048,0.048014224,0.25721905,0.39440256,0.5761707,0.77165717,0.823101,0.9568549,1.0323058,0.96714365,0.8093826,0.7442205,0.9774324,0.84367853,0.7339317,0.7682276,0.7922347,0.90198153,0.83681935,0.84367853,0.9294182,0.8711152,0.922559,0.7476501,0.5453044,0.4355576,0.4355576,0.39097297,0.36010668,0.3806842,0.4389872,0.45956472,0.5418748,0.6173257,0.607037,0.52815646,0.52472687,0.6893471,0.9842916,1.4267083,1.8691251,1.9823016,2.4212887,2.5001693,2.2326615,1.7216529,1.1351935,0.61389613,0.6173257,0.7613684,0.805953,0.66876954,0.72364295,0.8676856,0.8745448,0.7476501,0.7133542,0.7373613,0.91227025,1.1866373,1.4404267,1.5158776,1.3649758,1.2620882,1.2243627,1.2312219,1.214074,1.1454822,1.0323058,0.9842916,0.97400284,0.85396725,0.70649505,0.6344737,0.5624523,0.48014224,0.432128,0.7305021,0.8779744,0.90198153,0.805953,0.5693115,0.5007198,0.37382504,0.26407823,0.216064,0.2194936,0.16462019,0.16119061,0.216064,0.3566771,0.6036074,0.8162418,1.0185875,1.1934965,1.3032433,1.3238207,1.0940384,1.0528834,1.1008976,1.2003556,1.3546871,1.2860953,1.2037852,1.0666018,0.90198153,0.8093826,0.83338976,0.84367853,0.805953,0.7339317,0.70649505,0.6824879,0.6790583,0.7510797,0.85739684,0.86082643,0.77508676,0.69963586,0.65162164,0.66533995,0.77165717,0.7510797,0.7476501,0.7305021,0.6790583,0.5796003,0.6756287,0.86082643,0.9431366,0.8779744,0.78537554,0.939707,1.0117283,1.0323058,1.0768905,1.2860953,1.4815818,1.5981878,1.8245405,2.0508933,1.8691251,1.4678634,1.4164196,1.3101025,1.0666018,0.9328478,0.7990939,0.72707254,0.72707254,0.7305021,0.59674823,0.52815646,0.4355576,0.36696586,0.36353627,0.42869842,0.48357183,0.4698535,0.4046913,0.33609957,0.32581082,0.28122616,0.30523327,0.37382504,0.4698535,0.6001778,0.89855194,0.9328478,0.94999576,1.0837497,1.3306799,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.048014224,0.072021335,0.09945804,0.1371835,0.08916927,0.07545093,0.06859175,0.058302987,0.044584636,0.38754338,0.5658819,0.5453044,0.48357183,0.70306545,0.5555932,0.47328308,0.41840968,0.34295875,0.18176813,0.14747226,0.09259886,0.0548734,0.072021335,0.18176813,0.53844523,1.7799559,3.3678548,4.3761535,3.508468,3.8274195,6.166398,9.335337,11.825217,11.825217,13.279363,19.637817,29.477304,40.23592,48.22,71.08163,70.83127,55.96058,37.114994,27.069735,23.736176,15.505165,8.621983,5.4084597,4.273266,3.3198407,3.0454736,3.083199,3.0729103,2.6716487,2.8534167,3.1449318,3.6456516,4.671098,6.759717,6.5642304,5.5833683,4.7088237,4.0606318,2.976882,2.620205,2.4795918,2.369845,2.253239,2.2292318,1.6427724,1.0734608,0.72707254,0.6276145,0.64133286,1.0666018,1.4850113,1.7010754,1.605047,1.1900668,0.97057325,0.8711152,0.8025235,0.6927767,0.47328308,0.71678376,0.70649505,0.52815646,0.34638834,0.3806842,0.3806842,0.39097297,0.3841138,0.432128,0.70306545,1.762808,2.935727,3.8514268,4.5270553,5.3707337,6.2144127,7.366754,9.345626,12.343085,16.249386,13.491997,9.294182,7.829748,10.010965,13.502286,14.723219,15.268523,14.407697,12.600305,11.489118,11.111863,11.465111,12.531713,14.095605,15.731518,13.3033695,9.115844,9.983529,15.553179,18.324286,16.993607,13.3033695,10.604284,9.956093,10.100135,12.202472,13.869251,16.263103,17.88873,14.616901,9.493098,9.884071,9.3593445,9.342196,19.11995,22.78275,29.583622,43.096195,53.738205,38.77149,15.724659,13.1593275,13.365103,9.873782,7.431916,7.795452,8.182996,13.437123,23.791048,34.851467,11.986408,6.7665763,7.425057,8.745448,12.055,15.398848,18.62609,22.806757,28.811964,37.307053,28.444998,25.660173,28.986874,34.371326,33.675117,29.35384,24.802776,22.258022,20.670124,15.700651,12.905538,11.262765,10.323058,8.344186,2.287535,12.579727,16.990177,13.975569,8.827758,13.687484,12.404818,9.009526,10.185875,13.834956,9.047252,9.146709,10.55284,12.109874,13.790371,16.70895,31.099499,32.608517,30.252392,29.031458,29.936869,16.729528,12.010415,10.611144,8.971801,5.127233,4.297273,3.9611735,3.9543142,4.2835546,5.113515,7.3839016,10.422516,12.13731,11.31078,7.599966,7.610255,10.113853,10.786053,10.268185,14.174485,22.11055,24.597002,25.19375,27.652763,35.90435,60.058937,77.66987,77.64586,58.567066,28.68507,26.01342,32.67711,39.00127,41.864975,44.708103,31.027477,17.223389,13.437123,18.766703,21.270302,42.98645,64.7026,82.51244,89.60826,76.27746,35.08125,19.95677,14.033872,9.06097,5.3878818,7.191845,5.2266912,8.285883,15.9921665,18.814716,15.748666,14.352823,10.086417,7.2604365,19.027351,12.80265,5.5147767,7.956643,17.027903,15.745236,7.0546613,5.360445,8.093826,11.605724,11.153018,6.138962,5.2506986,4.0229063,2.4624438,5.051782,12.960411,8.903209,4.2423997,5.861165,16.173935,14.0750265,12.312219,8.656279,5.535354,10.038403,13.996146,19.397747,20.941061,17.974468,14.496866,26.178041,23.201159,19.833303,21.078245,22.690151,17.905876,28.33525,26.7645,14.637479,22.03167,12.768354,12.082437,27.073164,42.81497,22.36777,17.1205,12.538571,11.567999,12.538571,9.170717,3.8377085,3.7005248,7.2707253,10.851214,8.543102,4.297273,3.5564823,5.171818,7.6033955,8.89635,7.5039372,6.1492505,4.763697,3.2958336,1.7079345,1.8176813,1.8999915,2.2978237,3.0969174,4.1360826,3.7794054,4.0846386,4.280125,3.799983,2.2738166,2.3595562,3.0660512,3.2066643,2.9151495,3.6456516,2.6819375,3.1655092,3.2306714,2.386993,1.4953002,1.704505,2.452155,2.5721905,2.3835633,3.6765177,3.690236,2.9700227,3.1723683,4.5339146,5.888602,5.0003386,4.3281393,2.8808534,1.646202,3.5873485,5.2335505,5.562791,4.307562,2.2463799,1.2209331,1.2689474,2.352697,3.40901,3.6147852,2.3972816,2.1160555,2.8945718,2.5721905,1.4198492,2.1503513,7.4627824,7.2775846,6.0703697,5.051782,2.1812177,2.9871707,2.5756202,1.7936742,1.2106444,1.1146159,0.7476501,0.4081209,0.18176813,0.10288762,0.15090185,0.116605975,0.09602845,0.09259886,0.07888051,0.030866288,0.06859175,0.15090185,0.22292319,0.216064,0.044584636,0.010288762,0.0,0.0,0.01371835,0.07545093,0.12346515,0.082310095,0.13032432,0.2709374,0.31895164,0.3806842,0.5144381,0.77165717,0.96371406,0.67219913,0.37725464,0.19548649,0.09259886,0.048014224,0.061732575,0.061732575,0.06859175,0.2777966,0.4972902,0.16804978,0.29151493,0.5658819,0.548734,0.22635277,0.030866288,0.32238123,0.7442205,0.6962063,0.23664154,0.07545093,0.4046913,0.26750782,0.12346515,0.28465575,0.9294182,1.2346514,0.89169276,0.805953,1.1351935,1.2826657,1.0871792,0.7990939,0.7682276,0.9534253,0.91569984,0.64819205,0.53501564,0.51100856,0.4664239,0.26064864,0.16119061,0.072021335,0.037725464,0.08916927,0.26064864,0.34638834,0.51100856,0.5418748,0.36010668,0.030866288,0.0548734,0.061732575,0.10288762,0.22635277,0.45613512,0.64133286,0.8162418,0.764798,0.4972902,0.22978236,0.5693115,0.42869842,0.21263443,0.11317638,0.07545093,0.17490897,0.17833854,0.17490897,0.15090185,0.030866288,0.030866288,0.030866288,0.024007112,0.017147938,0.030866288,0.030866288,0.06859175,0.12346515,0.16804978,0.16804978,0.20577525,0.17833854,0.17833854,0.20920484,0.18176813,0.12346515,0.06859175,0.034295876,0.024007112,0.061732575,0.28122616,0.5007198,0.64133286,0.66533995,0.5796003,0.8471081,0.980862,0.94999576,0.805953,0.67219913,0.5624523,0.45956472,0.4972902,0.65848076,0.7922347,0.9877212,0.9911508,0.99801,1.08032,1.1900668,1.0940384,0.8676856,0.59674823,0.38754338,0.34981793,0.32581082,0.31895164,0.34981793,0.38754338,0.34981793,0.36353627,0.5041494,0.61389613,0.6241849,0.548734,0.548734,0.66876954,0.91227025,1.2620882,1.6633499,1.8108221,1.8005334,1.6221949,1.2826657,0.7922347,0.58645946,0.5796003,0.65162164,0.71678376,0.71678376,0.99801,0.9774324,0.84367853,0.7510797,0.823101,0.83681935,1.0048691,1.1934965,1.3203912,1.3581166,1.430138,1.3409687,1.2792361,1.2758065,1.1900668,0.9945804,0.8711152,0.84367853,0.8676856,0.85396725,0.7579388,0.6962063,0.65162164,0.59331864,0.45613512,0.48357183,0.6344737,0.823101,0.9362774,0.84024894,0.6927767,0.5727411,0.4698535,0.39097297,0.36696586,0.29151493,0.20234565,0.17147937,0.20234565,0.21263443,0.44584638,0.7407909,0.8711152,0.86082643,1.0082988,1.0323058,0.96371406,0.8676856,0.8162418,0.91569984,0.91569984,0.84367853,0.8128122,0.83338976,0.8093826,0.78537554,0.805953,0.78194594,0.67219913,0.48700142,0.548734,0.6276145,0.6962063,0.72707254,0.70306545,0.66533995,0.6379033,0.6241849,0.6379033,0.6859175,0.72364295,0.70649505,0.6756287,0.65162164,0.64133286,0.6790583,0.7339317,0.77508676,0.8093826,0.8711152,1.0151579,1.1454822,1.1866373,1.1763484,1.2346514,1.3341095,1.3752645,1.4850113,1.7113642,2.0303159,1.821111,1.6496316,1.5055889,1.3615463,1.1900668,0.86082643,0.7339317,0.70306545,0.66876954,0.53501564,0.5453044,0.5590228,0.5212973,0.4664239,0.5041494,0.42869842,0.37382504,0.37382504,0.4115505,0.4115505,0.42526886,0.42869842,0.42183927,0.42869842,0.5041494,0.72364295,0.823101,0.89855194,0.9534253,0.91569984,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.030866288,0.106317215,0.17490897,0.12346515,0.06516216,0.05144381,0.044584636,0.044584636,0.06859175,0.26407823,0.44927597,0.5693115,0.59331864,0.53158605,0.5212973,0.40126175,0.32924038,0.3018037,0.13375391,0.08916927,0.06859175,0.06859175,0.116605975,0.25721905,0.66876954,1.6976458,2.9048605,3.6525106,3.1072063,3.4433057,5.919468,8.80718,10.762046,10.847785,12.830087,18.228258,25.320644,34.127827,46.446903,64.89809,62.126976,48.840755,34.655983,28.09518,17.78927,10.415657,6.258997,4.4687524,3.0386145,2.633923,2.5550427,2.5619018,2.4658735,2.1194851,2.3252604,2.8054025,3.4227283,4.184097,5.2472687,5.1580997,4.6402316,4.2389703,3.882293,2.901431,2.2052248,1.6976458,1.3341095,1.1146159,1.08032,0.91569984,0.78194594,0.78537554,0.91227025,1.0323058,1.3992717,1.4953002,1.3786942,1.1729189,1.08032,0.8128122,0.66191036,0.6276145,0.64819205,0.59674823,0.66191036,0.5796003,0.42183927,0.29837412,0.34638834,0.4115505,0.36010668,0.36696586,0.59331864,1.1660597,2.2669573,3.2889743,4.40702,5.785714,7.5553813,9.091836,11.55428,18.008764,28.894274,42.015877,40.517147,28.009441,16.907866,12.555719,13.224489,12.531713,11.619442,9.798331,7.747438,7.534804,11.197603,11.941824,12.315649,13.042721,13.008426,11.293632,9.877212,9.993818,11.516555,12.9809885,12.908967,12.994707,13.982429,15.443433,15.765814,17.034761,15.817257,15.563468,15.80011,12.127021,9.314759,15.481158,15.9750185,11.187314,16.530611,22.350622,33.397324,53.498135,69.08904,49.22144,18.46147,9.445084,9.105555,9.205012,6.3447366,9.338767,19.253704,41.549454,64.44538,58.94432,22.645567,8.549961,7.623973,10.799771,8.992378,13.409687,15.103903,16.05733,18.588364,25.344652,22.470657,20.858751,22.628418,26.42497,27.44013,22.5221,21.338894,20.824455,18.842154,14.188204,8.872343,11.05356,12.867812,10.14129,2.3972816,9.328478,16.345413,15.786391,10.563129,14.150477,13.375391,8.958082,7.73029,10.415657,11.63659,10.991828,13.810948,15.1862135,16.317978,24.507832,52.071426,59.139805,51.88966,38.445675,28.853119,27.302946,30.622786,30.83542,24.487255,12.644889,9.3936405,7.6857057,8.519095,9.47938,4.7328305,6.2727156,7.6788464,9.208443,10.508256,10.6145735,8.525954,10.247607,11.427385,11.756626,14.980438,22.155134,25.93797,28.211786,32.738842,45.167667,77.604706,94.44741,86.346725,57.35985,24.93996,17.638369,20.954779,27.337242,31.027477,28.071173,15.4914465,9.287323,11.008976,19.312008,29.950588,54.86654,65.93039,68.59175,63.728596,47.64383,26.033998,20.61868,17.388008,11.571428,7.6445503,9.73317,7.517656,8.97523,13.999576,14.407697,13.190193,12.706621,11.163307,10.97468,18.746124,12.80608,6.90033,9.770895,19.154245,21.77788,7.363324,5.686256,11.026124,15.031882,6.697984,2.7470996,2.2841053,2.551613,5.703404,18.807858,24.27462,11.869802,2.7951138,4.290414,9.595985,7.8777623,6.5539417,4.6127954,3.1449318,5.353586,7.6685576,10.477389,12.411677,14.016724,17.741257,26.593021,18.677534,15.614912,22.659285,28.695358,14.455711,28.455288,35.50995,25.032558,11.036412,11.214751,14.102464,22.61127,30.430729,22.062536,11.05356,6.036074,8.570539,13.927555,11.074138,5.7308407,10.288762,14.658057,13.701202,7.2158523,4.1189346,3.8205605,4.8014226,5.7239814,5.4187484,3.9268777,3.0523329,2.311542,1.5947582,1.1592005,1.2998136,1.5364552,1.7113642,1.9754424,2.7813954,3.1963756,5.020916,6.807731,7.164408,4.73969,2.5584722,2.503599,3.1106358,3.8617156,5.161529,3.7382503,3.9646032,3.9543142,3.07634,1.9720128,2.452155,3.40901,3.1826572,2.0303159,2.1023371,2.6922262,2.9803114,4.0880685,5.892031,7.0135064,5.3981705,3.433017,2.1194851,2.1812177,4.0606318,6.5196457,6.715132,5.439326,3.4535947,1.488441,1.6359133,2.2909644,3.1895163,3.6387923,2.5070283,1.862266,3.2443898,3.3815732,2.1332035,2.4452958,10.079557,7.723431,4.1155047,2.942586,2.8156912,3.8377085,2.644212,1.6084765,1.3821237,0.89512235,0.607037,0.44927597,0.29151493,0.14061308,0.14061308,0.11317638,0.12003556,0.10288762,0.06859175,0.06859175,0.044584636,0.07545093,0.13375391,0.16804978,0.09602845,0.0274367,0.0034295875,0.0,0.006859175,0.041155048,0.14747226,0.08916927,0.12003556,0.23664154,0.18519773,0.6962063,0.86082643,0.8128122,0.7510797,0.96371406,0.4938606,0.19548649,0.058302987,0.037725464,0.061732575,0.05144381,0.07888051,0.1371835,0.19548649,0.216064,1.0323058,0.9911508,0.5453044,0.10288762,0.041155048,0.2469303,1.1592005,1.4232788,0.84024894,0.37039545,0.97057325,0.6310441,0.25721905,0.18862732,0.20920484,1.0528834,0.83338976,0.91912943,1.6016173,2.0989075,1.3855534,0.8745448,0.78194594,0.97057325,0.96371406,0.51100856,0.44584638,0.48014224,0.4389872,0.26064864,0.14061308,0.06516216,0.0548734,0.10288762,0.1371835,0.14404267,0.24007112,0.32924038,0.37382504,0.3841138,0.23321195,0.14404267,0.09259886,0.08573969,0.15090185,0.22978236,0.41840968,0.47671264,0.38754338,0.36353627,0.7339317,0.71678376,0.45613512,0.16804978,0.09945804,0.1097468,0.12346515,0.11317638,0.08573969,0.07888051,0.06859175,0.037725464,0.017147938,0.01371835,0.006859175,0.017147938,0.034295876,0.06859175,0.11317638,0.13032432,0.08916927,0.116605975,0.116605975,0.082310095,0.09602845,0.0548734,0.037725464,0.0274367,0.0274367,0.072021335,0.18519773,0.26750782,0.31552204,0.34638834,0.39783216,0.548734,0.66533995,0.6241849,0.45270553,0.31895164,0.31552204,0.29837412,0.40126175,0.64133286,0.939707,1.039165,1.0666018,1.0631721,1.0837497,1.214074,0.97057325,0.7373613,0.51100856,0.33266997,0.26407823,0.32924038,0.3806842,0.39097297,0.38754338,0.44927597,0.4115505,0.39440256,0.4115505,0.45956472,0.51100856,0.53158605,0.64133286,0.72364295,0.8093826,1.0666018,1.3581166,1.2826657,0.9945804,0.6927767,0.6344737,0.58302987,0.5418748,0.5761707,0.7099246,0.9259886,1.097468,1.1008976,1.097468,1.1249046,1.08032,1.0151579,1.0323058,1.2037852,1.4850113,1.6873571,1.605047,1.605047,1.587899,1.4918705,1.2895249,1.0425946,0.89512235,0.78537554,0.7339317,0.82996017,0.82996017,0.84367853,0.84024894,0.7888051,0.66533995,0.5727411,0.5796003,0.6893471,0.83681935,0.8745448,0.8162418,0.7990939,0.71678376,0.59674823,0.61046654,0.52815646,0.3806842,0.31895164,0.36353627,0.432128,0.53844523,0.66191036,0.71678376,0.70306545,0.7133542,0.7888051,0.9294182,0.9602845,0.8676856,0.82996017,0.7407909,0.6756287,0.7682276,0.9568549,0.9911508,1.0048691,1.0460242,0.9328478,0.6962063,0.5624523,0.6036074,0.5590228,0.52815646,0.5658819,0.6790583,0.72707254,0.7613684,0.7510797,0.72707254,0.7339317,0.7339317,0.70649505,0.66876954,0.6173257,0.5178677,0.5555932,0.6756287,0.8025235,0.89855194,0.980862,1.039165,1.0563129,1.0460242,1.0323058,1.0528834,1.0220171,1.0700313,1.2346514,1.4541451,1.5638919,1.6907866,1.762808,1.7525192,1.6667795,1.5433143,1.3409687,1.039165,0.83338976,0.7682276,0.7407909,0.65505123,0.6001778,0.53501564,0.47671264,0.5041494,0.5761707,0.5658819,0.4938606,0.4081209,0.38754338,0.33952916,0.3806842,0.41840968,0.44584638,0.53844523,0.69963586,0.8162418,0.91569984,1.0048691,1.0871792,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.09945804,0.26750782,0.45270553,0.22292319,0.07545093,0.024007112,0.037725464,0.058302987,0.2469303,0.4389872,0.548734,0.53501564,0.42526886,0.39783216,0.31209245,0.28465575,0.2777966,0.12346515,0.08916927,0.09602845,0.16804978,0.3018037,0.47671264,0.764798,1.5570327,2.5447538,3.2272418,2.9220085,3.3232703,5.4153185,7.9257765,9.815479,10.285333,11.818358,16.13621,22.319756,30.92802,44.008465,60.09666,59.86345,48.20971,32.522778,22.666143,12.38424,7.373613,5.0929375,3.7965534,2.5207467,2.435007,2.4384367,2.2429502,1.8999915,1.8176813,2.253239,2.7299516,3.117495,3.2512488,2.8980014,2.8019729,2.7711067,2.8328393,2.8019729,2.287535,1.7696671,1.4095604,1.1214751,0.91912943,0.90198153,0.9945804,1.1694894,1.313532,1.3375391,1.1832076,1.2380811,1.255229,1.1351935,0.9294182,0.8505377,0.70306545,0.7339317,0.7613684,0.71678376,0.65162164,0.72707254,0.65848076,0.47328308,0.30866286,0.4081209,0.4424168,0.4081209,0.6790583,1.2380811,1.704505,2.6304936,3.5393343,4.5647807,6.0703697,8.652849,11.574858,16.914726,29.168642,47.739857,66.95241,61.98979,44.361713,28.863409,21.215427,18.04992,12.922686,10.628291,9.129561,8.220721,9.5205345,12.71691,13.828096,13.536582,11.952112,8.632272,7.716572,7.459353,7.1541195,6.835168,7.3118806,9.856634,13.7526455,15.597764,14.562028,12.401388,13.193623,12.823228,14.819247,17.78927,15.422854,10.971251,14.640909,16.94902,16.29397,18.931322,18.180243,27.546446,50.775043,72.10708,56.300106,23.640146,15.560039,16.822126,18.557497,18.259123,14.658057,19.198832,42.657207,69.1199,55.981155,22.144846,7.6857057,10.151579,17.069057,5.953764,13.6086035,16.993607,14.743796,10.261326,11.698323,13.138749,13.214201,13.673765,15.21022,17.4566,16.63007,16.173935,14.321958,10.827208,6.9620624,4.9488945,9.866923,13.039291,10.388221,2.435007,6.15268,13.046151,16.554619,16.46545,18.917604,20.989075,14.009865,7.675417,6.759717,11.122152,17.61436,26.208908,29.43272,26.647894,24.061985,38.377083,41.31624,35.39334,26.088871,21.849901,26.147175,30.070623,29.59391,23.098272,11.348505,9.534253,8.635701,8.100685,7.8126,8.073249,12.079007,12.617453,11.173596,10.600855,15.110763,9.877212,9.057541,10.199594,11.753197,13.066729,17.158226,20.86561,24.09971,28.400414,36.946945,62.823185,73.605804,64.13672,40.102165,18.015623,11.585147,13.073587,17.600643,20.886189,19.233126,13.190193,12.116733,14.599753,20.872469,32.82458,49.684433,48.885338,43.024174,37.951817,32.773136,18.924463,16.88043,16.225378,12.566009,7.5039372,10.076128,9.122703,8.320179,9.712592,13.725209,12.9707,15.63206,13.63261,10.271614,20.224277,14.572317,10.213311,11.948683,18.54378,22.755312,7.407909,5.761707,11.698323,15.827546,5.4736214,1.6873571,2.760818,5.3501563,9.0369625,16.341984,17.562918,9.115844,4.187526,9.146709,23.547548,12.133881,5.8817425,3.1209247,2.6407824,3.7039545,4.355576,6.5882373,11.207891,16.62321,18.866161,19.143957,11.159878,13.104454,26.610168,36.76861,14.424845,22.347193,30.876575,25.372087,6.2075534,9.719451,11.598865,14.428274,18.108221,19.86417,8.30646,4.650521,10.30934,17.909306,11.276484,7.160979,16.54433,20.574095,14.222499,6.2864337,4.417309,5.802862,6.210983,4.6265135,3.2375305,2.170929,1.587899,1.1900668,0.91912943,0.9842916,1.1832076,1.4610043,1.3546871,1.0734608,1.488441,2.1812177,3.4707425,5.0174866,6.0223556,5.219832,3.059192,2.6236343,3.0626216,3.865145,4.852866,4.389872,4.4721823,3.8342788,2.603057,2.301253,2.5138876,3.1620796,2.6716487,1.6153357,2.7162333,3.4398763,2.952875,3.8034124,5.861165,6.324159,5.90575,4.396731,3.1655092,3.0557625,4.383013,6.509357,7.06495,6.5196457,4.8288593,1.4472859,1.4644338,2.0268862,2.9460156,3.566771,2.7711067,1.3855534,2.9940298,4.180667,3.9028704,3.4776018,8.368194,7.517656,4.852866,2.767677,2.1057668,3.0489032,2.2086544,1.3341095,1.039165,0.8196714,0.82996017,0.6927767,0.4389872,0.18176813,0.1097468,0.11317638,0.15090185,0.18862732,0.18519773,0.10288762,0.037725464,0.048014224,0.10288762,0.14747226,0.106317215,0.0548734,0.024007112,0.010288762,0.010288762,0.020577524,0.12003556,0.10288762,0.08573969,0.09602845,0.08916927,0.41840968,0.5693115,0.6001778,0.764798,1.4953002,0.89512235,0.39440256,0.14061308,0.106317215,0.08916927,0.06859175,0.06859175,0.07888051,0.11317638,0.1920569,0.78537554,0.70649505,0.38754338,0.13375391,0.09945804,0.26064864,0.96714365,1.762808,1.9548649,0.607037,0.8745448,0.8745448,0.6790583,0.36696586,0.020577524,0.4629943,0.78537554,0.90198153,0.94999576,1.2895249,1.6256244,1.3752645,1.0906088,0.9431366,0.6927767,0.4698535,0.5693115,0.58645946,0.4081209,0.22292319,0.1371835,0.09602845,0.17490897,0.37382504,0.6276145,0.29494452,0.22292319,0.28122616,0.38754338,0.490431,0.34638834,0.18519773,0.08573969,0.058302987,0.06859175,0.17490897,0.3018037,0.33266997,0.32238123,0.4972902,0.53158605,0.5418748,0.45956472,0.29494452,0.12346515,0.106317215,0.09259886,0.07888051,0.07545093,0.09945804,0.10288762,0.061732575,0.0274367,0.01371835,0.0,0.0034295875,0.01371835,0.030866288,0.05144381,0.07545093,0.10288762,0.14747226,0.14061308,0.08573969,0.058302987,0.0274367,0.020577524,0.020577524,0.020577524,0.048014224,0.15776102,0.22635277,0.28122616,0.32924038,0.37725464,0.3018037,0.29494452,0.25721905,0.16804978,0.09945804,0.10288762,0.1097468,0.15776102,0.26750782,0.41840968,0.50757897,0.65162164,0.8025235,0.9534253,1.138623,1.1420527,0.881404,0.6310441,0.490431,0.3806842,0.29837412,0.274367,0.274367,0.31552204,0.47328308,0.607037,0.48357183,0.38754338,0.40126175,0.42183927,0.432128,0.5007198,0.5761707,0.6756287,0.88826317,1.2243627,1.1180456,0.8779744,0.6893471,0.61389613,0.44584638,0.4972902,0.65505123,0.8265306,0.939707,0.94656616,1.0082988,1.1523414,1.3341095,1.4369972,1.2415106,1.1866373,1.2586586,1.4369972,1.6976458,1.5158776,1.587899,1.6221949,1.4781522,1.1660597,1.0048691,0.922559,0.823101,0.7407909,0.83338976,0.9602845,1.0528834,1.08032,1.0151579,0.8265306,0.70649505,0.6310441,0.6379033,0.71678376,0.8128122,0.8196714,0.83338976,0.805953,0.77165717,0.85396725,0.9294182,0.77851635,0.6173257,0.58645946,0.7442205,0.8162418,0.7682276,0.69963586,0.65505123,0.6241849,0.71678376,0.7682276,0.72707254,0.6310441,0.6173257,0.5796003,0.61046654,0.7305021,0.88826317,0.97400284,0.99801,1.0460242,1.0185875,0.89169276,0.72707254,0.6893471,0.6241849,0.6241849,0.70649505,0.8093826,0.85396725,0.85739684,0.8265306,0.78194594,0.77508676,0.8128122,0.8128122,0.8025235,0.764798,0.64476246,0.72364295,0.84024894,0.91569984,0.9774324,1.1454822,1.2689474,1.2106444,1.1351935,1.1180456,1.1454822,1.0837497,1.039165,1.0871792,1.2072148,1.2758065,1.4095604,1.5055889,1.546744,1.5673214,1.6324836,1.5193073,1.4918705,1.3341095,1.0563129,0.89512235,0.7922347,0.7133542,0.67219913,0.65505123,0.65848076,0.64476246,0.6173257,0.5693115,0.5041494,0.47328308,0.4698535,0.53501564,0.59331864,0.61046654,0.5761707,0.607037,0.7407909,0.91569984,1.0597426,1.0837497,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058302987,0.19891608,0.42869842,0.30523327,0.11317638,0.010288762,0.020577524,0.034295876,0.1920569,0.39440256,0.490431,0.4664239,0.4115505,0.39097297,0.32924038,0.28465575,0.25721905,0.18176813,0.12346515,0.14061308,0.25378948,0.4355576,0.61046654,0.8505377,1.5193073,2.503599,3.426158,3.649081,4.1292233,5.9983487,8.357904,10.439664,11.592006,12.253916,15.001016,20.080235,28.17749,40.414257,58.237823,58.340714,45.24312,26.973705,15.042171,8.2310095,5.7754254,4.623084,3.3678548,2.2566686,2.3424082,2.2292318,1.937717,1.6873571,1.879414,2.153781,2.3492675,2.4247184,2.2120838,1.4095604,1.2243627,1.3341095,1.6770682,2.0440342,2.0886188,1.8005334,1.6221949,1.3786942,1.08032,0.939707,1.0220171,1.2346514,1.3512574,1.2860953,1.0666018,1.0185875,1.0117283,0.881404,0.6790583,0.65505123,0.6241849,0.72021335,0.77508676,0.72707254,0.64133286,0.6859175,0.66876954,0.53844523,0.39440256,0.4938606,0.5761707,0.7682276,1.2483698,1.845118,2.0268862,2.7333813,3.5359046,4.715683,6.543653,9.280463,12.9707,21.139977,38.10272,60.720844,78.41752,66.57515,47.99365,36.233593,33.040646,28.3524,16.20137,9.990388,7.891481,8.604835,11.341646,12.171606,12.994707,13.505715,12.634601,8.543102,7.4696417,7.9737906,7.846896,6.8454566,6.701414,8.299602,11.519984,13.783512,15.422854,19.675543,22.991955,18.03277,14.915276,15.645778,14.13676,10.508256,11.962401,17.641798,24.85765,29.082901,22.94051,25.049707,46.741848,73.780716,66.3728,33.222412,20.882757,20.70785,26.661613,35.304173,29.906002,21.386908,29.59391,46.693832,37.15958,15.885849,6.327589,10.429376,17.53548,4.396731,14.2533655,17.562918,13.601744,6.1561093,3.5187566,8.285883,9.287323,7.9909387,7.2467184,11.297061,17.741257,16.990177,11.489118,4.897451,2.061182,4.7808447,10.419086,13.406258,10.765475,2.1194851,6.4887795,13.337666,19.161106,21.963078,21.260014,20.598103,15.63206,10.1481495,7.4627824,10.429376,22.707298,41.590607,50.37378,42.664066,22.422644,19.325726,17.394867,15.415996,13.560589,13.371962,16.770683,19.188541,18.70497,14.479718,6.7357097,8.279024,9.801761,9.242738,7.301592,7.431916,11.852654,13.893259,12.38767,9.949233,12.956982,10.604284,8.868914,9.788043,11.89038,10.206452,12.147599,16.156786,19.716698,22.234016,25.029129,39.690617,43.56948,36.789185,23.749893,13.125031,7.73372,7.4353456,9.318189,11.101575,11.125582,10.930096,13.625751,16.828985,21.503513,31.956896,40.270218,35.482513,31.991192,34.33703,37.214455,26.205479,17.885298,14.109323,13.22106,10.048691,10.179015,8.546532,7.1849856,8.368194,14.606613,13.056439,15.354263,14.153908,11.026124,16.45859,12.72034,10.041832,10.302481,12.826657,14.3974085,5.0929375,8.093826,13.88297,14.695783,4.5167665,4.887162,10.8958,12.792361,9.472521,8.48137,7.630832,5.2266912,4.431027,9.3764925,25.169743,13.210771,5.8337283,2.7985435,2.760818,3.2581081,3.234101,5.7411294,11.074138,16.074476,14.143619,11.814929,7.373613,11.691463,24.981115,36.796043,14.102464,19.744135,25.049707,18.183672,4.15666,8.337327,8.608265,7.846896,9.794902,19.058218,9.925226,8.172707,13.937843,19.486916,9.225591,7.6445503,17.532051,19.486916,10.751757,5.2301207,5.2026844,6.375603,6.012067,3.998899,2.860276,1.4129901,0.8779744,0.6893471,0.64819205,0.91912943,0.9842916,1.1763484,1.0631721,0.8711152,1.4953002,1.7525192,1.8691251,2.393852,3.2992632,4.0023284,3.0797696,2.6613598,2.633923,3.0420442,4.108646,4.1189346,4.3109913,3.5530527,2.2498093,2.311542,2.2292318,2.7333813,2.8396983,2.8328393,4.2595477,4.448175,3.0077481,3.223812,5.195825,5.8405876,5.7377,4.7534084,3.8720043,3.7553983,4.7499785,4.8014226,5.5490727,6.2898636,5.689686,1.8176813,1.4610043,1.728512,2.5996273,3.391862,2.7539587,1.2072148,2.277246,3.806842,4.434457,3.5839188,4.5510626,6.060081,5.675967,3.3952916,1.6290541,2.6853669,2.393852,1.8519772,1.4575747,0.89855194,0.8848336,0.7442205,0.5624523,0.3841138,0.19548649,0.16119061,0.19891608,0.23664154,0.22292319,0.1097468,0.044584636,0.06859175,0.16462019,0.2503599,0.17833854,0.09945804,0.05144381,0.0274367,0.01371835,0.01371835,0.08573969,0.09259886,0.05144381,0.010288762,0.034295876,0.32581082,0.4046913,0.6276145,1.0906088,1.6530612,1.2209331,0.65505123,0.29151493,0.18862732,0.14404267,0.09945804,0.06859175,0.072021335,0.09945804,0.12346515,0.38754338,0.3566771,0.22978236,0.16119061,0.26407823,0.4081209,0.607037,1.2243627,1.7113642,0.58988905,0.67219913,0.8025235,0.9842916,0.9294182,0.041155048,0.09259886,0.7339317,0.8196714,0.36353627,0.5418748,1.6256244,1.529596,1.0666018,0.6790583,0.42869842,0.41840968,0.5453044,0.5453044,0.37039545,0.20920484,0.37382504,0.26750782,0.2503599,0.4664239,0.85396725,0.4115505,0.20920484,0.274367,0.44927597,0.39440256,0.33609957,0.16804978,0.058302987,0.05144381,0.061732575,0.1920569,0.24007112,0.21263443,0.20234565,0.3566771,0.274367,0.4698535,0.70649505,0.7373613,0.29151493,0.12003556,0.07888051,0.08573969,0.09259886,0.07545093,0.082310095,0.082310095,0.0548734,0.01371835,0.0,0.0,0.006859175,0.010288762,0.01371835,0.034295876,0.10288762,0.14747226,0.14404267,0.09945804,0.041155048,0.020577524,0.010288762,0.010288762,0.01371835,0.024007112,0.106317215,0.17490897,0.24350071,0.30866286,0.34295875,0.14404267,0.06859175,0.048014224,0.037725464,0.034295876,0.017147938,0.017147938,0.020577524,0.024007112,0.0274367,0.08573969,0.2194936,0.39440256,0.6001778,0.8711152,1.1008976,0.96714365,0.7442205,0.5693115,0.42869842,0.274367,0.20920484,0.20234565,0.2469303,0.3566771,0.5212973,0.4389872,0.3566771,0.34638834,0.31209245,0.32238123,0.36696586,0.45270553,0.607037,0.88826317,1.1283343,1.0014396,0.8196714,0.6962063,0.5453044,0.41498008,0.6001778,0.83338976,0.922559,0.77508676,0.70306545,0.8196714,1.0220171,1.2380811,1.4507155,1.5810398,1.3375391,1.2209331,1.3786942,1.5913286,1.5638919,1.5501735,1.5673214,1.529596,1.2517995,1.1934965,1.1283343,0.980862,0.823101,0.88826317,1.0048691,1.1763484,1.2860953,1.2689474,1.0940384,0.99801,0.8711152,0.7579388,0.6859175,0.65848076,0.66533995,0.8162418,0.90541106,0.89512235,0.91569984,1.0940384,0.9945804,0.8162418,0.71678376,0.8128122,0.8128122,0.70649505,0.607037,0.5658819,0.59674823,0.6824879,0.6859175,0.6001778,0.48700142,0.47671264,0.5521636,0.6276145,0.7099246,0.7990939,0.88826317,0.94656616,0.9945804,1.0151579,0.96714365,0.77508676,0.72021335,0.7442205,0.7956643,0.8471081,0.90198153,0.90541106,0.864256,0.85396725,0.8779744,0.8676856,0.90541106,1.0185875,1.1351935,1.1866373,1.1077567,1.0940384,1.1454822,1.1420527,1.1454822,1.3649758,1.5570327,1.5536032,1.5090185,1.5227368,1.6016173,1.488441,1.3032433,1.1866373,1.1626302,1.1763484,1.2243627,1.2792361,1.3169615,1.3752645,1.5227368,1.4918705,1.6599203,1.6290541,1.3512574,1.1008976,1.0563129,1.0048691,0.94999576,0.90541106,0.89855194,0.7956643,0.7613684,0.7407909,0.6893471,0.5693115,0.548734,0.58988905,0.6379033,0.64476246,0.5693115,0.5761707,0.66876954,0.7990939,0.91227025,0.980862,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.048014224,0.216064,0.1097468,0.006859175,0.0034295875,0.01371835,0.09259886,0.28808534,0.42183927,0.44927597,0.4698535,0.5007198,0.42183927,0.31552204,0.25378948,0.32238123,0.19548649,0.18862732,0.29494452,0.4698535,0.6276145,0.9431366,1.5844694,2.6750782,3.974892,4.897451,5.675967,7.6685576,10.134431,12.442543,14.088745,13.96185,15.165636,18.187103,24.302057,35.57511,55.95372,53.35409,37.612286,19.11309,8.779744,5.693115,4.9248877,4.290414,3.069481,2.0097382,2.1880767,1.8999915,1.6633499,1.7319417,2.0749004,1.920569,1.7422304,1.5776103,1.3924125,1.0734608,0.805953,0.75450927,1.1111864,1.7319417,2.153781,2.0303159,1.8279701,1.4918705,1.0871792,0.7956643,0.7442205,0.7922347,0.8265306,0.823101,0.864256,0.9259886,0.84024894,0.6379033,0.45956472,0.5796003,0.5453044,0.53158605,0.5693115,0.6173257,0.5727411,0.58988905,0.6173257,0.6001778,0.5727411,0.6379033,0.8779744,1.2963841,1.7730967,2.1297739,2.1469216,2.7230926,3.4055803,4.9214582,7.4284863,10.528833,14.404267,22.62156,39.049282,58.838,68.413414,51.831356,38.77149,37.711742,43.98789,39.8278,21.1194,10.031544,6.8866115,9.3764925,12.566009,9.956093,9.3079,11.489118,14.157337,11.784062,10.63858,11.207891,10.837497,9.383351,9.22902,8.056101,8.882631,13.471419,23.719027,41.635193,48.178844,31.929459,16.383139,10.81006,10.230459,9.270175,10.9369545,19.071936,31.003471,37.533405,31.26069,25.252052,40.846386,69.00673,70.33741,40.537724,21.829325,18.44775,29.377846,48.336605,49.101402,29.542467,16.938732,18.03963,19.082224,10.81006,8.484799,12.596875,16.067617,4.262977,14.239647,16.074476,12.332796,6.39961,2.4795918,9.427936,9.932085,6.5470824,4.396731,11.153018,22.43979,21.407484,12.710052,3.3061223,2.4384367,8.7283,13.886399,14.839825,10.422516,1.3992717,9.719451,17.442883,23.009102,24.171732,18.019053,11.008976,12.010415,13.282792,12.295071,11.739478,22.628418,46.124523,59.633667,51.172874,19.377169,8.347616,5.586798,7.449064,9.942374,8.7283,9.253027,9.3079,8.296172,6.0497923,2.8019729,7.6514096,13.22106,15.755525,13.056439,4.5030484,5.4153185,10.909517,15.247946,16.088194,14.496866,13.673765,10.521975,10.796341,13.183334,9.290752,9.901219,13.924125,17.04848,17.703531,17.03819,22.11055,21.554956,18.691252,15.127911,10.751757,5.470192,3.7965534,3.8274195,4.314421,4.647091,7.2124224,12.298501,16.438013,20.11453,27.76937,32.40274,31.360147,35.81518,45.767845,50.034252,40.366245,23.232025,14.016724,14.994157,15.333686,11.633161,7.589677,7.023795,10.868362,17.189093,14.990726,12.874671,12.363663,12.445972,9.561689,8.81747,7.6205435,6.9860697,6.183546,2.726522,3.590778,12.106443,15.721229,10.97468,3.4981792,10.930096,19.853882,17.7927,6.6122446,2.5241764,3.5187566,5.007198,4.7808447,4.633373,10.353925,8.553391,4.9351764,2.8980014,3.1586502,3.7519686,3.9200184,6.433906,9.407358,10.621432,7.5450926,9.856634,9.098696,10.9198065,17.730967,28.736513,13.834956,22.254593,22.755312,9.695444,3.0283258,8.056101,7.5279446,5.144381,6.0326443,16.739817,13.245067,13.790371,16.444872,16.403717,5.9812007,7.0443726,14.390549,14.438563,6.8145905,4.3761535,6.111525,5.672538,4.7979927,4.184097,3.4776018,1.2758065,0.64133286,0.5178677,0.490431,0.7613684,0.65162164,0.6824879,0.7373613,1.1489118,2.6853669,2.6236343,1.762808,1.2003556,1.4232788,2.277246,2.4898806,2.3835633,2.16064,2.318401,3.6627994,3.4810312,3.9543142,3.6970954,2.7128036,2.4007113,1.903421,2.469303,3.673088,4.99005,5.778855,5.1752477,3.474172,3.1552205,4.5442033,5.7994323,5.521636,4.290414,3.5599117,3.9028704,5.003768,2.6545007,3.2958336,5.1855364,6.0737996,3.1963756,1.8897027,1.5707511,2.277246,3.1449318,2.386993,1.3032433,1.4438564,2.5241764,3.6319332,3.199805,1.8142518,3.8960114,5.0449233,3.8548563,1.9239986,2.9391565,3.3129816,3.3026927,2.784825,1.2415106,0.7579388,0.6241849,0.67219913,0.6824879,0.40126175,0.24007112,0.2469303,0.22635277,0.1371835,0.07545093,0.048014224,0.11317638,0.28465575,0.432128,0.29837412,0.15090185,0.07888051,0.037725464,0.01371835,0.01371835,0.0548734,0.0548734,0.037725464,0.020577524,0.01371835,0.5555932,0.5658819,0.89169276,1.4987297,1.4987297,1.4610043,1.0082988,0.5555932,0.29494452,0.20920484,0.12003556,0.07888051,0.07545093,0.08916927,0.061732575,0.2503599,0.31209245,0.22978236,0.17833854,0.5555932,0.78537554,0.5041494,0.37382504,0.51100856,0.4938606,0.5624523,0.5453044,0.97400284,1.3409687,0.09602845,0.072021335,0.607037,0.67219913,0.28465575,0.53501564,1.3821237,1.1934965,0.70306545,0.39440256,0.48700142,0.39783216,0.35324752,0.34638834,0.32924038,0.22292319,0.6344737,0.41840968,0.216064,0.29837412,0.5693115,0.36353627,0.16804978,0.25721905,0.4664239,0.1920569,0.23321195,0.12003556,0.058302987,0.09259886,0.10288762,0.17833854,0.15433143,0.09945804,0.061732575,0.06859175,0.11317638,0.5178677,1.0323058,1.2380811,0.548734,0.14061308,0.07545093,0.1097468,0.10288762,0.041155048,0.034295876,0.082310095,0.07545093,0.01371835,0.0,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0548734,0.082310095,0.09602845,0.082310095,0.030866288,0.017147938,0.0034295875,0.0,0.0034295875,0.01371835,0.034295876,0.072021335,0.12346515,0.17833854,0.21263443,0.06859175,0.024007112,0.020577524,0.030866288,0.05144381,0.030866288,0.0274367,0.0274367,0.020577524,0.0,0.0,0.006859175,0.05144381,0.18176813,0.48357183,0.7922347,0.90541106,0.7579388,0.4698535,0.34981793,0.29837412,0.26750782,0.23664154,0.20234565,0.16804978,0.19548649,0.24350071,0.274367,0.26750782,0.20920484,0.23664154,0.274367,0.33266997,0.47328308,0.8196714,0.9259886,0.78537554,0.6276145,0.53158605,0.432128,0.5624523,0.8265306,0.9877212,0.9259886,0.607037,0.5590228,0.66191036,0.823101,0.97400284,1.0837497,1.6976458,1.3203912,1.08032,1.2860953,1.3992717,1.6976458,1.5707511,1.5055889,1.5844694,1.471293,1.471293,1.3821237,1.1660597,0.9362774,0.9534253,0.97057325,1.1866373,1.3855534,1.4678634,1.4129901,1.4061309,1.2689474,1.0734608,0.8505377,0.5693115,0.5178677,0.8162418,1.0151579,0.96371406,0.83338976,0.980862,0.9602845,0.8676856,0.7613684,0.67219913,0.5624523,0.52815646,0.490431,0.45613512,0.5144381,0.6173257,0.6893471,0.65848076,0.5453044,0.48357183,0.61046654,0.64819205,0.6790583,0.7339317,0.7888051,0.90198153,0.9328478,0.90884066,0.83681935,0.70306545,0.6893471,0.8265306,0.90541106,0.88826317,0.922559,0.90541106,0.83338976,0.86082643,0.96714365,0.96714365,1.0048691,1.2895249,1.5536032,1.6804979,1.6770682,1.5330256,1.5158776,1.4781522,1.4541451,1.6256244,1.8039631,1.9274281,1.9891608,2.0303159,2.1434922,1.9823016,1.7113642,1.471293,1.3203912,1.2277923,1.2346514,1.2449403,1.2380811,1.2517995,1.3443983,1.4095604,1.5501735,1.6187652,1.5570327,1.3821237,1.4232788,1.3958421,1.2689474,1.1214751,1.1214751,1.0220171,1.0082988,0.9842916,0.8848336,0.67219913,0.61046654,0.58988905,0.5796003,0.5521636,0.490431,0.53501564,0.5521636,0.5453044,0.5727411,0.7579388,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.22292319,0.37039545,0.45613512,0.5178677,0.5178677,0.42869842,0.32924038,0.32238123,0.5178677,0.31209245,0.2503599,0.32238123,0.4938606,0.70306545,1.0563129,1.5741806,2.5996273,4.0057583,5.2026844,6.9380555,9.081548,11.640019,14.003006,14.970149,14.579176,15.6697855,16.20137,18.605513,29.799686,44.924168,42.20793,29.49788,14.894698,6.728851,4.7774153,4.0023284,3.4673128,2.7059445,1.7559488,2.0097382,1.8656956,1.6221949,1.5364552,1.8313997,1.8416885,1.6187652,1.3546871,1.1111864,0.7922347,0.5727411,0.52815646,0.64476246,0.89855194,1.2517995,1.4575747,0.980862,0.5693115,0.48014224,0.4424168,0.5144381,0.48700142,0.53158605,0.70649505,0.9602845,0.8745448,0.65162164,0.51100856,0.53158605,0.64133286,0.42183927,0.33952916,0.34981793,0.41498008,0.48700142,0.7579388,0.7956643,0.7956643,0.85739684,0.9911508,1.371835,1.4918705,1.6942163,2.0508933,2.3801336,3.0146074,3.5599117,4.9008803,8.014946,13.944703,18.828436,20.460918,25.207468,32.24498,33.58595,24.212887,26.781649,38.1473,48.923065,43.50089,24.912523,13.735497,12.240198,16.911295,18.46147,10.347065,6.64997,8.707723,12.857523,10.4533825,12.490558,10.621432,7.2467184,4.7842746,5.675967,8.31332,15.076467,26.1849,42.736088,66.70891,69.919,42.307392,19.394318,14.359683,18.019053,13.893259,13.934414,17.919594,22.789608,22.628418,19.723558,13.790371,20.11796,36.586838,43.641502,30.286688,21.846472,21.232576,29.710516,46.920185,54.1086,37.725464,20.989075,16.005884,23.756752,15.395418,20.004784,29.508171,30.444448,3.981751,13.101024,17.78927,15.608052,8.899779,4.7602673,11.780633,10.285333,5.425607,3.8788633,13.838386,17.820137,16.983316,10.007536,2.2909644,5.967482,13.876111,19.919044,16.523752,5.9880595,0.45613512,11.163307,19.569225,24.027689,21.897917,9.582268,4.4687524,8.069819,13.227919,16.160215,16.46545,16.417435,18.272842,24.92624,27.909983,7.4010496,2.9460156,4.0366244,7.7851634,11.780633,14.099034,20.251715,14.246507,6.800872,2.9494452,2.0440342,8.134981,19.984205,28.712505,27.258362,10.374502,5.360445,13.855534,30.224955,45.733547,48.566387,26.082012,13.347955,11.7257595,15.9921665,14.342535,10.960961,11.626302,13.214201,14.157337,14.448852,13.88983,13.557159,12.843805,10.899229,6.636252,3.673088,3.2409601,4.2835546,6.1629686,8.652849,12.240198,17.20281,18.269413,16.45173,19.027351,24.76505,25.85223,28.966295,35.948936,43.80955,33.946056,22.974806,18.348293,19.60695,18.386019,15.6526375,11.351934,9.856634,13.773223,23.94195,23.880217,17.96761,10.875222,7.058091,10.7586155,11.379372,10.840926,10.504827,9.369633,4.057202,11.345076,14.1299,9.72288,2.668219,4.729401,15.0456,11.746337,5.802862,2.6579304,2.2429502,8.48137,13.4645605,11.7257595,5.312431,3.799983,6.7048435,4.712253,3.2889743,4.396731,6.48535,6.495639,7.6616983,7.2364297,6.495639,10.741467,15.758954,13.197053,10.497967,12.744347,22.645567,18.015623,23.341772,21.256582,9.815479,2.503599,10.803201,9.105555,5.535354,3.9200184,3.799983,11.869802,16.074476,14.675205,9.156999,4.2115335,5.5662203,14.328816,17.024471,11.101575,4.914599,6.4133286,7.0752387,7.14726,6.1766872,2.9906003,1.8416885,1.2003556,0.78537554,0.490431,0.3806842,0.5658819,0.4629943,0.36010668,1.0014396,3.6010668,5.1992545,3.7794054,2.4898806,2.3252604,2.1057668,1.8005334,2.0714707,2.7368107,3.4295874,3.6010668,4.1120753,4.746549,4.746549,4.098357,3.525616,1.8142518,2.0474637,3.340418,5.0243454,6.6225333,6.036074,4.8837323,4.297273,4.4687524,4.6402316,7.3118806,5.0243454,3.0077481,3.2821152,4.6402316,2.9906003,3.5942078,5.3330083,6.7494283,6.042933,2.5756202,1.7456601,2.3081124,2.8877127,1.9823016,1.1180456,1.0734608,2.0131679,3.5804894,4.897451,4.3109913,2.719663,2.4830213,3.350707,2.4727325,2.1297739,4.0777793,5.0826488,4.0606318,2.061182,0.9602845,0.805953,0.8676856,0.7888051,0.59674823,0.29151493,0.26064864,0.20920484,0.07545093,0.01371835,0.01371835,0.13375391,0.34638834,0.50757897,0.33609957,0.17833854,0.072021335,0.017147938,0.0034295875,0.01371835,0.01371835,0.041155048,0.0548734,0.037725464,0.0,0.61046654,0.66191036,0.91227025,1.4610043,1.7559488,1.9514352,1.6599203,1.097468,0.52815646,0.26064864,0.09945804,0.034295876,0.05144381,0.09602845,0.061732575,0.37725464,0.64133286,0.53158605,0.33609957,0.94656616,1.5570327,1.0768905,0.8162418,1.0185875,0.8848336,0.39783216,0.548734,0.64133286,0.4389872,0.18176813,0.048014224,0.28122616,0.40126175,0.4355576,0.89855194,1.0357354,0.8196714,0.6207553,0.6824879,1.1592005,0.61046654,0.32581082,0.26407823,0.29494452,0.19891608,0.2469303,0.14061308,0.08573969,0.13032432,0.16804978,0.25378948,0.2469303,0.22978236,0.1920569,0.044584636,0.15433143,0.1097468,0.17147937,0.32238123,0.274367,0.21263443,0.12346515,0.06859175,0.082310095,0.16804978,0.044584636,0.14404267,0.58988905,1.039165,0.67219913,0.18176813,0.07888051,0.09602845,0.09945804,0.07545093,0.05144381,0.037725464,0.030866288,0.024007112,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.01371835,0.034295876,0.044584636,0.041155048,0.030866288,0.006859175,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.037725464,0.041155048,0.030866288,0.030866288,0.030866288,0.024007112,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.017147938,0.082310095,0.22978236,0.64476246,0.8471081,0.67219913,0.3018037,0.29151493,0.4115505,0.39783216,0.274367,0.13032432,0.106317215,0.14404267,0.216064,0.25378948,0.22292319,0.1371835,0.17490897,0.1920569,0.20577525,0.26064864,0.4424168,0.6241849,0.4972902,0.38754338,0.4081209,0.45613512,0.8128122,0.9568549,0.91912943,0.8025235,0.77851635,0.7305021,0.67219913,0.7888051,0.94999576,0.71678376,0.864256,0.94656616,0.9534253,0.922559,0.94656616,1.4232788,1.5124481,1.3924125,1.2380811,1.2517995,1.2517995,1.2517995,1.1729189,1.0254467,0.91569984,1.0117283,1.1660597,1.3169615,1.4369972,1.5090185,1.7182233,1.6770682,1.5364552,1.3032433,0.84024894,0.71678376,0.823101,0.9568549,0.9911508,0.8711152,0.91912943,0.94999576,0.94999576,0.89169276,0.7339317,0.6241849,0.6790583,0.66533995,0.5041494,0.26064864,0.5144381,0.607037,0.64476246,0.65505123,0.59674823,0.53501564,0.5178677,0.5555932,0.6207553,0.65505123,0.764798,0.7476501,0.6790583,0.64133286,0.70306545,0.6893471,0.7682276,0.8676856,0.94656616,1.0082988,1.0185875,0.94999576,0.88826317,0.881404,0.9294182,1.1763484,1.5741806,1.7833855,1.762808,1.8005334,1.862266,1.8862731,1.903421,1.920569,1.9068506,1.9685832,2.085189,2.1469216,2.1297739,2.1057668,2.0817597,1.9102802,1.6907866,1.4815818,1.313532,1.3992717,1.3101025,1.2175035,1.2106444,1.2963841,1.4678634,1.6221949,1.6804979,1.6633499,1.6633499,1.7250825,1.6187652,1.4061309,1.2072148,1.2209331,1.1489118,1.155771,1.0906088,0.939707,0.85396725,0.9877212,0.922559,0.7922347,0.6241849,0.31895164,0.19891608,0.20577525,0.24007112,0.26750782,0.30523327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.116605975,0.23664154,0.34981793,0.42183927,0.432128,0.37039545,0.3018037,0.274367,0.32238123,0.29151493,0.26064864,0.30523327,0.44584638,0.65162164,1.0837497,1.7833855,2.5550427,3.2306714,3.666229,4.557922,6.756287,9.39021,11.753197,13.334236,13.858963,14.208781,14.099034,16.70895,28.664492,38.449104,35.33161,24.322634,11.873232,5.874883,4.400161,3.6079261,2.9631636,2.2052248,1.3512574,1.3546871,1.3924125,1.4781522,1.5604624,1.5501735,1.5124481,1.5913286,1.4198492,1.0768905,1.0631721,0.7922347,0.5658819,0.45270553,0.44927597,0.48357183,0.53501564,0.4698535,0.432128,0.4389872,0.39440256,0.42869842,0.3841138,0.40126175,0.5144381,0.64476246,0.58645946,0.52472687,0.5453044,0.61389613,0.5693115,0.45613512,0.41498008,0.39097297,0.4115505,0.5624523,0.7922347,0.922559,0.99801,1.0288762,1.0151579,1.0837497,1.3032433,1.4678634,1.903421,3.4433057,2.7573884,3.6970954,6.866034,12.758065,21.747015,27.09717,24.11,21.891056,24.53184,31.120077,34.820602,39.0047,43.34313,44.200523,34.64226,21.225718,13.358243,13.663476,18.663815,18.766703,9.860064,5.586798,5.439326,7.4799304,8.327039,7.740579,7.922347,8.868914,11.664027,18.492336,28.901134,37.16987,40.757217,43.692944,56.605343,48.772163,27.090311,21.3629,32.461044,32.32729,24.185452,17.247395,13.876111,15.271953,21.469217,18.934752,12.593445,13.954991,24.19231,34.16898,22.494663,13.392539,13.399398,22.793037,35.58197,40.194763,27.560165,13.1593275,6.941485,13.296511,11.917816,14.027013,16.952452,15.608052,2.49331,6.807731,9.928656,9.280463,6.9860697,9.849775,10.659158,7.7885933,5.305572,7.1369715,17.04848,15.981877,11.8115,6.509357,4.537344,12.850664,17.147938,17.182234,12.017275,4.5167665,1.3478279,7.6788464,12.445972,14.88441,13.786942,7.4936485,2.9288676,8.004657,15.549749,20.649546,20.649546,18.11165,11.825217,10.734609,12.9707,5.8508763,4.822,7.1232533,10.645439,12.627741,9.657719,10.048691,10.655728,7.8091707,2.6956558,1.3615463,6.3790326,15.426285,21.572105,20.906765,12.548861,9.89436,18.132229,39.687187,64.23274,68.69463,34.532516,14.068168,9.619993,14.325387,12.120162,11.163307,12.257345,12.867812,12.542002,12.912396,10.652299,9.088407,9.2153015,9.914937,7.98065,7.514226,7.3358874,6.451054,5.645101,7.4799304,9.407358,11.910957,15.7795315,20.656404,25.056566,46.477768,43.31912,33.877464,27.594461,25.035988,22.817045,29.223515,38.07871,42.8184,36.5011,24.696459,15.673215,10.765475,10.803201,16.12935,15.988737,13.238208,11.900668,13.642899,17.751545,10.161868,6.3447366,5.0826488,5.161529,5.3878818,16.756964,14.0750265,6.7940125,4.2355404,15.54632,17.422304,11.89038,7.4524937,7.48336,10.199594,19.222837,18.646667,11.14273,6.0395036,19.349733,9.3079,5.871454,5.1821065,5.456474,6.9963584,7.7920227,8.820899,7.8537555,6.327589,9.3764925,15.6526375,12.130451,8.128122,8.742019,14.843254,18.468328,30.969175,28.410702,10.998687,3.0523329,22.573545,16.942162,8.303031,5.871454,5.936616,8.182996,11.688034,14.020154,13.176475,7.5690994,10.679735,15.6697855,14.2362175,7.0306544,3.642222,5.2335505,7.431916,10.408798,11.698323,6.186976,3.40901,2.8054025,2.3218307,1.4061309,1.0048691,0.5727411,0.64819205,1.4918705,2.6613598,3.0146074,3.6387923,2.9460156,2.037175,1.6187652,1.9823016,1.3066728,1.7216529,2.294394,2.9288676,4.3692946,4.5990767,5.0346346,4.928317,4.2252517,3.57363,1.903421,2.3664153,3.1723683,3.6868064,4.437886,4.417309,4.3590055,5.3741636,6.543653,4.9077396,4.5922174,2.867135,2.5138876,4.184097,6.4098988,4.5956473,3.8171308,5.0620713,7.2947326,7.4456344,3.8034124,2.3595562,2.435007,2.8396983,1.8485477,1.1180456,0.8848336,1.5158776,2.8122618,3.981751,3.923448,3.4604537,3.5187566,3.9268777,3.3987212,6.327589,5.4839106,3.8137012,2.6613598,1.7422304,1.1214751,0.8162418,0.7510797,0.78194594,0.70649505,0.39097297,0.37039545,0.30866286,0.13032432,0.041155048,0.07888051,0.106317215,0.21263443,0.36696586,0.42183927,0.23321195,0.09945804,0.024007112,0.0,0.0034295875,0.01371835,0.09259886,0.17833854,0.19891608,0.072021335,0.28465575,0.50757897,0.7476501,0.9259886,0.88826317,1.3855534,1.3101025,1.097468,0.8676856,0.4424168,0.19548649,0.06859175,0.048014224,0.082310095,0.08573969,0.36353627,0.4115505,0.42869842,0.6173257,1.1763484,1.6907866,1.1214751,0.6927767,0.89512235,1.4815818,0.8676856,0.8711152,0.7579388,0.39440256,0.25721905,0.15090185,0.23664154,0.4355576,0.6790583,0.90198153,1.0837497,0.72021335,0.6859175,1.1317638,1.5021594,1.430138,1.0254467,0.6276145,0.38754338,0.26064864,0.2503599,0.28808534,0.2777966,0.20577525,0.14404267,0.22978236,0.16462019,0.09259886,0.1371835,0.40126175,0.274367,0.28808534,0.33609957,0.5761707,1.4335675,0.7476501,0.2777966,0.07545093,0.1097468,0.25378948,0.11317638,0.16804978,0.64133286,1.2072148,0.9774324,0.4115505,0.15433143,0.07545093,0.06516216,0.05144381,0.058302987,0.034295876,0.017147938,0.01371835,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.030866288,0.017147938,0.0034295875,0.006859175,0.006859175,0.0034295875,0.01371835,0.01371835,0.030866288,0.044584636,0.037725464,0.006859175,0.017147938,0.024007112,0.024007112,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.006859175,0.034295876,0.1097468,0.26407823,0.58302987,0.7133542,0.6173257,0.39783216,0.2777966,0.32238123,0.24350071,0.14061308,0.07888051,0.082310095,0.09945804,0.14747226,0.16462019,0.1371835,0.09945804,0.1371835,0.14061308,0.15776102,0.22292319,0.3566771,0.34638834,0.28465575,0.28122616,0.3841138,0.5796003,0.805953,0.91912943,1.1249046,1.4438564,1.6942163,1.4404267,1.1763484,1.1420527,1.2998136,1.3409687,1.0666018,1.0288762,1.1214751,1.1592005,0.86082643,1.3066728,1.4198492,1.2689474,1.0323058,0.9945804,1.0323058,1.2037852,1.214074,1.0220171,0.84367853,1.0666018,1.2380811,1.3101025,1.3169615,1.3409687,1.5261664,1.5570327,1.5570327,1.4918705,1.1454822,0.89512235,0.8162418,0.7613684,0.71678376,0.8093826,1.0425946,1.0460242,1.0220171,1.0151579,0.91569984,0.7682276,0.7888051,0.8711152,0.7990939,0.2709374,0.25378948,0.32924038,0.3841138,0.3841138,0.36353627,0.3806842,0.39783216,0.5007198,0.65505123,0.7305021,0.67219913,0.65162164,0.69963586,0.8025235,0.8711152,0.7442205,0.6893471,0.6859175,0.7305021,0.86082643,0.90198153,0.90541106,0.94656616,1.0357354,1.1146159,1.2689474,1.546744,1.7490896,1.8485477,1.9720128,2.0337453,2.1229146,2.1572106,2.1846473,2.4075704,2.352697,2.2566686,2.136633,2.0406046,2.0440342,1.9720128,1.8691251,1.7559488,1.6530612,1.5810398,1.4129901,1.2586586,1.1454822,1.1008976,1.1866373,1.2895249,1.3821237,1.4678634,1.5913286,1.8348293,1.9239986,1.7388009,1.5261664,1.4198492,1.4404267,1.3478279,1.3443983,1.2963841,1.1934965,1.1489118,1.2037852,1.0871792,1.0185875,0.99801,0.8093826,0.5590228,0.38754338,0.2777966,0.2194936,0.20920484,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.006859175,0.05144381,0.12689474,0.21263443,0.28808534,0.31209245,0.29151493,0.26064864,0.24350071,0.25721905,0.25378948,0.23664154,0.25721905,0.36696586,0.6036074,0.97400284,1.920569,2.8019729,3.3232703,3.5016088,3.758828,5.8371577,8.7317295,11.382801,12.668896,14.860402,14.479718,13.797231,16.341984,26.898254,34.08667,32.51592,23.19087,11.087856,5.137522,3.9440255,3.1620796,2.750529,2.4212887,1.6256244,1.2003556,1.2312219,1.488441,1.6770682,1.4438564,1.2037852,1.1763484,1.0528834,0.8196714,0.77165717,0.6756287,0.58645946,0.51100856,0.4424168,0.36353627,0.39783216,0.4355576,0.45613512,0.41840968,0.29151493,0.28465575,0.29494452,0.37039545,0.490431,0.5658819,0.44927597,0.47671264,0.5418748,0.5555932,0.44927597,0.4938606,0.5041494,0.48700142,0.490431,0.5796003,0.7476501,0.94656616,1.0528834,1.0631721,1.0871792,1.2586586,1.4644338,1.546744,1.920569,3.5804894,2.8156912,4.180667,8.255017,14.860402,23.046827,29.467016,26.232914,24.500973,30.18723,43.950165,49.938225,46.254845,39.546574,32.296425,22.813616,14.21564,11.101575,13.361672,17.741257,17.87501,10.151579,6.358455,5.377593,6.23156,8.080108,9.297611,12.271064,14.040731,16.986746,28.829113,40.5,43.65865,38.4251,29.954018,28.444998,21.356041,14.843254,20.656404,34.59768,36.545685,32.807434,18.091074,10.360784,13.80409,18.807858,19.675543,13.54687,10.943813,14.730078,20.080235,15.350834,11.396519,9.619993,12.600305,24.075705,31.915741,22.717587,9.966381,2.6373527,5.178677,4.996909,5.8543057,7.7268605,8.477941,3.841138,4.1943855,5.1821065,5.3570156,5.610805,9.201583,8.594546,6.090947,5.5490727,9.06097,16.945591,13.7938,7.9189177,4.3692946,4.945465,8.189855,11.2421875,14.030442,12.312219,6.9517736,3.9508848,7.870903,10.203023,10.950673,9.668007,5.453044,2.7882545,9.338767,15.265094,16.259674,13.577737,14.29795,10.14472,8.196714,8.735159,5.2438393,4.7499785,7.058091,8.9100685,8.594546,5.953764,5.3673043,12.912396,14.764374,8.255017,1.8862731,6.4064693,12.2093315,14.829536,15.309678,20.186552,22.494663,19.86417,31.226395,52.438393,56.289818,25.351511,10.316199,7.874333,11.180455,9.863494,10.916377,12.363663,11.513125,9.122703,9.424506,8.364764,7.500508,7.431916,7.764586,7.0889573,9.057541,9.585697,8.354475,6.989499,9.071259,10.710602,12.120162,15.316538,22.422644,35.67457,54.979717,49.89364,36.610847,26.212337,24.662163,35.846046,55.861122,82.14548,99.68439,81.01714,43.281395,23.19773,14.198492,11.201033,10.6145735,12.902108,13.066729,14.973578,18.972477,21.908205,9.328478,7.034084,8.296172,8.399059,4.650521,22.892496,19.637817,9.640571,6.6293926,23.310905,15.484588,10.659158,8.594546,8.570539,9.373062,13.258785,11.177026,8.632272,11.362224,25.327503,8.381912,3.8205605,5.874883,9.561689,10.659158,11.348505,9.342196,7.3393173,7.4799304,11.369082,13.821238,8.584257,6.2418494,10.460241,17.984756,17.154797,29.158352,30.92116,19.432043,11.756626,23.259462,16.760393,7.64798,3.4055803,3.5942078,5.501058,6.725421,9.31133,13.663476,18.560926,15.63206,15.436573,12.195613,6.5985265,5.8165803,8.790032,10.618003,11.763485,11.705182,8.947794,8.001227,6.2555676,4.290414,2.7745364,2.4590142,1.1111864,0.64133286,1.2792361,2.6956558,3.974892,4.3624353,3.625074,2.287535,1.1351935,1.1934965,0.9294182,1.2072148,1.5673214,2.0303159,3.117495,4.07435,4.8185706,5.0895076,5.003768,5.079219,3.0214665,3.333559,3.7965534,3.5804894,3.223812,3.5873485,4.32128,5.6656785,6.8283086,6.0086374,3.7382503,2.5619018,3.0660512,4.5030484,4.791134,4.057202,4.1635194,5.470192,7.085528,6.8728933,4.5270553,3.3712845,3.3061223,3.4021509,1.9068506,1.371835,1.0425946,1.2380811,2.0817597,3.4776018,4.057202,4.5270553,5.0929375,5.164959,3.3472774,5.7274113,5.1066556,3.5050385,2.2463799,1.9754424,1.5193073,0.881404,0.5796003,0.6344737,0.5761707,0.39097297,0.39097297,0.33952916,0.18519773,0.06516216,0.12003556,0.12003556,0.14404267,0.2194936,0.31552204,0.24350071,0.14061308,0.048014224,0.0,0.0,0.020577524,0.09259886,0.17833854,0.2194936,0.14747226,0.1920569,0.33609957,0.61046654,0.8093826,0.48700142,0.90884066,0.8711152,0.7305021,0.61046654,0.39783216,0.216064,0.09259886,0.05144381,0.06859175,0.082310095,0.19548649,0.26750782,0.5144381,0.84367853,0.84367853,1.2929544,0.89512235,0.7133542,1.0117283,1.2758065,0.75450927,0.6173257,0.4972902,0.29151493,0.18176813,0.1371835,0.19891608,0.4046913,0.72707254,1.0837497,1.7113642,1.3958421,1.039165,1.1043272,1.6221949,1.7525192,1.4644338,0.90541106,0.3806842,0.34638834,0.5590228,0.6824879,0.5796003,0.31209245,0.1371835,0.42869842,0.33266997,0.20234565,0.31895164,0.91912943,0.5453044,0.4081209,0.31895164,0.40126175,1.0940384,0.6824879,0.26750782,0.0548734,0.06859175,0.14747226,0.1097468,0.23664154,0.6001778,0.97057325,0.83338976,0.41498008,0.19891608,0.1371835,0.15433143,0.12689474,0.09602845,0.061732575,0.037725464,0.030866288,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.030866288,0.024007112,0.0034295875,0.010288762,0.010288762,0.0034295875,0.01371835,0.006859175,0.024007112,0.044584636,0.048014224,0.017147938,0.006859175,0.01371835,0.01371835,0.006859175,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.15433143,0.39440256,0.66533995,0.7133542,0.6173257,0.4389872,0.2194936,0.18519773,0.12003556,0.06516216,0.041155048,0.041155048,0.05144381,0.07545093,0.09259886,0.09259886,0.082310095,0.082310095,0.09602845,0.12346515,0.18519773,0.30866286,0.22635277,0.16119061,0.15433143,0.2503599,0.48357183,0.72707254,1.0425946,1.3581166,1.6153357,1.7593783,1.7662375,1.6187652,1.3924125,1.2277923,1.3306799,1.0117283,1.155771,1.4472859,1.6359133,1.5433143,1.6016173,1.488441,1.3238207,1.138623,0.8745448,0.9602845,1.0631721,1.0940384,1.0460242,0.9877212,1.155771,1.3546871,1.3958421,1.3101025,1.3066728,1.4438564,1.5398848,1.6221949,1.6221949,1.3855534,1.0768905,0.8779744,0.7305021,0.6310441,0.64819205,0.78194594,0.82996017,0.90198153,0.96714365,0.8505377,0.7510797,0.78537554,0.8745448,0.8711152,0.5590228,0.22978236,0.18519773,0.20577525,0.19548649,0.17833854,0.2194936,0.2709374,0.34295875,0.45270553,0.6207553,0.6241849,0.64819205,0.72021335,0.7990939,0.7682276,0.66876954,0.66533995,0.69963586,0.7613684,0.8779744,0.91912943,0.94999576,1.0597426,1.255229,1.471293,1.5673214,1.7388009,1.9274281,2.0920484,2.1880767,2.0646117,2.1263442,2.2120838,2.2909644,2.4795918,2.335549,2.1640697,2.037175,1.9651536,1.920569,1.7971039,1.6530612,1.5536032,1.5124481,1.5021594,1.4678634,1.4198492,1.3684053,1.3203912,1.2895249,1.4095604,1.3924125,1.4232788,1.5776103,1.8039631,1.8931323,1.7799559,1.6290541,1.5570327,1.6324836,1.6599203,1.5433143,1.3992717,1.3169615,1.3409687,1.4129901,1.3821237,1.313532,1.196926,0.94999576,0.7407909,0.6207553,0.52472687,0.4355576,0.36696586,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.0034295875,0.020577524,0.061732575,0.116605975,0.16462019,0.19548649,0.34981793,0.41498008,0.33952916,0.22635277,0.23321195,0.22978236,0.2469303,0.31895164,0.48357183,0.8676856,1.9548649,2.9974594,3.6765177,4.098357,3.7519686,5.48734,8.117833,10.710602,12.614022,16.143068,15.13134,13.906977,16.088194,24.579853,30.862858,30.482174,22.758743,11.571428,5.346727,3.9954693,3.1072063,2.726522,2.5173173,1.7799559,1.1420527,1.1249046,1.371835,1.5398848,1.2963841,1.0837497,1.1043272,1.1008976,0.9602845,0.7339317,0.61389613,0.6036074,0.5624523,0.45613512,0.36353627,0.4424168,0.432128,0.39783216,0.3806842,0.41840968,0.4629943,0.4355576,0.5041494,0.66191036,0.75450927,0.5418748,0.58645946,0.58988905,0.48014224,0.3806842,0.53158605,0.53844523,0.548734,0.6173257,0.7133542,1.0288762,1.2758065,1.3203912,1.2243627,1.2209331,1.5193073,1.6942163,1.7593783,2.0234566,3.0969174,3.5942078,6.2658563,10.247607,15.107333,20.879328,26.061436,25.636166,29.26124,41.41913,61.423912,61.447918,49.900497,35.715725,23.712168,14.589465,10.659158,9.719451,12.435684,16.53404,16.79469,12.939834,9.822338,7.4456344,6.327589,7.5210853,13.629181,16.11906,17.339994,19.404606,24.216316,30.845709,31.867727,26.908543,18.595222,12.524854,8.844906,10.659158,18.097933,27.639046,32.1078,31.065203,14.977009,6.6636887,10.549411,12.644889,14.928994,10.381361,6.869464,6.8728933,7.500508,8.457363,11.06042,9.047252,5.329579,12.0138445,19.744135,14.754086,6.416758,0.85739684,0.9259886,0.6036074,0.89169276,2.9185789,5.3673043,4.48933,3.5873485,3.6627994,4.1120753,4.8254294,6.217842,5.8543057,4.4104495,5.5319247,9.458802,13.035862,8.824328,5.3330083,4.9351764,6.108095,3.474172,5.4496145,10.429376,11.571428,8.134981,5.4770513,7.31531,8.704293,9.084977,7.6857057,3.5359046,2.3149714,8.64599,12.583157,11.008976,7.613684,9.112414,8.608265,7.8091707,7.1884155,5.994919,6.1801167,6.948344,6.2898636,4.245829,2.901431,4.057202,11.9040985,15.71437,12.010415,4.540774,7.2707253,11.166737,10.875222,9.997248,21.091963,28.883986,22.463799,22.504953,31.555634,34.01122,15.275383,6.8591747,5.4839106,7.2878733,7.829748,10.377932,10.168727,8.203573,6.39961,7.579388,6.756287,7.689135,8.690575,8.676856,7.174697,9.942374,10.360784,9.040393,8.114404,11.22161,12.6929035,13.13532,15.385129,22.769032,39.117874,48.19599,41.199635,30.42044,23.338343,22.642136,39.31679,58.855152,83.544754,100.89846,83.671646,42.866413,22.727877,14.520873,11.166737,7.2707253,11.231899,12.5145645,15.697222,20.749004,23.03311,9.187865,11.784062,15.121051,12.082437,4.1326528,20.989075,18.903887,10.655728,8.038953,21.877338,11.664027,7.4627824,6.5024977,6.4373355,5.360445,7.257007,7.2467184,8.97523,13.776653,20.663265,5.936616,2.3904223,7.7783046,14.819247,11.190743,11.074138,9.702303,8.388771,8.275595,10.329918,10.515115,6.355026,5.888602,12.291641,23.880217,14.490007,20.94792,28.18435,27.553307,16.818697,17.484037,11.873232,5.7308407,2.6545007,4.0880685,7.6651278,7.9429245,7.349606,9.177576,17.61436,13.54687,11.540562,8.824328,6.4716315,9.403929,15.769243,16.719238,14.579176,11.190743,7.9292064,7.4970784,6.866034,5.3570156,3.3678548,2.3561265,1.3169615,0.7888051,1.2003556,2.4761622,4.0366244,4.2869844,3.590778,2.2258022,0.91227025,0.8162418,1.1729189,1.5604624,1.7593783,1.7936742,1.9308578,2.9391565,3.8548563,4.5510626,4.955754,5.0414934,3.7622573,4.0880685,4.4927597,4.3349986,3.8445675,4.190956,4.6676683,5.4496145,6.2864337,6.495639,4.513337,3.7965534,3.875434,3.9303071,2.8088322,2.702515,3.340418,4.763697,6.0703697,5.4324665,3.9783216,3.525616,3.8891523,3.9954693,1.8588364,1.4987297,1.8073926,1.7113642,1.587899,3.2958336,4.6402316,6.166398,6.90033,6.2555676,4.0434837,3.7313912,5.6142344,5.209543,2.6064866,2.4795918,1.7422304,0.88826317,0.4424168,0.45270553,0.47328308,0.41498008,0.41840968,0.39097297,0.28808534,0.09602845,0.13032432,0.13032432,0.12346515,0.15090185,0.23664154,0.22635277,0.16119061,0.07545093,0.010288762,0.0,0.020577524,0.072021335,0.1371835,0.19891608,0.26407823,0.16462019,0.28465575,0.6756287,1.0357354,0.72707254,0.91227025,0.66533995,0.4046913,0.3018037,0.29151493,0.20920484,0.116605975,0.06859175,0.072021335,0.08916927,0.09259886,0.25721905,0.47671264,0.59331864,0.40126175,1.1626302,0.7922347,0.53501564,0.6893471,0.6344737,0.5624523,0.34295875,0.18862732,0.14404267,0.072021335,0.14061308,0.15433143,0.32238123,0.65505123,0.9911508,2.253239,2.2463799,1.670209,1.3101025,2.0028791,2.1572106,1.7902447,1.2380811,0.7510797,0.52472687,0.77508676,0.9945804,0.8265306,0.36010668,0.14404267,0.61046654,0.52472687,0.37725464,0.48357183,0.9602845,1.4267083,0.90198153,0.34295875,0.216064,0.48357183,0.52472687,0.3806842,0.19548649,0.06859175,0.048014224,0.072021335,0.19891608,0.39783216,0.58645946,0.6310441,0.33952916,0.2469303,0.20577525,0.16119061,0.12689474,0.09602845,0.07545093,0.061732575,0.048014224,0.041155048,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.006859175,0.01371835,0.020577524,0.024007112,0.0034295875,0.006859175,0.006859175,0.0034295875,0.01371835,0.006859175,0.020577524,0.034295876,0.037725464,0.024007112,0.010288762,0.010288762,0.010288762,0.006859175,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.044584636,0.18519773,0.52815646,0.6756287,0.7099246,0.70649505,0.607037,0.23321195,0.14747226,0.106317215,0.082310095,0.05144381,0.01371835,0.017147938,0.0274367,0.041155048,0.0548734,0.06516216,0.048014224,0.061732575,0.08573969,0.116605975,0.18176813,0.12003556,0.07888051,0.07888051,0.15090185,0.32924038,0.67219913,1.1592005,1.471293,1.5604624,1.6187652,1.862266,1.9582944,1.7147937,1.3615463,1.5638919,1.1489118,1.1351935,1.5021594,1.978872,2.0508933,1.6942163,1.4644338,1.2963841,1.1180456,0.8505377,0.9945804,0.9568549,0.9328478,1.0048691,1.1523414,1.1900668,1.3409687,1.3992717,1.3203912,1.2449403,1.3203912,1.371835,1.3992717,1.3855534,1.2758065,1.0425946,0.89855194,0.7956643,0.70306545,0.6173257,0.6824879,0.764798,0.8505377,0.88826317,0.78537554,0.8162418,0.85396725,0.89512235,0.8779744,0.69963586,0.28808534,0.16119061,0.15090185,0.15090185,0.12346515,0.1371835,0.17833854,0.20920484,0.26064864,0.42869842,0.490431,0.6036074,0.69963586,0.72021335,0.6276145,0.5761707,0.6276145,0.72364295,0.8093826,0.85396725,0.9602845,1.0323058,1.1866373,1.4438564,1.7388009,1.9137098,2.095478,2.3149714,2.4624438,2.2978237,2.0131679,2.0028791,2.1503513,2.3081124,2.2841053,2.1194851,1.9342873,1.8245405,1.7971039,1.7662375,1.6016173,1.5090185,1.4987297,1.5261664,1.4815818,1.5124481,1.5981878,1.5981878,1.5055889,1.4335675,1.4747226,1.4267083,1.4610043,1.5947582,1.7182233,1.7730967,1.6804979,1.5536032,1.4918705,1.5844694,1.7147937,1.7147937,1.6324836,1.5193073,1.4438564,1.4815818,1.5227368,1.4918705,1.3306799,1.0151579,0.922559,0.82996017,0.7373613,0.6310441,0.52472687,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.06859175,0.07545093,0.09602845,0.4046913,0.5590228,0.42869842,0.20920484,0.24350071,0.24350071,0.2469303,0.274367,0.29837412,0.823101,1.8519772,2.9117198,3.8102717,4.6676683,3.8034124,4.8322887,6.776865,9.297611,12.6757555,16.324837,15.141628,13.7526455,15.477728,22.340332,28.252941,27.717926,21.287449,12.103014,5.892031,4.3041325,3.2958336,2.7093742,2.2738166,1.587899,1.08032,1.0700313,1.2072148,1.2689474,1.138623,1.0906088,1.2723769,1.3615463,1.2209331,0.9328478,0.6927767,0.64133286,0.5693115,0.42183927,0.31895164,0.41498008,0.35324752,0.28808534,0.36010668,0.6756287,0.7956643,0.70649505,0.71678376,0.881404,0.9945804,0.7579388,0.7682276,0.69963586,0.5178677,0.4629943,0.61389613,0.59674823,0.6859175,0.9328478,1.1694894,1.5536032,1.7936742,1.7696671,1.605047,1.6496316,2.0714707,2.3664153,2.6064866,3.0386145,4.064061,6.464772,10.113853,12.8197975,15.0250225,19.805868,22.515242,25.711617,34.75887,51.251755,73.0022,63.882927,49.314037,34.659412,22.638706,13.310229,11.513125,9.836057,11.509696,15.244516,15.261664,16.403717,14.102464,10.155008,7.14726,8.450503,17.689812,17.027903,17.583494,19.644676,12.655178,13.094165,15.6252,17.528622,17.463459,15.46744,13.622321,12.843805,14.174485,17.662374,22.371199,20.364891,9.523964,3.642222,5.223262,5.4839106,6.0326443,3.8685746,1.9754424,1.2106444,0.29151493,3.0454736,9.589127,9.297611,2.9391565,2.668219,5.796003,4.537344,2.0028791,0.21263443,0.08573969,0.32924038,0.50757897,1.937717,3.8720043,3.4776018,3.4638834,3.957744,4.396731,4.3487167,3.508468,3.192946,2.7779658,4.938606,8.182996,6.869464,2.9151495,3.9611735,6.9963584,8.268735,3.2958336,3.542764,6.9963584,8.495089,6.8969,5.1100855,5.086078,6.468202,7.4284863,6.4304767,2.218943,1.3341095,5.686256,8.597976,8.004657,6.4579134,5.5593615,6.0497923,5.98463,5.6245236,7.4456344,8.56025,7.250148,4.7499785,2.452155,1.8965619,4.5099077,6.4544835,8.97866,10.998687,9.108984,9.098696,11.499407,10.134431,7.4010496,14.249936,25.114868,23.516682,18.571217,15.676644,16.53747,10.39508,5.4907694,3.806842,5.0174866,6.4990683,9.709162,6.8214493,4.623084,5.7308407,8.56368,6.7459984,9.071259,11.547421,11.780633,8.961512,11.273054,10.377932,8.261876,7.4044795,10.765475,11.893809,11.760056,14.003006,20.423193,31.01033,31.030907,22.991955,17.017612,15.724659,14.225929,28.530739,38.016975,44.92074,47.938774,42.23537,22.498095,14.836395,12.319078,10.268185,6.245279,9.170717,9.342196,12.079007,17.329706,19.661825,8.553391,15.29253,18.643238,12.247057,4.636802,13.437123,11.763485,8.330468,8.855195,16.084764,9.379922,4.588788,3.4055803,4.4104495,3.0557625,7.233,10.940384,12.000127,10.88894,10.7586155,5.7411294,5.1683884,11.170166,17.182234,7.9600725,7.284444,9.102125,9.325048,7.3839016,6.2212715,7.040943,6.6636887,7.795452,13.262215,26.02371,12.05843,12.812939,22.662714,29.477304,14.616901,10.388221,6.5367937,5.1066556,6.279575,8.39563,11.859513,12.6586075,9.06097,4.6676683,8.412778,10.100135,8.841476,6.9552035,7.0786686,12.1921835,20.237995,21.163984,18.262554,13.207341,6.029215,4.2698364,5.2987127,5.130663,3.083199,1.7593783,1.7250825,1.5364552,1.762808,2.4041407,2.8739944,2.9254382,2.5138876,1.6427724,0.8128122,1.0151579,1.6907866,2.3321195,2.551613,2.2669573,1.7113642,1.8897027,2.5996273,3.426158,3.9063,3.542764,3.8034124,4.413879,4.8151407,4.9523244,5.2747054,5.7136927,5.3981705,5.271276,5.7891436,6.910619,6.464772,5.5250654,4.139512,2.644212,1.6496316,1.6496316,2.0440342,3.2889743,4.698535,4.448175,2.8637056,2.9803114,4.0880685,4.5990767,2.0577524,1.5536032,2.609916,2.435007,1.4061309,3.059192,5.020916,7.1849856,7.606825,6.3447366,5.435896,2.8054025,6.334448,6.999788,3.7451096,3.5050385,1.7765263,0.7990939,0.41498008,0.41840968,0.53501564,0.51100856,0.5521636,0.6036074,0.53844523,0.15433143,0.12003556,0.12003556,0.13032432,0.16462019,0.24007112,0.22292319,0.17490897,0.09945804,0.0274367,0.0,0.01371835,0.048014224,0.09602845,0.20234565,0.432128,0.21263443,0.4046913,0.91569984,1.4061309,1.2860953,1.2072148,0.7579388,0.4046913,0.28808534,0.24350071,0.216064,0.16804978,0.13032432,0.1097468,0.09945804,0.08573969,0.28465575,0.274367,0.11317638,0.33266997,1.4953002,0.9294182,0.2469303,0.072021335,0.041155048,0.42183927,0.23664154,0.05144381,0.048014224,0.01371835,0.19891608,0.13032432,0.23664154,0.58988905,0.8848336,2.4487255,2.8534167,2.4727325,1.9891608,2.4212887,2.4555845,2.0749004,1.7147937,1.4678634,1.0494537,0.9362774,1.1214751,0.97057325,0.45613512,0.16119061,0.65162164,0.6036074,0.48357183,0.47328308,0.47671264,2.1572106,1.3409687,0.41840968,0.26064864,0.22635277,0.42183927,0.5007198,0.36353627,0.1097468,0.05144381,0.048014224,0.08573969,0.15433143,0.28465575,0.53158605,0.3018037,0.31209245,0.274367,0.1371835,0.082310095,0.10288762,0.08916927,0.06859175,0.0548734,0.034295876,0.0274367,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.0274367,0.017147938,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.048014224,0.20920484,0.6036074,0.58645946,0.65848076,0.83681935,0.8848336,0.31552204,0.22978236,0.22635277,0.20920484,0.14061308,0.041155048,0.010288762,0.006859175,0.01371835,0.024007112,0.05144381,0.05144381,0.05144381,0.05144381,0.048014224,0.020577524,0.020577524,0.030866288,0.06516216,0.13032432,0.23321195,0.61389613,1.1420527,1.4369972,1.488441,1.6393428,1.862266,2.0989075,1.9651536,1.6290541,1.8176813,1.313532,0.9774324,1.2380811,1.8313997,1.8005334,1.3581166,1.2792361,1.1489118,0.89855194,0.8162418,1.0048691,0.922559,0.83681935,0.89855194,1.1283343,1.0734608,1.1283343,1.2175035,1.2449403,1.1146159,1.1523414,1.097468,1.0082988,0.9431366,0.9362774,0.8745448,0.881404,0.89855194,0.881404,0.8128122,0.89512235,0.939707,0.90541106,0.8093826,0.7339317,0.8676856,0.94656616,0.97057325,0.90198153,0.65162164,0.37039545,0.216064,0.17147937,0.18519773,0.15776102,0.12689474,0.13375391,0.15776102,0.19891608,0.2777966,0.33609957,0.52815646,0.64476246,0.6241849,0.52472687,0.5041494,0.5761707,0.6962063,0.7956643,0.7888051,1.0597426,1.214074,1.4027013,1.6667795,1.9308578,2.2223728,2.411,2.5550427,2.5413244,2.1023371,1.8588364,1.7936742,1.9582944,2.1640697,1.961724,1.8759843,1.7422304,1.6427724,1.6221949,1.6667795,1.5604624,1.605047,1.7010754,1.7456601,1.605047,1.5604624,1.6804979,1.7010754,1.6016173,1.611906,1.4918705,1.4815818,1.5501735,1.6393428,1.670209,1.6633499,1.5158776,1.3821237,1.3375391,1.3958421,1.5330256,1.762808,1.8313997,1.6907866,1.4815818,1.4335675,1.471293,1.4987297,1.4369972,1.1866373,1.1420527,1.0048691,0.8745448,0.78194594,0.7099246,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.0274367,0.01371835,0.01371835,0.034295876,0.06859175,0.13375391,0.24350071,0.28122616,0.23664154,0.16804978,0.12689474,0.15090185,0.8128122,1.5638919,2.428148,3.3644254,4.2423997,3.2272418,2.9391565,4.73969,8.429926,12.236768,14.068168,13.831526,13.37882,14.990726,21.3629,26.1849,24.497543,18.660385,11.190743,4.746549,3.782835,2.9734523,2.4418662,2.0508933,1.4027013,1.2209331,1.3032433,1.4369972,1.4541451,1.2346514,0.9431366,0.7510797,0.5727411,0.44584638,0.5178677,0.6790583,0.7339317,0.7099246,0.61389613,0.4424168,0.42869842,0.42869842,0.42869842,0.45613512,0.5658819,0.58988905,0.6962063,0.7682276,0.7888051,0.823101,0.8128122,0.7888051,0.7956643,0.8162418,0.7922347,0.85396725,0.88826317,1.1934965,1.7422304,2.1812177,1.7662375,1.8554068,1.9582944,2.1023371,2.8225505,3.7005248,4.506478,5.2506986,6.6876955,10.31277,13.7697935,14.750656,14.757515,16.901007,25.910534,29.984882,34.43992,41.957573,53.494705,68.25222,54.44813,41.840965,33.002922,26.93598,19.071936,11.88352,9.966381,10.707172,11.893809,11.732618,15.199932,14.586036,11.598865,10.220171,16.678083,18.924463,17.662374,17.864721,20.515793,22.628418,25.8488,25.282919,25.18003,25.159454,20.217419,19.277712,12.926115,9.033533,9.966381,12.603734,12.202472,6.4716315,3.74168,5.0929375,4.3487167,2.702515,1.7936742,1.0014396,0.25721905,0.061732575,2.0028791,6.1766872,6.4579134,3.1449318,2.959734,3.8514268,2.2600982,0.6790583,0.14747226,0.24350071,1.3684053,2.0063086,2.5481834,2.8911421,2.4247184,2.4624438,3.1209247,3.6353626,3.5839188,2.8980014,1.8485477,2.037175,3.7519686,5.113515,2.061182,2.2052248,3.5873485,6.800872,9.290752,5.3707337,3.7725463,5.0277753,6.310441,6.060081,3.998899,3.74168,4.6848164,5.435896,4.9180284,2.3664153,1.2037852,3.433017,5.2781353,5.446185,5.127233,5.518206,4.763697,5.06893,6.677407,7.874333,7.3358874,5.7822843,4.5201964,4.400161,5.826869,5.658819,3.3541365,3.1517909,6.9380555,14.2362175,13.114742,10.772334,11.084427,12.857523,9.8429165,17.580065,14.802099,11.821788,11.763485,10.545981,6.1492505,5.0140567,6.526505,8.378482,6.560801,9.088407,6.4133286,5.079219,7.3290286,11.1393,10.4533825,11.585147,11.931535,11.06042,10.679735,13.612033,10.700313,6.468202,3.7313912,3.5873485,4.8425775,6.3035817,8.7145815,11.821788,14.359683,15.385129,11.173596,6.5950966,5.3501563,9.962952,27.834532,37.025826,38.603436,33.10238,20.556948,8.834618,11.856084,14.4145565,11.434244,7.98065,6.492209,4.012617,4.513337,7.7131424,9.078118,4.756838,8.080108,10.05898,7.9943686,5.4770513,13.790371,9.945804,7.2467184,11.653738,21.77445,13.046151,7.191845,6.509357,8.64599,6.6053853,8.546532,14.232788,12.590015,5.435896,7.4627824,13.330807,15.505165,14.212211,10.449953,5.9812007,6.701414,5.4736214,4.07435,3.782835,5.3570156,5.7822843,8.186425,12.373952,17.000465,19.576086,12.607163,14.682064,19.857311,20.989075,9.736599,7.6342616,5.919468,8.697433,13.471419,11.153018,8.601405,8.735159,9.496528,11.478829,17.899017,23.499533,19.143957,14.315098,12.617453,11.763485,11.667457,14.7369375,18.28313,18.883308,12.3911,11.204462,7.5588107,4.1360826,2.9220085,5.2026844,4.3007026,3.415869,2.5241764,1.9342873,2.287535,2.3972816,1.9411465,1.1283343,0.52815646,1.0528834,1.2963841,1.605047,2.0920484,2.49331,2.1503513,1.920569,2.2292318,2.5927682,2.9700227,3.7382503,3.9097297,4.7499785,4.6093655,3.7965534,4.5784993,6.495639,6.632822,5.926327,6.1149545,9.764035,8.9100685,5.9434752,3.0489032,1.3101025,0.6859175,1.8108221,2.959734,3.5393343,3.923448,5.4633327,3.3369887,3.3301294,4.746549,5.778855,3.508468,2.020027,2.0234566,1.8828435,1.4575747,2.1057668,3.9611735,4.945465,4.8734436,4.530485,5.693115,4.4584637,3.2615378,3.9646032,5.885172,5.813151,2.0063086,0.65848076,0.5555932,0.7888051,0.77851635,0.66876954,0.90541106,1.1626302,1.0837497,0.29151493,0.12003556,0.10288762,0.14747226,0.1920569,0.22978236,0.29151493,0.22292319,0.12003556,0.037725464,0.0,0.01371835,0.024007112,0.08573969,0.26407823,0.64133286,0.5178677,0.66191036,1.1214751,1.5776103,1.3581166,1.0151579,0.94999576,0.90541106,0.72021335,0.30523327,0.26750782,0.26750782,0.26750782,0.22292319,0.07545093,0.05144381,0.09945804,0.12346515,0.30866286,1.1146159,1.8965619,1.138623,0.36353627,0.14061308,0.09259886,0.07888051,0.14061308,0.20234565,0.19548649,0.061732575,0.25721905,0.16804978,0.22292319,0.70306545,1.7388009,2.4247184,3.0043187,3.2443898,2.9460156,1.9685832,1.7113642,2.287535,2.3801336,1.978872,2.3801336,1.5261664,1.1660597,1.0631721,0.881404,0.19891608,0.5521636,0.5590228,0.41840968,0.23321195,0.0,0.7339317,0.45613512,0.36010668,0.6036074,0.33609957,0.14061308,0.09945804,0.08916927,0.07545093,0.1371835,0.12346515,0.12346515,0.15090185,0.2503599,0.45613512,0.3841138,0.37382504,0.4115505,0.4115505,0.22978236,0.29151493,0.15776102,0.061732575,0.058302987,0.044584636,0.058302987,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0274367,0.041155048,0.0274367,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09259886,0.26407823,0.5796003,0.5418748,0.6241849,0.90198153,1.0460242,0.34981793,0.32581082,0.42869842,0.4664239,0.3566771,0.1371835,0.041155048,0.006859175,0.01371835,0.041155048,0.07545093,0.07545093,0.06859175,0.072021335,0.082310095,0.044584636,0.044584636,0.0548734,0.07888051,0.13375391,0.24350071,0.40126175,0.90884066,1.3375391,1.5913286,1.9068506,1.9068506,1.8897027,1.6770682,1.2586586,0.7922347,0.70649505,0.8779744,0.9877212,0.8848336,0.5796003,0.7613684,1.039165,1.039165,0.764798,0.59674823,0.764798,0.881404,0.89855194,0.823101,0.70306545,0.7133542,0.7339317,0.83338976,0.96714365,0.9911508,1.0906088,1.0768905,1.0048691,0.9259886,0.90198153,0.9362774,0.94656616,1.0014396,1.1043272,1.1900668,1.1660597,1.0666018,0.8711152,0.6344737,0.48700142,0.48700142,0.78194594,0.9774324,0.9294182,0.7476501,0.52815646,0.29837412,0.15090185,0.1097468,0.12346515,0.1097468,0.14404267,0.216064,0.29151493,0.29151493,0.4355576,0.58302987,0.61389613,0.51100856,0.36696586,0.41498008,0.5555932,0.6824879,0.77851635,0.89855194,1.4267083,1.6942163,1.8999915,2.1263442,2.335549,2.469303,2.318401,1.9582944,1.5536032,1.3581166,1.5055889,1.4850113,1.5364552,1.6564908,1.6324836,1.7319417,1.8176813,1.8005334,1.7147937,1.7388009,1.9823016,2.037175,1.9685832,1.8245405,1.6187652,1.6770682,1.6290541,1.6839274,1.8554068,1.9514352,1.8416885,1.7696671,1.7456601,1.7422304,1.6942163,1.6084765,1.4953002,1.4267083,1.430138,1.4815818,1.529596,1.4953002,1.4335675,1.4095604,1.4953002,1.4472859,1.4164196,1.4232788,1.4678634,1.5398848,1.3101025,1.1866373,1.1146159,1.1008976,1.2346514,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0034295875,0.01371835,0.05144381,0.1097468,0.17147937,0.18862732,0.29151493,0.2777966,0.16119061,0.16462019,0.6001778,1.039165,1.7593783,2.8534167,4.2286816,3.5290456,2.7299516,4.064061,7.274155,9.637141,11.8115,12.068718,12.343085,14.747226,21.568676,25.317215,23.743034,17.693241,9.815479,4.5613513,3.7725463,3.2203827,2.7230926,2.2120838,1.7216529,1.529596,1.4404267,1.2655178,1.0837497,1.2243627,0.8711152,0.70306545,0.65505123,0.65505123,0.59331864,0.5178677,0.6036074,0.71678376,0.7682276,0.72364295,0.58302987,0.490431,0.45613512,0.45613512,0.42869842,0.4046913,0.50757897,0.6344737,0.7339317,0.7990939,0.91569984,1.1146159,1.2380811,1.2758065,1.3786942,1.4095604,1.3992717,1.4953002,1.6770682,1.7559488,1.7388009,2.177788,3.0866287,4.1326528,4.616225,4.6745276,5.2747054,9.208443,14.5414505,14.610043,13.320518,13.519434,16.352274,22.679861,33.07494,32.65996,36.17186,47.99022,63.666862,69.94987,49.163136,31.830002,24.69303,24.284908,16.914726,11.382801,12.055,13.262215,12.291641,9.39021,12.72034,14.829536,17.137648,19.62753,20.841602,15.734947,12.569438,11.115293,13.077017,22.093403,23.887077,20.262003,17.586924,17.312557,15.971589,12.764925,8.930646,6.2967224,5.675967,6.866034,7.548522,4.870014,3.5290456,4.386442,4.4721823,1.7765263,0.6893471,0.4972902,0.6962063,0.9877212,4.6676683,5.2918534,3.707384,1.9651536,3.3129816,3.2375305,2.153781,1.1626302,0.8265306,1.1592005,2.2429502,2.6579304,2.2566686,1.5981878,1.9754424,1.7182233,1.9239986,2.1297739,2.085189,1.7525192,1.6393428,2.3252604,3.3026927,3.5873485,1.704505,2.2120838,2.843128,4.955754,6.944915,4.2355404,2.1194851,1.7319417,1.8279701,1.7799559,1.5810398,1.9102802,2.4144297,3.1106358,3.3026927,1.5707511,0.75450927,1.6153357,3.4364467,4.945465,4.3452873,5.079219,4.064061,3.625074,4.623084,6.495639,6.835168,5.5902276,5.113515,6.728851,10.72432,8.344186,3.9440255,4.091498,10.22703,18.680964,11.122152,8.886061,9.925226,10.978109,7.582818,6.924337,6.042933,5.5113473,5.504488,5.796003,4.2423997,7.641121,10.463672,10.556271,9.136421,9.702303,7.3873315,10.096705,15.584045,11.444533,9.647429,8.381912,7.73029,7.7748747,8.604835,6.8385973,6.210983,6.5950966,7.040943,5.7822843,7.1952744,10.707172,14.486577,15.570327,9.866923,10.823778,11.986408,12.377381,11.1393,7.5245147,21.486366,29.607628,29.569902,21.829325,9.592556,6.9552035,12.349944,14.164196,10.2236,7.7851634,4.8425775,4.3349986,4.9591837,6.121814,7.966932,6.917478,8.004657,6.608815,4.547633,10.079557,15.05246,8.30646,5.8645945,11.856084,18.526632,10.172156,10.81006,13.725209,14.270514,9.877212,5.5902276,7.133542,8.23444,7.8366075,10.096705,24.11343,19.922474,11.269625,5.826869,5.188966,13.077017,10.803201,6.0566516,3.2992632,3.7691166,3.923448,5.645101,9.054111,12.298501,11.543991,10.960961,22.717587,25.399525,15.645778,8.158989,8.412778,7.4044795,5.8988905,4.7191124,4.7328305,4.976331,5.103226,4.3521466,5.761707,16.163645,18.224829,16.62664,14.918706,14.956431,16.904436,14.79524,17.425734,21.294308,21.263443,10.569988,7.4353456,4.280125,2.959734,4.197815,7.582818,5.672538,3.0523329,1.5638919,1.6599203,2.3732746,2.6613598,2.085189,2.0097382,2.3767042,1.7010754,1.3272504,1.6153357,2.3046827,2.8808534,2.5790498,2.435007,2.2463799,2.3561265,2.8945718,3.7622573,5.2918534,6.0875177,5.2609873,3.7039545,4.1155047,6.8900414,6.90033,6.948344,7.9429245,8.886061,7.250148,5.120374,3.5359046,2.9185789,3.0660512,3.9646032,4.633373,4.3795834,3.4776018,3.1792276,2.1880767,2.836269,4.180667,5.0174866,3.899441,2.3046827,2.294394,2.4624438,2.270387,2.0577524,2.534465,3.806842,3.8788633,3.2512488,4.897451,3.3232703,2.8980014,3.566771,4.1635194,2.4212887,1.1592005,0.61389613,0.9568549,1.5741806,1.0357354,0.7099246,0.7407909,0.8196714,0.7476501,0.42526886,0.22292319,0.12003556,0.09602845,0.1371835,0.25378948,0.274367,0.22635277,0.1371835,0.048014224,0.0,0.0034295875,0.01371835,0.0548734,0.13032432,0.22635277,0.38754338,0.6962063,1.2312219,1.7525192,1.7010754,1.786815,1.4335675,0.99801,0.65848076,0.39097297,0.274367,0.26407823,0.274367,0.2503599,0.16119061,0.09945804,0.116605975,0.14404267,0.4115505,1.4438564,1.6290541,0.9945804,0.47671264,0.34638834,0.18862732,0.06859175,0.044584636,0.05144381,0.06859175,0.1097468,0.14061308,0.14747226,0.16462019,0.2709374,0.6173257,0.8711152,0.9568549,1.2723769,1.903421,2.6167753,1.5090185,1.3684053,1.313532,1.3409687,2.318401,3.4673128,3.2478194,2.5721905,1.7799559,0.6379033,1.7936742,1.9411465,1.4335675,0.70649505,0.26750782,0.34638834,0.34638834,0.28465575,0.17833854,0.06859175,0.037725464,0.13375391,0.31895164,0.4115505,0.09945804,0.23664154,0.25378948,0.24007112,0.25378948,0.32238123,0.2709374,0.29494452,0.33952916,0.32924038,0.15433143,0.13032432,0.2469303,0.22635277,0.061732575,0.020577524,0.024007112,0.0274367,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.020577524,0.0274367,0.017147938,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.07545093,0.22978236,0.5178677,0.5796003,0.6001778,0.65848076,0.66191036,0.32581082,0.37039545,0.5418748,0.7510797,0.8025235,0.4046913,0.14061308,0.030866288,0.01371835,0.0548734,0.15090185,0.2194936,0.18176813,0.14061308,0.116605975,0.06859175,0.06859175,0.07888051,0.11317638,0.16462019,0.19548649,0.4698535,1.0494537,1.5124481,1.7250825,1.8588364,1.9171394,2.0165975,1.6564908,0.9362774,0.548734,0.5212973,0.58988905,0.6173257,0.5521636,0.42183927,0.5761707,1.8313997,2.1091962,1.1420527,0.47328308,0.5658819,0.64133286,0.7510797,0.88826317,0.9842916,0.96714365,0.8779744,0.8196714,0.8196714,0.83338976,0.78537554,0.8162418,0.8025235,0.7510797,0.8162418,0.881404,0.88826317,0.881404,0.94656616,1.2277923,1.2998136,1.2860953,1.2380811,1.1489118,0.96371406,0.7990939,0.7407909,0.7682276,0.805953,0.7613684,0.77508676,0.4664239,0.19548649,0.1097468,0.12346515,0.13032432,0.16804978,0.216064,0.25721905,0.2777966,0.34638834,0.4938606,0.5693115,0.51100856,0.35324752,0.35324752,0.5178677,0.7442205,1.0014396,1.3409687,1.6393428,1.8656956,2.0097382,2.1057668,2.2258022,2.2429502,2.1503513,1.9068506,1.6016173,1.4541451,1.4850113,1.5776103,1.6530612,1.728512,1.8897027,1.879414,1.903421,2.0097382,2.1400626,2.153781,2.0749004,2.054323,2.1194851,2.2223728,2.2395205,2.153781,2.0234566,1.9137098,1.8108221,1.6359133,1.5741806,1.5124481,1.5364552,1.670209,1.8656956,1.7696671,1.6599203,1.6187652,1.6667795,1.7730967,1.6839274,1.7353712,1.6839274,1.5261664,1.4815818,1.5227368,1.4918705,1.4404267,1.4061309,1.4198492,1.2758065,1.1832076,1.1763484,1.3032433,1.6016173,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.030866288,0.072021335,0.106317215,0.18519773,0.28808534,0.28465575,0.21263443,0.28808534,0.44584638,0.84367853,1.6667795,2.8294096,3.9783216,3.4878905,3.0248961,4.1772375,6.8866115,9.445084,12.055,12.788932,13.780083,16.101913,19.764713,23.321196,23.153145,17.556059,9.177576,4.9831905,3.8788633,3.0283258,2.4075704,1.9925903,1.7559488,1.6770682,1.6187652,1.3512574,1.0117283,1.1214751,0.90198153,0.70649505,0.6036074,0.61389613,0.7305021,0.7476501,0.7339317,0.66876954,0.6036074,0.66533995,0.66876954,0.70306545,0.66876954,0.5761707,0.5521636,0.65505123,0.70649505,0.7682276,0.864256,1.0048691,1.2826657,1.5604624,1.7319417,1.7696671,1.7353712,1.8931323,1.937717,2.0165975,2.1640697,2.2978237,2.9391565,3.7519686,4.4104495,5.0655007,6.355026,7.380472,6.341307,8.790032,14.466,17.278261,17.518333,18.70154,23.081123,29.463587,33.191547,33.16754,37.74947,48.833897,62.319035,68.08417,49.756454,38.040985,30.122066,23.791048,17.463459,11.036412,12.836946,15.556609,18.842154,29.292107,61.691418,76.19858,81.14747,78.0094,61.393044,41.05902,33.613388,25.10115,15.086755,16.674654,18.475187,14.613472,10.618003,10.127572,14.88098,9.623423,5.717122,3.426158,2.8019729,3.683377,4.314421,3.1209247,2.2841053,2.4658735,2.8156912,1.1900668,0.64133286,1.1694894,2.0680413,1.9239986,4.2526884,4.73969,3.2478194,1.4369972,2.7882545,2.6476414,1.821111,1.0220171,0.72364295,1.1592005,1.5021594,2.085189,2.153781,1.762808,1.7696671,1.6907866,1.529596,1.4438564,1.5261664,1.8313997,1.7422304,2.1297739,2.9391565,3.309552,1.5536032,1.7765263,2.2463799,3.7005248,4.8494368,2.3767042,1.0254467,0.77165717,0.77851635,0.69963586,0.6756287,2.0646117,3.9886103,4.6848164,3.7039545,1.9137098,2.1983654,2.5961976,3.6970954,4.8322887,4.057202,4.122364,3.1037767,2.9906003,4.197815,5.562791,6.7459984,5.888602,5.411889,6.5127864,9.146709,7.1849856,3.7176728,4.262977,9.31133,14.363112,7.1884155,5.5902276,8.529384,11.650309,7.2947326,5.429037,7.466212,8.292743,6.3721733,3.7553983,4.437886,9.1981535,11.976119,11.080997,9.177576,11.293632,10.2236,12.363663,16.530611,13.954991,8.351046,6.2898636,6.540223,7.4936485,7.160979,4.1189346,5.161529,7.881192,9.781183,8.2653055,7.5862474,14.750656,22.03167,24.247183,18.766703,11.396519,11.417097,12.823228,11.399949,4.698535,15.553179,21.02337,20.752434,15.443433,6.852316,5.137522,6.8763227,8.683716,8.886061,7.534804,6.0635104,6.351596,6.200694,5.8062916,7.7714453,9.729739,9.246168,5.675967,3.199805,10.81006,13.118172,7.291303,5.844017,11.067279,15.031882,7.15069,12.432255,17.772121,16.979887,10.762046,3.8514268,6.108095,9.692014,10.271614,7.0306544,19.582945,15.9613,8.412778,6.15268,15.350834,15.234227,10.031544,5.192395,3.3232703,4.1772375,3.3472774,4.4721823,8.344186,12.295071,10.196163,12.315649,22.089973,21.69557,10.703742,6.0737996,6.783724,5.7651367,3.5393343,2.1434922,5.1066556,8.1041155,7.8434668,6.358455,7.0272245,14.568888,14.387119,11.876661,10.971251,13.13532,17.364002,15.717799,19.987637,24.250612,22.738165,9.860064,5.435896,4.8254294,4.5442033,4.3041325,7.006647,4.386442,2.2566686,1.728512,2.644212,3.566771,3.4124396,2.9734523,2.6167753,2.386993,2.0268862,1.8759843,2.6990852,3.5221863,3.6970954,2.9151495,2.6750782,2.5961976,2.6785078,2.942586,3.4295874,4.763697,5.4324665,4.7534084,3.542764,4.1155047,6.464772,6.800872,7.4936485,8.707723,8.419638,6.2144127,4.4584637,3.5599117,3.7108135,4.887162,5.7377,5.312431,4.2286816,3.1963756,3.0111778,2.1880767,2.644212,3.858286,4.715683,3.5050385,2.7368107,2.9665933,3.1826572,2.9563043,2.4487255,2.0337453,2.6990852,3.2478194,3.474172,4.1600895,3.5187566,3.74168,3.923448,3.4295874,1.9274281,1.4541451,1.7079345,1.8588364,1.6016173,1.1729189,0.99801,0.72707254,0.64819205,0.70649505,0.48357183,0.28465575,0.16804978,0.1097468,0.12003556,0.23321195,0.25721905,0.19891608,0.12346515,0.06859175,0.0274367,0.01371835,0.017147938,0.037725464,0.07545093,0.15090185,0.2709374,0.78194594,1.704505,2.6476414,2.8122618,2.49331,1.6530612,0.9534253,0.6344737,0.5041494,0.3018037,0.26064864,0.25378948,0.22292319,0.16462019,0.11317638,0.12346515,0.15090185,0.39097297,1.2895249,1.4472859,1.0631721,0.72707254,0.5521636,0.14061308,0.13375391,0.12689474,0.08573969,0.030866288,0.058302987,0.06859175,0.116605975,0.12689474,0.14061308,0.32581082,0.45270553,0.38754338,0.45613512,0.78537554,1.313532,0.70306545,0.58302987,0.5521636,0.6379033,1.3066728,2.2429502,2.4487255,2.386993,2.386993,2.6613598,3.6353626,3.216953,2.1674993,1.0940384,0.44584638,0.39097297,0.29494452,0.16804978,0.044584636,0.010288762,0.034295876,0.23664154,0.5624523,0.78194594,0.47671264,0.39783216,0.30523327,0.21263443,0.15776102,0.216064,0.21263443,0.26064864,0.33609957,0.35324752,0.18176813,0.11317638,0.2194936,0.29151493,0.22635277,0.061732575,0.024007112,0.020577524,0.020577524,0.01371835,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.010288762,0.006859175,0.0,0.0,0.006859175,0.010288762,0.010288762,0.006859175,0.01371835,0.006859175,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.05144381,0.18176813,0.4389872,0.5624523,0.64476246,0.6893471,0.64133286,0.4115505,0.4938606,0.64133286,0.86082643,0.9602845,0.53844523,0.23321195,0.09602845,0.041155048,0.037725464,0.10288762,0.22635277,0.25721905,0.23321195,0.17147937,0.09602845,0.116605975,0.12689474,0.15090185,0.20234565,0.274367,0.5212973,1.1660597,1.6427724,1.786815,1.8279701,1.6084765,1.5261664,1.2998136,0.91569984,0.607037,0.50757897,0.51100856,0.48014224,0.3806842,0.28122616,0.3018037,1.8656956,2.5173173,1.6839274,0.66191036,0.66876954,0.71678376,0.83338976,0.9842916,1.0700313,1.0254467,0.9568549,0.91227025,0.90541106,0.9294182,0.8745448,0.8196714,0.7922347,0.805953,0.8848336,0.89169276,0.864256,0.823101,0.85739684,1.1077567,1.2998136,1.313532,1.2792361,1.2380811,1.138623,1.1934965,1.0357354,0.83681935,0.6962063,0.6241849,0.70649505,0.5007198,0.28122616,0.17833854,0.16804978,0.15776102,0.18176813,0.22635277,0.28122616,0.31895164,0.37725464,0.45270553,0.5144381,0.53844523,0.4972902,0.5144381,0.65848076,0.8779744,1.1351935,1.4232788,1.6736387,1.7936742,1.8005334,1.7833855,1.903421,1.8554068,1.8691251,1.7971039,1.6667795,1.6736387,1.5844694,1.6633499,1.762808,1.8142518,1.862266,1.9068506,1.9445761,1.9582944,1.9582944,1.9823016,1.9480057,2.0440342,2.1503513,2.194936,2.1674993,2.1674993,2.1057668,2.0131679,1.8965619,1.7388009,1.6599203,1.646202,1.7010754,1.8279701,2.0268862,1.920569,1.8176813,1.7765263,1.8073926,1.8554068,1.7696671,1.937717,2.037175,1.9720128,1.8554068,1.8862731,1.7730967,1.6496316,1.5913286,1.5981878,1.4987297,1.4027013,1.3855534,1.4918705,1.7319417,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.041155048,0.06859175,0.18862732,0.23321195,0.23321195,0.2503599,0.36696586,0.36696586,0.764798,1.7010754,2.935727,3.8342788,3.4433057,3.3644254,4.4687524,6.989499,10.518545,13.279363,14.376831,15.590904,17.391438,18.921034,22.789608,22.786179,17.254255,8.8929205,4.763697,3.8548563,2.7745364,2.0337453,1.762808,1.7010754,1.7250825,1.6393428,1.3649758,1.0185875,0.9259886,0.90198153,0.7510797,0.607037,0.5624523,0.65505123,0.78194594,0.7922347,0.65848076,0.51100856,0.6241849,0.6756287,0.77165717,0.77165717,0.6962063,0.7407909,0.9568549,1.0528834,1.1454822,1.3203912,1.6153357,1.8828435,2.061182,2.136633,2.0920484,1.8828435,2.0097382,2.0337453,2.1846473,2.702515,3.8102717,4.400161,4.6127954,4.887162,5.754848,7.857185,8.128122,7.346176,9.983529,16.780972,24.754763,29.202938,27.621897,27.93399,33.00635,40.63718,49.509525,52.96655,52.153736,49.825047,50.336056,37.872936,35.92836,31.054914,20.670124,13.066729,13.639469,16.990177,18.166525,22.823904,47.225418,100.209114,127.37831,135.3281,122.05216,76.966805,50.034252,44.900158,35.098396,17.418875,11.900668,14.356253,13.279363,9.383351,6.166398,9.901219,6.090947,2.959734,1.3375391,1.3924125,2.620205,2.5790498,1.862266,1.3169615,1.2895249,1.6324836,1.2792361,1.1763484,1.6976458,2.4247184,2.1469216,3.0351849,4.173808,3.5976372,1.879414,2.0989075,2.1332035,1.488441,0.84024894,0.6756287,1.2826657,1.9514352,2.3732746,2.3801336,2.0508933,1.7147937,1.6839274,1.6016173,1.6599203,1.8554068,1.9891608,1.7490896,1.7079345,2.2292318,2.760818,1.8588364,1.845118,2.1126258,3.0386145,3.6696587,1.704505,1.6564908,1.7113642,1.5947582,1.4129901,1.6564908,3.3369887,5.0243454,4.931747,3.3369887,2.5961976,4.4756117,3.74168,3.1552205,3.7725463,4.9488945,4.554492,3.525616,3.6216443,4.6676683,4.5613513,5.161529,5.3878818,5.8508763,6.2692857,5.4736214,4.2355404,2.976882,3.3781435,5.3227196,6.8797526,4.029765,4.976331,9.602845,14.160767,11.266195,11.814929,14.229359,12.785502,7.1061053,2.1743584,3.3266997,7.98065,11.914387,12.655178,9.506817,12.542002,12.394529,12.476839,13.4474125,13.234778,6.4990683,4.911169,5.693115,6.478491,5.336438,3.0900583,4.8151407,7.8263187,9.908078,9.294182,7.2192817,13.954991,22.69358,27.165762,21.637268,10.88894,9.421077,10.521975,9.352485,2.9700227,11.297061,14.404267,14.613472,12.325937,6.046363,3.566771,3.806842,6.420188,8.954653,6.8557453,7.6376915,8.64599,7.4113383,5.2472687,7.2364297,12.850664,10.31277,5.4496145,4.3007026,13.13532,10.988399,6.0497923,6.4098988,11.993267,14.582606,5.7068334,11.633161,17.562918,16.266533,8.1041155,3.2615378,9.091836,13.337666,11.067279,4.695105,12.415107,10.796341,6.8969,7.6857057,20.015072,13.214201,6.893471,3.9646032,4.3658648,5.051782,3.4398763,3.998899,7.0032177,10.628291,10.947243,13.279363,17.051908,14.359683,6.694555,4.9488945,7.8194594,5.672538,2.6956558,2.2909644,7.06495,10.984968,10.220171,9.211872,10.329918,13.834956,12.284782,9.849775,9.472521,11.640019,14.366542,15.46058,19.94305,24.000254,22.673002,9.873782,5.8337283,7.596536,7.949784,5.909179,6.715132,3.6044965,2.6304936,2.6133456,2.9322972,3.5359046,4.8082814,3.3781435,1.937717,1.5055889,1.4267083,1.9274281,2.877424,3.3266997,3.0077481,2.3149714,2.2292318,2.3424082,2.4967396,2.6922262,3.1072063,4.314421,4.32128,3.6216443,3.117495,4.1155047,5.627953,6.2144127,7.0889573,8.182996,8.107545,5.994919,4.2286816,3.5016088,4.190956,6.355026,6.210983,5.2301207,4.125794,3.6525106,4.605936,2.417859,2.4487255,3.9440255,5.0586414,2.8259802,3.3541365,3.4844608,3.4535947,3.5804894,4.2835546,2.7470996,2.3389788,3.0523329,4.2389703,4.5922174,3.642222,4.506478,4.623084,3.3781435,2.0749004,1.6667795,3.3747141,4.262977,3.357566,1.6221949,1.3443983,0.8025235,0.59674823,0.70306545,0.4664239,0.2469303,0.16462019,0.13375391,0.13032432,0.18862732,0.20234565,0.15776102,0.12003556,0.09602845,0.06859175,0.041155048,0.037725464,0.037725464,0.0548734,0.15090185,0.31209245,0.8676856,1.7799559,2.719663,3.0797696,2.8499873,2.0131679,1.2277923,0.77851635,0.5658819,0.34638834,0.3018037,0.29494452,0.25721905,0.18862732,0.12689474,0.12003556,0.14061308,0.30866286,0.8676856,1.1317638,0.99801,0.7510797,0.490431,0.10288762,0.13032432,0.13032432,0.1371835,0.16119061,0.17490897,0.09945804,0.09945804,0.09259886,0.09259886,0.22978236,0.32924038,0.24350071,0.19891608,0.23664154,0.22635277,0.1371835,0.14404267,0.16119061,0.216064,0.4629943,0.85396725,1.5433143,2.177788,2.8739944,4.180667,4.9351764,4.4550343,3.3815732,2.311542,1.8176813,1.4747226,0.8779744,0.39097297,0.15776102,0.11317638,0.07545093,0.25721905,0.5418748,0.72364295,0.5007198,0.30866286,0.20920484,0.1371835,0.10288762,0.16119061,0.17147937,0.20577525,0.28122616,0.33609957,0.23321195,0.106317215,0.13375391,0.216064,0.2503599,0.13375391,0.058302987,0.024007112,0.01371835,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.010288762,0.0,0.0,0.006859175,0.0034295875,0.0034295875,0.006859175,0.010288762,0.0034295875,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.034295876,0.13375391,0.34638834,0.5418748,0.6344737,0.65848076,0.64133286,0.58988905,0.64819205,0.7099246,0.84367853,0.91912943,0.59331864,0.28122616,0.14404267,0.07545093,0.034295876,0.037725464,0.13375391,0.20234565,0.20577525,0.16462019,0.12346515,0.16804978,0.20920484,0.2469303,0.2777966,0.32238123,0.5453044,1.1043272,1.5193073,1.6496316,1.6804979,1.3821237,1.2346514,1.0940384,0.89169276,0.64476246,0.548734,0.5555932,0.59674823,0.59674823,0.45613512,0.274367,1.255229,2.253239,2.585909,2.061182,1.2826657,0.94656616,0.90541106,0.9877212,0.99801,0.9945804,1.0460242,1.1180456,1.1729189,1.1694894,1.0528834,0.96714365,0.97400284,1.0528834,1.0871792,0.9774324,0.8711152,0.84024894,0.91569984,1.0940384,1.3752645,1.4438564,1.3546871,1.2106444,1.1626302,1.4438564,1.2929544,1.0597426,0.8779744,0.65505123,0.6344737,0.548734,0.4424168,0.33609957,0.22292319,0.16804978,0.17147937,0.22292319,0.3018037,0.37382504,0.39783216,0.37382504,0.4081209,0.4972902,0.53501564,0.5418748,0.64819205,0.8265306,1.0254467,1.1763484,1.4815818,1.546744,1.4644338,1.3821237,1.4953002,1.587899,1.6873571,1.6907866,1.6290541,1.6736387,1.5844694,1.646202,1.6907866,1.670209,1.6736387,1.7216529,1.7593783,1.7353712,1.6873571,1.728512,1.903421,2.0817597,2.1674993,2.136633,2.037175,2.1880767,2.1640697,2.095478,2.0337453,1.9411465,1.8382589,1.8588364,1.8965619,1.903421,1.8931323,1.845118,1.8348293,1.821111,1.786815,1.7319417,1.7113642,1.961724,2.1812177,2.2463799,2.201795,2.153781,1.9925903,1.8897027,1.903421,1.9823016,1.9137098,1.8382589,1.7696671,1.7490896,1.845118,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.061732575,0.15776102,0.16119061,0.17490897,0.24007112,0.32924038,0.34638834,0.6756287,1.6187652,2.942586,3.8720043,3.4467354,3.3129816,4.3041325,7.0306544,11.862943,14.579176,15.930434,16.732958,17.864721,20.255144,24.051697,22.271742,16.194511,8.656279,4.0229063,3.6525106,2.6167753,1.8691251,1.6770682,1.5913286,1.5913286,1.4815818,1.3375391,1.1797781,0.9568549,0.84367853,0.764798,0.7579388,0.764798,0.64476246,0.64476246,0.70649505,0.6790583,0.6001778,0.70649505,0.6824879,0.75450927,0.88826317,1.0323058,1.1249046,1.2586586,1.4061309,1.5741806,1.8108221,2.2086544,2.301253,2.4247184,2.4144297,2.2635276,2.1469216,2.5619018,3.2649672,4.064061,4.9831905,6.279575,5.4736214,4.3281393,4.8254294,7.0615206,9.263316,7.1678376,9.139851,15.103903,25.60873,41.840965,52.393806,41.840965,30.880005,31.991192,49.427216,67.83724,67.96071,53.36438,33.671688,24.538698,16.70895,21.404055,22.566685,15.189643,5.3330083,17.322845,21.85676,19.219408,20.073376,45.424885,92.31421,123.67778,134.74506,116.14641,53.923405,33.133244,35.719154,31.202387,15.004445,8.47451,11.7257595,13.862392,10.947243,4.7088237,2.527606,2.177788,1.0940384,0.78537554,1.6633499,3.0386145,2.1743584,1.4129901,1.1592005,1.3581166,1.4987297,1.6496316,1.728512,1.8656956,2.0268862,2.020027,2.2120838,3.625074,4.057202,2.959734,1.4541451,1.5433143,1.3341095,1.1043272,1.1146159,1.5844694,3.3061223,3.2718265,2.5619018,1.937717,1.8073926,1.6187652,1.9685832,2.3458378,2.393852,1.8931323,1.4953002,1.2483698,1.3101025,1.6804979,2.1983654,2.3767042,2.3218307,2.6545007,3.0729103,2.3286898,3.566771,3.5530527,2.8980014,2.4041407,3.0386145,4.190956,4.0537724,3.0248961,2.287535,3.8102717,7.0203657,4.773986,2.1023371,2.136633,6.101236,6.1629686,4.9488945,4.506478,4.8185706,3.8171308,2.7230926,3.875434,5.8371577,6.5813785,3.5016088,2.2360911,2.5378947,2.3218307,1.4027013,1.4850113,2.942586,6.8043017,11.348505,14.592895,14.321958,17.010754,17.446312,13.056439,5.6142344,1.2312219,1.214074,5.662249,11.856084,15.62863,11.379372,11.965831,12.22648,11.413667,9.801761,8.687145,5.1066556,5.195825,5.6519604,5.0140567,3.6353626,3.2683969,4.2115335,6.0154963,8.035523,9.448513,8.069819,10.041832,16.602633,22.405495,15.549749,8.457363,6.7357097,7.5039372,7.3530354,2.3424082,8.004657,10.542552,12.312219,12.22305,5.7479887,3.690236,5.552502,8.471081,9.568549,5.9400454,8.217292,9.918367,7.9017696,4.4241676,7.1232533,15.333686,10.6317215,5.6073756,7.2707253,17.03819,9.517105,4.7019644,7.160979,14.222499,15.96816,5.3878818,9.194724,14.750656,14.315098,5.06893,3.5118976,13.13532,16.324837,9.750318,4.383013,8.48137,7.5039372,6.15268,8.073249,15.858413,8.81061,3.806842,3.117495,5.2266912,4.7979927,3.6147852,4.972902,6.4098988,7.6925645,10.81006,13.111313,12.6586075,9.170717,4.787704,4.0846386,10.117283,7.8949103,4.245829,3.4810312,7.377043,10.439664,9.1810055,8.851766,11.039842,13.663476,11.413667,10.528833,11.129011,12.21619,11.650309,14.939283,18.965618,22.210009,21.270302,10.847785,9.719451,12.096155,11.369082,7.3873315,6.475061,3.9303071,3.957744,3.8445675,2.860276,2.2738166,5.305572,2.7128036,0.5418748,0.5796003,0.37039545,1.3409687,1.8519772,1.6736387,1.1763484,1.3306799,1.430138,1.5227368,1.7182233,2.0886188,2.6750782,4.396731,4.15666,3.234101,2.8225505,4.0023284,4.7328305,5.381023,6.138962,6.927767,7.4044795,6.279575,4.4104495,3.8514268,5.079219,6.9792104,5.3981705,5.3090014,5.096367,4.7499785,5.8508763,2.4795918,2.4795918,4.355576,5.6073756,2.726522,3.6010668,3.2443898,3.0626216,3.9646032,6.358455,4.32128,3.0523329,3.2889743,4.5922174,5.3227196,3.858286,4.972902,5.0895076,3.4810312,2.287535,1.6873571,4.1943855,5.9640527,5.2266912,2.311542,1.529596,0.8711152,0.6207553,0.65162164,0.4424168,0.18862732,0.13375391,0.15090185,0.17490897,0.17147937,0.13032432,0.12346515,0.12003556,0.11317638,0.09945804,0.06859175,0.061732575,0.05144381,0.0548734,0.13032432,0.5418748,0.9602845,1.3958421,1.8519772,2.3424082,2.6887965,2.3801336,1.7593783,1.1180456,0.6859175,0.5144381,0.45956472,0.42183927,0.34295875,0.22292319,0.14061308,0.116605975,0.13375391,0.216064,0.41840968,0.70649505,0.7339317,0.5418748,0.274367,0.19548649,0.13032432,0.082310095,0.19891608,0.42526886,0.490431,0.26407823,0.13375391,0.08573969,0.09259886,0.1097468,0.15090185,0.082310095,0.12003556,0.2194936,0.0548734,0.06859175,0.106317215,0.1371835,0.1920569,0.36010668,0.66191036,1.5673214,2.4761622,3.3129816,4.537344,5.079219,4.99005,4.280125,3.4192986,3.340418,2.8911421,1.7422304,0.77508676,0.33952916,0.23664154,0.12689474,0.18176813,0.2709374,0.29151493,0.17147937,0.106317215,0.274367,0.37382504,0.30523327,0.17833854,0.1371835,0.12003556,0.15776102,0.2194936,0.22635277,0.06859175,0.041155048,0.06516216,0.10288762,0.16804978,0.082310095,0.034295876,0.010288762,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.010288762,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.08573969,0.23664154,0.53844523,0.5624523,0.5178677,0.5453044,0.75450927,0.78537554,0.77851635,0.8128122,0.84367853,0.6859175,0.36010668,0.18176813,0.09945804,0.061732575,0.010288762,0.020577524,0.0548734,0.07545093,0.09259886,0.15090185,0.20577525,0.30866286,0.39097297,0.4115505,0.34638834,0.6207553,0.9945804,1.3341095,1.546744,1.5741806,1.4369972,1.371835,1.1729189,0.8505377,0.65505123,0.65505123,0.70306545,0.85396725,1.0151579,0.9568549,0.70306545,0.7339317,1.6427724,3.0043187,3.3952916,2.0063086,1.1626302,0.85739684,0.8848336,0.84024894,0.9431366,1.1008976,1.2586586,1.3649758,1.3615463,1.2003556,1.155771,1.2003556,1.2689474,1.2483698,1.1180456,0.94656616,0.9294182,1.0700313,1.2037852,1.4507155,1.5947582,1.488441,1.2277923,1.1489118,1.5261664,1.4404267,1.3375391,1.2792361,0.97057325,0.7305021,0.6893471,0.7133542,0.65505123,0.34981793,0.20234565,0.17147937,0.216064,0.3018037,0.4046913,0.37039545,0.3018037,0.32581082,0.42869842,0.47328308,0.4424168,0.5212973,0.6824879,0.84024894,0.8745448,1.1454822,1.2106444,1.1900668,1.1729189,1.2072148,1.4953002,1.6599203,1.6496316,1.5330256,1.5158776,1.5193073,1.6221949,1.5844694,1.4404267,1.5193073,1.4747226,1.4953002,1.5330256,1.587899,1.6873571,2.0131679,2.1091962,2.0989075,2.0577524,2.0097382,2.318401,2.2566686,2.1469216,2.1263442,2.1469216,2.020027,2.0508933,2.0303159,1.8828435,1.6667795,1.704505,1.7799559,1.7902447,1.7182233,1.6393428,1.6496316,1.8554068,2.054323,2.1674993,2.2498093,2.177788,2.1091962,2.1160555,2.218943,2.369845,2.3458378,2.2909644,2.1846473,2.0680413,2.020027,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.048014224,0.061732575,0.09602845,0.116605975,0.14061308,0.17147937,0.18176813,0.31895164,0.5418748,1.3786942,2.7368107,3.9200184,3.2615378,2.4384367,3.0317552,6.186976,12.617453,15.659496,17.250826,17.21653,17.703531,23.20802,25.19718,20.797018,14.205351,8.220721,4.2423997,3.4124396,2.4795918,1.9068506,1.6770682,1.2963841,1.0528834,1.2860953,1.6496316,1.8965619,1.845118,0.7956643,0.6173257,1.0185875,1.5364552,1.5090185,0.9842916,0.6790583,0.607037,0.6927767,0.77851635,0.864256,1.0494537,1.5433143,2.1263442,2.1503513,1.845118,1.7525192,1.6839274,1.6359133,1.7696671,1.7456601,2.352697,2.609916,2.534465,3.1586502,5.429037,9.263316,12.3533745,12.908967,9.674867,5.830299,4.0057583,5.8817425,9.849775,11.046701,8.7145815,13.773223,22.786179,38.874374,71.69896,92.2902,67.1376,38.870945,28.064314,33.205265,42.434284,41.168766,35.633415,28.458717,18.691252,11.026124,10.858074,13.025573,12.644889,5.127233,15.553179,17.415445,14.376831,10.960961,12.576297,28.01973,47.04365,57.870857,52.438393,26.383816,16.191082,20.591244,18.331144,6.852316,2.2738166,6.217842,6.615674,4.3281393,1.7456601,2.8088322,1.6496316,1.313532,2.3629858,4.0023284,4.0880685,2.6990852,1.7833855,1.5570327,1.6942163,1.3272504,1.155771,1.6187652,2.5447538,3.350707,3.0214665,1.8725548,3.508468,4.6676683,3.6970954,0.548734,0.5144381,1.5021594,2.2223728,2.0714707,1.1454822,2.1812177,2.1674993,1.8313997,1.7079345,2.136633,2.0268862,2.6304936,2.5447538,1.8313997,2.0131679,1.0631721,0.8505377,0.91912943,1.0871792,1.4644338,2.369845,2.3389788,1.9102802,1.7319417,2.5481834,4.6848164,4.7328305,3.525616,2.0508933,1.4644338,2.4418662,2.5378947,2.5447538,3.5050385,6.728851,9.791472,7.747438,4.0366244,2.0234566,4.99005,6.6122446,4.9420357,3.1655092,2.9631636,4.4996185,2.633923,2.194936,3.7519686,6.138962,6.468202,4.5784993,3.7553983,3.1723683,2.7299516,3.0969174,3.7931237,6.5127864,7.438775,5.7891436,3.799983,4.15323,4.1600895,4.605936,4.99005,3.525616,2.1332035,7.267296,14.112752,18.008764,14.479718,7.939495,8.8929205,10.539123,9.249598,4.5613513,6.2830043,9.431366,10.041832,7.407909,4.07435,6.0497923,4.184097,4.1120753,7.4113383,11.595435,12.864383,10.957532,12.6929035,16.832415,14.085316,8.601405,4.852866,5.254128,6.8557453,1.3272504,2.9871707,7.881192,13.697772,16.235666,9.400499,8.237869,8.580828,8.580828,7.466212,5.5250654,7.64798,8.985519,7.1061053,4.8288593,10.2236,15.63206,10.528833,7.3427467,10.618003,17.014183,7.3839016,4.32471,8.107545,14.246507,13.488567,3.5633414,7.0889573,13.742357,15.995596,9.108984,4.057202,14.411126,16.582056,7.0306544,2.2600982,6.835168,5.079219,3.789694,6.3481665,12.696333,5.5902276,1.8725548,1.6667795,2.9906003,1.7696671,3.333559,9.571979,12.562579,10.63858,8.3922,13.701202,14.764374,12.085866,6.7802944,0.5796003,5.7925735,9.283894,8.868914,5.802862,4.7774153,7.0958166,5.360445,3.450165,4.863155,12.710052,10.4533825,8.927217,10.347065,13.848674,15.470869,14.973578,22.875349,25.35494,19.565796,13.656617,18.650097,18.962189,12.144169,2.8019729,2.5927682,3.3884325,4.2081037,5.099797,5.06893,2.0920484,1.6770682,1.039165,0.5521636,0.3566771,0.3806842,0.8471081,1.0254467,0.89169276,0.8779744,1.8931323,1.3684053,1.1351935,1.2037852,1.430138,1.5398848,3.9474552,6.2041235,5.7994323,3.6387923,4.029765,4.0537724,4.938606,5.919468,6.3035817,5.4633327,6.245279,4.681387,5.212973,7.332458,5.6005163,4.245829,7.157549,8.169277,5.7274113,2.884283,2.49331,3.5221863,4.773986,5.302142,4.4104495,2.3458378,1.5844694,2.1640697,3.6696587,5.2335505,5.7582774,4.7808447,3.8720043,3.5873485,3.4776018,5.871454,6.012067,4.557922,3.0077481,3.6936657,2.4830213,1.8897027,1.5055889,1.5055889,2.6407824,1.3203912,0.8093826,0.66876954,0.6241849,0.5658819,0.31895164,0.18519773,0.18519773,0.25721905,0.24350071,0.14747226,0.08573969,0.072021335,0.08916927,0.07545093,0.06516216,0.06859175,0.06859175,0.082310095,0.16804978,0.90198153,1.1283343,1.1763484,1.3409687,1.8759843,1.961724,2.085189,1.961724,1.5776103,1.1763484,1.039165,0.8505377,0.607037,0.34638834,0.1371835,0.11317638,0.12346515,0.14404267,0.16119061,0.19891608,0.4664239,0.4972902,0.4355576,0.40126175,0.48700142,0.40126175,0.29837412,0.40126175,0.6756287,0.8093826,0.5521636,0.26064864,0.1920569,0.29151493,0.18176813,0.048014224,0.05144381,0.05144381,0.017147938,0.030866288,0.20234565,0.3806842,0.4115505,0.45613512,1.0082988,1.3992717,1.8348293,2.633923,3.6970954,4.5030484,3.9886103,3.4295874,2.5378947,1.6324836,1.6324836,2.5961976,1.611906,0.59674823,0.274367,0.15090185,0.17833854,0.12689474,0.061732575,0.061732575,0.24350071,0.36696586,1.2037852,1.5433143,1.0563129,0.274367,0.116605975,0.048014224,0.041155048,0.06859175,0.09259886,0.030866288,0.006859175,0.006859175,0.020577524,0.044584636,0.010288762,0.010288762,0.010288762,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09259886,0.5178677,0.5624523,0.4698535,0.45956472,0.71678376,0.8745448,0.91569984,0.94656616,0.9911508,0.9911508,0.6241849,0.26750782,0.1097468,0.12003556,0.044584636,0.010288762,0.0,0.006859175,0.041155048,0.1371835,0.22292319,0.36353627,0.53501564,0.6379033,0.5041494,0.90541106,1.255229,1.6804979,2.0508933,1.9514352,1.7456601,1.5913286,1.3478279,1.0597426,0.9602845,0.94999576,1.0117283,1.0117283,1.0563129,1.4953002,1.6770682,1.6599203,1.3615463,1.0288762,1.2346514,1.8588364,1.2175035,0.7099246,0.7407909,0.71678376,0.90198153,0.97400284,0.9842916,1.0323058,1.2517995,1.371835,1.3032433,1.1694894,1.0666018,1.0528834,1.2860953,1.1592005,1.0871792,1.1694894,1.2037852,1.1694894,1.3169615,1.3958421,1.3203912,1.1763484,1.6393428,1.7010754,1.5913286,1.4815818,1.4953002,1.0323058,0.9328478,1.1283343,1.2655178,0.71678376,0.36353627,0.26407823,0.2709374,0.30866286,0.3806842,0.34638834,0.37382504,0.4389872,0.5212973,0.59674823,0.59674823,0.6962063,0.8779744,1.0460242,1.0220171,0.864256,0.8779744,1.1729189,1.5124481,1.3443983,1.4027013,1.6770682,1.7353712,1.5913286,1.6633499,1.6770682,1.8965619,1.8965619,1.6770682,1.6770682,1.5570327,1.6359133,1.6599203,1.6633499,1.9685832,2.1263442,1.9480057,1.704505,1.5947582,1.7559488,2.3149714,2.201795,1.9925903,2.0508933,2.503599,2.294394,2.3081124,2.2326615,2.0577524,2.0440342,2.0337453,1.9274281,1.862266,1.8965619,2.0303159,1.9308578,1.862266,1.8554068,1.8828435,1.845118,2.07833,2.311542,2.4247184,2.4315774,2.4555845,2.5173173,2.369845,2.311542,2.3492675,2.1674993,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.0548734,0.08573969,0.082310095,0.14404267,0.23664154,0.29837412,0.23321195,0.28808534,0.4664239,1.1317638,2.2429502,3.3609958,2.8088322,2.201795,3.673088,7.7542973,13.375391,16.444872,16.86671,15.875561,15.145059,16.763824,20.227707,18.005335,12.88839,7.7097125,5.3398676,3.981751,3.0900583,2.6236343,2.311542,1.6393428,1.4438564,1.4747226,1.4267083,1.3615463,1.7113642,1.5604624,1.1660597,1.0014396,1.1180456,1.1317638,0.99801,1.1214751,1.1454822,1.0323058,1.0597426,1.2312219,1.3512574,1.4918705,1.6187652,1.6153357,1.6221949,1.7216529,1.845118,1.9411465,1.978872,3.6147852,4.664239,4.955754,5.305572,7.5279446,9.877212,11.345076,10.545981,8.076678,6.5127864,7.8434668,8.4264965,10.257896,12.751206,12.754636,16.04018,21.11597,25.142305,30.701668,45.812428,65.33021,52.987125,33.42819,21.541239,22.46037,23.331484,22.161995,22.46037,22.302607,14.335675,7.8983397,7.0786686,7.795452,7.5210853,5.284994,8.279024,6.9963584,4.7328305,3.5942078,4.4927597,10.844356,23.221737,29.26467,24.638157,13.042721,7.010077,8.032094,6.9346256,2.5001693,1.4678634,2.5790498,2.5653315,2.0440342,1.5707511,1.6496316,0.84024894,0.84024894,1.8142518,3.2683969,4.0777793,2.6853669,2.6545007,2.767677,2.5619018,2.3389788,1.6324836,1.5501735,2.7779658,4.3761535,3.7519686,1.9514352,2.7882545,3.82399,3.4913201,1.0734608,0.8128122,0.8093826,0.9294182,1.0700313,1.155771,1.8313997,1.9102802,1.6153357,1.3203912,1.5638919,1.4438564,1.9651536,2.8054025,3.1106358,1.4781522,1.2003556,0.89169276,0.6962063,0.70649505,0.9877212,1.7079345,2.054323,2.1674993,2.1880767,2.2429502,3.8137012,3.5221863,2.9871707,2.8705647,2.8808534,3.8479972,3.9440255,3.4398763,3.4776018,6.046363,7.7611566,7.5107965,5.4839106,3.0900583,2.952875,2.767677,2.2258022,1.9342873,2.4830213,4.4413157,4.0091877,3.275256,2.8465576,2.8465576,2.942586,2.750529,1.9582944,1.5604624,2.085189,3.5873485,4.7499785,5.3158607,4.7191124,3.8788633,5.178677,6.2830043,7.805741,8.189855,6.7459984,3.6216443,4.0846386,9.619993,13.612033,13.584596,11.207891,9.589127,9.97324,10.134431,8.872343,6.001778,6.8145905,9.956093,12.703192,12.926115,9.115844,5.6828265,3.4227283,3.391862,5.8508763,10.254466,11.670886,12.092726,14.894698,17.4566,11.166737,8.64599,6.526505,5.5250654,4.5990767,0.97400284,1.7833855,3.3301294,5.0586414,7.1849856,10.679735,9.884071,9.554831,8.1041155,5.892031,5.2301207,7.48336,8.800322,7.2158523,7.0443726,18.866161,20.570665,11.4033785,6.684266,10.374502,15.073037,6.3310184,4.8494368,9.067829,13.450842,8.484799,2.603057,7.582818,15.278812,18.612371,11.598865,6.077229,10.052121,10.47396,5.0757895,2.393852,6.2384195,5.878313,3.923448,4.2218223,11.876661,5.874883,6.6533995,7.4113383,5.8508763,4.149801,2.7745364,5.693115,8.659708,9.89436,10.089847,15.848124,15.258235,9.770895,3.0248961,0.83681935,15.285671,21.760733,18.845583,11.499407,11.050131,12.792361,11.417097,9.22902,9.249598,15.223939,12.332796,8.553391,8.011517,11.396519,15.947581,16.726099,18.8593,19.994495,20.299728,22.456938,31.34643,29.991743,21.990515,12.037852,5.9126086,5.2609873,4.4104495,4.389872,4.3624353,1.6256244,1.1729189,0.7099246,0.4081209,0.32924038,0.4424168,1.2277923,1.3272504,1.1592005,1.4953002,3.4673128,2.0337453,1.0837497,0.7888051,1.1523414,2.0063086,2.8465576,5.7411294,6.557371,4.9660425,4.417309,5.312431,5.4633327,5.377593,5.5250654,6.341307,5.90232,6.0395036,7.1026754,8.004657,6.2212715,4.8082814,6.5779486,7.1369715,5.6965446,5.06893,4.804852,4.040054,4.170378,5.3261495,6.39961,3.673088,3.3301294,3.875434,4.4927597,5.051782,4.746549,3.9200184,3.309552,3.0626216,2.7470996,3.333559,3.532475,3.1415021,2.3492675,1.762808,1.961724,2.5241764,2.568761,2.2978237,2.9940298,2.4075704,1.4335675,0.7373613,0.5212973,0.52815646,0.32238123,0.18519773,0.12346515,0.12689474,0.13375391,0.12346515,0.09945804,0.08916927,0.08916927,0.07545093,0.044584636,0.044584636,0.061732575,0.07888051,0.106317215,0.6344737,1.1694894,1.4404267,1.6564908,2.534465,2.201795,1.9171394,1.6221949,1.2998136,1.0048691,0.8025235,0.72707254,0.6379033,0.4664239,0.20920484,0.12689474,0.082310095,0.06859175,0.09602845,0.16119061,0.23664154,0.34981793,0.40126175,0.42869842,0.6241849,0.72364295,0.45956472,0.4081209,0.5761707,0.41840968,0.20234565,0.09945804,0.106317215,0.14061308,0.061732575,0.09259886,0.23321195,0.33609957,0.32238123,0.18862732,0.5761707,1.1146159,1.4850113,1.4747226,1.0082988,1.3786942,1.430138,1.7456601,2.352697,2.719663,2.8705647,2.836269,2.6304936,2.2463799,1.6804979,1.3375391,0.90198153,0.91569984,1.3203912,1.4815818,1.155771,1.5741806,1.605047,1.0220171,0.5007198,1.1008976,1.6324836,1.7936742,1.4061309,0.4081209,0.30866286,0.44584638,0.4355576,0.26407823,0.29837412,0.082310095,0.010288762,0.0,0.006859175,0.020577524,0.0034295875,0.017147938,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0548734,0.36353627,0.5041494,0.5178677,0.5178677,0.66876954,0.91569984,0.9259886,0.9259886,0.9911508,1.039165,0.7613684,0.44927597,0.30523327,0.3018037,0.17833854,0.0548734,0.017147938,0.006859175,0.020577524,0.08916927,0.21263443,0.3566771,0.47328308,0.5555932,0.6241849,0.922559,1.2792361,1.8073926,2.2635276,2.037175,1.7525192,1.7353712,1.7388009,1.6736387,1.5947582,1.4678634,1.4027013,1.3169615,1.2415106,1.3478279,1.1111864,1.0768905,1.0117283,0.8779744,0.8196714,0.9362774,0.9362774,0.864256,0.7613684,0.66876954,0.8025235,0.7613684,0.67219913,0.64476246,0.77508676,0.9568549,1.155771,1.2860953,1.3066728,1.2346514,1.2826657,1.1694894,1.1043272,1.1694894,1.3032433,1.2483698,1.4335675,1.4781522,1.2826657,1.0288762,1.2380811,1.3684053,1.471293,1.5844694,1.704505,1.4541451,1.2998136,1.2106444,1.1351935,0.9842916,0.5453044,0.5041494,0.4972902,0.4081209,0.39440256,0.32924038,0.31209245,0.34981793,0.4389872,0.5693115,0.58988905,0.6241849,0.7373613,0.91912943,1.0700313,1.196926,1.1146159,1.3272504,1.728512,1.587899,1.4541451,1.4781522,1.5330256,1.6016173,1.7730967,2.1846473,2.4727325,2.2806756,1.7765263,1.6290541,1.6839274,1.7765263,1.8176813,1.786815,1.7490896,1.7010754,1.6976458,1.728512,1.7593783,1.7422304,1.8656956,1.879414,1.8931323,1.9891608,2.2463799,2.428148,2.335549,2.1674993,2.0337453,1.9239986,1.9582944,1.9925903,2.037175,2.095478,2.1503513,2.0920484,2.061182,2.061182,2.085189,2.1263442,2.311542,2.4555845,2.5447538,2.5481834,2.4555845,2.527606,2.644212,2.585909,2.3629858,2.2292318,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.044584636,0.1097468,0.20920484,0.823101,1.1214751,0.8471081,0.30866286,0.2503599,0.3841138,0.9259886,1.8313997,2.7985435,2.2223728,2.2395205,4.184097,7.9737906,12.127021,14.932424,15.717799,15.343974,15.2033615,17.21996,20.481497,18.903887,14.2190695,8.851766,5.888602,4.7088237,4.0091877,3.4638834,2.8294096,1.9514352,1.6393428,1.5776103,1.3821237,1.1489118,1.430138,1.6221949,1.6153357,1.5090185,1.3615463,1.1763484,1.2346514,1.3889829,1.3752645,1.2346514,1.313532,1.670209,1.7319417,1.7147937,1.7559488,1.920569,2.393852,2.9700227,3.865145,4.938606,5.6828265,7.6445503,6.7357097,5.7274113,5.9434752,7.257007,7.5588107,9.551401,11.502836,12.5145645,12.531713,14.160767,13.203912,12.740917,13.7697935,15.206791,17.302269,24.305487,28.475864,29.67279,35.34533,47.04708,44.598354,36.309044,29.480734,30.393003,27.138325,22.20315,18.921034,17.583494,15.422854,9.054111,5.3741636,3.7382503,3.2203827,2.5961976,4.2526884,2.6647894,1.2655178,1.5021594,2.8294096,5.0757895,11.705182,14.373401,11.005547,5.8062916,2.6716487,2.9665933,2.5927682,1.039165,1.3752645,1.7936742,1.6667795,1.430138,1.2860953,1.2106444,0.90884066,1.2037852,1.8656956,2.633923,3.2032347,2.8877127,3.1963756,3.2306714,2.8294096,2.5584722,2.9665933,3.2683969,3.940596,4.770556,4.852866,3.7211025,3.8137012,3.8617156,3.3198407,2.3595562,2.3286898,1.5741806,0.99801,0.91912943,1.0871792,2.4624438,3.642222,3.4776018,2.3904223,2.3424082,2.0028791,1.978872,2.9734523,4.4859004,4.822,2.1057668,1.0906088,0.9362774,1.0254467,0.9534253,1.1763484,1.5673214,1.7971039,1.8588364,2.085189,3.8274195,3.4810312,2.8019729,2.5413244,2.4658735,2.9117198,2.983741,2.585909,2.287535,3.3301294,4.2115335,4.57164,3.8342788,2.452155,1.8999915,2.8328393,3.6696587,4.1155047,4.122364,3.8925817,3.6147852,3.6044965,3.5702004,3.333559,2.8294096,3.1106358,2.901431,2.9460156,3.357566,3.6147852,5.0449233,5.267846,4.3487167,3.3781435,4.4721823,5.5662203,6.23499,6.3481665,6.029215,5.6519604,4.4413157,6.975781,9.078118,10.333347,14.099034,12.682614,10.707172,9.517105,8.700864,6.0703697,5.5422134,8.916927,14.352823,18.118511,14.568888,9.506817,6.324159,4.15323,3.683377,7.1712675,9.14328,7.9017696,8.299602,10.302481,8.961512,8.213862,6.893471,5.4633327,4.372724,4.0709205,5.329579,5.161529,4.2081037,4.139512,7.6685576,10.542552,11.47197,10.381361,8.207003,6.9071894,7.4970784,7.298162,5.8680243,6.416758,15.806969,14.898128,7.8194594,5.8165803,10.30934,12.902108,6.046363,5.209543,9.084977,13.275933,10.288762,6.042933,6.6053853,14.006435,21.009653,11.132441,5.861165,6.667118,6.608815,4.081209,2.8294096,10.065839,8.663138,5.56965,5.425607,10.573419,4.396731,7.8366075,9.942374,7.233,3.7005248,2.0303159,4.928317,8.296172,10.062409,10.155008,11.091286,15.642348,14.277372,7.116394,3.9474552,19.53836,28.76052,23.376068,9.716022,8.690575,9.009526,9.057541,9.366203,10.6317215,13.72178,13.145609,10.580277,10.38479,13.673765,18.327715,19.12681,19.308577,19.260563,19.761284,21.993944,30.657082,28.2598,20.21399,11.509696,6.7185616,6.684266,4.8254294,3.8685746,3.9371665,2.5447538,1.5090185,0.7510797,0.40126175,0.4424168,0.72364295,1.3409687,1.3684053,1.3786942,1.8519772,3.1826572,1.6907866,0.97400284,0.77851635,1.0631721,1.9823016,3.3061223,6.773435,8.056101,6.4407654,4.856296,5.4016004,5.3707337,5.4976287,6.135532,7.267296,6.375603,5.936616,7.274155,9.287323,8.429926,6.2384195,6.7357097,6.7494283,5.645101,5.3330083,5.288424,4.383013,4.033195,4.8905916,6.842027,4.616225,4.434457,5.086078,5.4770513,4.6402316,4.1120753,3.974892,3.642222,3.0351849,2.5824795,2.201795,2.1332035,2.2463799,2.2086544,1.4644338,2.335549,2.2635276,1.961724,1.9137098,2.369845,2.7642474,2.417859,1.7388009,1.0563129,0.6207553,0.34295875,0.19891608,0.12346515,0.082310095,0.07888051,0.11317638,0.09259886,0.07545093,0.08573969,0.09602845,0.072021335,0.048014224,0.048014224,0.07545093,0.09945804,0.4389872,1.1489118,1.5364552,1.6016173,2.0234566,2.585909,2.726522,2.2155135,1.3924125,1.1797781,0.764798,0.805953,0.97400284,0.97400284,0.5590228,0.29837412,0.16119061,0.082310095,0.05144381,0.07888051,0.19891608,0.23664154,0.30866286,0.4424168,0.58302987,0.5693115,0.3841138,0.41840968,0.5796003,0.31209245,0.16119061,0.08573969,0.07888051,0.09945804,0.08573969,0.30523327,0.8711152,1.4267083,1.4987297,0.5212973,0.8505377,1.5433143,1.7696671,1.3992717,1.0082988,1.4987297,1.587899,1.8039631,2.1023371,1.862266,2.2360911,2.7711067,3.457024,3.8548563,3.093488,2.767677,2.1297739,3.0454736,5.0620713,5.40503,3.5187566,4.1326528,4.6745276,3.7279615,1.0323058,1.0768905,1.1489118,1.1317638,0.89512235,0.30523327,0.19891608,0.4355576,0.4664239,0.274367,0.37039545,0.09259886,0.006859175,0.0,0.0,0.006859175,0.0,0.017147938,0.024007112,0.01371835,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.24007112,0.45956472,0.5624523,0.58645946,0.6927767,0.94656616,0.9294182,0.89512235,0.922559,0.9259886,0.7407909,0.5727411,0.5007198,0.490431,0.37725464,0.12346515,0.030866288,0.01371835,0.01371835,0.041155048,0.13032432,0.274367,0.4081209,0.5178677,0.64819205,0.85739684,1.2723769,1.7010754,1.937717,1.7765263,1.4781522,1.5433143,1.6976458,1.7422304,1.5913286,1.5261664,1.5536032,1.646202,1.7147937,1.6221949,1.4438564,1.3546871,1.4095604,1.4541451,1.155771,0.7990939,0.8162418,0.864256,0.805953,0.70306545,0.6859175,0.5590228,0.45613512,0.45613512,0.5658819,0.78194594,1.0734608,1.3546871,1.5158776,1.4095604,1.4815818,1.3306799,1.155771,1.0940384,1.2072148,1.2998136,1.3443983,1.2655178,1.1317638,1.138623,1.1763484,1.2655178,1.3889829,1.4987297,1.5364552,1.4267083,1.4129901,1.3786942,1.2792361,1.1351935,0.78194594,0.70306545,0.66191036,0.5658819,0.48014224,0.37039545,0.33266997,0.3566771,0.41840968,0.490431,0.5521636,0.66876954,0.823101,0.9877212,1.1489118,1.430138,1.4541451,1.5090185,1.6290541,1.611906,1.2758065,1.2106444,1.3581166,1.6324836,1.9274281,2.2738166,2.4075704,2.3252604,2.1229146,1.9925903,1.7593783,1.7319417,1.7559488,1.7353712,1.6221949,1.5090185,1.471293,1.5021594,1.5433143,1.5090185,1.5364552,1.6667795,1.8005334,1.9102802,2.0440342,2.1503513,2.0920484,1.937717,1.7730967,1.7182233,1.8108221,1.9342873,2.0817597,2.2155135,2.2463799,2.0646117,2.0063086,2.037175,2.1229146,2.1983654,2.4418662,2.6236343,2.7779658,2.877424,2.8122618,2.6956558,2.750529,2.7539587,2.6716487,2.6373527,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.006859175,0.034295876,0.09259886,0.4664239,2.0886188,2.9048605,2.16064,0.40126175,0.24350071,0.34638834,0.86082643,1.6942163,2.5173173,1.9068506,2.3286898,4.3109913,7.589677,11.132441,14.13676,15.498305,15.158776,14.829536,17.991615,19.850452,17.88873,14.092175,10.072699,7.0375133,4.955754,4.2938433,4.016047,3.450165,2.294394,1.8965619,1.5844694,1.3169615,1.155771,1.2483698,1.3032433,1.5261664,1.6324836,1.5330256,1.3443983,1.4575747,1.5021594,1.4850113,1.4781522,1.605047,1.7525192,1.8382589,1.99602,2.1812177,2.170929,3.0969174,3.957744,5.271276,6.694555,7.0135064,7.6033955,6.1732574,5.295283,5.672538,6.121814,5.48734,9.815479,15.05246,18.482046,18.70497,19.03421,14.96672,11.948683,12.260776,14.994157,14.788382,20.340883,25.961977,29.871706,34.210136,41.281944,43.06533,38.946396,32.725124,32.618805,28.619907,22.762173,16.575195,12.05843,11.664027,10.436234,6.5024977,3.3541365,2.1400626,1.6873571,3.8891523,2.2395205,0.7133542,1.0357354,2.702515,3.6182148,5.6519604,6.121814,4.48933,2.3492675,1.2209331,1.5124481,1.4198492,0.8676856,1.5090185,1.9823016,1.9274281,1.7353712,1.5536032,1.2723769,1.1934965,1.6976458,2.0508933,2.1812177,2.6716487,3.0214665,3.1963756,3.1620796,2.9048605,2.4247184,3.4227283,4.1120753,4.32128,4.40702,5.2438393,5.693115,5.429037,4.722542,3.9680326,3.6696587,4.1017866,2.6750782,1.4507155,1.1351935,1.0563129,4.4241676,8.423067,8.783174,5.8200097,4.4241676,3.5770597,2.4418662,3.2786856,6.2075534,9.205012,3.391862,1.3169615,2.0234566,3.3438478,1.8965619,1.0082988,1.4095604,1.937717,2.1057668,2.0920484,3.4913201,3.7039545,3.292404,2.6167753,1.8416885,1.9685832,1.7662375,1.4267083,1.1934965,1.3512574,1.8965619,2.277246,2.1572106,1.7593783,1.8656956,3.5942078,5.0003386,5.562791,5.0106273,3.357566,3.1140654,4.0023284,4.4859004,4.15323,3.7451096,3.6216443,3.8102717,4.0434837,4.0229063,3.4227283,4.4687524,4.4516044,3.525616,2.7093742,3.8617156,4.0091877,3.7176728,3.99204,5.171818,6.9380555,3.858286,4.5682106,7.500508,12.9638405,23.163433,18.303709,11.595435,8.793462,9.205012,5.686256,4.729401,8.011517,12.864383,16.63007,16.664366,14.088745,10.367643,5.751418,2.469303,4.7191124,9.6645775,8.152129,5.435896,4.8940215,8.035523,8.1212635,8.086967,7.671987,7.274155,7.936065,8.207003,7.966932,6.9037595,5.6313825,5.6793966,11.814929,13.893259,12.723769,9.952662,8.073249,6.9723516,5.5559316,4.7431192,5.552502,9.074688,7.130112,4.383013,6.2658563,11.091286,10.065839,5.15467,4.623084,7.274155,11.369082,14.610043,12.082437,7.3118806,12.024134,20.697561,10.569988,6.40304,5.2575574,4.804852,3.8720043,2.4384367,10.086417,9.499957,6.917478,6.0635104,8.169277,2.8122618,8.47451,10.796341,6.2487082,2.1332035,1.6633499,7.6857057,11.859513,11.47197,9.448513,6.550512,14.088745,18.756414,15.971589,9.870353,21.712719,31.384155,25.557285,9.321619,6.193835,5.1100855,5.9640527,7.720001,9.616563,11.1393,16.602633,14.970149,13.481709,15.3302555,19.654966,21.304598,21.486366,20.361462,19.219408,20.467777,25.492125,23.849352,17.833855,11.423956,10.261326,8.282454,4.976331,3.5359046,4.180667,4.173808,2.6956558,1.3684053,0.6344737,0.5693115,0.88826317,1.5090185,1.4472859,1.6804979,2.2806756,2.4247184,1.3821237,0.9534253,0.91227025,1.1660597,1.7456601,4.1292233,7.610255,9.321619,8.351046,5.7651367,4.773986,4.15666,4.5956473,6.0737996,7.857185,7.1026754,5.5147767,6.0806584,8.2481575,7.9600725,5.7754254,6.0052075,6.1904054,5.4084597,4.256118,5.0757895,5.0449233,4.5510626,4.6093655,6.8557453,5.3398676,4.8837323,5.305572,5.576509,3.8274195,3.1277838,3.4535947,3.4844608,2.9117198,2.428148,1.6564908,1.3066728,1.4747226,1.7490896,1.2277923,2.3664153,1.7422304,1.1317638,1.2277923,1.6221949,2.020027,2.767677,2.5790498,1.4335675,0.5761707,0.34981793,0.22635277,0.14404267,0.08573969,0.06859175,0.09259886,0.07545093,0.06859175,0.09602845,0.14404267,0.14061308,0.106317215,0.09259886,0.12003556,0.18519773,0.44927597,1.2449403,1.7147937,1.7902447,2.194936,3.3061223,3.625074,2.959734,1.7936742,1.3101025,0.7099246,0.69963586,0.96714365,1.1454822,0.8025235,0.48014224,0.26407823,0.12003556,0.041155048,0.030866288,0.15090185,0.15090185,0.20920484,0.35324752,0.47328308,0.36010668,0.2777966,0.3566771,0.4629943,0.19548649,0.16804978,0.1097468,0.07545093,0.08573969,0.116605975,0.31209245,0.805953,1.3203912,1.4198492,0.5212973,0.72364295,1.2998136,1.4438564,1.2312219,1.6221949,2.0886188,2.095478,2.0680413,1.9685832,1.313532,1.4232788,1.99602,2.9906003,3.923448,3.865145,3.882293,3.018037,4.722542,8.224151,8.522525,4.996909,5.346727,6.1561093,5.2472687,1.6770682,1.4027013,1.08032,0.7888051,0.52815646,0.2194936,0.1371835,0.2503599,0.2709374,0.19548649,0.29494452,0.072021335,0.006859175,0.0034295875,0.006859175,0.01371835,0.0034295875,0.01371835,0.020577524,0.01371835,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.010288762,0.010288762,0.006859175,0.010288762,0.01371835,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.01371835,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13032432,0.36010668,0.52815646,0.6207553,0.77851635,0.91912943,0.881404,0.89855194,0.9911508,0.97400284,0.7990939,0.71678376,0.69963586,0.66876954,0.51100856,0.20920484,0.07545093,0.030866288,0.01371835,0.01371835,0.058302987,0.1920569,0.36010668,0.53158605,0.7133542,0.805953,1.1283343,1.4267083,1.5707511,1.5638919,1.2586586,1.3478279,1.6359133,1.8965619,1.8416885,1.4918705,1.4610043,1.6599203,1.8862731,1.8142518,1.7936742,1.6427724,1.6016173,1.5981878,1.2620882,0.8745448,0.764798,0.7990939,0.8505377,0.7888051,0.6001778,0.42183927,0.34638834,0.38754338,0.4664239,0.6859175,0.96371406,1.2689474,1.4953002,1.471293,1.529596,1.3341095,1.0940384,0.9328478,0.89855194,1.1626302,1.1283343,0.9911508,0.9568549,1.2483698,1.1283343,1.138623,1.2620882,1.4164196,1.4507155,1.4061309,1.3752645,1.3855534,1.3855534,1.2277923,0.97057325,0.8505377,0.8162418,0.805953,0.7305021,0.53158605,0.45270553,0.4389872,0.45613512,0.48357183,0.61046654,0.77165717,0.9259886,1.0768905,1.2929544,1.6359133,1.7147937,1.6016173,1.4335675,1.4164196,1.0700313,1.039165,1.2689474,1.6256244,1.9102802,2.0646117,2.0989075,2.1297739,2.1572106,2.07833,1.8759843,1.8519772,1.8382589,1.7388009,1.5158776,1.4438564,1.4644338,1.4747226,1.4472859,1.430138,1.4198492,1.5158776,1.6256244,1.6942163,1.7147937,1.7422304,1.786815,1.7388009,1.611906,1.5536032,1.670209,1.821111,2.0508933,2.2738166,2.2566686,1.9891608,1.9068506,1.9720128,2.1126258,2.2223728,2.4761622,2.620205,2.7882545,2.9906003,3.1072063,2.9803114,2.9906003,3.0283258,3.0283258,2.976882,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.006859175,0.01371835,0.037725464,0.061732575,0.94656616,3.3712845,4.461893,3.2066643,0.44927597,0.25721905,0.32581082,0.8162418,1.6393428,2.452155,1.9274281,2.836269,4.7842746,7.4936485,10.81006,14.514014,16.019604,14.654627,12.950122,16.61292,17.470318,15.165636,12.449403,10.326488,8.076678,5.0757895,4.3007026,4.2423997,3.8514268,2.534465,2.1743584,1.605047,1.2723769,1.2449403,1.2277923,1.0631721,1.214074,1.3889829,1.4575747,1.4507155,1.5570327,1.5193073,1.5844694,1.7696671,1.8588364,1.5501735,1.6976458,2.1263442,2.469303,2.16064,3.1552205,3.981751,5.3330083,6.608815,5.90575,5.212973,4.863155,4.979761,5.545643,6.4098988,7.0375133,12.521424,17.892159,20.467777,19.850452,19.720127,13.529722,9.239308,9.616563,12.236768,12.703192,13.96185,19.229696,27.52587,33.67855,39.88267,40.40397,34.179268,25.039417,21.699,18.451181,15.337115,10.875222,5.885172,3.5050385,9.129561,7.750868,4.9008803,3.350707,3.0866287,5.3981705,3.5702004,1.2929544,0.58302987,1.7730967,3.433017,2.651071,1.786815,1.6393428,1.4644338,1.2175035,1.4369972,1.4541451,1.3306799,1.8759843,2.534465,2.5961976,2.5619018,2.435007,1.7182233,1.5433143,1.9891608,2.2600982,2.3629858,3.1106358,3.450165,3.2992632,3.1586502,3.0111778,2.3149714,3.210094,3.940596,4.0057583,3.8205605,4.722542,6.728851,7.0958166,6.7185616,6.101236,5.3398676,6.2864337,5.1512403,3.4776018,2.1229146,1.2586586,6.0052075,12.758065,13.704632,8.80718,5.7925735,4.8082814,2.884283,3.3987212,6.848886,10.861504,3.99204,1.4369972,2.9631636,5.4153185,2.7402403,1.1111864,1.6839274,2.6304936,2.935727,2.417859,2.8019729,3.625074,3.9783216,3.5050385,2.393852,2.6956558,2.1434922,1.4335675,1.0151579,1.097468,1.6873571,2.0989075,2.2463799,2.253239,2.4315774,3.234101,4.07435,4.437886,4.064061,2.9563043,2.9220085,4.166949,4.5099077,3.7759757,3.799983,3.0351849,3.2375305,3.4467354,3.3266997,3.175798,3.3712845,2.651071,1.9445761,2.270387,4.729401,3.1380725,2.4007113,3.1037767,4.863155,6.3207297,3.100347,4.0057583,9.211872,18.488907,31.198957,22.659285,12.041282,8.124693,9.81205,6.142391,5.1752477,8.573969,10.525404,11.067279,16.105343,16.70895,12.682614,7.06495,3.1072063,4.262977,11.694893,12.109874,8.416207,5.0312047,7.8537555,8.128122,9.14328,10.179015,10.683165,10.268185,7.623973,8.289313,9.239308,8.694004,6.108095,13.011855,14.764374,12.576297,9.167287,8.766026,6.217842,4.5922174,5.1238036,6.3824625,4.2698364,2.3149714,3.1380725,7.658269,12.072148,7.870903,4.1017866,3.841138,4.712253,7.997798,18.629519,16.2974,9.156999,11.0981455,19.267422,14.081886,9.078118,5.6039457,4.32471,4.1326528,2.1503513,5.8200097,8.351046,8.515666,6.9380555,6.0806584,2.3081124,10.041832,11.47197,4.1155047,0.805953,3.1449318,11.149589,14.634049,11.7086115,8.779744,5.751418,11.989838,21.342323,26.287788,17.95389,22.223726,30.228384,27.42641,14.79867,8.848335,5.593657,6.042933,7.740579,9.211872,9.9801,20.131678,18.427174,14.953001,15.46401,21.383478,23.904224,23.623,21.44521,19.716698,22.210009,23.427511,22.216867,18.852442,15.5085945,16.280252,10.854645,6.217842,4.2869844,4.8734436,5.65539,3.9303071,2.1160555,0.96371406,0.6756287,0.89855194,1.6770682,1.6770682,1.9411465,2.3835633,1.7799559,1.255229,0.86082643,0.89169276,1.313532,1.762808,4.5682106,7.1987042,9.139851,9.595985,7.486789,4.856296,2.7985435,2.7299516,4.7259717,7.531374,7.1232533,5.295283,4.7534084,5.4907694,4.791134,3.6285036,4.5819287,5.576509,5.288424,3.1449318,4.880303,5.8371577,5.4667625,4.928317,7.0958166,5.9812007,5.2815647,5.3330083,5.2506986,2.9288676,2.136633,2.3835633,2.7470996,2.7299516,2.2395205,1.4644338,0.9842916,0.89855194,0.9911508,0.7099246,1.7216529,1.2929544,0.764798,0.78537554,1.2895249,0.9842916,2.2360911,2.4487255,1.2312219,0.39783216,0.33266997,0.2503599,0.16804978,0.10288762,0.06859175,0.06859175,0.07545093,0.082310095,0.106317215,0.18176813,0.216064,0.19548649,0.16804978,0.17833854,0.274367,0.58302987,1.4541451,1.9685832,2.1332035,2.884283,4.173808,4.482471,3.7279615,2.3801336,1.4575747,0.8471081,0.5453044,0.6173257,0.8745448,0.864256,0.6344737,0.36696586,0.16462019,0.06516216,0.037725464,0.061732575,0.09602845,0.12689474,0.19548649,0.39440256,0.34638834,0.2503599,0.22292319,0.22635277,0.058302987,0.12003556,0.10288762,0.07545093,0.06859175,0.09945804,0.12346515,0.12689474,0.15090185,0.20920484,0.29494452,0.36696586,0.607037,0.8025235,1.1214751,2.1263442,2.469303,2.2909644,2.0680413,1.8348293,1.2037852,0.7373613,0.86082643,1.5638919,2.5447538,3.2203827,3.4124396,2.8705647,4.856296,8.464222,8.628842,4.8151407,4.7534084,5.346727,4.7191124,2.2292318,1.9925903,1.5981878,1.2346514,0.881404,0.3018037,0.34981793,0.17833854,0.1097468,0.18519773,0.16119061,0.044584636,0.006859175,0.010288762,0.024007112,0.037725464,0.006859175,0.006859175,0.01371835,0.017147938,0.020577524,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.030866288,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.20577525,0.39440256,0.5727411,0.77165717,0.77851635,0.7613684,0.8745448,1.0597426,1.0666018,0.91227025,0.8745448,0.8505377,0.7579388,0.53158605,0.28122616,0.1371835,0.058302987,0.01371835,0.01371835,0.020577524,0.12346515,0.29837412,0.5212973,0.7888051,0.7990939,0.90884066,1.1249046,1.3615463,1.4610043,1.1797781,1.2037852,1.5741806,2.0680413,2.2258022,1.4095604,1.155771,1.3341095,1.6804979,1.7936742,1.8416885,1.670209,1.4507155,1.2826657,1.1832076,1.0563129,0.8265306,0.77165717,0.89512235,0.89169276,0.5796003,0.37382504,0.31209245,0.3566771,0.37382504,0.5624523,0.77165717,0.99801,1.214074,1.3992717,1.3649758,1.1420527,0.90198153,0.71678376,0.5590228,0.90198153,0.94656616,0.85739684,0.8471081,1.1832076,1.0563129,1.0288762,1.2380811,1.5673214,1.6599203,1.5981878,1.3889829,1.3066728,1.3581166,1.3101025,1.2106444,1.039165,0.9534253,0.9602845,0.91227025,0.65848076,0.5658819,0.53844523,0.53844523,0.58645946,0.764798,0.88826317,1.0048691,1.1866373,1.5330256,1.7113642,1.7250825,1.5570327,1.2998136,1.1454822,0.9842916,1.0494537,1.3101025,1.6359133,1.7799559,1.8108221,1.8656956,1.8965619,1.8931323,1.8656956,1.961724,2.0474637,2.020027,1.8279701,1.4815818,1.488441,1.6187652,1.6427724,1.5364552,1.5021594,1.4610043,1.4369972,1.4781522,1.5433143,1.529596,1.5433143,1.6153357,1.6633499,1.6324836,1.5021594,1.587899,1.7182233,1.9720128,2.218943,2.1297739,1.9068506,1.8862731,1.99602,2.153781,2.2669573,2.4624438,2.5173173,2.627064,2.8499873,3.117495,3.175798,3.2718265,3.292404,3.2032347,3.0557625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.048014224,0.12346515,1.8176813,3.5804894,3.4467354,1.5947582,0.34981793,0.216064,0.2194936,0.48357183,1.1111864,2.1983654,2.0131679,4.705394,7.3118806,8.735159,9.736599,13.958421,15.223939,12.97413,10.460241,14.771234,17.737827,16.767254,13.279363,9.098696,6.4407654,6.3893213,5.6999745,4.5030484,3.1826572,2.3664153,2.1194851,1.8588364,1.5364552,1.2517995,1.2517995,1.5090185,1.728512,1.7216529,1.5227368,1.3889829,1.5364552,1.5433143,1.704505,1.9445761,1.845118,1.6153357,1.6942163,1.8965619,2.1229146,2.3801336,2.4795918,3.1517909,5.051782,7.4181976,8.100685,10.1652975,8.985519,7.051232,6.4579134,8.9100685,11.948683,12.507706,13.560589,15.196502,14.647768,16.492886,11.907528,8.721441,9.3079,10.590566,17.168514,17.641798,18.392878,21.033659,22.402065,22.69358,19.52807,16.266533,13.128461,7.1712675,3.2409601,1.4815818,1.1626302,1.5981878,2.136633,3.3678548,2.9185789,2.417859,2.585909,3.2203827,4.770556,4.5167665,2.7093742,0.5658819,0.26064864,5.5319247,4.7534084,3.0077481,2.5996273,3.0523329,1.7696671,2.1640697,2.6579304,2.74367,2.976882,4.122364,4.170378,3.8548563,3.4021509,2.5481834,2.3046827,2.095478,2.74367,4.0023284,4.5613513,5.1855364,5.0003386,4.2081037,3.1963756,2.5481834,4.4756117,5.1512403,4.887162,4.2355404,3.9680326,6.029215,8.879202,10.515115,10.261326,8.759167,10.124143,12.21619,10.432805,5.2026844,1.9685832,3.4227283,8.580828,9.246168,4.852866,2.4727325,3.117495,2.6133456,2.4487255,3.316411,5.113515,2.1572106,1.2998136,1.3786942,1.4472859,0.764798,1.0563129,2.0817597,2.8088322,3.0283258,3.357566,2.9906003,3.0077481,3.5530527,4.4584637,5.2644167,6.0806584,5.717122,4.0949273,2.136633,1.7696671,2.5619018,3.6044965,4.5990767,4.7499785,2.760818,1.3581166,0.8711152,1.2175035,1.9925903,2.4555845,2.2258022,2.6613598,2.935727,2.603057,1.6016173,0.90541106,1.0528834,1.6016173,2.287535,3.0043187,2.6647894,1.371835,1.7902447,4.437886,7.658269,3.998899,2.3046827,2.719663,4.122364,4.1360826,3.0248961,3.2409601,7.8846216,16.245956,23.787619,17.075916,10.343636,7.723431,8.903209,9.108984,6.217842,11.543991,14.04759,13.018714,18.097933,15.350834,10.069269,6.492209,5.813151,6.1801167,7.7920227,8.515666,8.954653,8.793462,6.8043017,6.9517736,6.0086374,6.4236174,8.255017,9.170717,3.4227283,4.6573796,7.654839,8.868914,6.4407654,11.163307,10.422516,7.517656,6.375603,11.550851,6.5710897,5.3981705,7.888051,10.151579,4.5613513,2.0234566,3.5873485,7.716572,11.252477,9.383351,5.147811,5.1409516,4.4413157,6.0703697,21.009653,11.63659,7.891481,12.6586075,22.395206,27.145185,13.642899,6.2487082,3.858286,4.420738,4.9591837,4.557922,9.078118,13.3033695,13.564018,7.7680154,3.590778,12.425395,13.433694,4.197815,0.7339317,8.872343,9.253027,6.800872,5.6073756,8.927217,8.632272,13.978998,25.138876,34.553093,26.959988,18.722118,25.378946,29.950588,26.219196,18.735836,10.069269,9.424506,12.439114,14.812388,12.298501,14.863832,14.393978,14.064738,17.62465,29.401854,29.072613,24.936531,21.596113,22.052248,27.6802,30.68109,24.19917,20.237995,21.016512,18.965618,15.37827,11.7257595,7.939495,5.2026844,5.936616,3.6147852,1.8999915,0.99801,0.823101,1.0082988,1.3992717,1.9720128,1.7765263,1.0117283,1.0220171,0.5453044,0.216064,0.37039545,1.1900668,2.7162333,4.3281393,5.113515,6.036074,7.682276,10.268185,8.05953,3.7622573,1.6804979,2.942586,5.4941993,5.055212,5.15467,5.422178,5.120374,3.1449318,2.9974594,4.48933,5.9434752,6.077229,4.012617,5.0140567,5.9126086,6.0840883,6.108095,7.7680154,6.632822,6.852316,7.2604365,6.444195,2.7470996,2.5378947,2.294394,2.6304936,3.1552205,2.4727325,2.020027,1.5227368,1.0768905,0.7956643,0.8093826,0.980862,0.939707,0.77508676,0.7990939,1.5570327,1.6530612,1.313532,0.8128122,0.4081209,0.33609957,0.31209245,0.26064864,0.18519773,0.106317215,0.044584636,0.082310095,0.12689474,0.12346515,0.08573969,0.12346515,0.23321195,0.23321195,0.17147937,0.116605975,0.15090185,0.5178677,1.5810398,2.0577524,1.821111,1.9068506,4.6402316,5.919468,5.0586414,2.9734523,2.1674993,1.786815,0.9877212,0.5555932,0.6790583,0.9602845,0.84024894,0.53501564,0.25378948,0.09602845,0.061732575,0.08573969,0.082310095,0.06859175,0.1371835,0.4424168,0.58988905,0.32238123,0.09602845,0.082310095,0.16804978,0.082310095,0.05144381,0.05144381,0.06516216,0.07545093,0.1371835,0.17833854,0.17490897,0.22292319,0.5658819,0.42869842,0.26750782,0.23664154,0.34638834,0.4424168,0.9294182,1.0631721,1.6221949,2.4487255,2.411,1.4472859,1.3169615,1.8759843,2.4144297,1.6324836,1.8142518,2.5756202,3.5393343,4.355576,4.6848164,3.683377,3.8720043,3.9268777,3.340418,2.411,1.5673214,1.7319417,2.1674993,2.0714707,0.59674823,0.9259886,0.5761707,0.3806842,0.4424168,0.1371835,0.041155048,0.01371835,0.0274367,0.048014224,0.061732575,0.01371835,0.0,0.006859175,0.034295876,0.106317215,0.058302987,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.058302987,0.18519773,0.3566771,0.3806842,0.4664239,0.5796003,0.64819205,0.65162164,0.6241849,0.7956643,0.94999576,0.8745448,0.6173257,0.45613512,0.274367,0.16462019,0.07888051,0.01371835,0.0,0.0,0.0274367,0.13032432,0.33952916,0.65505123,0.7888051,0.86082643,1.0082988,1.1934965,1.2037852,1.0597426,0.922559,1.1043272,1.5055889,1.6016173,0.9911508,0.6927767,0.9568549,1.5638919,1.8313997,1.8313997,1.7490896,1.6324836,1.6359133,2.0131679,1.7216529,1.1626302,0.8745448,0.939707,0.9774324,0.6344737,0.3841138,0.28808534,0.29151493,0.22978236,0.37382504,0.4664239,0.58988905,0.823101,1.2517995,1.2380811,0.99801,0.69963586,0.51100856,0.59674823,0.84024894,1.039165,1.0563129,0.9294182,0.85396725,1.1832076,1.3032433,1.6873571,2.2086544,2.136633,1.9651536,1.7765263,1.5261664,1.3203912,1.4198492,1.8108221,1.4575747,0.9774324,0.65505123,0.47328308,0.37382504,0.45956472,0.5658819,0.6344737,0.7339317,0.89169276,0.9945804,1.1832076,1.4953002,1.862266,1.3992717,1.3375391,1.371835,1.3169615,1.0837497,1.1214751,1.2380811,1.4953002,1.7902447,1.8759843,1.8897027,1.937717,1.9548649,1.9514352,1.9994495,1.8039631,1.8108221,1.8588364,1.8348293,1.6633499,1.7010754,1.6256244,1.5227368,1.4267083,1.3443983,1.4781522,1.4918705,1.6633499,1.9925903,2.2120838,1.9445761,1.7765263,1.6976458,1.6599203,1.587899,1.587899,1.6873571,1.845118,1.9480057,1.8005334,1.762808,1.9651536,2.1983654,2.3286898,2.3046827,2.5001693,2.6476414,2.7539587,2.8122618,2.8225505,2.9322972,3.1072063,3.1312134,2.9940298,2.884283,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.034295876,0.05144381,0.2194936,0.82996017,4.040054,4.57507,3.1586502,1.0871792,0.25378948,0.274367,0.33266997,0.64476246,1.3889829,2.7093742,2.4384367,4.4859004,7.130112,9.071259,9.417647,11.80464,14.064738,13.728639,13.272504,20.093952,22.131128,19.164536,14.531162,10.556271,8.549961,6.8900414,5.219832,3.765687,2.7985435,2.633923,2.07833,1.6427724,1.4541451,1.4164196,1.2037852,1.5090185,1.879414,2.0234566,1.9445761,1.937717,1.9582944,1.8759843,1.8725548,1.8897027,1.6256244,1.471293,1.704505,2.1194851,2.527606,2.7470996,2.5413244,2.9940298,4.1600895,5.552502,6.138962,8.601405,12.377381,16.750105,20.954779,24.182022,22.19286,20.423193,21.479506,23.475527,20.056227,13.88297,15.062748,16.942162,16.019604,11.979549,16.79469,18.142517,17.257685,15.433144,14.027013,12.260776,10.933525,10.127572,9.126132,6.4407654,3.7965534,2.0646117,1.5055889,2.4144297,5.137522,5.2575574,4.822,4.190956,3.4055803,2.194936,3.1106358,4.835718,4.9831905,2.9803114,0.07545093,1.6873571,2.3664153,2.3972816,2.6476414,4.5647807,5.130663,3.683377,2.9631636,3.4776018,3.525616,2.867135,2.7573884,3.3747141,4.0606318,3.3061223,2.7779658,3.2821152,3.6113555,3.415869,3.1963756,4.314421,5.377593,5.1066556,3.7382503,3.0248961,4.180667,5.562791,6.557371,6.869464,6.543653,9.602845,10.628291,11.345076,11.602294,9.369633,7.181556,6.427047,6.910619,7.281014,5.0312047,2.568761,4.962613,6.3173003,4.8014226,2.6545007,4.6676683,3.7794054,2.510458,2.0817597,2.4007113,1.7422304,1.3272504,1.2209331,1.3443983,1.471293,1.6084765,2.5207467,3.57363,4.4687524,5.23698,9.870353,10.792912,8.31332,4.866585,5.007198,5.4941993,5.422178,4.633373,3.5976372,3.4055803,3.3198407,2.5893385,2.4590142,2.8294096,2.2360911,1.214074,1.2175035,2.5996273,4.091498,2.7985435,1.8828435,1.546744,1.4061309,1.1420527,0.490431,0.44927597,0.6927767,1.039165,1.488441,2.2498093,2.3561265,2.0474637,2.6956558,4.4756117,6.341307,3.4981792,2.0920484,2.867135,4.4516044,3.3301294,2.8534167,3.6765177,6.351596,10.316199,13.876111,15.189643,12.751206,8.597976,5.1340923,5.1066556,4.5956473,10.079557,17.20967,20.824455,14.946142,10.854645,8.330468,6.625963,6.64997,11.002116,7.4284863,7.4696417,8.738589,9.132992,6.8283086,7.953213,6.615674,5.4976287,5.470192,5.593657,5.7136927,7.301592,7.716572,7.48336,10.30934,16.828985,15.254805,8.694004,2.7711067,5.641671,4.3624353,6.8043017,9.870353,10.237319,4.341858,2.3321195,3.9508848,6.193835,7.010077,5.31929,3.8171308,11.019264,13.649758,10.443094,12.175035,13.893259,12.072148,12.2093315,15.944152,21.04395,11.05699,6.0052075,5.0826488,6.042933,5.2026844,4.605936,10.251037,15.827546,15.988737,6.3618846,4.588788,9.469091,9.794902,4.372724,2.037175,7.6616983,7.9943686,5.6142344,3.7005248,6.0326443,9.47938,17.034761,29.473875,38.023838,24.387796,14.534592,13.327377,15.367981,16.180794,12.181894,10.655728,14.668345,16.973028,16.311117,17.449741,18.3723,17.86815,18.941612,22.642136,28.074602,30.51647,27.93742,25.862518,27.618467,34.31988,34.031796,30.043186,24.254042,18.54035,14.791811,14.610043,12.586586,8.934075,5.429037,5.411889,3.7553983,2.3595562,1.6976458,1.4335675,0.44584638,2.7128036,2.0474637,1.1454822,1.1111864,1.4850113,0.70649505,0.274367,0.36696586,0.90198153,1.5193073,2.2909644,2.867135,3.3061223,4.355576,7.449064,7.016936,4.972902,4.1189346,5.3432975,7.641121,5.1821065,3.7862647,4.2355404,5.5250654,4.8768735,4.1635194,3.9543142,4.6402316,5.892031,6.660259,7.9086285,7.5862474,6.728851,6.1904054,6.667118,6.478491,7.449064,7.9017696,6.8969,4.2218223,4.1635194,4.249259,3.9783216,3.6044965,4.1326528,2.3732746,1.4095604,1.039165,0.939707,0.65162164,0.52815646,0.4972902,0.77851635,1.1729189,1.0323058,1.7147937,1.1694894,0.61046654,0.5041494,0.5693115,0.47328308,0.29494452,0.16462019,0.11317638,0.082310095,0.07888051,0.1097468,0.11317638,0.10288762,0.15776102,0.18176813,0.16462019,0.15776102,0.22978236,0.48357183,0.8779744,2.0714707,2.3561265,1.5947582,1.2106444,2.5584722,3.74168,3.7794054,3.0317552,3.192946,4.355576,3.357566,1.8897027,0.91569984,0.6790583,0.9602845,0.70306545,0.33952916,0.106317215,0.061732575,0.0548734,0.082310095,0.07888051,0.061732575,0.11317638,0.17147937,0.26407823,0.48700142,0.607037,0.058302987,0.041155048,0.034295876,0.041155048,0.061732575,0.11317638,0.24350071,0.30866286,0.33266997,0.34638834,0.39440256,0.2503599,0.15776102,0.12689474,0.15776102,0.2469303,0.48014224,0.83338976,1.6736387,2.7779658,3.3369887,2.8054025,2.6545007,2.8945718,3.2203827,3.0351849,2.8396983,5.0414934,5.8405876,5.051782,6.111525,6.0086374,6.2487082,6.025785,5.3501563,5.0483527,2.9048605,2.2841053,2.6304936,2.9460156,1.7902447,1.5055889,0.7339317,0.26064864,0.2194936,0.08916927,0.08916927,0.10288762,0.13032432,0.13032432,0.024007112,0.0034295875,0.0,0.006859175,0.020577524,0.034295876,0.024007112,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0034295875,0.010288762,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0274367,0.082310095,0.18519773,0.3566771,0.39440256,0.36353627,0.32238123,0.32238123,0.4046913,0.53844523,0.66533995,0.8128122,0.9431366,0.97057325,0.6001778,0.31209245,0.12689474,0.030866288,0.0,0.0,0.020577524,0.07545093,0.20234565,0.45956472,0.65505123,0.75450927,0.85739684,0.96714365,1.0117283,0.9328478,0.805953,0.7888051,0.9911508,1.4815818,1.0254467,0.6927767,0.6173257,0.7510797,0.84367853,1.2723769,1.3924125,1.2758065,1.1008976,1.1489118,1.371835,1.3238207,1.1866373,1.0871792,1.0871792,0.881404,0.70306545,0.53501564,0.40126175,0.34981793,0.4081209,0.42183927,0.4938606,0.7133542,1.1420527,1.1592005,1.0117283,0.8745448,0.77851635,0.6207553,0.70649505,0.7407909,0.805953,0.90198153,0.96371406,1.1763484,1.3238207,1.4850113,1.6496316,1.7216529,1.6667795,1.5810398,1.6221949,1.728512,1.6016173,1.2689474,0.7888051,0.4629943,0.37039545,0.36353627,0.34295875,0.42526886,0.5418748,0.6859175,0.939707,1.2758065,1.3203912,1.4404267,1.6427724,1.5673214,1.728512,1.5913286,1.4027013,1.2723769,1.1694894,1.1180456,1.3375391,1.6153357,1.7730967,1.6942163,1.8416885,2.1469216,2.3801336,2.503599,2.6716487,2.6785078,2.318401,1.8759843,1.5261664,1.3443983,1.3546871,1.3684053,1.3238207,1.2758065,1.4027013,1.3238207,1.3786942,1.546744,1.7559488,1.9068506,1.8039631,1.6564908,1.6256244,1.7079345,1.7216529,1.605047,1.7422304,2.037175,2.3458378,2.4830213,2.428148,2.4041407,2.3732746,2.3595562,2.4624438,2.7059445,3.0969174,3.4192986,3.5393343,3.3850029,3.1517909,3.0351849,3.069481,3.2066643,3.309552,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.034295876,0.10288762,0.19548649,0.5590228,1.7216529,4.9351764,4.6608095,2.8019729,0.9431366,0.31895164,0.3018037,0.33952916,0.61389613,1.2072148,2.1332035,2.1332035,3.8171308,6.341307,8.841476,10.446524,14.270514,15.21365,14.490007,14.946142,21.067955,21.45893,16.88729,12.367092,10.134431,9.647429,6.5813785,4.65395,3.3609958,2.5619018,2.4898806,2.0303159,1.7216529,1.5810398,1.5638919,1.5638919,2.0646117,2.311542,2.2360911,2.0749004,2.3767042,2.4384367,2.417859,2.5070283,2.719663,2.8980014,2.719663,3.5702004,5.7102633,8.944365,12.624311,9.962952,8.97523,10.069269,12.3533745,13.6086035,15.542891,19.764713,25.372087,30.379286,31.727114,27.76937,28.208357,29.947157,28.709076,19.027351,11.602294,11.434244,14.428274,16.990177,16.026463,15.21365,14.376831,13.282792,11.900668,10.39508,9.174147,9.201583,8.385342,6.375603,4.588788,4.6127954,4.4859004,4.256118,4.2698364,5.1752477,3.99204,3.9680326,4.262977,4.400161,4.245829,3.069481,3.3026927,6.5230756,8.7317295,0.37039545,0.6173257,1.2380811,1.7902447,2.2566686,3.0386145,4.7088237,5.1238036,5.0140567,4.746549,4.32128,4.0674906,4.389872,4.7945633,4.7774153,3.8342788,4.1943855,4.437886,4.57164,4.5339146,4.170378,4.0023284,4.431027,4.8494368,5.127233,5.586798,5.6965446,6.0395036,6.999788,8.261876,8.844906,9.55826,8.433355,7.9017696,8.40249,8.357904,7.0032177,6.138962,6.451054,7.431916,7.390761,3.6627994,5.271276,6.8591747,6.210983,4.256118,5.038064,4.2869844,3.4021509,2.901431,2.393852,2.0131679,2.428148,2.633923,2.4418662,2.4624438,4.105216,5.3501563,5.662249,5.552502,6.584808,9.626852,9.880642,7.7885933,5.209543,5.4187484,4.431027,5.2301207,5.576509,4.7534084,3.566771,2.6750782,1.5090185,1.1249046,1.5158776,1.5947582,1.3615463,1.99602,3.3266997,4.108646,2.0337453,1.4644338,1.4644338,1.4198492,1.1763484,1.0185875,2.6647894,3.391862,3.0969174,2.2738166,1.9857311,2.8739944,3.0900583,2.8739944,2.6133456,2.8808534,2.0303159,1.845118,2.2463799,2.6304936,1.8554068,1.6839274,2.2498093,4.3349986,7.623973,10.683165,12.723769,12.373952,8.964942,4.5270553,3.8205605,3.4364467,7.915488,15.6697855,21.493225,16.568336,13.601744,11.691463,9.328478,7.2604365,8.491658,6.3310184,6.636252,7.7885933,8.237869,6.5230756,7.1095347,5.7925735,4.897451,5.1855364,5.8543057,7.438775,8.405919,7.5519514,6.759717,10.957532,17.655516,15.261664,8.536243,2.5893385,2.8945718,5.2644167,9.887501,12.97413,11.64345,3.940596,2.644212,4.6573796,7.160979,7.7920227,4.6402316,3.7142432,12.103014,17.556059,15.621771,9.654288,14.143619,14.232788,11.499407,9.345626,12.987847,11.1393,9.14328,7.7097125,6.475061,4.0091877,3.4878905,7.016936,10.9369545,11.430815,4.537344,6.931196,11.441104,10.679735,5.5147767,5.0483527,9.153569,7.706283,5.6210938,5.2575574,6.4373355,5.669108,10.117283,17.305698,21.808746,15.265094,11.177026,12.38424,14.184773,13.251926,7.623973,7.1541195,14.13333,19.322296,19.596663,17.95046,17.117071,17.936743,20.762722,24.631298,27.244642,31.535057,29.916292,29.292107,33.356167,42.581757,35.75002,29.01431,22.985096,18.28656,15.525743,15.704081,12.356804,8.001227,4.6573796,3.8342788,3.0454736,1.821111,1.3203912,1.3684053,0.42526886,1.862266,1.7250825,1.2826657,1.138623,1.2072148,0.66191036,0.41498008,0.7682276,1.5124481,1.9239986,1.5947582,1.6599203,2.0268862,3.0043187,5.288424,5.717122,4.6402316,4.1189346,5.0414934,7.099246,4.7979927,3.4398763,3.8548563,5.295283,5.446185,4.2938433,3.7039545,3.7176728,4.437886,6.025785,7.98065,7.7680154,6.677407,6.125243,7.610255,7.366754,8.097256,8.357904,7.3255987,4.8117113,4.8837323,5.1580997,4.513337,3.1860867,2.7711067,1.9720128,1.2963841,1.0048691,0.9774324,0.7305021,0.490431,0.39440256,0.53158605,0.77508676,0.7888051,1.1283343,0.8162418,0.5418748,0.52472687,0.50757897,0.432128,0.29837412,0.17490897,0.09602845,0.072021335,0.082310095,0.13375391,0.13032432,0.07545093,0.08573969,0.13032432,0.15433143,0.18519773,0.31552204,0.6927767,1.1454822,1.6770682,1.6804979,1.214074,0.9911508,1.9994495,3.2786856,3.340418,2.5378947,3.0626216,4.341858,4.033195,2.7333813,1.2620882,0.64819205,1.0323058,0.99801,0.7099246,0.33266997,0.041155048,0.05144381,0.048014224,0.041155048,0.22978236,1.0014396,0.5693115,0.7339317,0.7339317,0.37382504,0.030866288,0.024007112,0.0274367,0.05144381,0.106317215,0.20577525,0.61389613,0.6207553,0.6173257,0.72364295,0.8162418,0.45270553,0.37382504,0.33952916,0.29151493,0.36353627,0.6962063,1.0734608,1.605047,2.2223728,2.6819375,2.942586,3.6319332,4.400161,4.938606,5.0003386,3.5770597,4.245829,4.4275975,3.8102717,4.338428,6.4887795,6.7357097,6.108095,5.3878818,5.103226,2.6133456,1.430138,1.5433143,2.2258022,2.0165975,1.862266,0.922559,0.22978236,0.09602845,0.12346515,0.32238123,0.24350071,0.14747226,0.11317638,0.024007112,0.0034295875,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.006859175,0.017147938,0.017147938,0.010288762,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.08916927,0.22292319,0.18862732,0.14061308,0.1097468,0.12346515,0.20577525,0.274367,0.4355576,0.77508676,1.1797781,1.3169615,0.939707,0.490431,0.17490897,0.044584636,0.0,0.0,0.006859175,0.030866288,0.1097468,0.3018037,0.5521636,0.70306545,0.823101,0.91912943,0.9534253,0.9431366,0.83681935,0.75450927,0.8196714,1.155771,1.0563129,0.83338976,0.61046654,0.4629943,0.40126175,0.6756287,0.84024894,0.8505377,0.77165717,0.8025235,1.1214751,1.2243627,1.1797781,1.0837497,1.039165,0.8265306,0.6962063,0.6310441,0.5727411,0.42869842,0.4698535,0.44584638,0.4629943,0.5693115,0.7476501,0.9911508,1.0666018,1.0563129,0.9568549,0.67219913,0.6241849,0.64476246,0.7373613,0.8779744,1.0288762,1.1008976,1.1146159,1.2072148,1.3649758,1.4267083,1.4678634,1.5055889,1.5707511,1.5741806,1.3169615,0.97400284,0.58645946,0.36353627,0.34981793,0.40126175,0.34981793,0.3841138,0.48357183,0.66533995,1.0014396,1.3512574,1.4129901,1.4541451,1.5604624,1.6324836,1.7079345,1.5707511,1.3889829,1.2723769,1.2620882,1.2929544,1.3992717,1.5090185,1.5604624,1.5090185,1.7662375,2.2326615,2.620205,2.7916842,2.784825,2.603057,2.201795,1.7662375,1.4267083,1.2655178,1.2449403,1.2003556,1.097468,0.9911508,1.0082988,0.9328478,0.96371406,1.0494537,1.1797781,1.4095604,1.4953002,1.4095604,1.3924125,1.488441,1.5638919,1.6221949,1.8588364,2.1812177,2.5447538,2.9665933,3.1826572,3.069481,2.8259802,2.644212,2.7128036,2.9322972,3.2992632,3.5770597,3.6319332,3.4433057,3.3952916,3.3850029,3.4878905,3.6113555,3.5016088,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0034295875,0.010288762,0.037725464,0.1371835,0.274367,0.64819205,1.6736387,4.623084,4.5030484,2.9631636,1.3272504,0.5761707,0.40126175,0.40126175,0.6001778,0.96371406,1.3958421,1.9137098,4.461893,6.756287,8.2481575,10.134431,14.112752,15.302819,15.896138,17.672665,22.011093,20.965069,15.337115,10.731179,9.338767,9.938945,6.5162163,4.664239,3.508468,2.6613598,2.2155135,2.0989075,1.961724,1.8005334,1.7353712,2.0406046,2.5481834,2.527606,2.3081124,2.2669573,2.8294096,2.8122618,3.018037,4.5784993,6.591667,6.138962,7.4113383,11.458252,16.503176,21.325174,25.27606,21.356041,20.220848,21.45207,23.184011,22.083115,25.084003,28.712505,33.157253,37.98954,42.180496,39.351086,41.000717,39.587727,31.826572,18.71526,13.704632,9.880642,10.010965,13.810948,17.981327,13.985858,10.491108,8.687145,8.48137,8.515666,8.3922,8.954653,8.656279,7.1849856,5.48734,5.120374,4.9934793,4.99005,5.144381,5.638242,4.722542,4.0846386,3.9680326,4.2389703,4.386442,2.8019729,2.095478,6.0840883,10.155008,1.2723769,0.67219913,0.89169276,1.5536032,2.1983654,2.2841053,3.806842,5.4667625,6.3001523,6.0875177,5.360445,5.6656785,6.2658563,6.111525,5.038064,3.7725463,4.4687524,5.0757895,5.4153185,5.439326,5.219832,4.5990767,4.40702,4.9214582,5.8817425,6.492209,6.540223,5.994919,6.307011,7.5588107,8.464222,7.5450926,6.0875177,5.1238036,5.2987127,6.883182,7.8263187,7.1952744,6.324159,6.3138704,8.032094,6.715132,6.543653,6.4887795,6.186976,5.960623,4.57507,4.2115335,4.3109913,4.1463714,2.843128,2.2463799,2.7711067,2.901431,2.4761622,2.7059445,4.40702,5.329579,5.2644167,4.787704,5.2747054,6.108095,5.6485305,4.9694724,4.7088237,5.0586414,3.216953,3.841138,4.307562,3.642222,2.5070283,1.961724,1.3032433,0.97057325,1.0871792,1.4815818,1.9308578,2.4967396,3.0386145,3.100347,1.9102802,1.8519772,1.8519772,1.7765263,1.7216529,1.99602,4.338428,4.8151407,4.249259,3.3266997,2.5961976,4.180667,3.882293,2.5961976,1.3375391,1.2312219,2.2326615,2.4590142,2.0063086,1.2826657,1.0117283,1.1214751,1.2826657,2.9906003,6.0566516,8.608265,8.669997,8.872343,7.4353456,4.9591837,4.40702,3.1243541,4.804852,9.921797,15.762384,16.420864,18.386019,15.824117,11.63659,8.1384115,7.0478024,5.9812007,5.686256,6.355026,7.1266828,6.0737996,5.2987127,4.40359,4.434457,5.7239814,7.874333,8.992378,9.544542,9.14328,8.296172,8.429926,12.161317,10.655728,6.636252,2.7539587,1.6187652,5.9571934,9.860064,11.712041,10.034973,3.4810312,3.0626216,5.2506986,7.1198235,7.0546613,4.746549,3.2375305,9.194724,14.71636,14.983868,8.237869,11.80464,13.927555,11.22161,6.427047,8.385342,10.563129,10.714031,8.690575,5.535354,3.4776018,2.8294096,3.9886103,5.9331865,6.6465406,3.1037767,9.619993,13.622321,11.245617,5.703404,7.298162,9.31133,6.7391396,5.206114,6.1046658,6.6122446,2.702515,7.606825,11.821788,11.382801,7.8606143,8.81404,13.344524,14.654627,11.050131,5.926327,5.2575574,10.916377,16.156786,18.255693,18.488907,17.309128,19.442331,22.988525,26.136887,27.162333,30.657082,29.199507,30.221525,36.81319,47.71585,36.33991,27.169191,21.60983,19.178253,17.501184,16.530611,11.849225,7.2158523,4.3590055,2.9906003,2.4590142,1.4644338,1.0871792,1.2106444,0.5144381,1.1523414,1.4987297,1.4095604,1.1111864,1.1832076,0.64819205,0.8265306,1.4815818,2.2086544,2.4555845,1.6427724,1.2380811,1.3649758,2.4384367,5.178677,5.8680243,5.192395,5.1683884,5.919468,5.689686,3.782835,3.309552,3.7862647,4.7774153,5.885172,4.420738,3.3198407,2.8705647,3.4604537,5.5902276,7.407909,8.045813,7.431916,6.5333643,7.3564653,7.281014,7.7920227,7.9429245,7.14726,5.171818,4.99005,5.8200097,5.4084597,3.673088,2.6922262,1.879414,1.2483698,1.0494537,1.1592005,1.0768905,0.84367853,0.53501564,0.35324752,0.36353627,0.5144381,0.5624523,0.5041494,0.50757897,0.5590228,0.48357183,0.3841138,0.31552204,0.2469303,0.16462019,0.08573969,0.08573969,0.15090185,0.14061308,0.058302987,0.030866288,0.07888051,0.12346515,0.16462019,0.28465575,0.6756287,1.4507155,1.3409687,1.0254467,0.9362774,1.2655178,1.903421,2.8877127,3.199805,2.9665933,3.4535947,3.275256,3.357566,2.7951138,1.5776103,0.5796003,0.6927767,0.7682276,0.64133286,0.32581082,0.037725464,0.07545093,0.041155048,0.020577524,0.33266997,1.5124481,1.0528834,0.91227025,0.6036074,0.15090185,0.10288762,0.072021335,0.05144381,0.06859175,0.1371835,0.26064864,0.82996017,0.7339317,0.65505123,0.8676856,1.2380811,1.0185875,0.7613684,0.53844523,0.45270553,0.6207553,1.0528834,1.4747226,1.8725548,2.2326615,2.534465,2.952875,3.5016088,4.307562,5.1409516,5.442755,3.8034124,3.6010668,3.8857226,3.9954693,3.5873485,6.56766,6.9380555,6.2555676,5.353586,4.3281393,2.4212887,1.1454822,0.8025235,1.2380811,1.8588364,1.5501735,0.91569984,0.34295875,0.106317215,0.36010668,0.7956643,0.75450927,0.4424168,0.106317215,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.0,0.006859175,0.017147938,0.017147938,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.082310095,0.044584636,0.024007112,0.020577524,0.037725464,0.08916927,0.12346515,0.3018037,0.72364295,1.2346514,1.4232788,1.0768905,0.58645946,0.21263443,0.05144381,0.006859175,0.006859175,0.0034295875,0.010288762,0.05144381,0.16119061,0.42869842,0.6824879,0.8471081,0.9259886,0.9877212,1.0082988,0.96714365,0.90541106,0.8848336,0.9842916,1.1249046,1.1008976,0.823101,0.4355576,0.28122616,0.33952916,0.42183927,0.5144381,0.61046654,0.7305021,0.8265306,0.91227025,0.97057325,0.980862,0.9259886,0.6893471,0.66876954,0.71678376,0.70649505,0.5418748,0.5007198,0.47328308,0.47671264,0.4972902,0.48014224,0.7579388,0.90541106,0.97057325,0.9362774,0.7133542,0.58988905,0.59331864,0.66191036,0.77165717,0.9259886,0.9431366,0.9431366,1.1111864,1.3409687,1.2312219,1.214074,1.2826657,1.3615463,1.3512574,1.1592005,1.039165,0.805953,0.5693115,0.42526886,0.47328308,0.45613512,0.52815646,0.66191036,0.83681935,1.0082988,1.2620882,1.3649758,1.4164196,1.5227368,1.7662375,1.5741806,1.4267083,1.2826657,1.1729189,1.1900668,1.3066728,1.3684053,1.4027013,1.4335675,1.4610043,1.7182233,2.1674993,2.5584722,2.7128036,2.5207467,2.153781,1.8245405,1.5501735,1.3478279,1.2346514,1.1180456,0.97400284,0.83338976,0.72707254,0.6790583,0.6344737,0.66533995,0.6927767,0.7510797,0.97057325,1.1180456,1.1660597,1.2449403,1.3889829,1.5433143,1.7388009,1.9514352,2.2120838,2.5996273,3.2272418,3.7725463,3.6285036,3.2649672,2.9185789,2.5653315,2.952875,3.292404,3.4638834,3.4398763,3.3026927,3.3472774,3.4981792,3.6593697,3.6970954,3.457024,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.05144381,0.0548734,0.024007112,0.061732575,0.13375391,0.28122616,0.6036074,1.2620882,4.201245,4.715683,3.6696587,2.0406046,0.9294182,0.58988905,0.607037,0.83681935,1.0906088,1.1180456,1.9857311,5.7239814,7.8606143,7.750868,8.584257,10.100135,13.965281,18.773561,22.652426,23.290329,20.718138,15.22051,10.772334,9.259886,10.463672,7.250148,5.254128,3.8891523,2.7985435,1.8691251,2.1915064,2.311542,2.2292318,2.1674993,2.5447538,2.668219,2.4452958,2.411,2.767677,3.4055803,3.5290456,4.712253,8.796892,13.649758,13.152468,20.505503,31.830002,39.879242,41.49458,37.59514,34.066093,34.728004,35.41392,33.805443,29.43272,37.128716,38.795494,39.718052,44.313698,56.132057,55.29181,55.161484,48.418915,35.053814,22.357481,19.668684,13.05301,8.39563,9.033533,15.721229,12.46312,7.829748,5.161529,5.6793966,8.491658,9.595985,9.517105,10.028113,10.635151,8.601405,5.6965446,4.0503426,3.7451096,4.6676683,6.5299344,7.4044795,6.1629686,4.5339146,3.2992632,2.318401,1.8588364,1.9068506,4.0503426,6.3035817,3.0797696,1.0871792,0.99801,1.7147937,2.5481834,3.216953,4.0777793,5.4804807,6.8454566,7.455923,6.468202,6.5367937,7.058091,6.756287,5.411889,3.8720043,3.9028704,5.3227196,6.001778,5.586798,5.5250654,5.6999745,5.562791,5.686256,5.9983487,5.813151,6.094377,5.161529,4.722542,5.223262,5.8680243,5.0483527,4.976331,4.5510626,4.1155047,5.453044,8.011517,7.1061053,5.4324665,5.051782,7.380472,9.80862,7.3084507,4.9934793,5.0620713,6.8111606,4.0880685,4.280125,5.3330083,5.422178,2.952875,2.2292318,2.1640697,1.7971039,1.3375391,2.1880767,2.4727325,2.5653315,2.9563043,3.3026927,2.4384367,2.7093742,2.0508933,2.5241764,4.0229063,4.2595477,2.5721905,2.2395205,2.2223728,2.0063086,1.5913286,2.393852,2.6750782,2.253239,1.6667795,2.1743584,2.7368107,2.5138876,2.16064,2.1126258,2.5961976,2.9082901,2.2429502,1.8759843,2.2841053,3.1517909,4.40702,4.122364,3.957744,4.266407,4.0846386,5.744559,4.190956,2.194936,1.4027013,2.3081124,3.7279615,3.391862,2.2360911,1.2483698,1.4850113,2.2120838,2.0577524,2.7333813,4.32128,5.2747054,3.882293,3.9783216,4.266407,4.513337,5.5730796,4.448175,2.9940298,3.7725463,7.3598948,12.325937,18.71183,16.002455,11.214751,8.388771,8.56368,7.3701835,5.9880595,5.73427,6.293293,5.7068334,4.4516044,4.064061,4.4275975,5.960623,9.602845,10.9541025,11.365653,11.38966,9.990388,4.547633,4.064061,4.4516044,4.0709205,3.0454736,3.2512488,6.358455,6.697984,6.5367937,6.0052075,3.093488,4.245829,6.701414,6.4716315,3.9646032,3.9714622,2.8088322,5.9983487,9.095266,9.410788,6.029215,8.162418,11.382801,10.600855,6.948344,7.7748747,8.522525,9.469091,7.98065,4.8597255,4.3349986,3.8548563,3.9097297,4.6608095,5.0174866,2.6613598,10.172156,12.3533745,9.030104,4.3521466,6.7940125,6.475061,4.3624353,4.1600895,5.960623,6.258997,2.8088322,13.584596,19.384027,14.160767,5.0414934,10.264755,17.21996,16.87014,10.124143,7.8331776,7.582818,9.626852,11.482259,13.581166,19.288,19.812727,22.336903,25.245193,27.234354,27.35096,28.27352,27.145185,29.8477,37.574562,46.855022,35.82547,27.652763,23.218307,21.3629,18.866161,16.427725,11.705182,7.613684,5.1238036,3.2546785,2.1194851,1.4027013,1.1763484,1.138623,0.5693115,1.2998136,1.5193073,1.2998136,1.039165,1.4644338,0.7579388,1.3409687,2.085189,2.5173173,2.7985435,2.0508933,1.3752645,1.0117283,1.8313997,5.3398676,6.166398,6.2212715,7.2638664,8.477941,6.4579134,3.6970954,3.6696587,4.040054,4.3624353,6.0737996,4.5956473,2.8877127,2.270387,3.3850029,6.1904054,6.9517736,8.258447,8.536243,7.3701835,5.5113473,6.1732574,6.759717,7.06495,6.790583,5.5662203,4.763697,6.1458206,6.433906,5.1855364,4.8082814,2.4007113,1.2723769,1.0871792,1.3786942,1.5638919,1.1797781,0.72021335,0.3841138,0.23321195,0.20920484,0.30866286,0.3566771,0.44927597,0.5521636,0.52472687,0.39440256,0.34638834,0.33952916,0.30866286,0.14404267,0.10288762,0.14061308,0.1371835,0.07545093,0.041155048,0.041155048,0.06516216,0.08573969,0.16462019,0.42869842,1.7696671,1.5261664,0.939707,0.8265306,1.5981878,1.7113642,2.1057668,2.935727,3.841138,3.9440255,2.1332035,2.1057668,2.3424082,1.9274281,0.5658819,0.15090185,0.14061308,0.15776102,0.082310095,0.048014224,0.09602845,0.06516216,0.0548734,0.28465575,1.0666018,1.255229,0.6927767,0.24350071,0.18519773,0.20920484,0.15776102,0.09945804,0.09602845,0.15776102,0.26407823,0.78194594,0.69963586,0.59674823,0.7922347,1.3443983,1.5947582,1.2415106,0.823101,0.7339317,1.2312219,1.5364552,1.9274281,2.4452958,2.9082901,2.9048605,3.2203827,2.719663,2.6647894,3.2992632,3.8479972,3.210094,3.6765177,4.8425775,5.703404,4.671098,6.324159,7.023795,6.8111606,5.8405876,4.383013,3.309552,2.1572106,1.1729189,0.7613684,1.4815818,0.85739684,0.77851635,0.53501564,0.19548649,0.6207553,1.2723769,1.2998136,0.83338976,0.2194936,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.020577524,0.048014224,0.07888051,0.22292319,0.5796003,1.0494537,1.3341095,1.0700313,0.65848076,0.30866286,0.10288762,0.020577524,0.017147938,0.006859175,0.006859175,0.024007112,0.058302987,0.2777966,0.6036074,0.8162418,0.89855194,1.0425946,1.0768905,1.1043272,1.0700313,1.0014396,0.9945804,1.2037852,1.4198492,1.1592005,0.548734,0.31895164,0.29837412,0.26750782,0.3566771,0.5453044,0.6756287,0.52815646,0.6241849,0.764798,0.8265306,0.7613684,0.58302987,0.70649505,0.7888051,0.72364295,0.6344737,0.48357183,0.5212973,0.58302987,0.58645946,0.5555932,0.59674823,0.59331864,0.65162164,0.7407909,0.69963586,0.58645946,0.5418748,0.5555932,0.6241849,0.70649505,0.7407909,0.8676856,1.1454822,1.3821237,1.1249046,0.96714365,0.980862,1.138623,1.3169615,1.3066728,1.313532,1.1351935,0.8196714,0.52815646,0.5521636,0.6344737,0.83338976,1.0494537,1.1660597,1.0254467,1.1694894,1.2998136,1.4061309,1.5193073,1.7010754,1.3615463,1.196926,1.0940384,1.0220171,1.0357354,1.1626302,1.3101025,1.4198492,1.4918705,1.5913286,1.7250825,1.9925903,2.253239,2.3664153,2.170929,1.7936742,1.5124481,1.3306799,1.2312219,1.1729189,0.9431366,0.7305021,0.59674823,0.548734,0.5658819,0.53501564,0.58988905,0.6001778,0.5796003,0.6756287,0.7682276,0.939707,1.155771,1.3992717,1.6496316,1.8039631,1.879414,2.0234566,2.3732746,3.0317552,3.6936657,3.542764,3.1655092,2.760818,2.1469216,2.8499873,3.2203827,3.333559,3.2958336,3.2512488,3.175798,3.333559,3.474172,3.4604537,3.2683969,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.09602845,0.2194936,0.28122616,0.12346515,0.15776102,0.18519773,0.38754338,1.0940384,2.7779658,5.744559,5.861165,4.417309,2.5310357,1.1763484,0.78537554,0.980862,1.5776103,2.0680413,1.6187652,1.9582944,4.4516044,6.807731,8.083538,8.683716,7.023795,13.838386,24.09971,30.063765,21.301168,15.614912,12.55229,10.847785,10.563129,13.077017,8.81747,5.7925735,3.673088,2.2258022,1.2963841,2.0303159,2.7985435,3.2306714,3.2786856,3.2032347,2.5070283,2.417859,2.9185789,3.7108135,4.2115335,5.662249,9.73317,15.63206,22.02824,27.069735,49.87992,73.4549,82.79367,73.16339,50.092556,46.175964,49.362053,47.48607,40.383392,39.868954,57.397575,51.601574,44.05305,47.149967,64.116135,61.615967,58.241253,51.8828,41.92328,29.26467,24.418663,17.357141,10.175586,6.1492505,9.750318,7.7748747,4.9248877,3.882293,6.4407654,13.533153,17.195951,14.915276,13.059869,12.583157,9.016385,7.6616983,6.327589,5.0140567,4.125794,4.4550343,6.773435,8.443645,7.1026754,3.6868064,2.4418662,1.1592005,1.9102802,2.435007,2.9700227,6.2418494,1.9925903,1.3615463,1.9411465,2.6785078,3.875434,5.5490727,7.73372,9.22902,9.22902,7.3255987,6.495639,6.9380555,7.596536,7.548522,5.994919,5.164959,5.9126086,6.2727156,5.830299,5.720552,6.1492505,6.1629686,6.3790326,6.924337,7.4627824,5.593657,3.5976372,2.633923,3.0489032,4.3795834,3.4021509,4.0846386,4.3521466,3.8548563,3.9508848,6.0532217,5.0312047,4.2835546,5.2301207,7.2947326,9.088407,7.5862474,6.358455,6.420188,6.2247014,4.870014,5.8508763,7.4970784,7.5931067,3.357566,2.270387,2.037175,1.5844694,1.0768905,1.9068506,2.3458378,2.503599,3.6970954,4.856296,2.486451,2.3767042,1.6084765,2.784825,5.2609873,5.127233,3.625074,3.724532,4.73969,5.2918534,3.3266997,5.0826488,6.0737996,5.113515,3.210094,3.5393343,3.2821152,2.3595562,1.9068506,2.2052248,2.6716487,3.4878905,2.2566686,1.7182233,2.9082901,5.1409516,3.9474552,3.9474552,4.695105,5.6245236,6.0875177,6.5162163,4.1772375,2.0474637,1.8313997,3.9680326,3.1140654,2.6716487,1.9548649,1.5604624,3.340418,5.4667625,4.8254294,3.2443898,1.9411465,1.5261664,1.0631721,1.5227368,1.3409687,1.5090185,5.5833683,8.611694,7.226141,4.338428,3.0111778,6.4544835,6.7974424,7.0923867,6.3618846,5.720552,8.3922,10.967821,10.6317215,8.268735,5.7068334,5.7068334,7.5382333,7.1061053,5.686256,5.3570156,9.016385,14.109323,13.5503,10.124143,6.036074,2.8980014,2.287535,2.4487255,3.4055803,6.094377,12.343085,9.623423,5.1512403,3.8342788,5.096367,2.8980014,7.438775,11.430815,9.527394,3.3712845,1.6016173,4.8734436,9.15014,10.072699,7.2878733,4.4550343,6.3721733,7.5107965,7.3873315,6.6053853,6.835168,6.7631464,7.870903,8.536243,7.9120584,5.936616,7.3873315,7.6788464,7.490219,6.543653,3.6010668,4.6265135,5.020916,3.981751,2.2292318,1.9823016,1.3752645,0.75450927,3.666229,8.457363,8.285883,4.9523244,21.843042,29.521889,19.507494,4.273266,21.009653,35.24244,32.769707,18.001905,13.96185,13.680624,16.383139,16.62321,14.586036,16.112202,20.104242,21.688711,23.34863,25.52985,26.641035,26.61703,28.139765,32.217545,37.24532,39.018417,33.729992,30.670801,28.84626,26.18833,19.562366,16.21852,12.377381,9.1810055,6.6225333,3.5702004,1.3238207,0.67219913,0.7510797,0.91227025,0.71678376,1.4267083,1.5741806,1.2826657,0.9294182,1.1592005,0.9534253,1.430138,1.8416885,2.2978237,3.799983,2.651071,1.862266,1.1832076,0.70306545,0.823101,2.3149714,4.4516044,6.914048,9.801761,13.670336,7.7748747,5.888602,5.1340923,4.4721823,4.729401,3.8891523,2.9906003,2.568761,3.2958336,5.9812007,5.9812007,6.475061,7.599966,7.939495,4.547633,5.950334,6.468202,7.205563,7.689135,5.857735,4.479041,5.1683884,5.9434752,6.1904054,6.6533995,3.100347,1.3512574,0.85739684,1.1626302,1.9068506,0.7099246,0.65162164,0.5761707,0.2194936,0.18176813,0.29151493,0.37382504,0.36353627,0.30523327,0.36696586,0.40126175,0.31895164,0.33952916,0.4115505,0.22978236,0.16804978,0.14404267,0.13032432,0.116605975,0.09259886,0.030866288,0.024007112,0.041155048,0.06516216,0.07545093,1.9308578,2.2292318,1.5364552,0.7442205,1.097468,1.3684053,1.6530612,2.2463799,2.7333813,2.0131679,1.3684053,1.4987297,2.2052248,2.5927682,1.0666018,0.21263443,0.017147938,0.030866288,0.037725464,0.061732575,0.061732575,0.05144381,0.13032432,0.22635277,0.09259886,1.1763484,0.66191036,0.15090185,0.17147937,0.18176813,0.18176813,0.1371835,0.15433143,0.24007112,0.29151493,0.6790583,0.99801,1.0906088,1.0254467,1.097468,1.4781522,1.8005334,1.7079345,1.6359133,2.8088322,2.6133456,2.5001693,2.7985435,2.9906003,1.7079345,3.4295874,2.935727,1.6599203,0.78537554,1.2346514,1.4198492,2.177788,3.974892,5.7582774,4.99005,4.465323,5.7239814,6.3721733,6.1286726,6.835168,5.528495,3.9303071,2.3081124,1.039165,0.6241849,0.83338976,0.90198153,0.6344737,0.25378948,0.4115505,1.2312219,0.8745448,0.58988905,0.5796003,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06859175,0.24007112,0.6001778,1.2346514,1.2346514,0.9431366,0.59674823,0.3018037,0.044584636,0.020577524,0.01371835,0.01371835,0.020577524,0.044584636,0.16804978,0.34638834,0.5521636,0.77508676,1.0082988,1.1180456,1.097468,1.0082988,0.90884066,0.8848336,1.2037852,1.6564908,1.5227368,0.84367853,0.4424168,0.33266997,0.32238123,0.39783216,0.4664239,0.3806842,0.42869842,0.77165717,0.864256,0.6379033,0.5041494,0.490431,0.67219913,0.6962063,0.53844523,0.48700142,0.4629943,0.7339317,0.90884066,0.922559,1.0082988,0.77508676,0.5418748,0.4629943,0.52815646,0.5658819,0.58988905,0.5418748,0.5521636,0.6241849,0.61046654,0.58645946,0.72707254,0.94656616,1.1249046,1.1146159,1.0048691,0.9842916,1.1866373,1.488441,1.5261664,1.3684053,0.980862,0.7099246,0.66191036,0.6859175,0.7613684,1.0700313,1.3032433,1.3066728,1.097468,1.2312219,1.3684053,1.3684053,1.2483698,1.1763484,0.90541106,0.82996017,0.89855194,1.0357354,1.1454822,1.1934965,1.4267083,1.5844694,1.6496316,1.845118,1.7971039,1.8416885,1.9514352,2.0714707,2.1194851,1.8519772,1.546744,1.2963841,1.1489118,1.097468,0.9294182,0.70306545,0.53844523,0.4664239,0.4424168,0.490431,0.51100856,0.4698535,0.4046913,0.4424168,0.52815646,0.6241849,0.82996017,1.1351935,1.4027013,1.4027013,1.430138,1.4541451,1.5536032,1.9068506,2.1880767,2.0749004,1.7525192,1.5947582,2.1812177,3.0111778,3.357566,3.4604537,3.4947495,3.5564823,3.532475,3.450165,3.4467354,3.426158,3.0969174,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.15776102,0.31552204,0.44584638,0.35324752,0.23321195,0.39097297,1.4027013,3.4638834,6.3790326,8.241299,7.257007,5.209543,3.2821152,2.054323,1.097468,0.8128122,1.1592005,1.8279701,2.2635276,4.852866,6.2727156,7.5450926,8.827758,9.427936,5.8234396,8.690575,16.177364,22.336903,17.12736,16.263103,15.776102,13.745787,10.81006,10.158438,7.64798,5.5662203,3.6765177,2.4384367,2.9940298,2.8945718,2.9803114,3.1723683,3.1860867,2.5584722,2.9151495,4.911169,7.0718093,9.129561,12.010415,11.101575,11.797781,19.919044,33.26357,41.607754,58.309845,89.258446,109.82225,104.506386,66.96269,56.931152,53.024853,47.79473,42.187355,45.520916,57.222668,50.44237,42.067318,42.434284,55.329536,51.265472,47.64726,42.458294,34.24786,22.12427,16.71238,12.46312,7.56224,3.8479972,6.783724,22.295748,17.302269,7.5416627,3.7039545,11.410237,16.928444,12.175035,6.6293926,4.149801,2.976882,2.568761,2.2806756,2.0714707,2.0714707,2.5893385,3.1586502,3.6010668,3.8685746,3.6044965,2.136633,1.6942163,2.2738166,3.7862647,5.895461,8.035523,4.2938433,2.9185789,3.1517909,4.057202,4.5099077,5.23698,6.252138,7.514226,8.697433,9.205012,7.006647,6.368744,6.691125,7.133542,6.6053853,7.641121,9.671436,10.2921915,9.321619,8.820899,9.006097,7.5690994,7.466212,9.163857,10.659158,7.689135,5.144381,3.6593697,3.74168,5.796003,3.82399,3.7108135,4.245829,4.6882463,4.804852,5.3741636,4.0194764,3.782835,5.1992545,6.3035817,7.6788464,5.8234396,4.372724,4.537344,5.103226,3.6387923,4.07435,5.3501563,5.6245236,2.2600982,2.294394,3.292404,3.5359046,2.7779658,2.2600982,2.7882545,4.190956,6.012067,6.7665763,3.940596,2.287535,1.7388009,2.4590142,3.4947495,2.784825,3.0283258,3.3850029,3.8445675,3.9063,2.5584722,4.170378,4.791134,3.6044965,1.6976458,2.0749004,1.9068506,1.6633499,1.8382589,2.3801336,2.7059445,2.3629858,2.0097382,2.085189,2.5893385,3.117495,3.3061223,2.7333813,2.5447538,3.1552205,4.245829,4.866585,3.7519686,3.1037767,3.799983,5.3707337,3.6182148,3.0248961,3.5804894,4.671098,5.086078,5.0243454,3.6970954,2.2738166,1.4027013,1.2209331,2.1126258,1.5433143,0.805953,1.1317638,3.7039545,12.579727,13.625751,9.990388,5.305572,3.673088,7.1095347,6.166398,4.623084,4.8117113,7.623973,10.628291,12.950122,10.7586155,6.0737996,6.7700057,8.501947,6.9620624,6.451054,8.303031,10.909517,14.455711,11.293632,6.574519,3.415869,2.8739944,4.6265135,6.2418494,7.2124224,8.543102,12.723769,10.635151,5.0140567,2.5756202,4.4413157,6.108095,10.816919,14.191633,11.334786,4.2252517,1.7250825,6.7940125,8.81061,7.2158523,4.4721823,6.042933,9.355915,7.8331776,6.5985265,9.448513,18.8593,16.811838,11.650309,7.963502,6.5299344,4.2869844,3.690236,6.615674,7.939495,6.046363,2.8328393,9.678296,14.7026415,13.711491,7.723431,2.9974594,1.2037852,1.6016173,4.835718,8.745448,8.371623,10.398509,20.598103,21.767591,11.88352,4.0880685,25.485264,45.349434,46.848164,31.192099,17.658945,13.649758,12.548861,11.7086115,10.906088,12.3533745,18.924463,22.930222,24.151155,23.588703,23.478956,25.125158,25.375517,27.772799,31.84372,33.09552,32.91718,30.482174,26.339231,21.493225,17.412016,14.448852,12.88839,11.746337,9.815479,5.669108,2.4761622,1.0220171,0.6241849,0.65505123,0.5453044,0.97057325,1.1729189,1.1111864,0.9842916,1.2449403,1.3786942,1.6359133,1.4198492,1.4541451,3.7862647,3.117495,2.0817597,1.2620882,0.7613684,0.20234565,0.881404,2.2909644,4.0846386,5.8234396,6.958633,7.2158523,5.9880595,6.3961806,7.922347,6.3893213,3.3712845,3.7965534,4.1429415,3.4776018,3.4776018,4.5339146,6.48535,7.438775,6.7494283,5.0346346,5.4153185,5.5559316,5.9812007,6.324159,5.3330083,4.149801,4.5819287,5.137522,5.23698,5.212973,3.6627994,2.7128036,1.5947582,0.5658819,0.91912943,0.64133286,0.5590228,0.4629943,0.29151493,0.15776102,0.17147937,0.22978236,0.26064864,0.28465575,0.41498008,0.42183927,0.3841138,0.3841138,0.40126175,0.32581082,0.14747226,0.09602845,0.116605975,0.15090185,0.12689474,0.058302987,0.041155048,0.05144381,0.15090185,0.5144381,2.3321195,2.7985435,1.9239986,0.5693115,0.41498008,0.96714365,1.8965619,2.1983654,1.8142518,1.611906,2.253239,1.2929544,0.6893471,0.8505377,0.65162164,0.17833854,0.10288762,0.1371835,0.13375391,0.061732575,0.030866288,0.01371835,0.0548734,0.17833854,0.3841138,0.33952916,0.16119061,0.09945804,0.18519773,0.25721905,0.15776102,0.17490897,0.23321195,0.53844523,1.5844694,3.4878905,2.469303,1.2689474,1.2895249,2.6133456,2.4727325,3.6113555,4.4859004,4.448175,3.7348208,3.6079261,2.4418662,1.9514352,3.2718265,6.9689217,5.7308407,3.9783216,2.2155135,1.1043272,1.4678634,0.7510797,2.7230926,4.787704,5.9640527,6.893471,5.754848,5.1169443,4.9488945,5.271276,6.1629686,3.7759757,2.2429502,2.1263442,2.702515,1.9548649,0.71678376,0.28122616,0.22292319,0.23664154,0.13032432,0.34295875,0.48357183,0.7613684,0.881404,0.017147938,0.061732575,0.07888051,0.05144381,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.020577524,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.07545093,0.28808534,0.89512235,1.762808,2.177788,1.6633499,0.5727411,0.082310095,0.0274367,0.01371835,0.010288762,0.010288762,0.034295876,0.09602845,0.28808534,0.490431,0.6859175,0.9568549,1.0871792,1.0528834,0.97057325,0.9259886,0.97057325,1.1523414,1.4850113,1.6633499,1.5536032,1.2003556,0.8265306,0.70649505,0.67219913,0.59331864,0.3806842,0.42183927,0.5178677,0.52815646,0.490431,0.65162164,0.764798,0.8745448,0.77508676,0.5693115,0.64819205,0.45613512,0.5007198,0.72021335,0.9328478,0.823101,0.6310441,0.5178677,0.4355576,0.36696586,0.34638834,0.37039545,0.40126175,0.4629943,0.53844523,0.58645946,0.6893471,0.65505123,0.70306545,0.90541106,1.1866373,1.1660597,1.2346514,1.3032433,1.3341095,1.3443983,1.1249046,0.9294182,0.78194594,0.64133286,0.39440256,0.6036074,0.89855194,1.0666018,1.0631721,1.0117283,1.3238207,1.3272504,1.2620882,1.2243627,1.1489118,0.9877212,0.9774324,1.1283343,1.3684053,1.546744,1.9685832,1.9342873,1.7490896,1.6804979,1.9445761,2.1983654,2.2292318,2.3629858,2.6064866,2.644212,2.6716487,2.3424082,1.7559488,1.1523414,0.9294182,0.8162418,0.72021335,0.6207553,0.52472687,0.490431,0.432128,0.4424168,0.432128,0.39783216,0.39440256,0.48014224,0.58988905,0.7373613,0.90198153,1.0254467,1.0254467,1.0906088,1.1077567,1.0563129,0.9911508,1.1180456,1.3821237,1.7113642,2.1160555,2.6819375,3.0454736,3.1826572,3.340418,3.666229,4.214963,3.6525106,3.357566,3.2443898,3.1792276,2.976882,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.13375391,0.21263443,0.24350071,0.24007112,0.2469303,0.34638834,1.5913286,3.7691166,6.3653145,8.577398,10.14472,9.496528,7.1987042,4.3590055,2.6579304,1.3032433,0.89169276,1.3889829,2.4624438,3.4776018,5.926327,7.939495,9.400499,10.028113,9.410788,6.807731,8.841476,14.30481,19.20912,16.777542,17.147938,15.902997,13.7938,11.880091,11.55428,7.81603,6.1904054,5.0106273,3.923448,3.875434,3.4467354,3.858286,3.9440255,3.6765177,4.15323,6.210983,8.285883,9.8429165,11.255906,13.797231,10.443094,14.407697,29.854559,50.274323,58.498474,60.892326,82.749084,99.660385,95.27737,61.324455,52.38352,47.424335,42.48916,37.9038,38.267338,44.985897,44.47832,41.796383,40.602886,43.171646,38.09929,37.24532,34.227283,26.699339,16.37628,14.095605,12.144169,8.124693,4.197815,7.085528,23.478956,25.132017,14.733508,2.3252604,5.284994,8.522525,8.2653055,6.7048435,5.055212,3.542764,2.7573884,2.294394,2.153781,2.287535,2.5790498,2.0749004,1.6976458,2.054323,2.843128,2.8465576,3.1723683,3.7931237,5.192395,7.3221693,9.599416,6.7940125,5.6793966,5.6348124,5.8988905,5.5662203,4.962613,5.1580997,5.926327,6.917478,7.6685576,6.001778,5.744559,5.9434752,6.1149545,6.2658563,7.0203657,9.054111,9.798331,9.283894,10.120712,10.388221,10.408798,10.288762,10.686595,12.823228,10.134431,8.608265,7.140401,5.844017,6.0497923,4.479041,3.8445675,4.5510626,6.138962,7.2707253,6.2247014,4.4413157,3.6147852,4.465323,6.7528577,5.7891436,4.197815,3.2512488,3.4433057,4.5030484,3.5016088,4.2286816,5.950334,6.6739774,3.1277838,2.1400626,2.5447538,3.9886103,4.938606,2.6785078,2.3629858,3.5187566,5.161529,6.001778,4.4584637,2.3389788,1.9754424,2.585909,3.1723683,2.534465,3.673088,3.0523329,2.8396983,3.3987212,3.2821152,3.0454736,4.0091877,3.5359046,2.0097382,2.8259802,2.8328393,1.903421,1.5330256,2.0337453,2.534465,1.7456601,1.7559488,1.9480057,2.0508933,2.1434922,2.5619018,2.16064,2.0508933,2.644212,3.6456516,3.1037767,2.3218307,2.3835633,3.4638834,4.835718,3.5221863,3.100347,3.2546785,3.5187566,3.2992632,2.702515,1.8142518,1.1523414,1.6427724,4.5956473,4.6127954,2.7402403,1.430138,2.085189,5.0655007,13.924125,12.912396,7.874333,3.450165,3.059192,6.7940125,7.006647,6.7665763,7.682276,9.911508,11.331357,10.796341,9.22216,8.179566,9.880642,11.187314,9.644,8.759167,9.911508,12.343085,12.435684,9.081548,5.4324665,3.1449318,2.3389788,5.40503,7.8331776,8.093826,7.56567,10.539123,7.716572,4.256118,4.232111,7.0272245,7.332458,8.032094,9.15014,7.473071,3.5770597,1.8279701,8.786603,10.017825,7.1232533,4.2423997,8.05953,10.762046,6.9620624,5.3673043,9.918367,19.78872,15.182784,8.419638,4.8082814,4.722542,3.5633414,8.018375,12.123591,10.72089,4.8734436,1.8519772,8.182996,11.694893,10.22703,5.429037,2.784825,3.1655092,4.139512,5.4941993,6.478491,5.802862,10.549411,18.45461,18.722118,11.30735,6.9380555,25.35837,42.24909,43.62778,30.495892,18.821575,15.433144,16.009314,16.595774,16.225378,16.942162,22.913074,25.492125,24.470106,21.561817,20.402617,22.758743,22.419212,22.919933,25.097721,27.09374,28.77081,28.959436,26.898254,23.256033,20.135109,16.46888,14.387119,13.145609,11.873232,9.56512,5.0655007,2.5173173,1.3512574,0.90541106,0.4389872,0.94656616,1.1763484,1.0871792,0.85739684,0.85396725,1.1043272,1.762808,1.9480057,1.8725548,2.860276,1.9891608,1.7319417,1.4644338,1.2620882,1.9137098,6.169828,4.2595477,2.277246,2.4658735,3.210094,4.170378,3.9474552,5.3158607,7.891481,8.131552,4.2081037,3.4810312,3.8034124,3.8857226,3.3026927,3.7553983,5.429037,6.3138704,5.9400454,5.3501563,5.422178,5.422178,5.768566,6.036074,4.9831905,4.420738,4.040054,3.858286,3.6970954,3.175798,3.0489032,2.7951138,1.879414,0.7990939,1.0940384,0.58302987,0.45956472,0.40126175,0.2777966,0.12346515,0.09945804,0.18519773,0.24350071,0.25721905,0.34638834,0.36010668,0.3806842,0.35324752,0.28122616,0.24007112,0.106317215,0.058302987,0.072021335,0.106317215,0.1097468,0.08916927,0.09945804,0.1097468,0.39440256,1.5501735,3.5976372,3.5187566,2.2498093,1.0666018,1.5638919,3.0557625,3.549623,3.4878905,3.4192986,4.0194764,4.029765,2.6304936,1.1866373,0.39783216,0.31209245,0.26407823,0.2194936,0.33952916,0.4629943,0.12346515,0.030866288,0.08573969,0.30523327,0.4972902,0.2469303,0.06516216,0.030866288,0.116605975,0.22635277,0.20234565,0.13032432,0.16119061,0.28465575,0.90884066,2.8396983,4.729401,3.6456516,1.8245405,0.8505377,1.6804979,2.7745364,4.0846386,4.7945633,4.400161,2.702515,2.5413244,2.3218307,1.8313997,2.0234566,4.99005,4.5510626,3.4707425,2.750529,2.8396983,3.6147852,3.0111778,4.5647807,6.2075534,6.8454566,6.355026,5.360445,4.1326528,4.3452873,5.9434752,7.140401,4.4927597,2.0406046,1.8382589,3.275256,3.0660512,1.2415106,0.32924038,0.07545093,0.14061308,0.07888051,0.58645946,0.6859175,0.66876954,0.53844523,0.024007112,0.06516216,0.09259886,0.06516216,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.106317215,0.39783216,0.96371406,1.3478279,1.1900668,0.6036074,0.20234565,0.082310095,0.030866288,0.01371835,0.010288762,0.01371835,0.0548734,0.1920569,0.37382504,0.5727411,0.77165717,0.9294182,0.97057325,0.9431366,0.90198153,0.9294182,1.0734608,1.2758065,1.4644338,1.529596,1.3341095,1.0837497,1.0014396,0.9362774,0.823101,0.66533995,0.6207553,0.45613512,0.3566771,0.45270553,0.823101,0.8745448,0.8676856,0.7888051,0.71678376,0.7956643,0.58645946,0.5418748,0.66876954,0.77508676,0.47671264,0.4115505,0.44584638,0.4424168,0.3841138,0.35324752,0.31209245,0.36353627,0.42869842,0.4629943,0.4424168,0.5041494,0.47328308,0.5212973,0.6790583,0.85739684,0.97400284,1.1111864,1.1866373,1.1866373,1.1866373,0.9328478,0.7682276,0.70306545,0.65848076,0.4664239,0.6001778,0.8265306,0.97400284,1.0323058,1.138623,1.2792361,1.3272504,1.2312219,1.0425946,0.9328478,1.0048691,1.2003556,1.4232788,1.605047,1.7216529,2.270387,2.3286898,2.2086544,2.1674993,2.3972816,2.7882545,2.9940298,3.07634,3.0351849,2.8225505,2.942586,2.7951138,2.194936,1.3478279,0.8676856,0.71678376,0.64819205,0.58988905,0.52472687,0.5041494,0.432128,0.4424168,0.45956472,0.48014224,0.5555932,0.59674823,0.65505123,0.7339317,0.8265306,0.90198153,0.9774324,1.0185875,1.0460242,1.0666018,1.1008976,1.2106444,1.5021594,2.0097382,2.5824795,2.9082901,2.836269,2.843128,2.884283,3.0077481,3.3266997,3.1072063,3.0111778,2.9391565,2.8499873,2.74367,0.017147938,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.17147937,0.25721905,0.28808534,0.28465575,0.2709374,0.5007198,2.5207467,5.5113473,8.515666,10.432805,11.701753,11.153018,8.327039,4.417309,2.2669573,1.2689474,1.1214751,1.762808,3.0111778,4.5647807,5.9469047,7.675417,9.386781,10.209882,8.783174,7.5862474,9.956093,14.246507,17.768692,16.79126,16.20137,14.946142,14.085316,13.63261,12.548861,7.8846216,6.341307,5.456474,4.3521466,3.7485392,5.1821065,5.9880595,5.1821065,3.8925817,5.3570156,8.1212635,9.914937,11.540562,13.495427,15.988737,13.9481325,18.752985,35.91464,57.8057,63.67029,56.70137,64.071556,71.04391,67.477135,47.822166,41.92671,38.373653,35.22872,31.799135,28.654203,30.489033,33.640823,35.791176,35.787746,33.647682,28.60276,28.619907,26.805656,20.752434,12.535142,11.910957,10.943813,7.98408,5.0174866,7.641121,19.6241,24.415234,16.894148,3.865145,4.033195,4.1635194,5.9880595,7.0958166,6.6225333,5.2335505,3.7313912,2.527606,2.0234566,2.1023371,2.1091962,1.7525192,1.2586586,1.313532,2.085189,3.2203827,4.2526884,4.897451,5.6005163,6.8043017,8.947794,8.292743,7.73029,7.486789,7.298162,6.3893213,4.746549,4.266407,4.3692946,4.602506,4.6402316,4.057202,4.3487167,4.530485,4.650521,5.7891436,6.358455,7.7680154,8.268735,8.200144,9.9801,11.55771,12.860953,12.744347,12.068718,13.697772,13.275933,13.677195,12.744347,10.100135,7.160979,5.7994323,4.770556,5.130663,6.560801,7.3839016,6.427047,4.8185706,3.9131594,4.4516044,6.5333643,4.32471,3.433017,3.1483612,3.216953,3.8548563,3.350707,4.396731,6.2247014,7.082098,4.2218223,2.1983654,1.9548649,3.57363,5.164959,2.867135,1.9445761,2.4041407,3.3815732,4.1120753,3.9165888,3.2855449,2.7882545,2.9288676,3.5153272,3.6765177,4.057202,2.651071,2.3424082,3.532475,4.1120753,3.059192,4.9180284,5.3090014,3.7313912,3.5461934,3.2958336,2.2429502,2.0063086,2.5893385,2.3801336,1.7730967,1.8862731,2.0920484,2.2635276,2.7882545,2.8396983,2.3561265,2.2566686,2.7333813,3.2615378,2.0234566,1.903421,2.6236343,3.649081,4.170378,3.5016088,3.2855449,2.8980014,2.1915064,1.4987297,1.138623,0.8779744,1.2277923,3.0523329,7.5690994,5.686256,3.3781435,2.568761,3.642222,5.4633327,11.084427,8.1384115,3.841138,1.9068506,2.5207467,4.3761535,6.368744,7.5039372,7.939495,8.964942,9.31133,7.274155,7.0478024,9.496528,12.147599,13.145609,11.938394,10.63858,10.607714,12.466551,10.117283,7.250148,4.804852,3.1346428,1.9823016,4.671098,6.557371,6.667118,5.90232,7.040943,4.671098,3.7794054,6.866034,11.156448,8.597976,5.6176643,6.852316,7.3084507,5.130663,1.5707511,9.1810055,10.179015,7.3530354,4.835718,8.090397,10.172156,5.926327,4.307562,8.351046,15.172495,10.813489,5.785714,3.3850029,3.7622573,3.9371665,13.485138,17.302269,13.042721,4.420738,1.2037852,5.552502,7.4113383,6.036074,3.117495,2.7642474,5.0243454,5.693115,5.103226,4.2218223,4.636802,8.841476,13.594885,14.260224,11.153018,9.517105,20.303158,29.298965,30.495892,24.888515,20.45406,15.933864,17.415445,19.658396,19.997925,18.3723,22.721018,23.667583,22.148275,20.066517,20.28601,22.12427,21.846472,22.919933,25.896814,28.43128,28.657633,28.218645,27.1932,25.293207,21.880768,18.067066,14.846684,13.214201,13.128461,13.512574,8.56368,4.7328305,2.3732746,1.3306799,0.922559,1.2723769,1.4129901,1.2243627,0.8196714,0.548734,0.86082643,1.7216529,2.1572106,2.07833,2.2669573,1.5673214,1.5947582,1.6393428,1.6427724,2.2052248,6.39961,4.372724,1.6084765,0.6859175,1.2998136,1.6736387,2.2909644,3.9851806,6.4887795,8.419638,5.6793966,3.649081,3.4776018,4.6402316,4.9180284,4.290414,4.513337,4.5853586,4.341858,4.4584637,4.7259717,4.9694724,5.3158607,5.521636,5.007198,4.6402316,4.125794,3.549623,2.8945718,2.0234566,2.1503513,2.1194851,1.6153357,0.9294182,0.9534253,0.53844523,0.44584638,0.37039545,0.216064,0.11317638,0.072021335,0.13375391,0.18862732,0.216064,0.28465575,0.33609957,0.39440256,0.35324752,0.23321195,0.16804978,0.10288762,0.07888051,0.07545093,0.082310095,0.09602845,0.106317215,0.116605975,0.1371835,0.67219913,2.7402403,4.5099077,4.046913,2.819121,2.1332035,3.1620796,4.496189,4.540774,4.166949,4.2286816,5.576509,5.3570156,3.6696587,1.7971039,0.53501564,0.19548649,0.2503599,0.2709374,0.42183927,0.548734,0.19891608,0.07888051,0.106317215,0.29837412,0.4629943,0.18519773,0.07545093,0.048014224,0.09602845,0.18519773,0.23664154,0.39097297,0.4115505,0.39440256,0.9568549,3.2135234,4.870014,4.122364,2.3458378,0.864256,0.9362774,2.0303159,2.8705647,3.2958336,2.9700227,1.3855534,1.5776103,1.9445761,1.7971039,1.4232788,2.085189,2.585909,2.5550427,3.4810312,5.1992545,5.895461,5.3261495,5.662249,6.5127864,6.9037595,5.2609873,5.4599032,4.448175,4.2526884,5.4633327,7.226141,5.206114,2.253239,1.3786942,2.5893385,2.8911421,1.3169615,0.4115505,0.072021335,0.106317215,0.20234565,0.94999576,0.88826317,0.5453044,0.23321195,0.048014224,0.044584636,0.06859175,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.116605975,0.29151493,0.5624523,0.7613684,0.7407909,0.37725464,0.16119061,0.061732575,0.0274367,0.017147938,0.0,0.020577524,0.09259886,0.23321195,0.41498008,0.5761707,0.7613684,0.83338976,0.8196714,0.77851635,0.7888051,0.9911508,1.1592005,1.3101025,1.4164196,1.4061309,1.3341095,1.2723769,1.2243627,1.1523414,0.9945804,0.7888051,0.48014224,0.34295875,0.4698535,0.7442205,0.7407909,0.78537554,0.8711152,0.9294182,0.84024894,0.6379033,0.5727411,0.6173257,0.6276145,0.35324752,0.4115505,0.48014224,0.5041494,0.48357183,0.45613512,0.40126175,0.4115505,0.4389872,0.42526886,0.33952916,0.3566771,0.36353627,0.4081209,0.48700142,0.5590228,0.7339317,0.89512235,0.9945804,1.0151579,0.9431366,0.78537554,0.7339317,0.72707254,0.69963586,0.5693115,0.6276145,0.7339317,0.8676856,1.0082988,1.1317638,1.2312219,1.2620882,1.1454822,0.9294182,0.823101,1.0460242,1.3272504,1.6221949,1.8965619,2.153781,2.527606,2.6922262,2.7573884,2.860276,3.1380725,3.5599117,3.9028704,3.9954693,3.7553983,3.1826572,3.07634,2.8911421,2.2635276,1.3443983,0.7922347,0.64819205,0.5796003,0.52472687,0.47671264,0.44927597,0.4355576,0.4698535,0.4972902,0.53844523,0.65848076,0.6824879,0.71678376,0.764798,0.8265306,0.91569984,1.1454822,1.2449403,1.2723769,1.3169615,1.4918705,1.6496316,1.8416885,2.2086544,2.6304936,2.7128036,2.5138876,2.5001693,2.4761622,2.3972816,2.3629858,2.4247184,2.49331,2.469303,2.3664153,2.335549,0.09945804,0.041155048,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.017147938,0.034295876,0.15776102,0.31552204,0.5007198,0.6173257,0.48700142,0.9259886,3.4295874,6.975781,10.350495,12.13731,12.22305,10.696883,7.250148,3.1449318,1.2037852,1.039165,1.2998136,1.9480057,3.1209247,5.130663,5.7102633,6.3790326,8.124693,9.770895,7.956643,7.157549,9.547972,13.248496,15.971589,15.0456,13.872682,14.808959,15.830976,15.237658,11.657167,8.282454,6.9620624,5.669108,4.1017866,3.6593697,6.9552035,7.459353,5.830299,4.2286816,6.341307,8.090397,10.779194,15.446862,20.4472,21.44521,21.009653,21.980227,33.781437,50.699593,51.86222,46.49492,44.780125,43.699802,41.2305,36.32276,32.553646,30.465025,28.619907,25.872808,21.35947,19.576086,21.44864,24.970827,27.892836,27.738503,23.184011,21.70929,20.111101,16.53747,10.449953,8.772884,7.5450926,5.9640527,4.8597255,6.711703,15.450292,16.564907,12.006986,6.5059276,7.596536,5.970912,5.579939,5.528495,5.3913116,5.223262,3.3438478,1.7216529,1.0288762,1.1317638,1.1180456,1.5227368,1.4232788,1.4918705,2.1263442,3.4467354,4.8322887,5.271276,5.2918534,5.56965,6.9552035,8.320179,8.124693,7.7714453,7.490219,6.3447366,4.554492,3.758828,3.2615378,2.719663,2.1469216,2.2806756,2.6990852,2.9185789,3.391862,5.4976287,6.8797526,7.390761,7.377043,7.6685576,9.547972,12.415107,13.694343,13.526293,12.761495,12.946692,14.898128,17.014183,17.477179,15.29253,10.30934,8.357904,6.660259,5.8234396,5.7136927,5.453044,5.9400454,4.9077396,4.5647807,5.2266912,5.302142,3.7211025,3.7862647,3.957744,3.6319332,3.1517909,2.8499873,3.9097297,5.3398676,5.9880595,4.530485,2.369845,2.0920484,2.8019729,3.415869,2.6545007,1.9754424,1.961724,2.2360911,2.6819375,3.4467354,4.434457,3.7039545,3.3266997,4.040054,5.24041,4.091498,2.4144297,2.3801336,3.8342788,4.3109913,3.8685746,6.046363,6.8797526,5.4804807,4.0434837,3.1415021,2.702515,3.2786856,4.0057583,2.6167753,2.3561265,2.411,2.6407824,3.1106358,4.0846386,3.7211025,3.0146074,2.6545007,2.6990852,2.5550427,1.6667795,2.3492675,3.5839188,4.420738,3.9954693,3.7794054,3.9337368,3.6593697,2.7402403,1.5741806,1.3752645,1.3101025,2.417859,4.9180284,8.224151,5.086078,3.5633414,3.7862647,4.629943,3.7348208,5.3673043,2.8294096,1.6084765,2.5756202,1.9823016,1.1866373,4.197815,6.355026,6.310441,6.0326443,5.8645945,5.113515,5.994919,8.7317295,11.540562,12.764925,12.38424,10.981539,9.777754,10.628291,7.966932,6.029215,4.273266,2.750529,2.0920484,4.420738,5.086078,5.2609873,5.038064,3.4364467,2.9185789,3.7108135,8.330468,13.128461,8.303031,5.099797,9.304471,11.8115,8.755736,1.5090185,9.187865,9.472521,7.4696417,6.420188,7.689135,9.280463,6.1972647,4.57507,6.3790326,9.379922,7.455923,5.4941993,4.173808,3.8171308,4.400161,14.2190695,16.7844,12.308789,4.698535,1.5638919,6.012067,7.9737906,6.660259,3.6765177,3.0214665,5.099797,4.856296,3.7108135,3.210094,5.0277753,6.8557453,7.380472,7.798882,8.721441,10.1652975,13.416546,14.243076,15.827546,18.900457,21.747015,14.695783,14.788382,17.384579,18.440891,14.534592,17.826996,18.927893,19.137098,19.86417,22.628418,22.885637,23.163433,26.579304,32.08722,34.477642,32.299854,29.151493,26.973705,25.296637,21.253153,18.073925,14.349394,12.634601,13.543441,15.748666,11.784062,6.9620624,3.3472774,1.8313997,2.1434922,1.9480057,1.8554068,1.546744,1.0288762,0.6241849,0.9534253,1.529596,1.7490896,1.7319417,2.3424082,2.5413244,2.201795,2.061182,1.978872,0.9294182,0.9774324,1.7525192,1.5055889,0.4389872,0.7339317,0.91227025,1.7422304,3.100347,4.8768735,6.9552035,6.7048435,4.5819287,3.9646032,5.453044,6.90033,5.669108,4.4996185,3.2855449,2.3561265,2.5001693,3.415869,4.2252517,4.5613513,4.5682106,4.9077396,4.647091,4.5647807,4.0537724,3.0351849,1.961724,1.646202,1.7250825,1.4507155,0.7922347,0.4424168,0.5590228,0.52815646,0.37039545,0.18862732,0.14747226,0.07888051,0.061732575,0.09945804,0.17833854,0.26750782,0.36010668,0.41840968,0.39097297,0.29151493,0.1920569,0.1371835,0.13375391,0.13375391,0.12346515,0.116605975,0.11317638,0.09259886,0.116605975,0.77851635,3.199805,4.2869844,4.0194764,3.2889743,2.9665933,3.8788633,4.0194764,4.1463714,3.8377085,3.7279615,5.4976287,5.7274113,3.9371665,2.037175,0.8848336,0.28122616,0.13375391,0.25378948,0.34981793,0.31895164,0.26750782,0.13032432,0.048014224,0.020577524,0.12689474,0.51100856,0.1920569,0.1371835,0.10288762,0.10288762,0.4081209,1.0220171,0.96714365,0.5796003,0.6962063,2.6579304,4.5201964,4.1772375,2.9288676,1.8656956,1.8691251,1.08032,1.1283343,1.646202,2.0165975,1.3581166,1.8965619,1.8176813,1.7936742,1.8279701,1.2895249,1.937717,2.5961976,4.5819287,7.0786686,7.130112,6.416758,5.9812007,5.936616,5.8543057,4.791134,6.2967224,5.830299,4.866585,4.698535,6.4407654,5.1238036,2.417859,0.9328478,1.214074,1.728512,1.0151579,0.39783216,0.09602845,0.13032432,0.3018037,0.8848336,0.7579388,0.41840968,0.15776102,0.06516216,0.024007112,0.034295876,0.044584636,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.030866288,0.01371835,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.11317638,0.24350071,0.5212973,0.8196714,0.91912943,0.51100856,0.24007112,0.1097468,0.05144381,0.024007112,0.0,0.0,0.024007112,0.10288762,0.24007112,0.4046913,0.59674823,0.66191036,0.65848076,0.64133286,0.65848076,0.939707,1.1249046,1.2449403,1.3478279,1.4781522,1.4678634,1.3992717,1.3889829,1.3786942,1.1351935,0.8093826,0.5521636,0.490431,0.5590228,0.5041494,0.59674823,0.8676856,1.1729189,1.2689474,0.8128122,0.6001778,0.548734,0.5693115,0.58302987,0.53158605,0.7305021,0.69963586,0.66533995,0.6927767,0.6824879,0.65505123,0.5624523,0.50757897,0.48357183,0.38754338,0.3566771,0.34981793,0.33609957,0.33952916,0.42183927,0.548734,0.6927767,0.8093826,0.82996017,0.6859175,0.71678376,0.8093826,0.8162418,0.70649505,0.5658819,0.65848076,0.6893471,0.805953,0.9774324,0.9842916,1.1592005,1.1214751,1.0357354,0.9774324,0.9362774,1.1797781,1.4061309,1.762808,2.2635276,2.7573884,2.8499873,2.9871707,3.1655092,3.40901,3.782835,4.2218223,4.557922,4.712253,4.530485,3.7553983,3.2032347,2.7642474,2.1023371,1.2826657,0.75450927,0.6207553,0.53844523,0.4698535,0.40126175,0.35324752,0.42869842,0.50757897,0.5521636,0.5796003,0.6310441,0.67219913,0.7407909,0.8128122,0.89169276,1.0117283,1.3581166,1.5638919,1.605047,1.5913286,1.7490896,1.9857311,2.0989075,2.2360911,2.3767042,2.3252604,2.2258022,2.2052248,2.1743584,2.0749004,1.8691251,1.8382589,1.8862731,1.8965619,1.862266,1.9068506,0.31895164,0.12346515,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06859175,0.08916927,0.058302987,0.044584636,0.13032432,0.45613512,0.6927767,0.70649505,0.548734,2.061182,6.0840883,10.827208,14.040731,13.015285,10.072699,6.509357,3.3232703,1.2655178,0.84024894,0.84024894,1.1043272,1.7833855,3.0420442,5.0826488,6.0326443,7.6342616,9.849775,10.971251,7.613684,5.9160385,6.9860697,10.048691,12.6757555,10.772334,13.166186,17.305698,18.338005,15.196502,10.621432,11.314209,11.269625,9.211872,6.258997,5.90575,4.9523244,3.8925817,4.1600895,6.327589,10.100135,9.283894,15.46058,27.837961,37.91066,29.463587,20.162544,17.189093,24.343212,33.904903,26.644464,32.711407,37.82492,38.34279,34.796593,31.891733,28.863409,27.062874,24.219748,19.833303,15.182784,14.119612,15.018164,18.632948,22.587263,21.37662,16.191082,14.812388,14.352823,12.854094,9.277034,6.5539417,4.804852,3.5839188,3.0248961,3.8308492,12.068718,8.4264965,4.5990767,5.0449233,6.9723516,5.98463,4.7019644,3.6353626,3.1209247,3.340418,1.8142518,1.2037852,1.0940384,1.2895249,1.8005334,1.8245405,1.9582944,2.6236343,3.8479972,5.2644167,6.046363,5.8645945,5.885172,6.5024977,7.3701835,7.1129646,6.9037595,6.5230756,5.844017,4.8082814,4.307562,4.190956,3.532475,2.486451,2.3046827,2.2909644,2.527606,2.8499873,3.5187566,5.2026844,7.9737906,7.3564653,7.010077,8.388771,10.7586155,11.513125,12.281353,12.133881,11.101575,10.161868,10.199594,12.250486,15.71094,18.255693,15.837835,12.871242,9.55826,6.475061,4.756838,6.0875177,6.869464,5.720552,5.1992545,5.5079174,4.4721823,3.9474552,5.051782,5.31929,4.1772375,2.9460156,2.4555845,3.3609958,4.7019644,5.312431,3.799983,2.07833,1.9308578,2.085189,2.020027,1.9823016,2.4830213,2.5173173,2.5961976,3.3369887,5.4633327,3.6559403,3.3061223,3.690236,4.530485,5.9983487,5.0826488,2.8945718,2.3732746,3.6044965,3.799983,3.4467354,3.2581081,3.7519686,4.911169,6.1801167,4.835718,4.180667,4.3933015,4.7774153,3.7382503,3.175798,2.935727,3.0626216,3.3884325,3.508468,3.2649672,3.415869,3.2066643,2.4452958,1.4815818,1.2963841,1.371835,2.0406046,3.0900583,3.7382503,4.1292233,5.381023,5.8988905,5.1752477,3.782835,2.8808534,2.2600982,3.2272418,5.4153185,6.8214493,5.1855364,5.2335505,4.8494368,3.4055803,1.7696671,0.939707,0.9877212,2.7539587,4.791134,3.3884325,1.3615463,3.6456516,7.6376915,10.6488695,9.901219,7.3530354,6.677407,6.2075534,5.8165803,6.927767,9.283894,11.273054,9.582268,5.796003,6.392751,4.8425775,5.535354,4.8940215,2.784825,2.5173173,8.597976,9.438225,7.8949103,5.1821065,0.8848336,1.471293,3.4124396,6.262427,7.2432885,1.2380811,2.9803114,10.000677,13.557159,10.4705305,3.0969174,12.922686,10.868362,9.0369625,11.118723,12.3911,11.900668,9.6645775,7.857185,6.927767,5.5833683,3.6696587,3.40901,3.8377085,3.9611735,2.7779658,5.377593,6.7322803,6.111525,4.32128,3.724532,12.596875,14.229359,10.635151,5.120374,2.287535,2.2292318,1.5090185,1.9582944,3.316411,3.2203827,4.307562,4.3658648,4.2938433,5.2815647,8.834618,11.228469,9.2153015,8.97866,12.603734,18.097933,13.896688,13.526293,14.38026,14.534592,12.740917,16.55119,19.929333,21.506943,21.87048,23.544119,21.750444,22.810186,26.26721,30.461596,32.563934,31.781986,31.42188,29.065754,24.816494,21.301168,18.348293,15.083325,12.950122,12.723769,14.479718,12.857523,8.213862,4.122364,2.5584722,3.875434,3.0454736,2.5824795,2.0920484,1.5124481,1.097468,1.2312219,1.3203912,1.3889829,1.6496316,2.503599,3.9783216,3.8274195,3.4192986,2.9700227,1.5398848,0.5041494,0.6276145,0.6962063,0.66191036,1.6633499,1.2243627,1.2346514,1.9582944,3.2821152,4.6848164,5.8680243,5.2506986,4.914599,5.641671,6.910619,6.327589,5.686256,4.122364,1.9754424,0.77851635,2.9151495,4.3349986,4.623084,4.029765,3.4776018,4.7602673,4.2389703,3.6113555,3.1963756,1.937717,2.0234566,3.1963756,2.7951138,1.0151579,0.9294182,0.7339317,0.59674823,0.44927597,0.30523327,0.24350071,0.09602845,0.06859175,0.11317638,0.18176813,0.24350071,0.31895164,0.36353627,0.37382504,0.34981793,0.29151493,0.16804978,0.14747226,0.17147937,0.18862732,0.15090185,0.14061308,0.1097468,0.10288762,0.41840968,1.6016173,2.5927682,3.0317552,2.6819375,2.061182,2.4247184,2.2566686,2.9906003,3.625074,4.214963,5.874883,5.4599032,4.32128,2.8396983,1.3924125,0.36696586,0.12346515,0.26407823,0.26750782,0.13375391,0.36696586,0.072021335,0.010288762,0.020577524,0.29151493,1.3272504,0.32581082,0.38754338,0.3806842,0.16462019,0.5796003,1.8862731,1.5810398,0.7922347,0.58302987,1.937717,4.417309,4.7602673,4.15666,3.782835,4.822,1.9514352,1.5090185,2.5001693,3.7862647,4.105216,3.7142432,3.1483612,2.3561265,1.7799559,2.3664153,4.0846386,5.164959,6.210983,7.0443726,6.715132,6.5779486,7.5245147,6.677407,4.619654,5.4016004,6.193835,6.1286726,6.8728933,8.076678,7.3701835,5.171818,2.702515,0.94999576,0.44584638,1.2517995,1.5570327,0.67219913,0.041155048,0.058302987,0.044584636,0.31552204,0.23664154,0.106317215,0.05144381,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.01371835,0.01371835,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.1371835,0.34638834,0.53501564,0.65505123,0.64819205,0.42869842,0.28122616,0.15090185,0.06859175,0.024007112,0.0,0.0,0.010288762,0.041155048,0.09945804,0.19891608,0.31895164,0.50757897,0.66533995,0.7442205,0.7339317,0.96371406,1.039165,0.9911508,0.939707,1.097468,1.0494537,1.0734608,1.1180456,1.0871792,0.85396725,0.6962063,0.72021335,0.7990939,0.7956643,0.5658819,0.980862,1.4507155,1.8759843,1.8965619,0.8848336,0.66533995,0.64819205,0.64133286,0.6276145,0.7613684,1.2758065,1.1008976,1.0048691,1.1729189,1.2209331,1.1214751,0.86082643,0.70649505,0.70649505,0.65505123,0.4115505,0.31552204,0.2469303,0.20234565,0.274367,0.32238123,0.4629943,0.59674823,0.6756287,0.6859175,0.7956643,0.7339317,0.64133286,0.5761707,0.5041494,0.77165717,0.94999576,1.0700313,1.1214751,1.0220171,0.91227025,0.9842916,1.0940384,1.1694894,1.2037852,1.4507155,1.704505,2.1057668,2.5893385,2.867135,3.0283258,3.059192,3.1620796,3.391862,3.6456516,4.197815,4.389872,4.4859004,4.4756117,4.07435,3.1723683,2.7162333,2.3629858,1.8416885,0.9602845,0.64476246,0.490431,0.4115505,0.35324752,0.30523327,0.42869842,0.5761707,0.6927767,0.71678376,0.59674823,0.65505123,0.77165717,0.90541106,1.0460242,1.2037852,1.3752645,1.5364552,1.6599203,1.7353712,1.786815,2.1400626,2.2841053,2.3629858,2.411,2.3492675,2.1434922,1.8897027,1.7182233,1.6256244,1.4815818,1.2620882,1.2415106,1.4061309,1.6633499,1.845118,0.6756287,0.37039545,0.12689474,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.024007112,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.024007112,0.07545093,0.12003556,0.17833854,0.20920484,0.12003556,0.14747226,0.26407823,0.6824879,1.8108221,4.2595477,9.033533,15.3817,19.726988,19.425184,12.734058,7.1369715,3.99204,2.253239,1.255229,0.7305021,0.9431366,1.4918705,2.5001693,3.8205605,5.007198,5.9812007,8.618553,11.592006,12.380811,7.298162,5.638242,5.785714,7.795452,10.117283,9.589127,14.030442,18.502625,18.269413,13.917266,11.341646,12.88496,12.343085,9.167287,5.9400454,8.357904,7.915488,6.927767,10.000677,15.611482,16.143068,13.862392,13.711491,13.790371,14.30481,17.562918,20.018501,22.26831,24.473536,27.361248,32.207256,45.579216,49.10826,39.947834,25.913963,25.457829,25.368658,25.389236,23.873358,19.514353,11.348505,7.0375133,5.7719955,7.5931067,10.693454,11.417097,8.279024,7.2604365,7.7783046,8.309891,6.3721733,4.3933015,3.426158,2.7299516,4.2766957,12.775213,6.0669403,3.542764,4.2115335,6.012067,5.813151,3.9474552,2.3218307,1.529596,1.5364552,1.6564908,1.3341095,1.1043272,1.196926,1.5330256,1.704505,1.9239986,2.177788,2.4830213,2.8122618,3.117495,2.726522,3.1963756,4.232111,5.4839106,6.5642304,5.144381,4.0880685,3.9165888,4.4584637,4.866585,5.305572,5.6210938,4.6573796,2.7951138,1.937717,3.1277838,4.8494368,5.336438,5.1409516,7.1061053,8.1487,7.459353,9.163857,12.401388,11.341646,8.906639,9.80519,10.662587,9.640571,6.416758,5.31929,7.6959944,12.63803,17.892159,19.829874,16.767254,12.788932,9.794902,7.7680154,4.7808447,5.271276,5.4976287,5.4324665,5.6485305,7.3255987,5.288424,5.0106273,4.57164,3.7622573,4.091498,3.2443898,4.0777793,4.012617,2.884283,2.9322972,2.5996273,1.8691251,2.1880767,3.2786856,3.1415021,2.4418662,2.4967396,3.1723683,4.2869844,5.610805,3.059192,2.2086544,2.0303159,2.5961976,5.055212,4.835718,3.0557625,2.7128036,3.82399,3.433017,4.15323,5.662249,6.0875177,5.192395,4.372724,4.064061,3.2786856,2.7368107,2.6956558,2.9563043,2.9048605,2.3218307,2.1297739,2.6579304,3.6182148,3.7862647,3.1723683,2.5893385,2.1674993,1.371835,1.7250825,2.4590142,2.9151495,3.083199,3.6044965,4.307562,5.0277753,4.976331,4.180667,3.5050385,3.8514268,3.974892,4.8288593,6.4716315,8.090397,7.040943,6.262427,4.547633,2.1812177,0.91569984,1.1214751,1.605047,2.9734523,4.681387,5.0346346,2.7745364,2.760818,4.5167665,6.042933,3.82399,3.3712845,3.309552,3.7725463,4.9077396,6.8797526,9.945804,12.854094,10.882081,5.1066556,2.4144297,3.9200184,4.8425775,4.705394,4.098357,4.6916757,8.241299,8.875772,6.23156,2.177788,0.8128122,3.457024,3.9886103,3.8925817,3.2786856,0.84367853,1.605047,4.619654,5.4976287,3.549623,1.7902447,6.138962,6.4716315,6.615674,7.8949103,9.095266,7.630832,5.3330083,4.73969,5.830299,5.9983487,3.7691166,3.5942078,5.6245236,9.006097,11.893809,7.0752387,5.7239814,5.703404,5.7582774,5.5422134,7.658269,8.525954,6.0497923,1.8931323,1.4815818,1.4335675,1.1180456,1.0185875,1.4232788,2.4384367,2.627064,3.100347,3.8034124,4.619654,5.381023,7.010077,8.80718,9.72288,11.050131,16.424294,17.655516,15.789821,14.531162,14.417986,12.840376,13.903547,15.440002,16.414005,17.271402,19.932762,20.656404,21.548098,23.739605,26.394106,26.726774,30.08777,32.3513,31.034336,25.85223,18.71526,16.55119,13.21763,11.626302,12.682614,15.29939,12.71691,8.244728,4.3590055,2.5550427,3.3266997,3.1415021,2.976882,2.5996273,1.920569,0.9774324,1.4918705,1.7422304,1.8142518,1.961724,2.5996273,2.2498093,2.0817597,1.9411465,1.6633499,1.0666018,0.4664239,0.70306545,0.7305021,0.4972902,0.9431366,1.1008976,1.3443983,1.5330256,1.7216529,2.170929,3.6559403,4.2252517,4.8288593,5.3090014,4.420738,4.245829,7.157549,7.0443726,3.3747141,1.1934965,3.8171308,5.521636,5.130663,3.1792276,1.9171394,2.651071,2.5481834,2.3424082,2.2326615,1.9137098,1.8931323,2.1229146,1.9514352,1.3752645,1.0666018,0.490431,0.28122616,0.28122616,0.34295875,0.34295875,0.106317215,0.05144381,0.06859175,0.11317638,0.19548649,0.26750782,0.3566771,0.40126175,0.36696586,0.2777966,0.16462019,0.12346515,0.13032432,0.14747226,0.14061308,0.1371835,0.1097468,0.11317638,0.34981793,1.1626302,2.218943,2.9254382,3.4604537,3.6285036,2.8396983,3.1483612,5.2335505,6.9723516,7.301592,6.217842,5.254128,4.40359,3.1415021,1.5913286,0.53844523,0.3018037,0.2194936,0.15090185,0.08916927,0.14747226,0.058302987,0.030866288,0.09259886,0.23321195,0.4115505,0.2503599,0.1920569,0.11317638,0.09259886,0.42183927,1.728512,1.978872,1.4747226,1.0734608,2.194936,4.046913,5.950334,7.4456344,8.203573,8.018375,5.6793966,4.0949273,2.959734,2.5481834,3.7142432,4.4756117,6.3893213,5.8062916,3.3232703,3.7794054,4.5442033,4.338428,4.2835546,4.2183924,2.6990852,4.2423997,5.6313825,5.192395,3.8034124,4.8768735,7.936065,7.870903,7.3839016,7.2604365,6.358455,3.7108135,2.4727325,1.7799559,1.1420527,0.432128,1.2655178,0.7407909,0.18519773,0.16462019,0.48357183,0.16804978,0.05144381,0.5521636,1.1489118,0.37039545,0.07545093,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.07545093,0.14747226,0.14747226,0.08916927,0.09602845,0.106317215,0.10288762,0.072021335,0.030866288,0.01371835,0.0034295875,0.0,0.024007112,0.13375391,0.41840968,0.6756287,0.9259886,1.0288762,0.9431366,0.7442205,0.490431,0.2777966,0.12346515,0.048014224,0.061732575,0.05144381,0.020577524,0.017147938,0.058302987,0.12346515,0.2194936,0.4046913,0.69963586,0.91912943,0.6824879,0.7682276,0.8676856,0.881404,0.82996017,0.84367853,0.83338976,0.8676856,0.9431366,0.9294182,0.548734,0.48014224,0.5555932,0.71678376,0.88826317,0.980862,0.85739684,0.6962063,0.7407909,0.91912943,0.823101,0.58302987,0.5761707,0.5521636,0.490431,0.6173257,0.9842916,1.0940384,1.138623,1.1729189,1.1214751,1.3101025,1.08032,0.89512235,0.8779744,0.84024894,0.67219913,0.4355576,0.24350071,0.16119061,0.17833854,0.274367,0.32581082,0.41498008,0.53158605,0.5521636,0.5555932,0.59674823,0.64133286,0.6927767,0.78537554,0.8265306,0.9774324,1.0563129,1.0117283,0.9259886,1.039165,1.2346514,1.2415106,1.1420527,1.3649758,1.646202,1.7936742,2.1229146,2.6476414,3.0626216,3.40901,3.5359046,3.7313912,4.15323,4.8322887,5.0586414,5.0586414,4.938606,4.647091,4.0023284,3.4673128,2.6956558,1.8656956,1.1351935,0.65505123,0.4664239,0.36010668,0.33266997,0.3841138,0.5007198,0.4972902,0.6276145,0.69963586,0.6756287,0.6790583,0.7613684,0.8745448,1.0734608,1.2860953,1.3272504,1.4198492,1.488441,1.488441,1.5055889,1.7490896,2.0234566,2.177788,2.270387,2.3801336,2.5927682,2.287535,1.937717,1.7079345,1.646202,1.6770682,1.5433143,1.4438564,1.471293,1.5947582,1.6496316,0.607037,0.9431366,0.490431,0.07888051,0.0034295875,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.024007112,0.01371835,0.017147938,0.017147938,0.0034295875,0.0,0.006859175,0.024007112,0.030866288,0.048014224,0.08573969,0.12689474,0.15090185,0.12689474,0.22978236,0.4972902,1.6393428,4.5956473,10.55284,16.684942,22.117409,26.1849,26.486704,18.879879,8.992378,4.1155047,2.095478,1.3478279,0.8196714,1.0597426,1.5604624,2.620205,3.9611735,4.722542,6.944915,11.321068,14.315098,13.495427,7.5382333,7.0615206,6.8283086,7.7542973,9.342196,9.695444,14.452282,15.954441,14.373401,12.092726,13.670336,14.448852,11.314209,8.56025,7.8434668,8.203573,8.464222,8.992378,15.388559,23.461807,19.246845,13.399398,15.566897,16.163645,13.670336,14.613472,19.730417,18.37916,16.273392,16.911295,21.572105,33.465916,37.776905,30.7634,19.353163,21.12283,19.548649,17.53548,15.028452,11.790922,7.3873315,4.7088237,3.4604537,4.1326528,6.0840883,7.56224,6.036074,4.8254294,4.3521466,4.197815,3.1106358,2.6990852,4.0674906,4.396731,4.506478,8.855195,3.3987212,2.551613,3.865145,5.0483527,3.957744,2.5653315,1.8142518,1.3649758,1.0734608,0.980862,1.0494537,1.1592005,1.3581166,1.4953002,1.2312219,1.587899,1.9342873,2.3801336,2.942586,3.532475,4.091498,4.8082814,5.1992545,5.1752477,5.0449233,3.8205605,2.9048605,3.018037,4.15323,5.586798,6.9552035,7.7680154,7.1369715,5.435896,4.3007026,4.3761535,6.1321025,7.0752387,7.257007,9.259886,9.523964,9.400499,12.212761,14.870691,7.864044,6.958633,9.712592,10.72089,8.268735,4.32471,4.2938433,7.191845,11.753197,16.273392,18.602083,16.780972,14.181344,11.303921,8.196714,4.4447455,4.5030484,4.9351764,5.2472687,5.425607,5.9434752,5.0140567,5.3741636,5.3878818,4.8082814,4.7808447,3.8274195,4.0091877,3.6593697,2.7573884,2.9185789,3.1655092,2.7985435,2.9631636,3.590778,3.3952916,2.767677,3.2546785,4.0194764,4.513337,4.465323,3.07634,2.2566686,1.5913286,1.605047,3.7519686,3.7691166,2.819121,3.0077481,4.040054,3.2409601,3.0866287,3.6285036,3.707384,3.3438478,3.7279615,3.7108135,2.9974594,2.4590142,2.486451,2.9906003,2.8877127,2.136633,1.7833855,2.1332035,2.750529,2.9734523,2.9906003,2.719663,2.1812177,1.4987297,1.7216529,2.1469216,2.3081124,2.1469216,2.0131679,2.620205,3.0729103,3.2443898,3.4638834,4.4859004,4.7499785,4.197815,4.331569,5.926327,9.057541,9.201583,6.169828,2.9906003,1.1489118,0.59331864,1.6633499,2.9631636,4.338428,5.2987127,5.007198,3.2821152,3.1209247,3.9028704,4.5784993,3.6593697,4.2389703,4.400161,4.355576,4.523626,5.528495,8.052671,8.508806,7.0272245,4.8837323,4.5030484,4.6127954,4.290414,4.465323,4.8837323,4.098357,5.528495,5.439326,3.6079261,1.6907866,3.210094,5.8165803,4.770556,3.0283258,2.294394,3.0283258,2.6887965,2.6613598,2.534465,2.1674993,1.704505,3.6936657,4.5922174,5.453044,7.1095347,10.175586,8.100685,4.7499785,4.1120753,6.560801,8.868914,6.355026,5.2815647,7.5588107,11.633161,12.46312,5.98463,5.2747054,5.312431,4.6745276,5.5559316,7.023795,7.7440085,5.8371577,2.4590142,1.8142518,2.510458,2.218943,1.7662375,1.6221949,1.9137098,1.7662375,1.9480057,2.5996273,3.625074,4.6916757,6.2555676,8.992378,9.421077,8.327039,10.751757,12.922686,13.437123,14.778092,16.383139,14.637479,13.992717,13.728639,14.651197,17.089634,20.896477,19.994495,20.893047,23.046827,24.627867,22.511812,24.624437,26.987423,27.244642,24.648445,20.097382,16.62321,13.491997,12.833516,14.441993,15.7966795,14.345964,10.415657,6.4373355,4.012617,3.9303071,2.9254382,3.0969174,3.3884325,3.216953,2.4555845,2.9631636,2.1812177,1.6187652,1.920569,2.836269,2.0886188,1.7250825,1.3032433,0.8196714,0.70649505,1.2826657,1.4129901,1.903421,2.9082901,3.9303071,3.0797696,1.7799559,1.5604624,2.270387,2.0920484,2.2841053,4.1635194,5.627953,5.5079174,3.5976372,4.417309,7.1232533,6.660259,3.1312134,1.8005334,3.9097297,6.948344,7.6925645,5.3878818,1.7730967,1.6393428,1.4918705,1.6221949,1.9754424,2.153781,1.9137098,2.1880767,2.2223728,1.8176813,1.3169615,0.7407909,0.39440256,0.25721905,0.24007112,0.1920569,0.06859175,0.041155048,0.06859175,0.12346515,0.20234565,0.25378948,0.30866286,0.37382504,0.40126175,0.31209245,0.20920484,0.14747226,0.13032432,0.1371835,0.1371835,0.12346515,0.10288762,0.30523327,0.77165717,1.3443983,1.7456601,2.4384367,3.2512488,3.8479972,3.74168,4.2046742,5.9228973,6.56766,5.504488,3.7931237,3.2375305,2.983741,2.2086544,1.0151579,0.45270553,0.21263443,0.14747226,0.11317638,0.06516216,0.0548734,0.041155048,0.034295876,0.09259886,0.1920569,0.2194936,0.24007112,0.23664154,0.19891608,0.18519773,0.33609957,1.1454822,1.2380811,1.2003556,1.4918705,2.4590142,3.9165888,5.953764,7.332458,7.514226,6.667118,6.2692857,5.223262,3.7759757,2.6407824,3.0043187,3.532475,5.1066556,5.7822843,5.1409516,4.262977,4.1943855,4.386442,5.130663,6.0052075,5.885172,4.1155047,4.2081037,3.7553983,2.7299516,3.474172,6.042933,6.193835,5.171818,4.461893,5.7754254,4.9248877,4.437886,3.1723683,1.6256244,1.9239986,1.5981878,0.6893471,0.09945804,0.12346515,0.47671264,0.18862732,0.08916927,0.30866286,0.5693115,0.18176813,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.010288762,0.0034295875,0.0034295875,0.006859175,0.006859175,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.048014224,0.1920569,0.45956472,0.58645946,0.53158605,0.48014224,0.53501564,0.52472687,0.40126175,0.216064,0.09602845,0.041155048,0.017147938,0.048014224,0.18176813,0.48700142,0.69963586,1.0288762,1.2175035,1.1317638,0.7682276,0.53158605,0.36353627,0.2194936,0.09945804,0.058302987,0.030866288,0.010288762,0.0034295875,0.020577524,0.061732575,0.14061308,0.3018037,0.5624523,0.8265306,0.89169276,0.7990939,0.84367853,0.8025235,0.6893471,0.72364295,0.8025235,0.8711152,0.91569984,0.8265306,0.39097297,0.29837412,0.4355576,0.6001778,0.75450927,1.0288762,0.881404,0.48014224,1.0357354,2.2052248,2.0989075,0.72021335,0.5521636,0.59331864,0.4938606,0.5418748,0.84367853,0.96371406,1.0048691,1.0460242,1.1729189,1.5981878,1.6873571,1.6016173,1.4129901,1.1146159,0.97400284,0.6344737,0.32238123,0.14747226,0.12346515,0.23664154,0.28465575,0.3806842,0.5212973,0.58302987,0.5453044,0.6241849,0.6927767,0.7442205,0.89855194,0.9842916,1.2037852,1.3615463,1.3889829,1.3855534,1.2620882,1.2415106,1.2312219,1.2380811,1.3306799,1.6804979,1.8108221,2.0886188,2.6887965,3.5804894,3.8445675,4.012617,4.184097,4.40359,4.650521,4.6573796,4.945465,5.223262,5.2506986,4.8322887,4.547633,3.542764,2.3286898,1.2826657,0.67219913,0.48357183,0.39783216,0.42183927,0.548734,0.7510797,0.764798,0.7099246,0.6859175,0.7407909,0.85739684,0.8128122,0.8471081,0.9328478,1.0460242,1.1832076,1.2860953,1.2415106,1.2072148,1.2758065,1.4747226,1.5913286,1.7765263,1.937717,2.0337453,2.0886188,1.9994495,1.8931323,1.8073926,1.7250825,1.587899,1.3684053,1.2963841,1.3855534,1.5673214,1.6942163,0.5693115,1.2826657,0.7682276,0.22635277,0.106317215,0.08573969,0.017147938,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.01371835,0.020577524,0.01371835,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.01371835,0.041155048,0.08916927,0.10288762,0.07888051,0.034295876,0.006859175,0.01371835,0.037725464,0.048014224,0.08916927,0.14061308,0.19891608,0.26750782,0.38754338,0.65162164,2.0577524,5.456474,11.567999,17.71039,24.93996,31.432169,33.215553,24.168303,11.31078,4.8940215,2.2258022,1.3443983,1.0151579,1.3272504,2.0508933,3.3369887,4.650521,4.7671266,7.891481,13.522863,15.824117,13.4645605,9.599416,9.904649,8.621983,8.735159,10.213311,9.983529,13.193623,12.833516,11.228469,10.717461,13.642899,12.836946,10.460241,10.062409,11.478829,10.834066,12.22648,16.667795,21.575535,23.386356,17.549198,14.229359,19.047928,20.52951,16.139639,12.295071,15.937293,14.661487,13.457702,13.687484,13.090735,16.94902,20.676983,18.193962,12.521424,15.762384,16.146498,12.932974,9.139851,6.310441,4.5201964,3.7622573,3.0900583,3.3987212,4.5099077,5.1683884,4.6402316,3.6387923,2.668219,1.8931323,1.1214751,1.5261664,3.782835,4.962613,4.554492,4.4756117,2.469303,2.2909644,3.0420442,3.649081,2.884283,2.2086544,2.0440342,1.7250825,1.2963841,1.5158776,1.5055889,1.5227368,1.7490896,2.0577524,2.0165975,2.1503513,2.2052248,2.668219,3.7005248,5.147811,6.447624,6.800872,6.3447366,5.31929,4.07435,3.2135234,2.9494452,3.4398763,4.6127954,6.1629686,7.1026754,7.915488,7.9463544,7.2604365,6.632822,5.809721,6.831738,8.327039,9.671436,10.97468,10.357354,10.700313,12.80608,13.639469,6.3447366,7.0615206,9.72288,10.0041065,7.1781263,4.098357,4.6779575,6.800872,9.259886,11.379372,13.008426,13.090735,13.008426,11.547421,8.738589,5.885172,5.65539,5.693115,6.2487082,6.7048435,5.5730796,4.773986,5.2575574,6.0086374,6.3721733,6.0635104,4.9180284,4.0091877,3.3369887,3.0111778,3.2478194,3.9268777,3.6010668,3.350707,3.508468,3.642222,3.457024,4.465323,5.23698,4.9660425,3.4810312,2.7402403,2.393852,2.0028791,1.8176813,2.784825,3.0489032,2.4384367,2.819121,4.07435,4.1189346,2.867135,1.9891608,1.7593783,2.2566686,3.3438478,3.1689389,2.719663,2.3595562,2.287535,2.5070283,2.2806756,1.762808,1.4747226,1.5193073,1.6084765,1.978872,2.6476414,2.7642474,2.2120838,1.5947582,1.5810398,1.5844694,1.5364552,1.3992717,1.1729189,1.4404267,1.6187652,1.9068506,2.5447538,3.8102717,4.5270553,4.400161,4.383013,5.130663,7.006647,6.711703,3.7313912,1.3615463,0.8196714,1.2620882,2.253239,3.4913201,4.3658648,4.4721823,3.6044965,2.9734523,3.1895163,3.666229,4.1360826,4.6848164,5.7994323,5.3673043,4.5922174,4.125794,4.0777793,4.8185706,4.6916757,5.693115,7.7268605,8.628842,5.164959,3.3815732,3.3884325,4.016047,2.8156912,3.2512488,2.8328393,2.3732746,2.8465576,5.3878818,6.584808,5.0586414,3.7451096,3.7691166,4.437886,3.5873485,2.1674993,1.5741806,2.0920484,2.8877127,4.9008803,4.8837323,4.715683,6.183546,10.998687,10.714031,6.2830043,4.3007026,6.310441,8.790032,6.6465406,5.411889,6.7048435,9.177576,8.525954,4.8288593,5.2026844,5.079219,4.2595477,6.893471,10.871792,11.681175,8.539673,3.799983,2.952875,4.297273,3.4947495,2.4624438,1.9582944,1.5844694,1.4129901,1.3889829,1.8999915,3.07634,4.8014226,5.6073756,6.9380555,6.783724,5.7479887,7.0032177,8.515666,10.957532,14.359683,17.027903,15.529172,14.2533655,14.284232,15.642348,18.149376,21.462358,20.299728,21.404055,23.743034,25.080574,21.993944,21.980227,22.957659,23.341772,22.86163,22.559826,17.682953,14.678635,14.819247,16.931873,17.370861,16.187653,12.734058,9.074688,6.40304,5.0346346,3.3472774,3.0317552,3.4021509,3.7759757,3.4776018,3.4947495,2.294394,1.4335675,1.605047,2.633923,2.4761622,1.8416885,1.0220171,0.45613512,0.72021335,2.0131679,2.301253,2.7985435,3.6044965,3.7005248,3.74168,4.40702,4.0606318,2.702515,1.9823016,1.9137098,3.6285036,4.7602673,4.3658648,2.9082901,4.636802,6.8797526,6.5642304,3.8617156,2.1846473,3.9371665,6.420188,7.466212,6.0737996,2.3972816,1.488441,1.1249046,1.4335675,2.2841053,3.2718265,1.9445761,2.7230926,3.8720043,4.105216,2.5996273,1.1729189,0.5521636,0.29494452,0.15776102,0.07545093,0.044584636,0.048014224,0.082310095,0.1371835,0.2194936,0.274367,0.31209245,0.37382504,0.42183927,0.34295875,0.23321195,0.18176813,0.15433143,0.14061308,0.1371835,0.12346515,0.15433143,0.48357183,1.039165,1.4369972,1.3169615,1.6667795,2.2326615,2.952875,3.9783216,4.386442,5.4667625,5.5250654,4.2081037,2.49331,2.3664153,2.4041407,1.762808,0.65848076,0.35324752,0.19891608,0.13032432,0.12003556,0.11317638,0.037725464,0.0274367,0.024007112,0.082310095,0.20234565,0.32238123,0.34638834,0.33609957,0.29494452,0.24350071,0.2194936,0.5144381,0.52815646,0.6756287,1.1934965,2.1434922,3.6113555,5.267846,6.0806584,5.7651367,4.746549,6.0395036,6.200694,5.2266912,3.6525106,2.5584722,2.760818,3.707384,4.962613,5.669108,4.5510626,4.897451,6.341307,7.939495,8.958082,8.879202,6.029215,5.4187484,4.465323,3.0626216,3.5770597,4.249259,4.40702,4.0023284,3.9371665,6.0497923,7.0375133,6.680836,4.633373,2.318401,2.9494452,1.4472859,0.4389872,0.010288762,0.048014224,0.23664154,0.1371835,0.08916927,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.31552204,0.7099246,0.94656616,0.939707,0.8196714,0.83338976,0.77165717,0.6036074,0.3806842,0.23664154,0.16119061,0.106317215,0.11317638,0.23321195,0.53844523,0.5727411,0.77508676,0.9602845,0.97057325,0.66533995,0.51100856,0.42183927,0.31209245,0.17490897,0.09602845,0.024007112,0.0034295875,0.0,0.0034295875,0.017147938,0.07545093,0.26064864,0.53158605,0.82996017,1.0631721,0.89855194,0.9294182,0.9774324,1.0220171,1.1934965,1.0734608,1.0220171,1.0220171,0.9362774,0.4938606,0.40126175,0.5041494,0.5761707,0.6241849,0.8711152,0.8025235,0.4115505,0.939707,2.0577524,1.8691251,0.6310441,0.70649505,1.0494537,1.0768905,0.64133286,0.864256,0.97057325,1.0117283,1.0563129,1.2209331,1.5364552,1.7456601,1.7833855,1.6221949,1.2415106,1.0048691,0.6790583,0.37382504,0.16804978,0.106317215,0.1920569,0.29494452,0.432128,0.58988905,0.70649505,0.69963586,0.77851635,0.8711152,0.9602845,1.0837497,1.1900668,1.3992717,1.5810398,1.6599203,1.611906,1.4781522,1.4575747,1.4541451,1.4507155,1.4953002,1.8897027,2.2292318,2.668219,3.3026927,4.166949,4.396731,4.4927597,4.448175,4.383013,4.540774,4.866585,5.3981705,5.751418,5.7822843,5.579939,5.3570156,4.3487167,3.1380725,2.0714707,1.2689474,0.8711152,0.7339317,0.7613684,0.864256,0.9568549,0.96714365,0.86082643,0.8128122,0.8848336,1.0460242,0.89169276,0.83338976,0.7922347,0.78194594,0.90198153,0.94656616,0.88826317,0.89855194,1.0185875,1.1317638,1.1900668,1.3958421,1.5913286,1.6770682,1.6187652,1.6016173,1.5913286,1.5604624,1.4644338,1.2312219,1.0666018,1.1523414,1.2758065,1.3512574,1.4438564,0.58988905,1.1249046,0.7510797,0.36696586,0.274367,0.17490897,0.041155048,0.0034295875,0.006859175,0.010288762,0.0034295875,0.01371835,0.024007112,0.024007112,0.017147938,0.006859175,0.0,0.0034295875,0.0034295875,0.006859175,0.017147938,0.017147938,0.006859175,0.0548734,0.14747226,0.18519773,0.15776102,0.06859175,0.006859175,0.01371835,0.0548734,0.11317638,0.14404267,0.2469303,0.40126175,0.47671264,0.5521636,0.5693115,1.488441,3.6010668,6.5470824,12.435684,23.989964,33.122955,34.00779,23.091412,10.957532,4.846007,2.170929,1.2483698,1.3066728,1.9445761,3.3781435,4.962613,5.8474464,4.962613,8.344186,14.04759,15.443433,12.63803,12.46312,12.408247,9.633711,9.352485,11.372512,10.089847,10.864933,10.844356,10.350495,10.161868,11.499407,10.05898,11.80121,14.232788,16.108772,17.439453,21.091963,28.400414,27.09374,17.851004,14.321958,19.102802,24.161444,22.865059,15.522313,9.403929,13.293081,17.717249,19.569225,17.686382,12.840376,7.3839016,8.735159,8.549961,6.245279,8.992378,14.71636,12.950122,9.15014,5.98463,3.340418,3.0523329,2.4418662,2.6750782,3.4398763,2.9391565,2.5893385,2.1469216,1.7765263,1.3924125,0.65848076,1.0151579,2.3835633,4.091498,5.3501563,5.271276,3.0351849,2.3732746,2.7402403,3.3815732,3.3198407,2.8911421,2.3424082,1.8108221,1.7010754,2.6647894,2.6750782,2.510458,2.6887965,3.2066643,3.5599117,3.2409601,2.8911421,3.234101,4.4996185,6.4304767,7.3290286,6.999788,6.2418494,5.2644167,3.7005248,3.0866287,3.525616,4.3521466,5.171818,5.8474464,5.9331865,6.64997,7.281014,7.613684,7.953213,7.4113383,7.5107965,8.992378,11.019264,11.156448,9.767465,10.079557,10.281903,9.352485,7.0958166,7.9017696,8.333898,7.7131424,6.509357,6.324159,5.5730796,5.164959,4.852866,4.9214582,6.1766872,7.5039372,9.544542,10.31277,9.410788,8.052671,8.110974,7.4799304,8.035523,9.163857,7.7577267,5.610805,4.99005,5.844017,7.1095347,6.691125,5.3158607,3.9303071,3.1243541,3.0797696,3.5633414,4.307562,3.6765177,3.3369887,3.7142432,4.012617,3.882293,4.9214582,5.535354,4.8905916,2.935727,2.0920484,2.1503513,2.3561265,2.452155,2.6853669,3.0557625,2.452155,2.5790498,3.7794054,5.0483527,3.6559403,2.318401,2.0886188,2.7813954,3.000889,2.5481834,2.287535,2.0063086,1.6907866,1.5364552,1.4267083,1.3032433,1.1180456,0.90198153,0.7579388,1.3924125,2.2635276,2.585909,2.2086544,1.5981878,1.5810398,1.4335675,1.2826657,1.2449403,1.4267083,1.3203912,1.2517995,1.3272504,1.5227368,1.6839274,3.117495,4.15323,4.5030484,4.040054,2.8054025,1.1214751,0.48700142,0.52815646,1.0837497,2.1812177,2.3972816,2.8980014,2.9665933,2.5653315,2.3149714,2.901431,3.0660512,3.3644254,4.180667,5.7308407,6.914048,5.223262,3.7725463,3.5599117,3.474172,2.311542,3.998899,8.169277,12.05843,10.532263,4.5853586,2.633923,2.527606,2.6887965,2.1091962,2.3252604,2.3389788,2.8739944,4.064061,5.4804807,5.394741,4.6779575,5.038064,5.874883,4.280125,3.5530527,2.3081124,1.3238207,1.6084765,4.386442,8.371623,7.0923867,4.972902,5.4941993,11.177026,12.929544,7.932636,4.437886,4.791134,5.442755,4.2938433,3.7965534,4.0503426,4.557922,4.2183924,4.482471,5.7719955,5.641671,5.120374,8.7283,14.942713,15.4742985,10.429376,3.9543142,4.2526884,5.7411294,4.0777793,2.2978237,1.5810398,1.2483698,1.2655178,1.488441,1.99602,2.9082901,4.389872,3.9440255,3.3850029,3.3266997,4.266407,6.557371,7.805741,10.31277,13.169616,15.110763,14.507155,14.284232,15.80011,17.099922,17.96418,19.884748,21.067955,22.817045,25.077143,26.407824,23.986534,22.95423,22.422644,21.915064,21.969936,24.123718,19.483486,16.606062,17.04505,19.507494,19.850452,17.833855,14.555169,11.06042,7.939495,5.3090014,4.1463714,3.0660512,2.867135,3.4124396,3.6147852,2.9665933,2.8877127,2.5996273,2.1057668,2.177788,2.6133456,1.920569,0.97400284,0.50757897,1.1111864,2.3595562,2.9974594,3.3987212,3.1072063,0.8162418,2.5207467,6.7871537,6.7871537,2.627064,1.3443983,1.99602,2.4590142,2.74367,2.760818,2.3081124,4.420738,6.6293926,6.989499,5.144381,2.318401,4.32471,4.804852,4.887162,4.65395,3.1723683,1.9274281,1.2483698,1.7696671,3.199805,4.341858,1.8999915,3.3678548,5.7822843,6.728851,4.3624353,2.1572106,0.9774324,0.42183927,0.18862732,0.09259886,0.06859175,0.07545093,0.10288762,0.15090185,0.25378948,0.32238123,0.37725464,0.44927597,0.490431,0.3806842,0.24350071,0.20577525,0.18176813,0.14747226,0.1371835,0.14404267,0.25378948,0.5453044,0.94656616,1.214074,1.0357354,0.939707,1.0323058,1.6667795,3.4433057,3.6970954,4.4756117,4.996909,4.6848164,3.1826572,3.2718265,3.0523329,2.0817597,0.7682276,0.36696586,0.31209245,0.16804978,0.13375391,0.17833854,0.037725464,0.030866288,0.0274367,0.09602845,0.24007112,0.37382504,0.53501564,0.4355576,0.31552204,0.25378948,0.13375391,0.12346515,0.3018037,0.32924038,0.39440256,1.2346514,2.760818,3.9097297,4.4104495,4.180667,3.3301294,5.4736214,6.6705475,6.3721733,4.8151407,3.0043187,3.0077481,3.841138,4.7431192,5.1992545,4.9214582,6.6739774,9.438225,11.05356,10.576848,8.255017,7.73029,7.5862474,6.4407654,4.9077396,5.6005163,4.547633,4.314421,4.6436615,5.453044,6.8283086,8.423067,7.9017696,5.7136927,3.275256,2.9460156,1.2517995,0.4355576,0.106317215,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.01371835,0.058302987,0.39440256,0.8196714,1.1008976,1.1489118,1.0048691,0.96371406,0.8265306,0.6756287,0.548734,0.42869842,0.34638834,0.26750782,0.23321195,0.29494452,0.5418748,0.4389872,0.41840968,0.5212973,0.66191036,0.6276145,0.5178677,0.45613512,0.37382504,0.26750782,0.20234565,0.06859175,0.01371835,0.0,0.0,0.0034295875,0.048014224,0.28122616,0.6207553,0.939707,1.0940384,1.0151579,1.0768905,1.3272504,1.7147937,2.0714707,1.5776103,1.2895249,1.2277923,1.2037852,0.8025235,0.72364295,0.7099246,0.66191036,0.61046654,0.6859175,0.6276145,0.37725464,0.2709374,0.33609957,0.28808534,0.4046913,0.922559,1.5536032,1.7765263,0.8162418,0.89169276,1.0734608,1.2072148,1.2277923,1.1729189,1.1489118,1.2072148,1.2963841,1.3238207,1.1523414,0.85396725,0.6379033,0.4355576,0.23664154,0.12689474,0.15776102,0.3018037,0.48357183,0.65505123,0.7990939,0.88826317,0.980862,1.1420527,1.3238207,1.3443983,1.3512574,1.4781522,1.6187652,1.6873571,1.611906,1.8073926,1.9754424,1.8999915,1.6942163,1.8142518,2.2292318,2.8396983,3.5153272,4.1360826,4.5853586,4.8322887,4.8185706,4.6402316,4.5853586,5.1238036,5.844017,6.2692857,6.2658563,5.977771,5.8165803,5.6142344,4.863155,3.99204,3.1689389,2.311542,1.5913286,1.2415106,1.1317638,1.1077567,0.9877212,0.99801,1.0494537,1.0631721,1.0666018,1.1797781,1.0288762,0.88826317,0.7682276,0.66876954,0.6241849,0.548734,0.548734,0.6241849,0.7442205,0.83681935,0.922559,1.0906088,1.2415106,1.3272504,1.3341095,1.214074,1.1008976,1.0151579,0.939707,0.8025235,0.83338976,1.0597426,1.1283343,0.9945804,0.9568549,0.26064864,0.490431,0.39440256,0.33266997,0.3566771,0.19891608,0.06516216,0.020577524,0.010288762,0.0034295875,0.01371835,0.0274367,0.030866288,0.030866288,0.030866288,0.030866288,0.006859175,0.010288762,0.01371835,0.017147938,0.030866288,0.017147938,0.006859175,0.006859175,0.0274367,0.07545093,0.041155048,0.01371835,0.006859175,0.030866288,0.09259886,0.18862732,0.15090185,0.29494452,0.548734,0.42869842,0.5624523,0.44927597,0.5418748,1.0288762,1.845118,8.841476,20.899906,25.317215,19.696121,11.931535,6.012067,2.983741,1.6359133,1.2826657,1.7696671,3.1483612,5.6176643,6.9071894,6.2555676,4.4241676,8.405919,12.768354,14.013294,12.572867,12.816368,11.317638,8.275595,7.9943686,10.271614,10.405369,9.942374,10.209882,10.185875,10.155008,11.718901,13.306799,17.106783,19.500635,20.749004,25.008553,33.212124,34.50165,27.738503,18.276272,17.960749,27.17605,32.90346,29.583622,19.315437,11.856084,24.476965,31.5865,27.961426,17.772121,14.586036,6.8728933,6.948344,7.034084,4.7534084,3.1449318,9.599416,10.868362,9.4862385,6.9792104,3.8308492,3.6593697,2.095478,1.3821237,2.0474637,2.9151495,1.704505,1.1283343,1.1523414,1.2929544,0.61046654,1.4164196,2.452155,4.756838,7.9189177,10.055551,6.210983,5.1580997,5.4804807,5.895461,5.2472687,4.273266,2.5173173,1.4541451,1.7010754,3.0043187,3.981751,4.6093655,4.616225,4.033195,3.2032347,2.7882545,2.7951138,3.5050385,4.695105,5.662249,5.5147767,4.945465,4.4721823,3.981751,2.760818,2.860276,3.642222,4.4859004,4.7842746,3.9680326,5.9571934,7.846896,8.529384,8.344186,9.0644,9.379922,8.838047,8.611694,8.776315,8.299602,7.740579,7.4696417,6.691125,5.4599032,4.715683,5.4736214,4.835718,4.5510626,6.3481665,11.962401,7.630832,3.4981792,1.6976458,2.3424082,3.5393343,3.4776018,5.0655007,6.6533995,7.5519514,8.042382,9.554831,8.056101,8.196714,10.295622,10.343636,7.963502,6.0978065,5.470192,5.2644167,3.1277838,1.9068506,2.6167753,3.4776018,3.7348208,3.6627994,2.9803114,2.9460156,3.9474552,5.0277753,3.8925817,2.7916842,2.5001693,2.218943,1.8382589,1.9239986,2.1915064,1.6359133,1.196926,1.6839274,3.782835,3.3815732,3.683377,3.5873485,3.0454736,3.083199,3.1552205,2.952875,3.234101,3.7313912,3.1586502,2.6579304,2.020027,1.728512,1.7319417,1.4644338,1.8931323,1.587899,1.097468,0.7442205,0.61046654,1.2586586,2.287535,2.7333813,2.3561265,1.6496316,2.0028791,1.8519772,1.5844694,1.3924125,1.2826657,0.9877212,1.0357354,1.039165,1.039165,1.4644338,1.4541451,1.138623,1.0768905,1.2175035,0.90198153,0.4972902,0.7442205,1.0563129,1.2175035,1.3889829,1.4369972,2.1812177,2.4624438,2.486451,3.8308492,5.099797,4.482471,4.262977,5.7308407,9.184435,9.431366,6.560801,3.8514268,3.059192,4.4241676,3.4467354,5.15467,9.373062,12.144169,5.7239814,2.6476414,3.5804894,4.7808447,4.389872,2.4247184,1.7902447,2.8054025,3.4398763,3.0626216,2.4418662,3.4673128,3.9886103,4.8185706,5.501058,4.3178506,3.7553983,3.3781435,2.2738166,1.529596,4.2252517,12.003556,11.05356,8.203573,8.368194,14.555169,12.236768,7.346176,4.4413157,4.232111,3.5873485,3.3678548,3.100347,4.547633,6.293293,3.7553983,3.9611735,7.7131424,8.1212635,5.284994,6.2864337,10.545981,9.626852,5.5113473,2.0097382,4.729401,5.9126086,3.57363,1.4129901,0.7613684,0.5658819,1.039165,1.8931323,2.2566686,2.2155135,2.7779658,2.3629858,2.651071,3.3712845,4.496189,6.2418494,8.718011,10.940384,11.777204,11.578287,12.175035,15.851553,16.156786,15.0456,14.723219,17.638369,20.762722,24.027689,25.996273,25.989414,24.048267,22.546108,22.079683,22.477516,23.28347,23.756752,22.426073,20.172834,20.172834,21.976797,21.500084,20.011642,16.599203,11.262765,5.5902276,2.7470996,3.858286,3.6696587,3.2958336,3.3815732,4.0880685,3.2958336,5.888602,7.164408,5.5113473,2.411,1.8965619,1.862266,1.4027013,0.82996017,1.646202,2.6613598,3.2272418,5.099797,6.7459984,3.340418,1.7182233,2.1915064,3.2409601,3.4776018,1.6496316,1.2586586,1.762808,3.1449318,4.3349986,3.234101,5.003768,5.4667625,4.7808447,3.5050385,2.5619018,5.164959,6.0532217,5.641671,4.540774,3.5393343,2.6236343,1.4061309,2.6407824,4.9660425,2.9151495,1.7799559,4.057202,5.456474,4.911169,4.5922174,4.763697,2.5001693,0.7339317,0.34638834,0.15090185,0.12689474,0.12346515,0.15090185,0.22978236,0.34981793,0.34981793,0.432128,0.6241849,0.7613684,0.5041494,0.30866286,0.23321195,0.18176813,0.1371835,0.1371835,0.17490897,0.31209245,0.50757897,0.72707254,0.94656616,0.9842916,0.8093826,0.7099246,1.2072148,3.0523329,3.210094,3.782835,4.15323,4.0846386,3.707384,4.245829,3.3541365,1.9754424,0.84367853,0.48700142,0.31895164,0.16462019,0.09259886,0.072021335,0.0,0.072021335,0.072021335,0.12689474,0.20577525,0.106317215,0.66876954,0.607037,0.4355576,0.36696586,0.30523327,0.15776102,0.33266997,0.33266997,0.15776102,0.30523327,1.0117283,1.4369972,1.4918705,1.1797781,0.59674823,3.2066643,4.602506,5.07236,5.0312047,5.020916,4.105216,4.40702,5.2609873,5.8508763,5.2026844,7.716572,11.101575,11.962401,9.318189,4.5922174,4.897451,5.2026844,5.826869,6.8214493,7.98065,7.2124224,6.2144127,4.8597255,4.3041325,6.989499,7.6342616,7.4044795,6.018926,4.1772375,3.5564823,3.0043187,1.670209,0.53501564,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.020577524,0.044584636,0.36353627,0.864256,1.2003556,1.2483698,1.1146159,1.3101025,1.1489118,1.0082988,0.9431366,0.6859175,0.5041494,0.4389872,0.37725464,0.29494452,0.26064864,0.4424168,0.5418748,0.6824879,0.8471081,0.8848336,0.6276145,0.4629943,0.39097297,0.37382504,0.33609957,0.15090185,0.041155048,0.0,0.0034295875,0.01371835,0.09945804,0.31552204,0.5590228,0.7990939,1.0666018,1.214074,1.2243627,1.4815818,2.0234566,2.5481834,2.0714707,1.6770682,1.4815818,1.3889829,1.0837497,0.88826317,0.8196714,0.764798,0.69963586,0.6859175,0.6379033,0.5418748,0.47671264,0.4698535,0.5178677,0.66533995,0.84024894,1.0940384,1.2346514,0.7922347,0.6241849,0.9294182,1.2758065,1.3546871,0.9774324,0.91569984,0.91912943,0.90198153,0.8745448,0.94656616,1.0082988,0.91227025,0.66876954,0.37382504,0.21263443,0.16462019,0.25378948,0.42869842,0.6173257,0.70306545,0.90884066,1.1180456,1.3684053,1.5638919,1.4815818,1.3101025,1.4953002,1.6667795,1.7936742,2.1983654,2.5893385,2.5207467,2.16064,1.786815,1.8005334,2.277246,2.760818,3.2821152,3.875434,4.6093655,4.633373,4.6573796,5.0586414,5.7582774,6.210983,6.0532217,5.9126086,5.826869,5.778855,5.7068334,5.8165803,5.48734,4.887162,4.1326528,3.2649672,2.3972816,1.5501735,1.0254467,0.82996017,0.67219913,0.91569984,1.1420527,1.2380811,1.2175035,1.2037852,1.1694894,0.9945804,0.7922347,0.6241849,0.48700142,0.41498008,0.37039545,0.4115505,0.53158605,0.64133286,0.64133286,0.65848076,0.6824879,0.7099246,0.7476501,0.7339317,0.7133542,0.70649505,0.70649505,0.65505123,0.70649505,0.7613684,0.7990939,0.8196714,0.8711152,0.3566771,0.6379033,0.4629943,0.31209245,0.28808534,0.15090185,0.044584636,0.024007112,0.0274367,0.024007112,0.01371835,0.0274367,0.024007112,0.01371835,0.01371835,0.041155048,0.017147938,0.034295876,0.06516216,0.07545093,0.017147938,0.006859175,0.006859175,0.017147938,0.034295876,0.06516216,0.037725464,0.034295876,0.05144381,0.07888051,0.09259886,0.12003556,0.15776102,0.23664154,0.36010668,0.5007198,0.66533995,0.7922347,0.8128122,0.8779744,1.3958421,6.1149545,11.026124,12.061859,9.016385,5.5490727,3.2135234,2.0165975,1.587899,1.6736387,2.1743584,3.6113555,5.267846,6.433906,6.958633,7.257007,9.839486,13.049581,15.172495,15.577187,14.695783,9.6988735,7.0889573,7.116394,8.30646,7.466212,12.079007,11.609154,9.091836,7.442205,9.472521,13.509145,16.328266,17.662374,18.725548,22.213438,27.008001,32.10437,29.8477,20.95135,14.493437,19.569225,26.195189,25.835083,20.241425,21.472647,40.55144,39.00127,26.253492,12.459691,8.484799,3.6696587,5.312431,9.2153015,10.9541025,5.8645945,4.413879,4.1360826,3.9303071,3.6525106,4.0846386,5.6828265,3.4844608,1.546744,1.3649758,1.8999915,1.3375391,0.9945804,1.2209331,1.5638919,0.7922347,0.69963586,0.66191036,1.5227368,3.0626216,3.9783216,4.0194764,5.658819,6.416758,5.6005163,4.307562,4.0846386,3.6593697,3.8720043,4.434457,3.9337368,4.314421,5.1100855,5.2438393,4.822,5.1340923,4.465323,4.40702,4.3178506,4.149801,4.4413157,4.4413157,4.245829,4.0434837,3.7691166,3.117495,4.2183924,4.712253,5.0620713,5.0757895,3.9063,5.885172,8.899779,9.729739,8.1384115,6.866034,7.016936,7.1061053,7.1781263,7.0923867,6.5196457,6.992929,7.414768,6.2418494,4.8185706,7.377043,9.9698105,6.81802,4.705394,7.0478024,13.903547,11.015835,4.835718,1.8485477,3.4021509,5.7136927,3.923448,3.724532,4.588788,5.6793966,5.857735,6.5299344,5.5113473,5.909179,7.9257765,8.844906,9.225591,8.597976,7.1952744,5.40503,3.7862647,2.7128036,2.8088322,3.4055803,3.9371665,3.9303071,2.4658735,2.2360911,3.7519686,5.672538,4.8322887,3.0969174,2.6373527,2.1640697,1.5398848,1.8005334,2.136633,1.7765263,1.2929544,1.5638919,3.758828,3.199805,2.7299516,2.7470996,2.9082901,2.153781,2.277246,2.8054025,3.3850029,3.625074,3.1106358,2.5893385,2.2841053,2.0337453,1.9582944,2.4418662,2.2326615,1.7490896,1.3032433,1.0460242,0.939707,0.8265306,1.08032,1.9651536,2.6853669,1.3924125,1.920569,2.0577524,1.7456601,1.2380811,1.097468,1.0220171,1.3821237,1.5707511,1.3821237,1.039165,1.1420527,1.2963841,1.2175035,0.881404,0.53501564,0.30866286,0.29837412,0.36353627,0.41840968,0.42526886,0.5693115,1.1111864,2.0131679,3.2443898,4.7808447,5.212973,4.1292233,3.117495,2.9288676,3.474172,6.56766,6.001778,3.7622573,2.177788,3.9371665,3.8377085,3.6182148,3.8137012,3.998899,2.7916842,1.9137098,3.7759757,4.8734436,3.7622573,1.0837497,1.1111864,2.5173173,2.9940298,2.218943,1.879414,3.0420442,3.2478194,2.6133456,1.6804979,1.4267083,2.5824795,3.525616,2.959734,2.0028791,4.201245,6.773435,5.6656785,6.989499,12.010415,17.144508,12.960411,8.217292,5.3844523,4.5853586,3.5873485,3.7485392,4.2869844,4.835718,4.9180284,3.9611735,4.773986,8.4264965,8.64942,5.346727,4.588788,10.755186,14.760944,10.995257,2.9220085,3.1072063,3.4124396,2.3767042,1.3615463,0.85396725,0.4424168,0.8128122,2.3321195,3.0489032,2.6167753,2.287535,2.8225505,2.901431,3.0146074,3.350707,3.7862647,4.3109913,7.174697,8.64599,8.64256,10.734609,13.718349,16.396858,19.11309,21.050808,20.227707,20.598103,20.834743,22.083115,24.202599,25.76992,23.232025,23.02625,24.466677,26.26721,26.527859,22.94394,21.887627,23.544119,25.44068,22.463799,19.977346,19.517782,16.39,10.343636,5.5662203,6.1492505,6.108095,5.3673043,4.214963,3.2821152,3.457024,3.1723683,4.8254294,7.15069,5.2438393,2.7368107,2.2120838,2.5927682,3.2581081,4.016047,5.195825,4.125794,2.9665933,2.3492675,1.3752645,2.633923,2.9322972,3.5873485,4.8425775,5.8817425,2.867135,2.335549,2.411,2.0268862,0.9294182,2.318401,2.7916842,2.4418662,2.0474637,3.100347,3.3850029,4.170378,6.9071894,9.760606,7.6171136,3.1072063,1.3786942,2.3046827,4.0709205,3.1826572,2.8568463,4.513337,6.262427,7.301592,7.9017696,5.1512403,2.5447538,1.0220171,0.6310441,0.5418748,0.30523327,0.36696586,0.3841138,0.30866286,0.40126175,0.3806842,0.42183927,0.5041494,0.5727411,0.53844523,0.31552204,0.22292319,0.22292319,0.2503599,0.22292319,0.2503599,0.28808534,0.36353627,0.47328308,0.6036074,0.77851635,0.6001778,0.64133286,1.2483698,2.5756202,3.2718265,3.2443898,2.9288676,2.7642474,3.1963756,2.7368107,2.3149714,1.704505,1.0288762,0.7442205,0.77851635,0.50757897,0.31895164,0.33952916,0.45270553,0.64133286,0.48014224,0.37039545,0.34981793,0.106317215,0.37382504,0.48357183,0.48700142,0.4698535,0.53844523,0.4698535,0.50757897,0.47328308,0.40126175,0.548734,0.39783216,0.980862,1.039165,0.6207553,1.0597426,1.9823016,1.978872,2.6407824,4.0194764,4.6402316,4.722542,4.8425775,4.5784993,4.420738,5.7754254,7.8023114,10.100135,9.9698105,7.4765005,5.446185,6.0635104,6.1321025,6.355026,6.5333643,5.562791,6.619104,6.8111606,6.262427,5.4324665,5.120374,10.943813,11.602294,9.80519,7.4010496,5.3741636,3.5050385,4.0366244,3.0523329,0.51100856,0.24350071,0.058302987,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.017147938,0.06859175,0.31895164,0.7510797,1.0871792,1.2003556,1.1146159,1.3101025,1.0528834,0.84367853,0.86082643,0.96714365,0.922559,0.71678376,0.59674823,0.53158605,0.22292319,0.33609957,0.4081209,0.5658819,0.8471081,1.1660597,0.881404,0.69963586,0.5590228,0.41498008,0.26407823,0.12003556,0.041155048,0.017147938,0.034295876,0.07545093,0.14061308,0.30866286,0.66876954,1.0185875,0.8471081,1.3752645,1.3855534,1.4164196,1.7353712,2.3286898,2.1263442,1.8965619,1.5398848,1.2003556,1.2655178,1.1283343,1.0117283,0.85739684,0.72021335,0.7476501,0.7476501,0.66533995,0.6173257,0.6962063,0.9568549,1.0082988,0.7613684,0.5693115,0.66191036,1.1592005,0.72364295,0.7888051,1.0631721,1.2998136,1.2826657,1.3478279,1.2209331,1.0563129,0.9328478,0.86082643,1.0871792,1.0631721,0.8162418,0.4698535,0.26407823,0.19548649,0.25721905,0.38754338,0.5178677,0.5418748,0.64476246,0.9911508,1.1900668,1.255229,1.6393428,1.7593783,1.9171394,2.0886188,2.2395205,2.318401,2.301253,2.4727325,2.469303,2.3972816,2.8499873,3.4535947,3.7211025,4.0949273,4.671098,5.219832,5.693115,6.101236,6.375603,6.4887795,6.4407654,6.0875177,5.9812007,5.7582774,5.3570156,5.0106273,5.2781353,5.051782,4.9180284,4.822,4.0846386,2.3458378,1.3101025,0.82996017,0.7339317,0.82996017,1.2415106,1.5810398,1.704505,1.6599203,1.704505,1.4541451,1.0597426,0.71678376,0.4938606,0.32924038,0.26750782,0.28808534,0.3566771,0.44927597,0.5796003,0.5418748,0.45270553,0.40126175,0.4081209,0.45613512,0.5418748,0.6173257,0.64819205,0.64133286,0.6310441,0.65162164,0.65848076,0.6790583,0.7305021,0.8093826,0.4081209,2.1812177,1.4369972,0.5041494,0.29494452,0.28465575,0.15776102,0.06859175,0.0274367,0.020577524,0.024007112,0.030866288,0.017147938,0.01371835,0.05144381,0.15433143,0.058302987,0.082310095,0.09259886,0.05144381,0.01371835,0.0034295875,0.0034295875,0.01371835,0.024007112,0.041155048,0.024007112,0.030866288,0.061732575,0.09602845,0.072021335,0.14404267,0.19891608,0.24350071,0.32924038,0.5727411,1.155771,1.4644338,1.4987297,1.845118,3.6525106,8.615124,11.159878,9.904649,6.1766872,3.998899,2.4761622,1.7799559,1.611906,1.8999915,2.7951138,4.5853586,6.9723516,8.433355,8.776315,9.136421,9.825768,12.528283,15.594335,16.561478,12.164746,8.31332,7.3564653,7.363324,7.208993,6.5470824,11.640019,9.921797,6.619104,5.5902276,9.314759,12.024134,12.343085,16.050468,23.290329,28.554745,29.559614,30.729103,28.582182,24.562706,25.032558,19.133669,16.21852,14.061309,13.762935,19.723558,34.151833,30.93145,21.304598,12.449403,7.4627824,3.3129816,3.6970954,6.783724,9.379922,6.931196,3.6387923,2.585909,2.1400626,1.7936742,2.1640697,4.715683,3.1860867,1.5364552,1.2072148,1.1180456,0.89855194,1.3409687,1.7593783,2.0920484,2.9185789,2.6064866,1.3272504,0.7339317,1.0837497,1.2380811,1.9754424,3.4227283,4.1429415,4.0503426,4.413879,4.4927597,4.2115335,4.8082814,6.029215,6.125243,6.245279,6.3138704,5.501058,4.4756117,5.40503,5.456474,5.219832,5.1580997,5.1169443,4.3452873,5.267846,5.24041,4.856296,4.57164,4.695105,5.4084597,6.574519,6.601956,5.456474,4.6608095,6.5710897,8.069819,8.086967,7.0889573,7.06838,6.5196457,6.842027,7.5107965,8.213862,8.875772,10.463672,10.175586,7.5759587,5.055212,7.822889,9.818909,6.694555,4.5922174,6.8728933,14.105893,7.939495,3.433017,2.4967396,4.9214582,8.388771,6.475061,4.8185706,4.647091,5.56965,5.5559316,5.0757895,5.164959,5.693115,6.40304,6.893471,7.1198235,7.363324,6.989499,6.1492505,5.7651367,4.647091,3.690236,2.9117198,2.469303,2.633923,1.9342873,2.4727325,4.029765,5.346727,4.1326528,2.4452958,1.9308578,1.5536032,1.1043272,1.1832076,1.6633499,1.4404267,1.2998136,1.9308578,3.9200184,3.841138,3.3369887,2.877424,2.4967396,1.7936742,2.061182,2.7882545,3.1826572,2.9563043,2.3389788,2.1846473,2.1572106,2.0680413,1.937717,1.9823016,2.054323,1.5844694,1.2517995,1.214074,1.0871792,0.66533995,0.77165717,2.277246,3.758828,1.5193073,1.4987297,1.6324836,1.5570327,1.2758065,1.1454822,1.155771,1.3992717,1.5947582,1.5810398,1.3066728,1.138623,1.0357354,0.9431366,0.8848336,0.96371406,0.9568549,0.9842916,0.96714365,0.90198153,0.84367853,1.2929544,1.4678634,1.9171394,2.7402403,3.6010668,2.7882545,2.2429502,2.170929,2.301253,1.8965619,5.3844523,4.763697,2.884283,2.3424082,5.4804807,8.186425,6.0669403,3.6627994,3.4364467,5.7754254,5.768566,4.5510626,3.0626216,1.7422304,0.5178677,0.5453044,1.4815818,2.3801336,2.7230926,2.417859,4.0023284,3.590778,2.3321195,1.4747226,2.386993,5.0483527,5.381023,3.5599117,1.5981878,3.3438478,3.0111778,3.2512488,5.7719955,9.870353,12.456262,8.117833,4.9591837,3.8548563,3.998899,2.8980014,3.059192,4.5922174,6.279575,7.2775846,7.0889573,4.3041325,5.1340923,5.360445,3.974892,3.1689389,9.956093,15.433144,11.598865,1.9548649,1.5090185,2.6133456,2.4144297,1.471293,0.48014224,0.3018037,1.2826657,2.3801336,2.9906003,2.8877127,2.2566686,2.428148,2.2120838,2.49331,3.508468,4.839148,4.7431192,7.73372,9.448513,9.14328,9.6988735,10.981539,13.745787,17.785841,20.443771,16.599203,17.388008,19.346302,20.807306,21.325174,21.69557,21.301168,22.899355,25.577864,27.796806,27.395544,25.221186,25.19375,26.133457,26.860529,26.174612,24.617579,22.669573,18.948471,13.766364,9.126132,7.966932,7.6033955,7.3701835,6.5882373,4.5647807,3.316411,2.1023371,4.729401,9.126132,7.332458,4.856296,2.9288676,2.5481834,3.4124396,3.8857226,4.7534084,3.806842,2.2978237,1.2895249,1.6530612,2.07833,2.568761,2.6887965,2.6647894,3.3815732,2.393852,1.8313997,2.3218307,3.350707,3.2615378,6.9963584,4.6573796,2.07833,1.7319417,2.7299516,2.7470996,3.0626216,4.7808447,6.5196457,4.396731,2.952875,3.0111778,3.6627994,4.2286816,4.2286816,3.799983,5.4907694,7.7028537,9.023245,8.23444,5.641671,3.549623,1.7765263,0.6824879,1.1626302,0.7099246,0.4938606,0.39097297,0.36353627,0.44927597,0.4081209,0.41498008,0.4355576,0.4629943,0.4938606,0.34981793,0.2709374,0.25378948,0.28122616,0.31895164,0.34295875,0.33609957,0.32924038,0.33609957,0.33609957,0.5212973,0.6173257,0.85739684,1.4472859,2.5927682,3.2272418,3.1106358,2.8396983,2.8225505,3.2683969,2.9117198,2.7333813,2.5070283,2.1091962,1.5055889,1.5021594,1.4438564,1.3924125,1.3169615,1.0871792,1.5707511,1.3203912,0.84024894,0.44927597,0.2709374,0.36353627,0.53844523,0.6790583,0.7339317,0.7133542,0.59331864,0.45956472,0.33609957,0.3018037,0.5007198,0.5144381,0.6276145,0.66191036,0.7613684,1.4129901,1.7216529,1.2312219,1.3992717,2.3218307,2.7162333,4.0503426,4.7842746,5.31929,5.470192,4.4927597,5.099797,7.5588107,8.954653,8.131552,5.669108,5.312431,5.953764,7.579388,8.985519,7.7783046,9.167287,11.338216,10.185875,6.307011,5.0106273,12.435684,14.685493,13.718349,10.628291,5.65539,6.4887795,6.1904054,4.4721823,2.5721905,3.2512488,1.6736387,0.51100856,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.16462019,0.490431,0.86082643,1.1008976,1.0117283,1.3478279,1.3546871,1.1317638,0.91569984,1.0734608,1.0185875,0.9259886,0.82996017,0.66876954,0.26750782,0.33609957,0.36696586,0.6001778,0.96371406,1.097468,0.89512235,0.77508676,0.66876954,0.5521636,0.4629943,0.16804978,0.05144381,0.048014224,0.11317638,0.22978236,0.30523327,0.44584638,0.7133542,0.94999576,0.7579388,1.1660597,1.2758065,1.4541451,1.845118,2.3732746,2.386993,2.1194851,1.6667795,1.2998136,1.4507155,1.3203912,0.9842916,0.7305021,0.64819205,0.6241849,0.72707254,0.83338976,0.91912943,0.9842916,1.0597426,1.097468,0.71678376,0.3566771,0.39097297,1.1214751,0.6241849,0.6310441,0.90884066,1.2072148,1.2586586,1.1351935,1.0357354,1.0048691,0.96371406,0.7305021,0.8676856,0.7956643,0.6001778,0.3841138,0.274367,0.23664154,0.33609957,0.4664239,0.58302987,0.66876954,0.61046654,0.84024894,1.0563129,1.2517995,1.7250825,2.0234566,2.1091962,2.1983654,2.3252604,2.3321195,2.486451,2.6887965,2.8225505,3.0146074,3.6353626,4.8322887,5.3741636,5.871454,6.4544835,6.7802944,7.250148,7.723431,7.675417,7.0752387,6.39961,5.953764,5.874883,5.7754254,5.5387836,5.3227196,5.3570156,5.4187484,5.686256,5.7377,4.5613513,2.3595562,1.2243627,0.8676856,0.94999576,1.0700313,1.3752645,1.5398848,1.6290541,1.6393428,1.4747226,1.2415106,0.922559,0.6241849,0.39440256,0.25378948,0.23664154,0.23664154,0.26750782,0.32924038,0.41840968,0.4355576,0.42183927,0.39783216,0.432128,0.6276145,0.6344737,0.65505123,0.64476246,0.607037,0.607037,0.70649505,0.75450927,0.77851635,0.7888051,0.8025235,0.45613512,2.7779658,1.978872,0.88826317,0.607037,0.51100856,0.22978236,0.08916927,0.034295876,0.020577524,0.017147938,0.017147938,0.006859175,0.024007112,0.09259886,0.22292319,0.09602845,0.09945804,0.082310095,0.024007112,0.01371835,0.05144381,0.034295876,0.030866288,0.044584636,0.037725464,0.037725464,0.07888051,0.14747226,0.22978236,0.274367,0.39097297,0.42869842,0.38754338,0.4389872,0.922559,1.3821237,1.6804979,2.3081124,4.2835546,9.156999,15.782962,16.997036,13.179905,7.2124224,4.4859004,2.7539587,2.0646117,1.9548649,2.5310357,4.4687524,6.461343,8.347616,9.225591,9.122703,8.988949,9.14328,12.130451,16.239098,18.12537,12.809509,9.331907,8.447074,7.8503256,6.9620624,6.924337,9.191295,7.1026754,5.501058,6.9620624,11.780633,11.087856,11.650309,19.250275,32.491913,42.777245,41.92671,33.054363,25.660173,24.891945,31.538486,22.77589,13.680624,9.270175,10.103564,12.264205,17.583494,16.417435,13.872682,11.362224,6.608815,3.0489032,2.1640697,3.3884325,5.2335505,5.302142,2.7951138,2.0097382,1.9548649,1.8176813,0.94999576,2.568761,2.0268862,1.529596,1.6804979,1.5090185,1.7353712,2.867135,3.4055803,3.525616,5.079219,5.3158607,4.5167665,3.9337368,3.875434,3.7279615,3.4913201,3.4535947,3.3266997,3.2581081,3.8205605,3.9508848,3.9268777,4.996909,6.8385973,7.5519514,7.226141,6.711703,5.579939,4.7842746,6.6739774,6.691125,5.878313,5.8474464,6.385892,5.4324665,6.029215,6.1458206,5.953764,6.0395036,7.4113383,7.9875093,8.522525,7.870903,6.3790326,5.885172,6.636252,6.40304,6.0395036,6.2830043,7.7577267,6.9654922,7.1884155,7.8983397,8.927217,10.436234,13.437123,14.38026,11.598865,7.48336,8.48137,8.783174,6.427047,4.996909,7.284444,15.275383,5.2609873,2.6476414,3.5770597,5.717122,8.255017,6.7185616,5.144381,4.856296,5.5833683,5.4770513,4.5784993,6.0737996,6.8866115,6.1321025,5.0929375,4.7808447,4.870014,5.1752477,5.857735,7.4181976,8.128122,5.6210938,2.959734,1.7319417,2.0303159,1.879414,2.5584722,3.5873485,4.125794,2.9494452,1.7971039,1.3615463,1.1592005,1.0425946,1.2072148,1.2517995,1.0117283,1.1832076,2.0474637,3.4673128,3.2135234,3.3301294,3.508468,3.2478194,1.862266,2.5584722,3.3301294,3.649081,3.1483612,1.6187652,1.6084765,1.8108221,1.9994495,1.99602,1.6496316,1.6770682,1.3341095,1.1008976,1.0323058,0.7922347,0.4972902,0.66533995,2.136633,3.6456516,1.8142518,1.4472859,1.4129901,1.488441,1.546744,1.5707511,1.3992717,1.3478279,1.4129901,1.5364552,1.6221949,1.3684053,0.9842916,0.823101,1.0734608,1.7456601,1.5330256,1.4850113,1.4541451,1.3684053,1.2312219,1.7799559,2.095478,2.0989075,1.9754424,2.1434922,1.3992717,1.1523414,1.7525192,2.5893385,2.0749004,4.125794,3.1140654,1.786815,2.386993,6.6396813,10.436234,8.069819,5.178677,4.7945633,7.301592,6.557371,3.5804894,1.3478279,0.91227025,1.3992717,1.2792361,1.7490896,4.1943855,6.9826403,5.456474,4.2183924,3.0557625,2.5138876,3.1963756,5.754848,7.658269,6.0052075,3.2615378,1.6599203,3.1860867,2.9940298,4.972902,7.06495,7.740579,6.0154963,3.192946,2.620205,3.1209247,3.4673128,2.3561265,2.7059445,4.4550343,6.108095,6.842027,6.5024977,2.6647894,2.0646117,2.952875,3.525616,1.9239986,6.3481665,10.947243,8.587687,1.3684053,0.6001778,1.8279701,1.845118,1.0666018,0.28808534,0.7099246,2.760818,3.508468,3.1449318,2.287535,1.9651536,1.646202,1.8519772,3.450165,6.025785,7.915488,6.464772,8.440215,9.764035,9.345626,9.074688,12.548861,14.225929,17.63151,21.098822,17.799559,17.364002,19.017063,19.363451,18.169954,18.37916,19.648108,22.378057,25.111439,26.51757,25.392666,28.002583,29.058895,28.52731,27.700777,29.209797,29.449867,24.648445,19.45262,15.54632,11.63659,9.030104,8.587687,9.153569,9.239308,7.0306544,4.4584637,2.8877127,5.1580997,9.427936,9.156999,7.0135064,3.882293,2.503599,3.1483612,3.6285036,4.1120753,4.15323,3.309552,2.16064,2.301253,1.9685832,2.2429502,2.020027,1.5124481,2.2395205,2.4144297,2.2360911,2.8877127,4.0537724,3.9028704,11.074138,9.740028,5.8165803,2.9700227,2.609916,2.301253,2.3424082,2.9082901,3.5187566,3.0489032,3.7211025,3.7451096,3.8960114,4.5030484,5.470192,4.928317,6.8557453,8.724871,9.277034,8.556821,6.3824625,4.6676683,3.2203827,2.335549,2.7985435,1.5673214,0.7922347,0.4698535,0.4664239,0.4972902,0.4629943,0.4424168,0.4355576,0.432128,0.44584638,0.37382504,0.30866286,0.28122616,0.30866286,0.39097297,0.42526886,0.39440256,0.34981793,0.30866286,0.26750782,0.36696586,0.6207553,1.039165,1.6359133,2.4590142,2.9700227,2.9871707,3.1689389,3.7211025,4.40359,3.7382503,3.450165,3.4844608,3.5461934,3.0969174,2.8019729,2.3321195,2.2052248,2.4144297,2.4247184,2.6373527,2.3972816,1.7319417,1.0117283,0.94999576,1.1249046,0.939707,0.8711152,1.0528834,1.2586586,0.764798,0.4629943,0.33952916,0.34981793,0.39783216,0.6859175,0.4698535,0.432128,0.77851635,1.255229,1.5947582,1.2175035,1.3341095,1.9994495,2.1229146,2.6956558,3.9268777,5.1580997,5.6348124,4.5030484,4.8494368,6.279575,7.6342616,7.9600725,6.5196457,6.8145905,8.093826,10.360784,12.21619,10.854645,12.332796,13.848674,11.657167,7.2707253,7.4353456,12.569438,13.3033695,13.101024,12.295071,8.114404,8.567109,7.0923867,5.8200097,5.662249,6.279575,3.875434,1.9548649,0.97057325,0.65505123,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.082310095,0.29837412,0.64819205,0.97400284,1.0082988,1.3889829,1.6221949,1.4987297,1.2689474,1.646202,1.1900668,0.922559,0.7099246,0.48357183,0.2194936,0.26407823,0.36010668,0.6962063,1.1180456,1.1351935,0.9431366,0.82996017,0.7133542,0.59331864,0.5727411,0.1920569,0.06516216,0.09945804,0.216064,0.34638834,0.44584638,0.5178677,0.6859175,0.89169276,0.8779744,1.1180456,1.3615463,1.7456601,2.1983654,2.428148,2.3492675,2.1469216,1.7936742,1.4267083,1.3409687,1.3032433,0.9534253,0.71678376,0.6859175,0.6241849,0.6962063,0.86082643,0.96714365,0.9568549,0.881404,0.8093826,0.50757897,0.22292319,0.19548649,0.6344737,0.38754338,0.5212973,0.78537554,1.0048691,1.08032,0.9328478,0.8471081,0.86082643,0.89855194,0.77165717,0.7476501,0.5521636,0.36696586,0.274367,0.24350071,0.20920484,0.32238123,0.5418748,0.77851635,0.91912943,0.8025235,0.91569984,1.1351935,1.4678634,2.0406046,2.2258022,2.2978237,2.3424082,2.3629858,2.2635276,2.9322972,3.3026927,3.4433057,3.57363,4.0606318,5.0174866,5.5250654,6.111525,6.8111606,7.1952744,7.689135,7.9257765,7.6205435,6.9380555,6.492209,6.3721733,6.2487082,5.967482,5.6176643,5.5490727,5.562791,5.3673043,5.5319247,5.7651367,4.9420357,2.5173173,1.2655178,0.8779744,0.96371406,1.0768905,1.2346514,1.3409687,1.4369972,1.4815818,1.3341095,1.1317638,0.8779744,0.59331864,0.34295875,0.24007112,0.2777966,0.23321195,0.22292319,0.2777966,0.36353627,0.4081209,0.4424168,0.44584638,0.47328308,0.65848076,0.6379033,0.6207553,0.58988905,0.5555932,0.5658819,0.66533995,0.7133542,0.7442205,0.77165717,0.77851635,0.84367853,2.3286898,1.903421,1.2723769,1.0597426,0.7888051,0.2777966,0.106317215,0.06859175,0.044584636,0.0034295875,0.020577524,0.01371835,0.037725464,0.1097468,0.20920484,0.116605975,0.09945804,0.06859175,0.017147938,0.017147938,0.12689474,0.10288762,0.08573969,0.10288762,0.07888051,0.09259886,0.17490897,0.28465575,0.4081209,0.5693115,0.7305021,0.8025235,0.70649505,0.7099246,1.4061309,1.3889829,2.0749004,4.249259,9.091836,18.159666,25.697899,24.058556,17.072487,9.187865,5.4633327,3.4295874,2.767677,2.8019729,3.6799474,6.385892,8.385342,8.865483,8.9100685,8.718011,7.6033955,8.2310095,11.543991,16.45859,19.836735,16.489456,11.856084,9.781183,8.570539,7.7920227,8.282454,6.697984,5.669108,7.301592,11.218181,14.544881,11.05356,14.256795,25.59844,43.31226,62.442497,62.5934,42.23194,25.622448,22.319756,27.165762,23.451519,16.935303,13.121602,11.626302,6.169828,3.899441,4.5784993,6.715132,7.9463544,5.020916,2.3904223,1.1592005,1.1832076,1.8588364,2.1091962,0.864256,0.91227025,1.9720128,2.8156912,1.2689474,1.0048691,1.0220171,1.5364552,2.2738166,2.486451,3.450165,5.0277753,5.802862,5.909179,7.006647,8.056101,8.735159,9.050681,8.985519,8.505377,7.0615206,5.7274113,4.5030484,3.4467354,2.6545007,2.5138876,3.2032347,4.9831905,7.010077,7.3255987,6.4373355,5.953764,5.4324665,5.6005163,8.354475,7.6342616,6.478491,6.3447366,7.1129646,7.0958166,6.4544835,6.4819202,6.5813785,7.431916,10.978109,10.7586155,9.349055,8.309891,8.011517,7.630832,6.334448,5.24041,5.2472687,6.427047,8.018375,7.3530354,7.363324,7.548522,8.049242,9.661148,14.733508,18.849012,17.099922,11.2421875,9.674867,8.210432,6.5127864,5.8165803,8.128122,16.194511,6.0703697,4.0057583,4.7774153,5.703404,6.6431108,4.705394,4.1155047,4.4275975,4.945465,4.7191124,4.15666,6.2418494,7.2295704,5.9160385,3.666229,3.82399,3.3472774,3.2958336,4.4687524,7.3873315,10.182446,6.7631464,3.210094,2.1091962,2.527606,2.1743584,2.1400626,2.369845,2.5207467,1.9891608,1.5776103,1.2929544,1.2449403,1.4369972,1.7765263,1.1317638,0.7990939,0.9877212,1.6324836,2.3972816,1.6084765,2.335549,3.6696587,4.1943855,1.9720128,2.8980014,3.6525106,4.170378,3.7931237,1.2895249,1.1729189,1.4472859,1.8039631,1.9891608,1.7799559,1.3821237,1.2175035,1.0323058,0.72707254,0.34638834,0.31552204,0.5590228,1.4061309,2.3218307,1.8999915,1.7490896,1.6016173,1.6530612,1.9068506,2.1743584,1.6770682,1.4232788,1.3341095,1.4061309,1.6907866,1.7113642,1.4335675,1.255229,1.4644338,2.2429502,1.6084765,1.3409687,1.3306799,1.3684053,1.1420527,1.4644338,2.2600982,2.2909644,1.6427724,1.7113642,2.1194851,1.5536032,1.7971039,2.7779658,2.568761,2.5824795,1.670209,1.0666018,2.020027,5.796003,8.217292,7.157549,5.4633327,4.7019644,5.137522,3.1620796,1.1832076,0.6310441,1.6221949,2.9665933,2.452155,3.0111778,7.239859,12.020704,8.519095,3.2032347,1.728512,2.4247184,4.4447455,7.7714453,7.3118806,4.3109913,2.177788,2.2326615,3.7142432,4.773986,7.3839016,8.491658,6.56766,1.5844694,1.0871792,2.9494452,4.262977,3.9097297,2.551613,2.877424,3.9714622,4.232111,3.5187566,3.1586502,2.0131679,1.978872,3.4192986,4.4859004,1.1249046,1.6599203,4.523626,4.8425775,2.1915064,0.61389613,0.75450927,0.5658819,0.30866286,0.4355576,1.5604624,4.057202,4.540774,3.0557625,1.0151579,1.1934965,0.90198153,2.0714707,5.103226,8.707723,9.911508,6.6053853,7.5519514,8.484799,8.1041155,8.069819,15.395418,16.47231,18.341434,21.976797,22.299177,19.723558,18.571217,17.20967,16.321407,18.924463,19.45262,21.469217,23.35549,23.921373,22.422644,30.050045,31.631084,29.881996,28.17406,30.51647,31.09264,24.507832,18.862732,16.352274,13.251926,10.192734,10.182446,11.190743,11.4376745,9.403929,6.776865,4.8322887,5.2164025,7.689135,10.131001,8.656279,5.353586,3.216953,3.3541365,4.972902,4.9008803,5.2575574,4.7602673,3.4467354,2.668219,2.6579304,2.3081124,2.0028791,2.287535,3.8720043,3.0317552,3.0866287,3.3266997,3.1826572,2.201795,10.868362,14.445422,11.581717,5.2506986,2.7711067,1.7936742,1.9925903,2.8499873,4.0194764,5.3330083,6.012067,4.3487167,4.064061,5.552502,5.885172,6.0395036,8.06639,8.776315,8.124693,9.201583,7.3393173,5.8988905,5.127233,4.880303,4.6127954,2.4727325,1.2003556,0.65162164,0.5796003,0.6241849,0.5727411,0.53844523,0.5144381,0.48700142,0.42869842,0.3841138,0.33609957,0.33266997,0.37725464,0.44584638,0.48357183,0.4424168,0.37725464,0.33266997,0.34295875,0.36696586,0.5624523,1.0837497,1.7833855,2.1983654,2.5961976,2.767677,3.4433057,4.65395,5.7239814,4.297273,3.6182148,3.765687,4.389872,4.7019644,4.091498,2.7642474,2.4144297,3.2683969,4.0709205,3.7279615,3.4844608,2.8705647,2.0714707,1.9342873,2.3458378,1.7079345,1.255229,1.4507155,1.9925903,1.0117283,0.5624523,0.50757897,0.5658819,0.31552204,0.5761707,0.44927597,0.3806842,0.5144381,0.6824879,1.2003556,1.1283343,1.6530612,2.6716487,2.7813954,1.7799559,3.1415021,4.1463714,4.4447455,6.0806584,7.5553813,7.349606,7.133542,7.531374,8.097256,10.185875,11.787492,13.179905,13.732068,11.931535,13.296511,12.428825,9.993818,7.997798,9.798331,10.844356,8.354475,8.282454,10.947243,11.067279,7.8983397,6.5950966,7.1061053,8.258447,7.7611566,5.3913116,3.542764,2.5241764,1.8656956,0.34638834,0.12689474,0.05144381,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.08916927,0.23664154,0.52472687,0.8848336,1.1043272,1.3786942,1.5913286,1.605047,1.6187652,2.1846473,1.2483698,0.64819205,0.28808534,0.1097468,0.07888051,0.11317638,0.33266997,0.7407909,1.1763484,1.3101025,1.1214751,0.9911508,0.8093826,0.58988905,0.47328308,0.15433143,0.06859175,0.15090185,0.29837412,0.37382504,0.5007198,0.5007198,0.6207553,0.881404,1.0666018,1.3032433,1.7113642,2.1812177,2.5241764,2.49331,2.1229146,2.0097382,1.8485477,1.5433143,1.2312219,1.3992717,1.1729189,0.9328478,0.82996017,0.75450927,0.72364295,0.77851635,0.7613684,0.64476246,0.5453044,0.31552204,0.22635277,0.14061308,0.037725464,0.0274367,0.13375391,0.41498008,0.64133286,0.7510797,0.84367853,0.94999576,0.8196714,0.7099246,0.7339317,0.8676856,0.77851635,0.48357183,0.274367,0.22635277,0.1920569,0.12003556,0.22978236,0.5590228,0.96371406,1.1111864,1.097468,1.1832076,1.3581166,1.7147937,2.4555845,2.3458378,2.4727325,2.534465,2.4315774,2.277246,3.391862,3.9440255,4.040054,4.0229063,4.4550343,4.448175,4.530485,5.0174866,5.878313,6.711703,7.3084507,7.160979,6.756287,6.5127864,6.7665763,7.1026754,6.9346256,6.3721733,5.754848,5.6828265,5.813151,5.127233,4.938606,5.312431,5.07236,2.6613598,1.3786942,0.85739684,0.78194594,0.881404,1.0048691,1.2346514,1.3855534,1.4335675,1.4987297,1.2449403,1.0185875,0.7407909,0.45270553,0.32581082,0.34981793,0.28465575,0.25721905,0.32238123,0.432128,0.45270553,0.4664239,0.45956472,0.44584638,0.4664239,0.5041494,0.50757897,0.4972902,0.48357183,0.4972902,0.5007198,0.490431,0.53158605,0.6276145,0.71678376,2.2120838,2.9940298,2.1640697,1.3101025,1.0700313,1.1454822,0.48357183,0.20920484,0.14404267,0.12346515,0.01371835,0.09945804,0.06859175,0.06859175,0.13375391,0.18176813,0.12346515,0.17147937,0.13375391,0.017147938,0.030866288,0.12689474,0.15090185,0.16462019,0.18862732,0.21263443,0.17833854,0.23321195,0.29151493,0.34981793,0.47328308,0.77851635,1.0940384,1.2072148,1.2106444,1.4815818,1.9308578,4.681387,9.654288,17.71039,30.622786,35.10526,27.68363,17.63494,10.209882,6.6225333,4.314421,3.8925817,4.280125,4.9831905,6.118384,8.255017,9.860064,11.372512,11.585147,7.630832,7.1884155,9.239308,13.996146,18.235117,15.306249,11.910957,10.80663,10.39165,10.161868,10.710602,7.5245147,8.687145,12.418536,15.326826,12.421966,10.39508,13.687484,27.169191,51.666737,83.95287,87.4922,61.883476,35.81518,21.819035,16.266533,10.189304,11.962401,13.920695,12.836946,9.918367,6.914048,4.588788,4.5853586,6.0806584,5.813151,3.117495,1.5158776,0.83338976,0.71678376,0.65505123,0.29151493,0.52815646,1.529596,2.5378947,1.8931323,1.7319417,1.3546871,1.4027013,1.8416885,1.937717,3.865145,6.0154963,7.606825,8.680285,10.069269,11.118723,10.943813,10.419086,9.616563,7.798882,6.2487082,5.15467,4.0434837,3.0454736,2.8980014,1.8485477,3.0866287,5.1340923,6.495639,5.675967,4.8082814,4.8494368,4.7808447,4.863155,6.608815,6.2898636,6.6053853,6.7322803,6.8385973,8.073249,7.9875093,7.0786686,6.217842,7.630832,14.908417,9.767465,7.3393173,8.021805,10.216741,10.316199,7.5553813,6.2247014,6.6053853,7.8366075,7.936065,6.6053853,6.684266,6.550512,6.427047,8.3922,16.715809,22.587263,20.762722,13.310229,9.613133,7.0375133,5.9812007,6.0806584,7.64798,11.688034,9.661148,7.205563,5.545643,5.9126086,9.537683,4.972902,3.7485392,3.7725463,3.74168,3.1449318,2.6785078,2.6373527,2.8499873,2.9700227,2.4555845,4.32471,4.773986,4.1326528,3.4707425,4.5922174,4.448175,3.083199,2.0337453,1.9651536,2.6853669,2.037175,1.611906,1.4541451,1.488441,1.5261664,1.6599203,1.4541451,1.6016173,1.9582944,1.5570327,1.2620882,1.0254467,0.84367853,0.881404,1.4815818,1.7010754,1.7456601,1.8725548,1.9582944,1.4953002,1.2895249,1.7765263,2.4795918,2.644212,1.2517995,1.3615463,1.2895249,1.2517995,1.3272504,1.4507155,1.4129901,1.4027013,1.2620882,0.9568549,0.5796003,0.37382504,0.7682276,1.3443983,1.6564908,1.2655178,1.6804979,1.7388009,1.8005334,2.0303159,2.3972816,1.845118,1.728512,1.6839274,1.5913286,1.5570327,1.99602,2.3081124,2.4418662,2.2806756,1.6324836,1.2415106,0.9259886,0.99801,1.2758065,1.0666018,1.0323058,1.6530612,2.0028791,2.1263442,3.0660512,3.542764,2.5173173,1.8108221,2.0920484,2.8980014,2.0817597,1.3992717,1.3649758,1.8519772,2.1229146,2.8534167,2.836269,2.4555845,2.1091962,2.1812177,0.99801,0.31895164,0.7339317,2.0028791,3.0523329,1.1729189,2.5893385,6.5196457,9.469091,5.2335505,2.095478,1.7593783,2.0406046,2.085189,2.3664153,1.3272504,1.0700313,1.3375391,2.0646117,3.3712845,2.177788,2.428148,2.7745364,2.428148,1.1454822,2.1332035,4.3933015,6.159539,6.200694,3.8445675,2.551613,2.8877127,3.2581081,3.6456516,5.6005163,6.5642304,6.1629686,6.036074,5.470192,1.4198492,1.1626302,3.3232703,4.863155,4.2252517,1.3581166,0.5041494,0.22635277,0.19548649,0.58302987,2.061182,2.486451,1.670209,0.71678376,0.216064,0.22978236,0.5693115,2.0749004,4.249259,6.090947,6.1046658,2.9906003,5.7754254,7.805741,6.848886,5.0655007,8.594546,11.7086115,12.723769,12.80265,15.9750185,16.62321,16.005884,16.074476,18.156237,22.964518,20.19341,19.510923,21.561817,24.35007,23.238884,30.1838,30.245531,27.951138,27.234354,31.432169,27.27208,21.78131,18.588364,17.816708,16.081335,13.433694,14.208781,14.586036,12.9809885,10.041832,8.464222,6.3310184,4.835718,5.188966,8.604835,9.911508,8.021805,4.99005,3.923448,9.002667,7.610255,5.4324665,3.9474552,3.508468,3.3266997,2.935727,2.3149714,1.9857311,2.2120838,3.0077481,1.8828435,1.4918705,2.0646117,3.069481,3.2032347,6.975781,12.891819,13.066729,7.116394,2.136633,1.6496316,2.3492675,4.0949273,5.8337283,5.6142344,9.448513,8.89635,9.132992,9.606275,4.029765,6.420188,8.162418,7.8091707,6.478491,7.857185,8.261876,8.069819,6.8283086,5.038064,4.1360826,2.3767042,1.2895249,0.70306545,0.5727411,0.9774324,0.7682276,0.72707254,0.70649505,0.6241849,0.4424168,0.4046913,0.4424168,0.4664239,0.4698535,0.5178677,0.5178677,0.48357183,0.39783216,0.30523327,0.30523327,0.47671264,0.58302987,1.1249046,2.0028791,2.503599,2.4041407,2.627064,3.4638834,4.5784993,5.003768,3.7725463,2.6956558,2.510458,3.275256,4.3487167,3.8857226,2.5790498,2.469303,3.74168,4.729401,4.8288593,4.3109913,3.724532,3.2032347,2.4727325,2.9220085,2.7333813,2.3424082,2.07833,2.1503513,1.1489118,0.5693115,0.4424168,0.4972902,0.16804978,0.20577525,0.34981793,0.48014224,0.48700142,0.30523327,0.59674823,0.45956472,0.7956643,1.5364552,1.6324836,2.9391565,4.5099077,4.712253,4.3349986,6.6053853,8.999237,10.120712,10.998687,11.30735,9.352485,10.477389,12.05843,12.120162,10.542552,9.0644,8.940934,9.211872,8.779744,7.4936485,6.1492505,5.8062916,4.972902,4.5510626,5.219832,7.414768,4.170378,5.453044,7.301592,7.846896,7.3084507,4.636802,3.2615378,2.8945718,2.7882545,1.7388009,0.6276145,0.2503599,0.1097468,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.037725464,0.18176813,0.53158605,0.9568549,1.1283343,1.2277923,1.1694894,1.155771,1.1832076,1.039165,0.40126175,0.13375391,0.0548734,0.041155048,0.030866288,0.0548734,0.2709374,0.6001778,0.9568549,1.2346514,1.3203912,1.3615463,1.2072148,0.8265306,0.29151493,0.106317215,0.07888051,0.17147937,0.3018037,0.34981793,0.4972902,0.5418748,0.58645946,0.70306545,0.94656616,1.3375391,2.0097382,2.3767042,2.4452958,2.8225505,2.4452958,1.9823016,1.7525192,1.8142518,1.9994495,2.4007113,1.9239986,1.2792361,0.8505377,0.71678376,0.8162418,0.8196714,0.70649505,0.48357183,0.22978236,0.09602845,0.28122616,0.28808534,0.06516216,0.01371835,0.0034295875,0.14747226,0.40126175,0.6241849,0.5658819,0.9431366,0.7990939,0.59331864,0.52472687,0.548734,0.64819205,0.432128,0.26750782,0.24007112,0.16804978,0.106317215,0.23664154,0.5418748,0.89169276,1.039165,1.2586586,1.3306799,1.4232788,1.7113642,2.3972816,2.1743584,2.386993,2.452155,2.3629858,2.6545007,3.5942078,3.7279615,3.8034124,4.32128,5.552502,5.4187484,5.284994,5.5113473,6.3447366,7.9189177,8.323608,7.963502,7.531374,7.2535777,6.910619,6.9380555,6.9346256,6.9654922,6.975781,6.8043017,6.427047,6.368744,6.5470824,6.3035817,4.4241676,2.3732746,1.4678634,1.0906088,0.90541106,0.8711152,1.1489118,1.3958421,1.5913286,1.6804979,1.5707511,1.2312219,1.2449403,1.196926,0.9362774,0.59674823,0.42526886,0.3806842,0.37382504,0.3841138,0.45613512,0.45613512,0.5041494,0.5212973,0.5041494,0.5041494,0.5418748,0.53158605,0.4938606,0.44927597,0.4115505,0.37382504,0.3566771,0.39440256,0.4972902,0.65505123,2.3835633,3.6627994,2.4795918,1.3101025,1.0597426,1.0837497,0.5418748,0.35324752,0.34638834,0.33609957,0.1371835,0.106317215,0.072021335,0.048014224,0.041155048,0.061732575,0.16462019,0.116605975,0.048014224,0.024007112,0.06859175,0.21263443,0.26407823,0.23321195,0.15433143,0.09259886,0.30866286,0.41840968,0.4355576,0.53844523,1.0700313,1.728512,1.5947582,1.3169615,1.3101025,1.7730967,4.3041325,12.936404,24.085993,32.49877,31.246971,27.17262,20.087093,13.042721,7.963502,5.6348124,4.3624353,4.506478,5.6176643,7.3118806,9.266746,11.657167,12.154458,11.417097,9.657719,6.6396813,7.9600725,12.46312,17.851004,20.663265,16.269962,11.002116,11.454823,12.545431,11.63659,8.56368,8.158989,10.72089,12.452832,12.768354,14.287662,14.565458,15.536031,24.981115,43.758106,65.8035,58.838,46.70412,36.586838,29.830551,21.95279,14.21564,14.068168,13.810948,10.957532,8.244728,6.697984,4.400161,2.7642474,2.277246,2.5173173,3.940596,3.7691166,2.5173173,1.0323058,0.47328308,0.9842916,5.7068334,7.7028537,5.7822843,4.479041,4.4275975,4.619654,4.448175,3.8137012,3.1209247,3.1277838,4.2081037,6.3790326,8.875772,10.179015,7.8023114,6.7322803,6.433906,6.2830043,5.576509,4.386442,3.642222,3.2718265,3.3884325,4.266407,3.175798,4.0023284,5.2815647,5.7754254,4.479041,3.690236,4.190956,5.3913116,6.1801167,4.897451,4.8734436,6.924337,7.7268605,7.208993,8.56025,10.7586155,9.403929,7.579388,6.958633,7.7783046,4.972902,4.2046742,4.9420357,6.5162163,8.117833,7.857185,7.6959944,9.129561,10.624862,7.6171136,6.715132,7.891481,8.875772,8.745448,7.9292064,10.39508,11.190743,10.645439,9.5205345,9.016385,6.9963584,6.6053853,7.4181976,8.766026,9.760606,9.959522,8.916927,6.9963584,5.693115,7.606825,6.478491,6.8111606,5.977771,3.9646032,3.3884325,3.216953,2.9906003,3.1552205,4.149801,6.4098988,6.8145905,6.632822,5.3570156,3.724532,3.7279615,2.5927682,2.294394,2.1846473,2.0131679,1.903421,1.8142518,1.8931323,1.920569,1.8897027,2.0131679,1.9342873,1.704505,1.587899,1.5741806,1.3855534,1.2963841,1.1763484,1.1832076,1.471293,2.1743584,1.7422304,1.5501735,1.5021594,1.5536032,1.7147937,1.5844694,1.7422304,1.7799559,1.7456601,2.1297739,1.5673214,1.1043272,1.0254467,1.2415106,1.3169615,1.0837497,0.8196714,0.65505123,0.6241849,0.66533995,0.4972902,0.4938606,0.6859175,0.9774324,1.1454822,1.255229,1.2963841,1.371835,1.4781522,1.4918705,1.862266,1.786815,1.6564908,1.6221949,1.605047,1.2620882,1.430138,1.5981878,1.5021594,1.1214751,0.7682276,0.70306545,0.9431366,1.196926,0.8711152,1.255229,1.4129901,1.3992717,2.0817597,5.130663,7.14726,5.038064,3.0386145,2.726522,2.983741,2.568761,2.3321195,2.3149714,2.3149714,1.8999915,1.3341095,1.5398848,1.6256244,1.3512574,1.1317638,0.72021335,0.3566771,0.7339317,2.318401,5.3570156,3.4776018,3.292404,4.3761535,4.98662,2.061182,1.9411465,4.2423997,5.055212,3.5187566,1.8142518,1.762808,1.3341095,1.196926,1.5501735,2.1023371,2.5173173,3.99204,5.295283,5.06893,1.8142518,1.9925903,4.2218223,7.720001,10.1481495,7.6171136,4.6916757,3.000889,2.7230926,3.666229,5.2575574,7.1095347,6.2658563,4.0846386,1.7902447,0.490431,3.0386145,7.208993,7.140401,2.9117198,0.5521636,0.4389872,0.37039545,0.33609957,0.7133542,2.2806756,1.5844694,0.77165717,0.29151493,0.2194936,0.24007112,1.5021594,2.867135,4.07435,4.554492,3.4433057,2.8294096,5.813151,7.5931067,7.016936,6.591667,8.597976,11.931535,15.542891,17.693241,15.964729,17.665806,19.672113,19.425184,17.78927,19.03421,16.664366,16.444872,19.833303,24.548986,24.569565,27.628757,28.630196,29.127487,30.938309,36.14442,31.229824,25.303495,20.776442,18.45461,17.511473,17.343424,19.03078,19.301718,17.113642,13.653188,10.847785,8.035523,6.615674,6.8900414,8.032094,10.539123,9.705732,6.4990683,4.1017866,7.881192,9.523964,7.7097125,4.9420357,3.223812,4.046913,3.1689389,3.275256,3.117495,2.3458378,1.529596,1.862266,2.0165975,3.0043187,4.6779575,5.7308407,4.280125,5.994919,6.2898636,4.081209,1.8073926,2.1469216,2.3561265,2.1434922,1.8656956,2.5138876,3.5633414,4.2355404,5.3432975,5.909179,3.1620796,6.138962,6.3824625,5.9983487,6.3378778,7.98065,7.160979,6.893471,6.464772,5.813151,5.5250654,3.6525106,2.0063086,1.1351935,1.0631721,1.2826657,0.8196714,0.8025235,0.7990939,0.64476246,0.4424168,0.5041494,0.45613512,0.40126175,0.4389872,0.65162164,0.84024894,0.67219913,0.48357183,0.4081209,0.37725464,0.40126175,0.6790583,1.1317638,1.5776103,1.6976458,1.9514352,2.6990852,3.4295874,3.799983,3.649081,3.0111778,2.054323,1.3889829,1.196926,1.2346514,2.1091962,3.5118976,4.417309,4.40359,3.642222,3.340418,3.1655092,2.7299516,2.1023371,1.786815,2.7299516,3.4878905,3.0146074,1.8108221,1.9308578,1.4575747,1.3306799,1.1763484,0.9568549,0.99801,0.7613684,0.4664239,0.36353627,0.71678376,1.7833855,2.3767042,2.0508933,2.1332035,2.3321195,0.7305021,1.4987297,4.7808447,7.130112,7.5450926,7.4627824,10.089847,11.105004,11.036412,10.192734,8.669997,10.329918,11.482259,11.660598,10.628291,8.378482,8.083538,8.4264965,8.4093485,6.9620624,2.9631636,4.262977,4.297273,3.2718265,2.8225505,6.036074,5.2609873,4.4516044,3.7931237,4.0263357,6.468202,5.305572,4.1429415,3.5770597,3.2443898,1.8142518,1.4644338,0.881404,0.33952916,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.037725464,0.07888051,0.2777966,0.59331864,0.823101,0.980862,0.9877212,0.9911508,0.9602845,0.6962063,0.33609957,0.13375391,0.044584636,0.020577524,0.017147938,0.14061308,0.607037,0.980862,1.1111864,1.138623,0.823101,0.6310441,0.4938606,0.35324752,0.16804978,0.072021335,0.082310095,0.18176813,0.30866286,0.33952916,0.44584638,0.65848076,0.77851635,0.8745448,1.2758065,1.6564908,2.0714707,2.2086544,2.1160555,2.2120838,1.7559488,2.153781,2.609916,2.9082901,3.415869,3.0557625,2.4487255,1.7182233,1.0871792,0.8745448,0.7990939,0.607037,0.4081209,0.23664154,0.058302987,0.1097468,1.4335675,1.903421,1.0734608,0.18519773,0.037725464,0.030866288,0.216064,0.4629943,0.4424168,0.70306545,0.7579388,0.77165717,0.78537554,0.7339317,0.7613684,0.61046654,0.40126175,0.22292319,0.12003556,0.09602845,0.26750782,0.42183927,0.5418748,0.805953,1.1626302,1.4369972,1.6016173,1.862266,2.651071,2.5481834,2.627064,2.6990852,2.8294096,3.3369887,4.2389703,4.9488945,5.346727,5.6005163,6.1904054,6.375603,6.8797526,7.507367,8.028665,8.186425,7.507367,7.4044795,7.6857057,8.004657,7.888051,7.7680154,7.332458,7.133542,7.1987042,7.0375133,6.64997,6.478491,6.1732574,5.4770513,4.2423997,2.6785078,1.6976458,1.1283343,0.89512235,1.0151579,1.3169615,1.4781522,1.4678634,1.4507155,1.7799559,1.7799559,1.704505,1.4781522,1.1077567,0.66876954,0.45956472,0.4046913,0.4081209,0.432128,0.50757897,0.48700142,0.48357183,0.47671264,0.47328308,0.490431,0.5178677,0.48357183,0.41840968,0.34981793,0.31552204,0.3566771,0.40126175,0.4115505,0.4115505,0.47328308,3.223812,5.1683884,3.9200184,2.2360911,1.3821237,1.1214751,1.0631721,0.77165717,0.6379033,0.66876954,0.48014224,0.21263443,0.13375391,0.14061308,0.14747226,0.09602845,0.12346515,0.09259886,0.072021335,0.072021335,0.048014224,0.36696586,0.59331864,0.59331864,0.45613512,0.48357183,0.5212973,0.607037,0.64476246,0.77508676,1.4027013,1.8931323,1.9068506,1.8554068,1.920569,2.0749004,7.06838,18.674105,28.060884,30.77369,26.76107,21.705858,14.904987,9.06097,5.4839106,4.1155047,4.1120753,5.2987127,6.4819202,7.4799304,9.122703,12.21962,12.507706,11.149589,9.6817255,10.017825,12.47341,18.355152,23.664154,24.518122,17.178804,13.022143,14.856973,16.19794,14.29795,10.151579,10.340206,13.934414,14.321958,10.923236,9.1981535,9.9869585,13.797231,27.025148,45.620373,55.086033,43.915867,34.07981,28.071173,24.778769,19.476627,14.589465,13.46799,11.739478,8.388771,5.785714,5.188966,4.108646,3.059192,2.218943,1.4267083,2.16064,2.369845,2.4418662,3.07634,5.2781353,6.2075534,7.81603,7.5690994,6.142391,7.414768,8.344186,7.39762,5.9640527,4.9248877,4.664239,3.690236,4.273266,5.48734,6.420188,6.2075534,5.103226,4.99005,4.6436615,3.882293,3.57363,3.1620796,3.6593697,4.3795834,5.0174866,5.6245236,5.411889,5.6793966,5.9400454,5.6348124,4.1429415,3.4638834,4.3349986,5.744559,6.601956,5.73427,6.4716315,8.505377,9.551401,8.831187,7.0889573,8.357904,7.56567,7.7097125,8.477941,6.2247014,5.9160385,5.1100855,4.7019644,5.346727,7.4765005,7.8194594,7.473071,8.189855,10.045261,11.410237,6.9620624,7.548522,9.06097,9.438225,8.663138,7.658269,7.058091,7.301592,8.128122,8.591117,7.6342616,6.4819202,6.3618846,7.6342616,9.798331,11.955542,10.844356,7.7748747,4.7362604,4.417309,6.1904054,5.9160385,4.636802,3.3026927,2.7813954,2.6373527,2.6133456,2.7059445,3.4124396,5.751418,7.085528,6.2487082,4.7019644,3.234101,1.9445761,1.6839274,1.6942163,1.7593783,1.8279701,2.037175,2.0714707,2.0474637,1.9102802,1.8073926,2.0989075,1.8999915,1.7147937,1.9925903,2.4247184,1.9480057,1.9754424,1.5776103,1.2449403,1.3821237,2.3046827,1.7216529,1.6393428,1.5638919,1.4267083,1.5604624,1.1797781,1.1523414,1.1454822,1.2209331,1.845118,1.9411465,1.2312219,0.8745448,1.1008976,1.2277923,0.83681935,0.6207553,0.47328308,0.4115505,0.5590228,0.5178677,0.52472687,0.66533995,0.89855194,1.0597426,0.9842916,1.0117283,1.1420527,1.2963841,1.3032433,1.6221949,1.6804979,1.4747226,1.196926,1.2037852,1.0117283,0.96714365,0.94999576,0.89169276,0.77165717,0.58988905,0.8711152,1.1008976,1.0563129,0.7956643,1.2689474,1.1900668,1.138623,1.9068506,4.5099077,4.9660425,3.2958336,2.2223728,2.5138876,2.9494452,1.8999915,1.7730967,1.7730967,1.5981878,1.4541451,1.2792361,1.2655178,1.1249046,0.84367853,0.65848076,0.490431,0.4629943,1.9239986,5.1066556,9.122703,5.411889,3.7211025,3.0283258,2.3321195,0.65162164,4.0503426,10.412228,10.789482,4.9420357,1.3306799,1.7456601,1.371835,1.1180456,1.2758065,1.5021594,2.5173173,5.5593615,8.076678,7.9017696,3.2375305,1.7936742,2.6579304,5.130663,7.191845,5.501058,3.216953,2.170929,2.8054025,4.1463714,3.8102717,4.5442033,3.192946,1.5330256,0.6962063,1.1832076,7.6685576,13.4645605,12.13731,5.130663,1.7593783,2.4212887,1.5433143,0.59331864,0.4629943,1.4541451,1.1180456,0.9431366,0.78537554,0.6276145,0.5555932,5.099797,6.3721733,6.550512,6.4133286,5.3570156,4.822,6.2692857,6.7631464,5.888602,5.7274113,6.5985265,7.970361,10.377932,13.588025,16.602633,16.427725,20.27915,20.824455,17.638369,17.20967,16.527182,16.688372,19.634388,24.03455,25.269201,27.210346,26.514141,26.466127,28.863409,34.018078,32.035778,29.161781,26.548437,24.583282,22.892496,24.487255,23.324625,20.875898,18.519772,17.532051,12.713481,9.3079,7.613684,7.1987042,6.90033,9.078118,9.757176,7.473071,4.671098,7.699424,12.315649,12.754636,10.2236,6.660259,4.729401,2.836269,3.7485392,3.882293,2.4830213,1.6359133,1.9445761,1.6667795,3.3301294,6.9723516,10.14472,6.0532217,4.846007,4.90431,5.1752477,5.1580997,6.8797526,5.3261495,3.093488,2.6236343,6.2144127,6.2692857,3.9680326,4.016047,6.783724,8.327039,7.5725293,6.385892,5.73427,6.118384,7.56224,6.262427,5.4839106,5.120374,5.3330083,6.550512,5.754848,3.5359046,1.8279701,1.2517995,1.138623,0.9294182,0.8848336,0.78537554,0.6173257,0.5796003,0.548734,0.4664239,0.37725464,0.37039545,0.5693115,0.7613684,0.65505123,0.50757897,0.432128,0.38754338,0.4629943,0.69963586,0.9259886,1.0700313,1.138623,2.277246,3.9303071,4.866585,4.7259717,4.016047,3.3232703,2.1400626,1.5227368,1.529596,1.2346514,1.4850113,3.234101,4.201245,3.7313912,2.8054025,3.1346428,4.098357,3.690236,1.9411465,0.922559,2.5550427,4.2286816,4.122364,2.4315774,1.371835,1.2072148,1.430138,1.3992717,1.2723769,2.020027,0.89512235,0.3841138,0.22635277,0.39783216,1.08032,1.9720128,2.1640697,2.5310357,2.7128036,1.1249046,2.294394,5.9160385,9.067829,10.072699,8.471081,9.523964,10.079557,10.816919,11.612583,11.537132,11.070708,11.019264,10.930096,10.329918,8.7317295,8.460793,8.158989,7.407909,6.416758,5.994919,6.7048435,6.121814,6.451054,7.4181976,6.2864337,6.334448,5.086078,3.957744,4.0846386,6.3481665,6.39961,5.086078,3.6147852,2.7299516,2.719663,2.1297739,1.611906,0.823101,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.030866288,0.044584636,0.16119061,0.38754338,0.6379033,0.70649505,0.72707254,0.7442205,0.7407909,0.64819205,0.33952916,0.21263443,0.116605975,0.024007112,0.01371835,0.07545093,0.32924038,0.6927767,1.0151579,1.0940384,0.7476501,0.48014224,0.32581082,0.26750782,0.22978236,0.08916927,0.09259886,0.22978236,0.4115505,0.4629943,0.42869842,0.65162164,0.922559,1.2175035,1.6770682,2.0508933,2.2669573,2.2669573,2.2841053,2.867135,1.8554068,2.3081124,2.9151495,3.3815732,4.437886,3.9543142,3.07634,2.1846473,1.4781522,0.9877212,0.72021335,0.91912943,1.2277923,1.3341095,0.9842916,0.34981793,1.0288762,1.7765263,1.8931323,1.2277923,0.37725464,0.06516216,0.06859175,0.3018037,0.83338976,0.77851635,0.7510797,0.7476501,0.7922347,0.9259886,0.9602845,0.6824879,0.39097297,0.21263443,0.07888051,0.12003556,0.19548649,0.41498008,0.7099246,0.8471081,1.1214751,1.4472859,1.6393428,1.7490896,2.037175,2.5447538,2.6236343,2.8465576,3.4433057,4.297273,4.8494368,5.641671,6.392751,7.0272245,7.675417,8.025234,8.378482,8.549961,8.279024,7.2192817,7.798882,8.56368,9.067829,9.153569,8.947794,8.663138,8.272165,7.7748747,7.407909,7.6445503,6.8591747,6.169828,5.610805,5.0243454,4.0674906,2.6579304,1.9274281,1.4438564,1.08032,1.0254467,1.3752645,1.7182233,2.0165975,2.2635276,2.4898806,2.435007,2.2223728,1.8588364,1.3752645,0.8162418,0.58645946,0.52472687,0.52815646,0.548734,0.59331864,0.48700142,0.4698535,0.4629943,0.4389872,0.4046913,0.4081209,0.3841138,0.33952916,0.29494452,0.28122616,0.31209245,0.37039545,0.38754338,0.3566771,0.33609957,4.400161,6.186976,4.9351764,3.1655092,2.037175,1.371835,1.1832076,1.0837497,1.2003556,1.3238207,0.91227025,0.6173257,0.66876954,0.67219913,0.5453044,0.53844523,0.37039545,0.2709374,0.25721905,0.29494452,0.31209245,0.58645946,0.8265306,0.881404,0.83338976,0.9877212,1.0082988,1.0425946,1.1111864,1.2929544,1.7456601,1.920569,2.0234566,2.1297739,2.2223728,2.1915064,6.7871537,15.536031,20.882757,20.992504,19.768143,16.87014,11.334786,6.5985265,4.122364,3.391862,3.8685746,5.381023,6.5230756,7.366754,9.445084,11.914387,11.434244,10.690024,10.916377,11.924676,15.134769,25.344652,34.535946,36.024387,24.476965,20.96164,19.37031,17.326277,14.472859,12.493987,11.691463,14.112752,13.865822,9.873782,5.871454,6.7048435,12.898679,26.867388,42.609196,45.70954,35.197857,26.047716,21.19485,19.819586,17.333136,14.105893,12.2093315,9.97324,7.0752387,4.540774,3.6593697,3.3026927,3.1620796,2.8054025,1.6976458,1.3924125,1.6976458,2.2120838,3.426158,6.725421,8.261876,8.045813,6.917478,6.3790326,8.587687,8.196714,6.866034,5.675967,5.0346346,4.681387,5.0243454,5.3673043,5.1580997,4.3178506,3.223812,2.9185789,3.3712845,3.426158,3.0454736,3.2855449,3.5359046,4.5853586,5.3741636,5.5147767,5.2781353,5.610805,5.6828265,5.6519604,5.3673043,4.383013,3.9543142,4.7602673,5.744559,6.4098988,6.831738,8.543102,9.647429,9.743458,8.47451,5.5387836,5.288424,5.4839106,8.556821,11.622872,6.451054,7.0752387,7.14726,6.7357097,6.619104,8.299602,8.368194,7.1781263,6.883182,8.450503,11.667457,6.866034,6.1046658,7.1095347,8.337327,8.968371,6.094377,5.888602,6.636252,7.1061053,6.5813785,6.461343,5.284994,4.523626,5.3090014,8.433355,11.832077,10.038403,6.800872,4.3007026,3.1517909,6.0806584,4.9934793,3.4295874,2.8877127,2.860276,3.4535947,3.4295874,2.8808534,2.5619018,3.865145,5.48734,4.6848164,3.450165,2.6750782,2.1400626,1.8691251,1.6942163,1.7388009,1.9274281,1.9891608,1.9411465,1.8176813,1.7799559,1.9068506,2.2086544,1.8691251,1.9171394,2.5173173,3.1449318,2.5824795,2.4247184,1.6393428,1.0014396,0.9534253,1.6084765,1.4541451,1.6359133,1.6770682,1.5158776,1.5227368,1.1454822,1.0871792,1.0185875,0.9877212,1.4129901,1.6599203,1.08032,0.7099246,0.8162418,0.90198153,0.66876954,0.58988905,0.490431,0.36696586,0.4046913,0.4664239,0.5521636,0.70649505,0.881404,0.91912943,0.8848336,0.8711152,1.0014396,1.1763484,1.0940384,1.3375391,1.4541451,1.3478279,1.1283343,1.1077567,1.2072148,1.1763484,1.0014396,0.7956643,0.78537554,0.83681935,1.255229,1.4438564,1.2895249,1.155771,1.7525192,1.920569,1.8897027,2.0817597,3.07634,2.6476414,1.8759843,1.7353712,2.2395205,2.4247184,1.7388009,1.7388009,1.605047,1.2449403,1.2998136,1.6839274,1.5330256,1.3821237,1.3272504,1.039165,0.7510797,0.71678376,2.0165975,4.616225,7.332458,4.4275975,2.9391565,2.0063086,1.1454822,0.26750782,4.9180284,13.365103,13.344524,5.06893,1.2380811,1.9239986,1.5536032,1.155771,1.097468,1.1043272,1.7936742,4.2526884,6.2144127,6.0223556,2.633923,1.5947582,2.9871707,5.363875,6.464772,3.2203827,2.0337453,1.9754424,3.292404,4.695105,3.350707,2.194936,0.8779744,0.4664239,1.0597426,1.7833855,7.2604365,11.845795,11.588576,6.9620624,2.8465576,3.8960114,2.750529,1.1729189,0.28122616,0.5453044,1.6564908,2.534465,2.2120838,1.2243627,1.587899,7.3427467,8.772884,8.035523,6.725421,5.885172,4.8185706,4.9831905,4.9248877,4.2355404,3.542764,3.7725463,4.7534084,6.4544835,9.431366,14.850114,15.189643,19.03421,20.04251,17.504614,16.317978,16.62321,16.983316,19.500635,23.595562,26.03057,27.85854,25.968836,24.408375,25.663603,30.650223,31.864298,31.850578,31.116648,30.056904,28.956007,31.730543,29.665932,26.198618,23.681301,23.386356,16.369421,11.825217,9.801761,9.0644,7.082098,7.7851634,8.567109,7.3290286,5.329579,7.191845,11.201033,12.634601,11.4376745,8.309891,4.7362604,2.9700227,4.671098,4.4721823,2.1057668,2.411,3.2409601,2.428148,3.9131594,8.090397,11.797781,7.490219,5.6656785,5.785714,6.9860697,8.06296,7.81603,5.0586414,2.8877127,3.3644254,7.4936485,6.9552035,3.707384,2.9700227,5.9743414,9.959522,8.440215,7.116394,6.1149545,5.7411294,6.4887795,5.593657,4.232111,3.875434,5.020916,7.174697,7.2947326,4.7328305,2.503599,1.6256244,1.1146159,1.0597426,0.9602845,0.8265306,0.70306545,0.6824879,0.6276145,0.490431,0.33266997,0.26407823,0.45613512,0.6036074,0.58645946,0.53844523,0.52472687,0.53844523,0.66533995,0.7579388,0.91912943,1.0906088,1.0666018,2.633923,5.2781353,6.1904054,5.15467,4.540774,3.882293,2.726522,2.095478,1.9925903,1.4129901,1.08032,2.3835633,3.3198407,3.1072063,2.1503513,3.175798,5.7068334,5.9914894,3.4844608,0.8779744,2.8499873,4.506478,4.48933,2.9288676,1.4575747,1.0597426,0.9945804,1.0185875,1.2998136,2.417859,0.9842916,0.39097297,0.1920569,0.16119061,0.28808534,1.2620882,2.2841053,3.0111778,2.952875,1.4678634,3.0660512,5.950334,8.838047,10.230459,8.423067,8.30646,7.671987,7.56224,8.597976,10.988399,8.539673,8.186425,8.443645,8.457363,8.004657,7.747438,7.641121,7.5416627,7.414768,7.3427467,7.5725293,6.5882373,7.870903,10.343636,8.378482,7.438775,6.591667,5.597087,5.0757895,6.5127864,6.8591747,6.169828,4.698535,3.1552205,2.726522,1.8039631,1.2929544,0.66533995,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.024007112,0.034295876,0.09602845,0.22978236,0.42526886,0.4938606,0.6036074,0.6790583,0.70306545,0.7510797,0.4629943,0.29494452,0.15090185,0.0274367,0.01371835,0.058302987,0.14061308,0.4081209,0.77508676,0.89512235,0.61389613,0.3841138,0.26750782,0.2503599,0.26064864,0.13375391,0.09602845,0.2503599,0.51100856,0.6036074,0.4972902,0.5796003,0.8196714,1.2037852,1.704505,2.1846473,2.7985435,2.884283,2.609916,2.9563043,2.194936,2.4144297,2.9322972,3.4604537,4.0949273,3.724532,2.942586,2.0714707,1.371835,1.0323058,0.77165717,1.3375391,2.1023371,2.3492675,1.2792361,0.42526886,0.6173257,1.3478279,1.8965619,1.3615463,0.4664239,0.12346515,0.05144381,0.25378948,1.0288762,1.039165,0.9431366,0.83338976,0.8128122,0.980862,0.980862,0.71678376,0.4664239,0.30866286,0.10288762,0.12689474,0.216064,0.52472687,0.94656616,1.1043272,1.1008976,1.3615463,1.7079345,1.9308578,1.8005334,2.4144297,2.9391565,3.6113555,4.431027,5.1580997,5.48734,5.878313,6.660259,7.682276,8.31675,8.639131,8.903209,8.951223,8.64599,7.8537555,8.769455,9.606275,10.010965,10.05898,10.261326,10.045261,9.839486,9.318189,8.659708,8.56025,7.6616983,6.691125,5.8543057,5.0757895,3.974892,2.6476414,2.1263442,1.7113642,1.2243627,0.9945804,1.2072148,1.670209,2.1983654,2.644212,2.8980014,2.7230926,2.3904223,1.9239986,1.3821237,0.8505377,0.6379033,0.5727411,0.5590228,0.5521636,0.5693115,0.42869842,0.38754338,0.3841138,0.3841138,0.36353627,0.3566771,0.33266997,0.3018037,0.2709374,0.26407823,0.2503599,0.2777966,0.29494452,0.28465575,0.23664154,5.360445,6.461343,5.295283,3.8342788,2.8019729,1.6667795,0.85739684,1.2792361,1.9411465,2.1126258,1.3272504,1.1797781,1.5055889,1.605047,1.4541451,1.7010754,1.3272504,0.9362774,0.7305021,0.7510797,0.881404,0.88826317,0.9911508,1.1351935,1.3443983,1.7319417,2.0337453,2.0063086,1.9891608,2.095478,2.2223728,2.2360911,2.0920484,2.0097382,2.0680413,2.201795,3.974892,6.5230756,8.7317295,10.419086,12.315649,11.698323,8.635701,5.878313,4.4721823,3.7759757,3.7759757,4.787704,6.077229,7.7371492,10.679735,11.080997,9.695444,10.199594,12.212761,11.283342,17.412016,36.020958,51.481537,52.96312,34.43649,30.002031,23.091412,16.767254,13.368532,14.493437,11.808069,10.984968,10.556271,9.746887,8.433355,9.517105,14.836395,23.184011,31.370436,34.223854,27.68706,21.674994,18.8593,18.684393,17.357141,14.037301,11.509696,9.421077,7.56567,5.8817425,3.4913201,2.74367,2.8911421,3.1106358,2.4967396,2.5824795,2.942586,2.4967396,1.9239986,3.6353626,5.545643,6.6568294,6.807731,6.5127864,6.9620624,4.5784993,4.249259,4.434457,4.2938433,3.6970954,6.7940125,6.6876955,5.206114,3.5976372,2.5310357,1.6427724,1.7971039,2.4315774,3.2786856,4.3521466,5.020916,5.7068334,5.7411294,5.0895076,4.331569,4.5201964,4.7671266,4.9248877,4.945465,4.852866,4.887162,5.411889,5.861165,6.3138704,7.5245147,9.619993,9.325048,7.8194594,6.0154963,4.5510626,3.799983,4.383013,8.580828,12.596875,6.5710897,6.186976,7.8983397,8.937505,8.913498,9.825768,9.458802,7.596536,6.725421,7.3839016,8.158989,6.3721733,4.523626,4.4413157,6.258997,8.388771,5.099797,5.31929,6.018926,5.5559316,3.673088,4.201245,4.033195,3.4947495,3.6285036,6.2075534,9.325048,6.842027,4.804852,5.0414934,5.137522,6.999788,5.645101,4.0057583,3.5359046,4.197815,5.7068334,5.394741,3.9646032,2.5413244,2.668219,3.4776018,3.57363,3.175798,2.8877127,3.7039545,2.4315774,2.2360911,2.49331,2.5790498,1.8554068,1.4781522,1.4472859,1.8176813,2.3286898,2.3972816,2.037175,2.2841053,2.6956558,2.877424,2.5070283,2.095478,1.2758065,0.71678376,0.6241849,0.72021335,1.155771,1.471293,1.5981878,1.5947582,1.6427724,1.6016173,1.5536032,1.2312219,0.86082643,1.1283343,0.922559,0.72707254,0.5796003,0.4972902,0.490431,0.5624523,0.5453044,0.47671264,0.38754338,0.3018037,0.39783216,0.4698535,0.5761707,0.6893471,0.69963586,0.805953,0.7922347,0.8848336,1.0014396,0.72707254,1.0425946,1.1283343,1.2175035,1.3375391,1.3066728,1.4472859,1.6256244,1.5124481,1.1832076,1.1146159,1.313532,1.5776103,1.7353712,1.728512,1.6016173,2.2360911,2.7985435,2.784825,2.2463799,1.8245405,1.9925903,1.9411465,1.9925903,2.0749004,1.7250825,2.2498093,2.3424082,2.0063086,1.5330256,1.5090185,1.862266,1.7765263,1.9651536,2.2909644,1.7662375,1.2826657,0.9877212,0.96714365,1.2106444,1.6187652,2.1194851,1.9754424,1.5124481,0.9602845,0.45270553,3.433017,10.14129,10.220171,3.9508848,2.2395205,2.7539587,1.937717,1.2346514,1.1180456,1.1008976,0.97057325,1.1763484,1.3889829,1.3821237,1.0254467,1.8862731,5.610805,9.541112,10.220171,3.3987212,2.5653315,3.1860867,4.40359,5.0243454,3.525616,1.2449403,0.5555932,1.155771,2.1880767,2.2360911,2.4247184,3.5050385,5.31929,6.1972647,2.9665933,3.8548563,3.2581081,1.7559488,0.29837412,0.18862732,2.7882545,4.341858,3.450165,1.4987297,2.6304936,6.7391396,8.207003,6.914048,4.434457,4.0503426,3.683377,3.1037767,2.8980014,2.7402403,1.3889829,1.3341095,3.923448,6.601956,8.687145,11.372512,14.387119,16.95931,18.180243,17.837284,16.424294,16.081335,16.822126,19.548649,23.5304,26.373528,27.436699,26.208908,24.209457,23.732746,27.84482,31.634514,33.308155,33.356167,32.86231,33.50707,36.7446,36.57998,35.08125,33.109238,30.300406,21.479506,15.6252,13.004995,11.80464,8.114404,7.3187394,7.164408,6.543653,5.7274113,6.368744,7.5588107,8.303031,8.501947,7.64798,4.8494368,4.0674906,5.5079174,4.5030484,1.8313997,3.7039545,5.9400454,4.4927597,4.5784993,7.380472,10.041832,7.6171136,7.1198235,7.6651278,8.371623,8.357904,4.386442,2.1160555,1.9514352,3.309552,4.6127954,3.690236,2.4555845,1.9754424,3.1620796,6.800872,7.6651278,7.2467184,6.121814,5.07236,5.086078,5.284994,3.9131594,3.690236,5.2438393,7.1061053,7.3701835,4.852866,2.6887965,1.8759843,1.2689474,1.2346514,1.0700313,0.94656616,0.8745448,0.6927767,0.7305021,0.5212973,0.26750782,0.15776102,0.36010668,0.4698535,0.5178677,0.58302987,0.6893471,0.8025235,0.8779744,0.85396725,1.1077567,1.5021594,1.3684053,2.6236343,5.9400454,6.7802944,4.962613,4.664239,4.064061,3.4467354,2.6853669,1.8279701,1.08032,1.0494537,2.1091962,3.4364467,3.9200184,2.1640697,2.6750782,5.936616,7.517656,5.861165,2.318401,3.40901,3.9714622,3.6319332,2.620205,1.7902447,1.0323058,0.4629943,0.5144381,1.1317638,1.7902447,1.1043272,0.6344737,0.36010668,0.23321195,0.18176813,0.980862,2.386993,3.3369887,3.2546785,2.054323,3.5599117,5.1752477,7.130112,8.556821,7.48336,6.8111606,4.914599,2.767677,2.2600982,6.169828,4.1360826,4.73969,5.90575,6.495639,6.310441,6.1149545,6.7940125,8.200144,8.718011,5.2747054,6.6122446,6.1321025,6.9792104,9.256456,10.028113,8.549961,8.279024,7.431916,6.258997,7.0272245,6.584808,6.9037595,6.48535,4.6402316,1.5021594,0.71678376,0.23321195,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.01371835,0.0274367,0.0548734,0.10288762,0.18176813,0.32238123,0.53844523,0.6927767,0.7510797,0.78194594,0.53844523,0.28122616,0.10288762,0.0274367,0.020577524,0.14747226,0.24350071,0.36353627,0.48357183,0.4972902,0.29837412,0.17490897,0.14061308,0.16804978,0.19548649,0.16462019,0.09259886,0.2194936,0.52815646,0.75450927,0.764798,0.61389613,0.58645946,0.8196714,1.2826657,1.920569,3.2409601,3.7005248,3.117495,2.6887965,2.6476414,2.5447538,2.7882545,3.1792276,2.9254382,2.4830213,2.054323,1.4472859,0.89512235,1.0528834,1.0048691,1.6427724,2.6956558,3.0660512,0.8162418,0.31209245,0.8711152,1.4335675,1.4507155,0.89169276,0.6241849,0.5178677,0.36696586,0.30523327,0.8025235,1.2209331,1.2037852,1.0563129,0.9431366,0.90884066,0.82996017,0.7099246,0.59331864,0.44927597,0.16804978,0.116605975,0.29837412,0.61046654,0.9774324,1.3546871,1.138623,1.2312219,1.728512,2.287535,2.1400626,2.386993,3.6353626,4.804852,5.422178,5.6210938,5.8645945,5.844017,6.5024977,7.671987,8.086967,8.213862,8.604835,8.999237,9.352485,9.8429165,9.870353,10.062409,10.275044,10.6488695,11.622872,11.760056,11.547421,11.063849,10.38479,9.585697,8.913498,8.069819,7.0032177,5.6999745,4.1635194,2.8945718,2.318401,1.845118,1.3306799,1.0666018,1.0425946,1.4438564,1.920569,2.3321195,2.7573884,2.5447538,2.1263442,1.5947582,1.0700313,0.69963586,0.548734,0.490431,0.45270553,0.41840968,0.42869842,0.33952916,0.274367,0.274367,0.32238123,0.37382504,0.36696586,0.32924038,0.29494452,0.26750782,0.23664154,0.18519773,0.17147937,0.18862732,0.20920484,0.1920569,5.3261495,6.8145905,6.060081,4.6436615,3.2272418,1.5570327,0.8848336,1.7147937,2.5070283,2.486451,1.6324836,1.4369972,1.8828435,2.5481834,3.2272418,3.9200184,3.4810312,2.503599,1.7147937,1.4198492,1.4815818,1.3101025,1.4575747,1.8142518,2.3904223,3.340418,3.9268777,3.8171308,3.391862,2.9665933,2.8088322,3.0283258,2.4144297,1.9308578,1.99602,2.4727325,3.069481,4.0057583,4.6848164,5.113515,5.919468,6.090947,6.142391,6.416758,6.3618846,4.530485,3.799983,4.4687524,6.159539,8.261876,9.932085,8.433355,8.275595,9.877212,12.003556,11.794352,27.84482,57.154076,73.42061,64.64772,33.14353,27.52587,23.835632,20.227707,17.069057,16.921585,12.247057,8.213862,7.4970784,10.717461,16.417435,17.981327,19.178253,19.768143,19.843594,19.805868,18.914175,17.04505,15.933864,15.673215,14.7095,14.123041,11.787492,9.647429,9.006097,10.542552,6.1732574,4.3590055,4.2115335,4.3761535,3.0214665,3.998899,4.0846386,3.0420442,1.704505,1.9994495,2.5721905,2.9803114,3.542764,3.8102717,2.5790498,3.9474552,4.8185706,4.201245,3.1243541,4.6402316,8.838047,7.4970784,5.0277753,3.2992632,1.6633499,2.1503513,2.4761622,2.603057,2.983741,4.547633,5.693115,6.228131,6.461343,6.5882373,6.697984,6.5779486,6.8763227,6.23499,4.98662,5.1580997,5.8645945,6.691125,7.1198235,7.438775,8.759167,9.321619,7.191845,5.254128,4.40359,3.525616,3.8788633,2.8054025,2.7368107,4.3624353,6.6053853,4.2526884,5.446185,7.658269,9.472521,10.621432,10.096705,8.656279,7.64798,7.5725293,8.073249,5.8371577,4.262977,3.8857226,4.996909,7.6445503,5.8988905,4.9214582,4.2938433,3.7108135,2.9906003,4.7979927,5.103226,4.846007,5.206114,7.599966,7.7097125,4.897451,4.3178506,6.992929,9.81205,8.676856,7.130112,5.994919,5.7239814,6.4098988,6.958633,6.5196457,5.1340923,3.4227283,2.5927682,3.6182148,5.103226,5.744559,4.887162,2.534465,1.786815,2.7916842,3.7622573,3.806842,2.9288676,1.6736387,1.6770682,2.2395205,2.6785078,2.3492675,2.4967396,2.3218307,1.8828435,1.3101025,0.8093826,0.7613684,0.89512235,0.9431366,0.9294182,1.1592005,1.4267083,1.3581166,1.2415106,1.2620882,1.4953002,1.6907866,1.4644338,0.9877212,0.5555932,0.5796003,0.97057325,0.9294182,0.66876954,0.4424168,0.5658819,0.48014224,0.31895164,0.22292319,0.22978236,0.29151493,0.37382504,0.37725464,0.37382504,0.39440256,0.4424168,0.4424168,0.59674823,0.78194594,0.8471081,0.64133286,0.6173257,0.66533995,0.7442205,0.85396725,1.039165,0.96371406,1.1763484,1.4678634,1.6393428,1.4815818,1.5055889,1.4472859,1.5330256,1.6016173,1.1146159,1.1008976,1.2998136,1.3924125,1.2380811,0.8848336,0.9328478,1.2209331,1.4541451,1.5913286,1.845118,2.1263442,1.8313997,1.5124481,1.4610043,1.6942163,1.4507155,1.3238207,1.587899,1.9514352,1.5707511,1.1934965,0.9328478,0.9534253,1.3615463,2.2292318,4.1943855,3.8137012,2.435007,1.196926,1.039165,0.85396725,1.7250825,2.3458378,2.9734523,5.4016004,4.5099077,2.2738166,1.1694894,1.6873571,2.335549,1.6873571,1.4267083,1.8759843,2.7711067,3.234101,3.5873485,8.035523,12.912396,13.810948,5.5833683,3.7519686,5.768566,6.773435,4.9523244,1.5124481,0.70649505,0.7510797,2.0440342,3.82399,4.166949,2.1743584,1.0185875,1.2449403,2.3081124,2.5619018,2.8088322,2.5756202,1.5193073,0.32238123,0.70306545,3.1072063,3.5976372,2.2498093,0.64133286,1.862266,4.338428,4.7499785,3.5770597,2.4007113,3.8925817,7.284444,5.0757895,2.726522,1.9857311,0.90198153,0.5212973,3.8137012,7.250148,9.321619,10.528833,12.617453,14.915276,17.648657,19.744135,18.828436,16.338554,18.406595,21.479506,23.640146,24.627867,22.724447,23.60242,23.931662,23.180582,23.61957,30.993181,34.933777,35.804893,35.10869,35.461933,38.023838,38.510838,40.256496,41.371113,34.74515,25.063425,19.109661,14.874121,11.080997,7.1884155,6.7219915,7.191845,6.625963,5.453044,6.5162163,8.944365,9.595985,9.602845,9.108984,7.2775846,6.1046658,4.249259,3.0077481,3.3987212,6.135532,9.294182,6.2487082,4.1017866,5.4153185,8.210432,9.283894,10.347065,11.173596,10.456812,5.844017,3.4638834,3.8479972,5.195825,5.662249,3.357566,3.223812,2.6133456,2.7402403,3.9954693,5.936616,5.3741636,5.1683884,4.619654,3.9165888,4.1360826,5.562791,5.6999745,5.3878818,5.2781353,5.813151,5.56965,3.5770597,1.7147937,0.91569984,1.1592005,1.5261664,1.3169615,1.0666018,0.9259886,0.65505123,0.7407909,0.5144381,0.25378948,0.116605975,0.15090185,0.26407823,0.39097297,0.5727411,0.77851635,0.89855194,0.84024894,0.86082643,1.0871792,1.4267083,1.587899,2.1983654,5.353586,6.992929,6.1286726,4.822,3.4433057,3.7931237,3.2615378,1.7765263,1.8005334,2.6167753,4.105216,6.368744,7.5588107,3.8617156,1.0906088,2.0920484,4.6608095,6.56766,5.552502,3.3815732,2.352697,1.7490896,1.1797781,0.59674823,0.51100856,0.607037,0.9294182,1.0700313,0.16804978,1.0220171,1.1077567,0.8162418,0.45270553,0.24350071,0.72021335,0.9294182,1.9925903,3.7622573,4.835718,5.5319247,6.108095,7.023795,7.8366075,7.2021337,4.773986,3.2409601,2.2326615,1.786815,2.3492675,4.8288593,6.684266,8.210432,8.604835,5.9812007,6.2727156,6.210983,6.39961,6.3001523,4.2115335,8.899779,9.4862385,8.886061,8.1487,6.4407654,9.551401,9.534253,9.112414,9.115844,8.467651,6.4544835,6.2247014,6.591667,5.518206,0.12346515,0.15776102,0.18519773,0.12003556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.037725464,0.061732575,0.058302987,0.044584636,0.06859175,0.14061308,0.32924038,0.52472687,0.42869842,0.18176813,0.06859175,0.024007112,0.020577524,0.044584636,0.22978236,0.34638834,0.34638834,0.22978236,0.044584636,0.034295876,0.020577524,0.041155048,0.08573969,0.12346515,0.1097468,0.07888051,0.12689474,0.38754338,1.0220171,1.4267083,1.039165,0.64476246,0.5727411,0.7339317,1.2826657,2.5447538,3.642222,4.190956,4.2869844,3.4947495,2.8739944,2.452155,2.3904223,2.976882,1.8279701,1.313532,1.039165,0.91912943,1.1763484,1.3341095,1.821111,3.4021509,4.4756117,1.0837497,0.37382504,1.5707511,2.2292318,1.9171394,2.1983654,2.037175,2.0165975,1.3341095,0.31552204,0.4115505,0.94999576,1.1283343,1.1592005,1.1043272,0.8848336,0.7888051,0.5796003,0.45613512,0.40126175,0.16804978,0.106317215,0.18176813,0.37382504,0.6962063,1.2209331,1.3546871,1.1420527,1.3786942,2.0303159,2.2120838,2.6647894,4.280125,5.3398676,5.439326,5.4633327,5.353586,5.8474464,6.914048,8.124693,8.635701,8.440215,8.64942,8.954653,9.294182,9.8429165,10.429376,10.803201,11.046701,11.441104,12.466551,13.087306,12.319078,11.173596,10.377932,10.39165,9.719451,9.129561,8.268735,6.910619,4.945465,3.5290456,2.5790498,1.9754424,1.6187652,1.4335675,1.4472859,1.6976458,2.0268862,2.294394,2.3801336,2.1846473,1.670209,1.1146159,0.6756287,0.3806842,0.37039545,0.32924038,0.28808534,0.26750782,0.30523327,0.30523327,0.2777966,0.29151493,0.33952916,0.34981793,0.3018037,0.2709374,0.26407823,0.26064864,0.19891608,0.15090185,0.16462019,0.19548649,0.216064,0.22978236,5.545643,7.2295704,6.3035817,5.2438393,4.420738,2.0920484,1.2449403,1.5776103,2.2052248,2.568761,2.4247184,1.9754424,2.3081124,3.1586502,4.40359,6.0566516,5.5387836,4.5853586,3.3541365,2.3286898,2.311542,2.2360911,2.3801336,2.7539587,3.275256,3.7691166,4.32471,4.647091,4.307562,3.5187566,3.1243541,3.3541365,3.5770597,3.57363,3.3198407,2.983741,3.6010668,4.170378,4.2766957,3.9097297,3.4673128,4.3590055,5.9914894,6.848886,6.1801167,4.0057583,4.1155047,4.8322887,5.892031,7.0375133,8.018375,7.0615206,8.875772,12.003556,15.028452,16.578627,35.139553,64.243034,76.037384,63.40964,39.978703,35.59226,28.949148,22.53925,17.429163,13.258785,13.975569,12.092726,9.342196,9.122703,16.492886,28.667921,31.771698,28.239223,22.223726,19.600092,21.969936,20.37175,16.681513,12.88496,11.070708,10.593996,9.561689,8.080108,6.6225333,6.001778,4.90431,4.629943,4.3178506,3.457024,1.8862731,2.6579304,2.2566686,2.3835633,3.3232703,3.940596,2.9700227,3.923448,4.8597255,4.945465,4.4447455,5.442755,4.866585,4.314421,4.7259717,6.3961806,6.0566516,5.3741636,4.557922,3.9303071,3.9440255,4.979761,4.650521,3.9474552,3.549623,3.8034124,4.3349986,4.863155,5.7479887,6.4819202,5.672538,5.425607,6.9517736,7.6342616,7.1061053,7.257007,6.540223,6.64997,6.159539,5.2026844,5.48734,7.922347,6.90033,5.6965446,4.9831905,2.8054025,5.4839106,5.137522,5.3913116,7.963502,12.662037,7.1232533,5.5147767,6.6122446,8.1212635,6.701414,7.514226,8.165848,8.06639,7.6857057,8.546532,8.179566,6.4716315,5.9126086,7.0375133,8.4264965,7.548522,5.970912,5.15467,5.254128,5.0895076,5.3330083,4.1943855,3.7622573,5.188966,8.683716,8.666568,5.6656785,4.108646,5.751418,9.6645775,9.078118,7.56224,5.953764,4.681387,3.782835,4.420738,6.0978065,6.135532,4.431027,3.474172,3.6765177,4.2595477,4.945465,5.0140567,3.3026927,4.0229063,5.751418,6.39961,5.885172,6.1286726,4.256118,4.0263357,3.8445675,3.059192,1.9582944,2.1057668,2.0714707,2.1229146,2.1743584,1.7593783,1.3203912,1.2860953,1.255229,1.1592005,1.2449403,1.0940384,1.2277923,1.3443983,1.4575747,1.8725548,1.2792361,1.214074,1.1489118,0.91569984,0.72707254,0.75450927,0.6756287,0.53501564,0.42183927,0.4664239,0.4972902,0.5007198,0.490431,0.47671264,0.44927597,0.5521636,0.5178677,0.4081209,0.30523327,0.29494452,0.2194936,0.23664154,0.4046913,0.66191036,0.83681935,0.8025235,0.6859175,0.607037,0.6379033,0.82996017,0.91227025,1.0906088,1.4472859,1.7216529,1.3101025,1.0597426,1.1763484,1.5193073,1.7216529,1.1763484,1.1523414,1.371835,1.6427724,1.8073926,1.728512,1.6393428,1.5638919,1.6393428,1.8073926,1.8108221,1.5810398,1.3512574,1.3101025,1.3615463,1.0940384,0.96714365,1.2243627,1.6290541,1.786815,1.1454822,1.214074,1.0906088,1.0357354,1.2346514,1.786815,2.2806756,1.8897027,1.7525192,2.0646117,2.1126258,1.646202,1.6770682,1.6187652,1.4335675,1.6187652,1.762808,1.2689474,1.0014396,1.1763484,1.3821237,1.2517995,1.3101025,3.3781435,6.8626046,8.752307,3.9028704,3.1586502,3.8617156,3.8445675,1.4472859,1.1694894,4.149801,5.020916,2.7573884,0.6927767,1.1180456,1.5364552,1.879414,2.469303,4.029765,6.4544835,5.48734,3.666229,2.860276,4.249259,3.457024,2.6304936,1.3992717,0.31552204,0.86082643,3.6765177,6.0703697,6.060081,4.4104495,4.6436615,4.0091877,2.627064,2.0406046,2.74367,4.184097,5.3227196,4.057202,2.8499873,2.3389788,1.3512574,1.4335675,3.7279615,6.3961806,8.539673,10.199594,15.059319,15.889278,16.540901,18.173384,19.267422,19.03421,21.074816,22.875349,23.705309,24.61415,24.147726,23.489244,22.659285,22.155134,22.923363,27.553307,31.929459,33.966633,34.463924,37.07384,39.83123,40.38682,40.63032,40.31823,37.08756,30.17008,26.527859,22.666143,17.508043,12.373952,10.504827,9.129561,8.189855,7.7611566,8.052671,9.97667,13.766364,14.836395,11.921246,7.082098,6.6225333,4.7671266,3.6593697,3.9371665,4.7191124,6.2692857,5.4633327,5.127233,6.111525,7.3050213,8.820899,9.386781,9.386781,8.1041155,3.7313912,3.100347,3.6147852,4.479041,4.7362604,3.2581081,2.1194851,4.0194764,4.2869844,2.767677,3.8102717,4.2183924,3.4707425,2.8534167,3.1277838,4.5510626,8.244728,6.2384195,4.139512,4.2081037,5.3501563,4.5682106,3.1586502,1.6530612,0.5521636,0.31895164,1.0151579,1.2380811,1.0323058,0.7339317,0.97400284,0.764798,0.34981793,0.09602845,0.09259886,0.12689474,0.16119061,0.29151493,0.7682276,1.2998136,1.0597426,0.96714365,1.3546871,1.9274281,2.2669573,1.8313997,1.9445761,6.4304767,8.971801,7.610255,4.7602673,3.5359046,3.391862,2.8877127,2.5207467,4.7431192,3.666229,3.3815732,4.619654,6.4133286,6.0806584,2.6373527,1.6324836,2.4144297,3.6559403,3.3438478,2.9185789,2.6956558,2.3492675,1.7147937,0.764798,0.37725464,0.274367,0.36353627,0.51100856,0.5453044,0.97057325,0.7442205,0.72021335,0.9842916,0.85396725,0.9774324,0.6241849,1.4198492,3.391862,4.9831905,7.8091707,8.361334,8.210432,7.9086285,6.9826403,4.856296,3.882293,3.4364467,3.3644254,3.9851806,7.517656,7.1987042,7.099246,8.491658,9.849775,8.64942,7.596536,6.142391,4.7671266,4.9934793,17.473747,28.112328,27.964857,17.189093,5.0586414,5.456474,7.682276,8.64256,8.611694,11.228469,9.163857,4.513337,1.7696671,1.8108221,1.8931323,2.054323,1.5364552,0.70649505,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.010288762,0.0274367,0.041155048,0.05144381,0.06859175,0.0548734,0.058302987,0.08916927,0.13032432,0.1097468,0.05144381,0.017147938,0.020577524,0.072021335,0.20577525,0.30866286,0.30523327,0.22292319,0.11317638,0.058302987,0.09602845,0.072021335,0.09259886,0.16119061,0.20920484,0.09602845,0.08573969,0.16462019,0.34638834,0.66876954,1.0425946,1.039165,0.8711152,0.72707254,0.7682276,0.9294182,1.4267083,1.9754424,2.386993,2.603057,2.5138876,2.5070283,2.301253,1.9068506,1.6324836,1.2277923,0.84024894,0.6379033,0.5761707,0.39440256,0.4629943,0.8711152,2.3767042,3.8445675,2.2669573,1.0906088,0.9774324,1.2449403,1.5124481,1.6976458,1.5776103,1.6324836,1.1729189,0.33609957,0.082310095,0.53158605,0.823101,0.89169276,0.864256,1.0563129,0.99801,0.823101,0.6790583,0.61046654,0.53501564,0.4046913,0.32581082,0.31209245,0.44927597,0.8676856,1.2175035,1.3341095,1.5810398,2.1400626,3.0043187,3.5359046,4.15323,4.5647807,4.822,5.305572,5.3501563,5.7891436,6.4133286,7.051232,7.56224,7.15069,7.891481,8.779744,9.294182,9.414218,10.2921915,12.017275,13.22106,13.807519,14.932424,14.647768,14.105893,13.697772,13.423406,12.867812,11.094715,9.767465,8.567109,7.1987042,5.4187484,3.7794054,2.9117198,2.4830213,2.2360911,1.99602,1.8416885,1.903421,1.99602,1.9994495,1.879414,1.6256244,1.4267083,1.1832076,0.8779744,0.5761707,0.47671264,0.39440256,0.32581082,0.28808534,0.30523327,0.33609957,0.29837412,0.2777966,0.29151493,0.3018037,0.29151493,0.30866286,0.28808534,0.22292319,0.16119061,0.14061308,0.16462019,0.18519773,0.19548649,0.22978236,5.3330083,10.460241,7.531374,4.616225,4.0674906,2.5310357,2.1229146,2.0817597,2.2292318,2.4315774,2.6167753,2.6064866,2.8328393,3.8891523,5.8543057,8.296172,8.176137,6.9071894,4.955754,3.1586502,2.719663,2.6990852,3.069481,3.5461934,3.9303071,4.105216,4.389872,4.5682106,4.3452873,3.9680326,4.2115335,4.180667,4.2286816,4.32128,4.3624353,4.1943855,4.6608095,4.955754,4.619654,3.7313912,2.9082901,5.0655007,6.615674,6.64997,5.4667625,4.5613513,5.597087,6.694555,8.049242,9.427936,10.1481495,8.735159,10.127572,13.361672,16.925014,18.746124,39.68033,63.978954,71.836136,61.26615,48.13083,38.795494,25.77335,16.510035,12.902108,11.255906,13.71492,16.53404,16.05733,14.023583,17.573206,30.410152,39.025276,36.25074,25.416672,20.344313,21.098822,19.78872,16.729528,12.977559,10.336777,9.033533,8.05953,7.010077,5.7651367,4.465323,3.474172,2.8911421,2.270387,1.4815818,0.72364295,1.0631721,0.89855194,1.1043272,1.8108221,2.411,2.7333813,6.121814,7.2364297,5.425607,4.722542,4.2389703,3.875434,4.863155,6.0737996,3.998899,4.6436615,4.3795834,3.6285036,3.2032347,4.297273,5.020916,5.689686,5.720552,5.07236,4.2389703,4.513337,5.4153185,6.6396813,7.3084507,5.9571934,6.166398,7.5519514,7.7577267,6.680836,6.492209,6.118384,6.293293,6.4236174,6.1972647,5.5833683,6.8043017,6.4819202,5.751418,5.0106273,3.9165888,10.792912,10.350495,9.270175,10.398509,12.758065,7.864044,6.725421,8.663138,10.371073,5.90575,6.7459984,7.8606143,7.8023114,6.9552035,7.548522,8.371623,7.1952744,6.584808,7.1541195,7.5759587,7.284444,6.711703,6.81802,7.682276,8.498518,8.872343,7.2535777,5.501058,5.06893,7.016936,7.085528,5.703404,5.7102633,7.932636,11.204462,8.81747,8.193284,7.720001,6.5642304,4.6573796,5.7479887,7.689135,7.671987,6.1732574,6.9346256,6.077229,4.9180284,4.671098,5.0620713,4.307562,5.936616,8.344186,9.613133,9.47595,9.325048,7.130112,7.0752387,5.919468,3.5839188,3.1620796,2.6133456,2.1846473,2.2258022,2.5721905,2.5481834,1.9582944,1.7730967,1.6839274,1.5193073,1.2380811,1.0700313,1.0837497,1.2243627,1.3546871,1.255229,1.0528834,1.1660597,1.2792361,1.2243627,0.97400284,0.823101,0.6756287,0.5727411,0.53501564,0.5418748,0.42183927,0.39783216,0.41498008,0.4938606,0.71678376,0.6893471,0.6344737,0.52815646,0.42526886,0.45270553,0.35324752,0.32238123,0.5007198,0.85396725,1.1592005,1.1077567,0.8676856,0.64819205,0.6036074,0.8162418,0.96714365,1.0220171,1.2209331,1.4953002,1.4575747,0.97400284,1.1489118,1.4815818,1.5741806,1.1454822,0.96714365,1.2003556,1.6221949,1.99602,2.0577524,1.8245405,1.903421,1.9891608,1.9754424,1.9754424,1.7319417,1.2346514,0.9259886,0.91227025,0.9568549,1.0906088,1.4678634,1.605047,1.3272504,0.77165717,0.99801,1.605047,1.9685832,1.8519772,1.4129901,1.4335675,1.2312219,1.3169615,1.646202,1.6221949,1.4061309,1.2723769,1.0597426,0.77851635,0.6344737,0.9431366,1.2106444,1.8519772,2.8122618,3.5702004,3.0351849,2.2223728,2.9082901,5.147811,7.239859,2.4555845,1.0597426,1.08032,1.2175035,0.83338976,0.7442205,1.8416885,2.2463799,1.7319417,1.7250825,2.1263442,1.8554068,1.4747226,1.5124481,2.4418662,4.8768735,4.2835546,2.585909,1.4232788,2.1503513,1.6290541,1.1866373,0.6241849,0.20234565,0.6241849,4.2252517,6.3378778,6.324159,5.113515,5.2026844,3.4433057,1.9685832,2.5138876,4.1326528,3.1963756,3.6010668,3.6387923,3.1072063,2.1572106,1.3169615,1.529596,3.6868064,7.1541195,10.515115,11.592006,13.4474125,14.332246,15.700651,17.514904,18.235117,19.888178,21.966507,22.306036,21.705858,23.952238,24.672453,23.382927,22.292318,22.491234,23.969387,26.380386,28.84969,30.276398,31.469894,35.139553,38.74748,38.915527,38.48683,38.538273,38.40795,35.10869,32.24155,27.309805,20.430052,14.339106,12.79922,10.590566,9.050681,8.663138,9.033533,9.458802,11.077567,12.600305,12.9638405,11.365653,8.337327,5.521636,4.386442,4.8837323,5.425607,5.284994,4.8117113,4.341858,4.3658648,5.5250654,6.025785,6.4579134,6.728851,5.9914894,2.6167753,2.4144297,2.9494452,4.081209,5.0586414,4.506478,2.5721905,4.7842746,5.586798,3.9543142,3.3815732,3.457024,2.411,1.9308578,2.8225505,5.020916,6.591667,4.856296,3.0626216,2.5893385,2.952875,2.0749004,1.4404267,0.9534253,0.5693115,0.31895164,0.59331864,0.8162418,0.7442205,0.65848076,1.3443983,0.8162418,0.32924038,0.11317638,0.17833854,0.28808534,0.6790583,0.53844523,0.7990939,1.4438564,1.5021594,1.1249046,1.0940384,1.2998136,1.6324836,1.9925903,2.1400626,4.619654,6.3481665,6.094377,4.4721823,3.3747141,3.841138,3.974892,3.7313912,4.928317,4.623084,4.108646,4.331569,5.65539,7.874333,5.658819,4.746549,4.57507,4.506478,3.8342788,3.5839188,3.5393343,2.8122618,1.6736387,1.5604624,0.58302987,0.33952916,0.30523327,0.35324752,0.7682276,0.5590228,0.490431,0.72021335,0.980862,0.5761707,0.5761707,0.85739684,1.3546871,2.1812177,3.6387923,5.919468,7.0786686,7.390761,6.9689217,5.7925735,3.4707425,4.482471,5.0312047,4.479041,5.3090014,7.5245147,6.090947,5.9297566,8.604835,12.291641,10.988399,9.657719,8.001227,7.4696417,11.249047,27.056015,42.372555,41.004147,23.43094,6.800872,5.24041,6.210983,7.222711,7.407909,7.5519514,4.523626,2.136633,1.6256244,2.5447538,2.784825,1.9239986,1.3169615,0.6379033,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.010288762,0.01371835,0.01371835,0.01371835,0.024007112,0.048014224,0.048014224,0.037725464,0.030866288,0.030866288,0.041155048,0.048014224,0.041155048,0.041155048,0.07888051,0.216064,0.25721905,0.22292319,0.15776102,0.08916927,0.041155048,0.048014224,0.034295876,0.041155048,0.07545093,0.09945804,0.07545093,0.1097468,0.1920569,0.29494452,0.37039545,0.50757897,0.6790583,0.72364295,0.64476246,0.6036074,0.6859175,0.89169276,1.0906088,1.2072148,1.1934965,1.2277923,1.529596,1.7696671,1.6907866,1.1214751,1.1900668,0.8265306,0.5555932,0.44927597,0.13375391,0.16804978,0.6893471,2.3732746,4.249259,3.690236,1.9411465,1.5227368,1.6427724,1.7490896,1.5261664,1.5536032,1.2826657,0.78537554,0.25378948,0.0,0.17147937,0.6001778,0.881404,0.9294182,0.9877212,1.0631721,0.91569984,0.77851635,0.71678376,0.64476246,0.59331864,0.5796003,0.58302987,0.6756287,1.0082988,0.88826317,1.1043272,1.4850113,1.9925903,2.6922262,3.1826572,3.9954693,4.4687524,4.5339146,4.715683,5.5250654,6.4064693,6.999788,7.3084507,7.706283,7.658269,8.258447,9.132992,9.692014,9.132992,9.777754,11.931535,13.176475,13.200482,13.790371,13.841815,14.376831,15.0250225,15.3302555,14.750656,12.860953,10.991828,9.246168,7.699424,6.39961,4.9660425,3.8342788,3.1517909,2.7779658,2.311542,1.8965619,1.762808,1.7250825,1.6667795,1.5261664,1.3958421,1.1832076,0.90884066,0.64133286,0.4972902,0.44927597,0.37725464,0.3018037,0.2503599,0.2777966,0.2777966,0.25378948,0.22635277,0.20920484,0.19891608,0.21263443,0.24007112,0.22978236,0.18862732,0.17833854,0.14747226,0.16462019,0.18176813,0.18862732,0.20920484,6.2692857,12.157887,9.445084,6.200694,5.1238036,3.5564823,3.216953,3.292404,3.216953,2.959734,3.0248961,3.4433057,3.5804894,4.2115335,5.675967,7.874333,8.525954,7.846896,6.2555676,4.4687524,3.4810312,3.2958336,3.549623,3.8171308,3.9028704,3.8171308,4.15323,4.4447455,4.3487167,4.1189346,4.6093655,4.8117113,5.3432975,6.001778,6.557371,6.7322803,6.989499,6.550512,5.3330083,4.0434837,4.1943855,6.0086374,6.1561093,5.40503,4.65395,4.9420357,6.1321025,7.9292064,9.877212,11.38623,11.72233,10.021255,9.97667,12.586586,17.689812,23.952238,46.282284,61.307304,62.205856,51.88623,42.976162,35.300743,23.890507,15.8138275,12.768354,11.084427,14.448852,20.920483,22.494663,19.586374,20.995934,28.321533,36.696587,35.17728,24.967398,19.421753,17.71039,16.317978,14.4145565,11.859513,9.194724,7.56567,6.7357097,6.5710897,6.2384195,4.197815,2.644212,1.6736387,0.9431366,0.37725464,0.17490897,0.48357183,0.59674823,0.5727411,0.5658819,0.823101,2.435007,6.6122446,7.414768,4.7431192,4.3624353,2.7230926,3.9165888,5.7479887,5.970912,2.294394,3.4981792,3.4055803,3.4638834,4.2526884,5.48734,5.439326,6.6396813,7.3118806,6.715132,5.1409516,5.007198,6.025785,7.2158523,7.579388,6.108095,6.3138704,6.9963584,6.725421,5.717122,5.813151,6.1492505,6.3893213,6.835168,7.250148,6.848886,6.7802944,6.1492505,5.0174866,4.1326528,4.9214582,10.744898,11.852654,11.063849,10.100135,9.589127,7.5759587,8.186425,10.525404,11.646879,6.5813785,6.715132,7.531374,7.6274023,7.1061053,7.5931067,7.332458,6.111525,5.470192,5.693115,5.8062916,6.018926,6.23156,6.677407,7.534804,8.944365,9.640571,8.687145,6.7322803,5.0312047,5.470192,6.334448,6.252138,7.3050213,9.729739,11.948683,8.546532,8.042382,8.285883,8.467651,9.112414,10.021255,9.208443,7.5553813,6.3824625,7.4524937,6.697984,5.0483527,4.6265135,5.5079174,5.720552,8.875772,10.844356,11.458252,10.964391,10.034973,9.239308,9.712592,7.966932,4.4996185,3.7794054,2.719663,2.3492675,2.3561265,2.4144297,2.170929,1.8005334,1.6599203,1.6187652,1.5673214,1.4095604,1.4850113,1.2346514,1.1489118,1.2003556,0.83338976,0.881404,1.0014396,1.138623,1.1934965,1.0117283,0.8848336,0.7305021,0.6824879,0.7373613,0.7613684,0.59674823,0.5144381,0.50757897,0.64476246,1.0700313,0.805953,0.64819205,0.5007198,0.3806842,0.42183927,0.37725464,0.4664239,0.67219913,0.9294182,1.1214751,0.94999576,0.7305021,0.5761707,0.61389613,0.97400284,0.9328478,0.90884066,0.9294182,1.0597426,1.371835,1.0768905,1.2758065,1.4953002,1.4438564,1.0357354,0.9431366,1.2449403,1.5638919,1.7662375,1.9342873,1.9925903,2.0165975,1.8588364,1.611906,1.6084765,1.3752645,0.9774324,0.823101,0.9431366,1.0048691,1.1180456,1.3478279,1.2929544,0.939707,0.66191036,0.8196714,1.8073926,2.4315774,2.1915064,1.3101025,1.4472859,1.3203912,1.1626302,1.1008976,1.1489118,1.3169615,1.2346514,0.94656616,0.6790583,0.84367853,1.2998136,1.4987297,2.0097382,3.0146074,4.307562,3.3678548,2.2463799,1.821111,2.386993,3.6627994,1.5707511,1.3958421,2.4144297,3.2581081,1.920569,1.2277923,0.8711152,1.6221949,3.1243541,3.9097297,2.3972816,1.9754424,2.1400626,2.270387,1.6427724,2.1091962,2.0028791,1.3066728,0.48357183,0.48014224,0.32238123,0.26750782,0.19548649,0.19548649,0.5453044,3.2581081,4.0229063,3.724532,3.2203827,3.3541365,3.0111778,3.350707,4.763697,5.885172,3.6147852,2.9974594,3.7211025,4.2526884,3.99204,3.2649672,2.7882545,3.9954693,7.3255987,11.519984,13.622321,13.7938,12.63117,12.936404,15.069608,16.976458,19.03764,21.181131,21.301168,20.738716,24.257473,25.300066,23.290329,21.969936,22.53239,23.640146,23.904224,25.6053,27.470995,29.326403,32.07693,35.623123,36.669147,37.293335,38.692604,41.17563,40.277077,37.142433,31.113218,23.540688,17.79613,17.069057,13.869251,11.303921,10.515115,10.669447,8.961512,7.822889,9.89436,14.174485,16.047039,9.674867,5.3741636,4.0949273,4.897451,4.931747,5.2506986,6.574519,6.2658563,4.5442033,4.4927597,4.537344,4.3007026,4.7019644,4.8905916,2.2463799,1.8485477,2.6922262,4.1017866,5.1340923,4.5819287,2.6990852,4.506478,5.518206,4.602506,3.9851806,3.275256,2.5138876,2.4555845,3.532475,5.885172,4.8905916,3.4844608,2.5481834,2.510458,3.3438478,1.9857311,1.1592005,1.1454822,1.5021594,1.08032,0.9259886,0.77508676,0.7099246,0.823101,1.2312219,0.6756287,0.2777966,0.16119061,0.274367,0.39097297,0.939707,0.805953,1.0288762,1.7388009,2.153781,1.4267083,1.1214751,1.1592005,1.4095604,1.704505,1.7971039,2.4830213,3.7313912,4.914599,4.8185706,3.7211025,4.5682106,5.0174866,4.48933,4.1463714,5.593657,5.5559316,4.746549,4.6779575,7.6616983,7.1095347,5.9640527,4.835718,4.1155047,3.981751,3.5118976,3.316411,2.469303,1.3203912,1.4815818,0.6756287,0.3806842,0.490431,0.7613684,0.8128122,0.64133286,0.5590228,0.65848076,0.7407909,0.30866286,0.26407823,1.1111864,1.4644338,1.4918705,2.8980014,4.1772375,5.6245236,7.2707253,8.117833,6.121814,4.098357,5.65539,6.9689217,6.8866115,6.9346256,5.662249,3.7553983,4.3041325,7.3564653,9.918367,9.551401,9.132992,8.831187,9.8429165,14.373401,27.227495,38.191887,35.33161,20.495214,9.328478,8.64599,6.3893213,5.1992545,5.1066556,3.5599117,1.4129901,1.5844694,2.7470996,3.6010668,2.8637056,1.7696671,1.4815818,0.94999576,0.1371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.024007112,0.030866288,0.030866288,0.034295876,0.037725464,0.044584636,0.061732575,0.058302987,0.048014224,0.05144381,0.13032432,0.1371835,0.11317638,0.08573969,0.058302987,0.017147938,0.01371835,0.020577524,0.020577524,0.020577524,0.034295876,0.058302987,0.106317215,0.1920569,0.2709374,0.23664154,0.18862732,0.31209245,0.39440256,0.37725464,0.35324752,0.51100856,0.6790583,0.7339317,0.64476246,0.45956472,0.42526886,0.6859175,1.1111864,1.4232788,1.1763484,1.1111864,0.823101,0.66533995,0.6036074,0.19548649,0.106317215,0.6173257,2.1297739,3.9200184,4.1292233,3.0900583,3.2409601,3.192946,2.5207467,1.7936742,1.4918705,0.97400284,0.48357183,0.15090185,0.0,0.0,0.3018037,0.6824879,0.9362774,0.8711152,1.0597426,0.9945804,0.84367853,0.72364295,0.71678376,0.7682276,0.78194594,0.78537554,0.8711152,1.1763484,1.1180456,1.3032433,1.546744,1.8348293,2.318401,2.8019729,3.415869,4.029765,4.4447455,4.4104495,5.4976287,6.5127864,7.1849856,7.490219,7.6514096,7.798882,7.7714453,8.519095,9.609704,9.23245,10.072699,11.499407,12.175035,11.965831,11.97269,11.852654,13.173045,14.784951,15.724659,15.2033615,12.946692,11.303921,9.877212,8.457363,7.010077,6.001778,4.602506,3.5118976,2.884283,2.3149714,1.9102802,1.670209,1.4953002,1.3443983,1.2312219,1.155771,0.97400284,0.72364295,0.48700142,0.4115505,0.3841138,0.33952916,0.2777966,0.22292319,0.22978236,0.20577525,0.21263443,0.19548649,0.15776102,0.1371835,0.16804978,0.19891608,0.22292319,0.22978236,0.22978236,0.17833854,0.20234565,0.22635277,0.22292319,0.20577525,8.433355,11.393089,10.542552,8.793462,7.1952744,4.928317,4.2286816,4.448175,4.3658648,3.789694,3.5393343,4.0194764,4.098357,3.9646032,4.15323,5.535354,7.006647,7.56567,7.1095347,5.960623,4.870014,4.290414,3.9371665,3.7519686,3.6525106,3.5050385,3.9371665,4.5030484,4.4927597,4.07435,4.2869844,5.1512403,6.8043017,8.210432,8.930646,9.122703,9.174147,7.864044,6.025785,4.9351764,6.310441,5.926327,4.6127954,4.0674906,4.557922,4.897451,5.2506986,7.3393173,9.671436,11.190743,11.2593355,10.14129,9.89436,12.812939,20.484926,33.781437,53.076294,57.572483,51.745617,40.729782,30.34156,30.146074,25.752771,21.524092,19.514353,19.480057,23.739605,27.241213,26.10945,22.415783,24.18888,25.351511,27.625326,26.088871,20.810738,16.852993,13.540011,11.657167,10.216741,8.64942,6.807731,5.6176643,5.288424,6.1286726,6.8591747,4.616225,2.5756202,1.7182233,1.3032433,0.9431366,0.58302987,0.97057325,1.1077567,1.0254467,0.8196714,0.67219913,2.6476414,5.4187484,5.874883,4.2423997,4.0674906,2.2806756,4.911169,6.4133286,5.1169443,3.2306714,3.3884325,3.981751,5.3981705,6.9517736,6.8900414,6.464772,7.281014,7.8983397,7.4936485,5.8680243,5.206114,5.895461,6.7357097,6.790583,5.3913116,5.212973,5.305572,5.1169443,4.8768735,5.5902276,6.276145,6.711703,7.006647,7.2707253,7.630832,7.449064,6.23499,4.2218223,2.843128,4.698535,5.579939,8.419638,9.136421,7.377043,6.5470824,7.164408,8.354475,9.575408,9.73317,7.157549,6.927767,7.332458,7.7851634,8.14527,8.690575,6.475061,4.705394,3.974892,4.098357,4.1120753,4.6093655,4.928317,5.0929375,5.5593615,7.2158523,7.881192,7.98408,7.164408,5.960623,5.809721,7.3598948,7.671987,8.635701,10.528833,12.037852,9.194724,7.9737906,7.8194594,9.091836,13.056439,13.152468,9.033533,5.8234396,5.1100855,4.9248877,5.9983487,5.751418,5.638242,6.1972647,7.034084,10.861504,11.441104,10.566559,9.3593445,8.2653055,9.544542,10.2236,8.371623,4.804852,3.0660512,2.2429502,2.2909644,2.3424082,1.961724,1.1454822,1.1729189,1.2209331,1.2689474,1.371835,1.6427724,1.9274281,1.5021594,1.1660597,1.1283343,1.0014396,0.8093826,0.764798,0.805953,0.8505377,0.77851635,0.8162418,0.764798,0.7990939,0.9294182,0.980862,0.94999576,0.89169276,0.8505377,0.91569984,1.2346514,0.84024894,0.58645946,0.37382504,0.20577525,0.1920569,0.20920484,0.4424168,0.65848076,0.7613684,0.78537554,0.4629943,0.34981793,0.36353627,0.53844523,1.0014396,0.7888051,0.8025235,0.7407909,0.65505123,0.94656616,1.08032,1.2860953,1.3992717,1.3066728,0.9362774,1.0700313,1.4095604,1.471293,1.3101025,1.5021594,2.0028791,1.7490896,1.2517995,0.864256,0.78537554,0.548734,0.6276145,0.9911508,1.3238207,1.0425946,0.8745448,0.85396725,0.83338976,0.77508676,0.7510797,0.77165717,1.4541451,1.9274281,1.8245405,1.313532,1.6359133,1.5261664,1.255229,1.0837497,1.2586586,1.6084765,1.546744,1.1729189,0.8711152,1.3101025,1.8965619,1.6873571,1.3443983,1.471293,2.5893385,1.7936742,1.3684053,1.1832076,1.1489118,1.196926,1.5913286,2.3904223,4.15323,5.40503,2.6407824,1.5021594,1.5673214,3.4638834,5.8165803,5.24041,1.7319417,2.201795,3.4981792,3.6319332,1.7593783,0.91569984,1.4987297,1.6324836,1.0082988,0.8711152,1.0837497,1.1489118,0.88826317,0.5178677,0.64476246,1.196926,0.78194594,0.50757897,0.7099246,0.94999576,3.0729103,5.7308407,7.346176,7.1884155,5.3844523,3.340418,3.5359046,4.7602673,5.7994323,5.446185,4.7362604,5.456474,8.272165,13.128461,19.28457,20.419764,14.009865,9.938945,11.513125,15.443433,16.952452,19.404606,20.742146,21.486366,24.723896,25.838512,23.869928,22.384918,22.20315,21.400625,20.234566,22.480946,25.485264,27.738503,28.883986,31.528198,34.25815,37.060123,40.170757,44.094208,43.590057,39.947834,33.952915,27.639046,24.302057,23.585274,19.45262,15.810398,13.96185,12.624311,9.294182,7.366754,9.654288,15.021593,18.37916,10.868362,6.15268,4.98662,5.627953,3.8514268,5.926327,9.294182,9.424506,6.262427,4.2355404,4.5510626,3.4398763,3.6525106,4.6882463,2.8054025,2.1194851,4.0194764,6.433906,7.431916,5.2164025,2.726522,4.122364,5.6039457,5.8165803,5.8337283,4.616225,4.4687524,4.6779575,5.103226,6.200694,4.619654,3.2855449,3.2855449,4.671098,6.464772,4.266407,2.4452958,2.136633,2.843128,2.4212887,1.8999915,1.2449403,0.9842916,1.0357354,0.7339317,0.4389872,0.24007112,0.2777966,0.45270553,0.42183927,0.8848336,1.1008976,1.4164196,1.8999915,2.3595562,1.5913286,1.4953002,1.7216529,1.7936742,1.1214751,1.0082988,1.4987297,3.0077481,4.8940215,5.439326,4.2835546,5.096367,5.586798,5.007198,4.139512,6.632822,7.4353456,6.2727156,4.681387,5.994919,6.138962,4.5510626,3.1072063,2.7573884,3.532475,2.9974594,2.49331,1.8691251,1.2792361,1.1420527,0.7613684,0.4938606,0.77851635,1.2312219,0.64476246,1.0048691,0.8848336,0.84024894,0.90541106,0.61046654,0.7339317,1.8313997,2.3732746,2.4247184,3.642222,4.105216,5.192395,8.217292,11.238758,9.057541,7.630832,7.7371492,8.940934,10.103564,9.386781,4.8597255,2.8877127,3.865145,6.2144127,6.3721733,7.058091,7.720001,8.999237,10.964391,13.114742,19.37031,21.356041,17.576635,11.149589,9.822338,10.738038,6.2898636,3.0660512,2.8396983,2.5584722,2.5653315,3.1072063,3.5804894,3.5873485,2.9151495,2.435007,2.3972816,1.6084765,0.274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.0034295875,0.006859175,0.01371835,0.017147938,0.0274367,0.030866288,0.024007112,0.017147938,0.020577524,0.024007112,0.030866288,0.041155048,0.041155048,0.041155048,0.041155048,0.030866288,0.017147938,0.030866288,0.030866288,0.024007112,0.017147938,0.01371835,0.0034295875,0.020577524,0.041155048,0.048014224,0.044584636,0.06516216,0.0548734,0.09602845,0.18176813,0.25721905,0.22978236,0.14747226,0.12003556,0.11317638,0.11317638,0.14747226,0.34295875,0.5212973,0.5624523,0.45270553,0.3018037,0.22978236,0.26750782,0.5521636,0.9911508,1.2620882,0.88826317,0.69963586,0.7133542,0.72364295,0.28465575,0.09259886,0.52815646,1.605047,2.877424,3.4364467,3.9851806,4.962613,4.695105,3.2409601,2.393852,1.5330256,0.8848336,0.4046913,0.08916927,0.0,0.0,0.058302987,0.3841138,0.7990939,0.7339317,0.96714365,1.1249046,1.0631721,0.8676856,0.86082643,0.91569984,0.8711152,0.8676856,0.9877212,1.2620882,1.6942163,1.9068506,1.9445761,1.99602,2.4007113,3.0214665,2.9254382,3.4364467,4.48933,4.605936,5.24041,5.861165,6.427047,6.824879,6.8557453,7.3290286,7.0375133,7.6274023,9.0644,9.633711,10.755186,11.132441,11.533703,11.965831,11.670886,10.943813,12.13731,14.150477,15.693792,15.278812,12.133881,10.97468,10.353925,9.249598,7.06838,6.3721733,4.8768735,3.5530527,2.767677,2.2978237,1.978872,1.6873571,1.3821237,1.1146159,1.0357354,0.8848336,0.805953,0.6893471,0.53158605,0.39440256,0.33609957,0.31895164,0.29151493,0.24007112,0.20577525,0.17833854,0.20234565,0.1920569,0.14061308,0.12346515,0.15433143,0.1920569,0.24007112,0.2709374,0.2503599,0.21263443,0.24007112,0.25721905,0.2469303,0.216064,10.422516,10.628291,8.107545,6.5710897,6.5642304,5.4770513,4.866585,3.9646032,3.433017,3.333559,3.1140654,3.309552,3.3747141,3.350707,3.74168,5.5250654,7.3187394,8.021805,7.4936485,6.4819202,6.6533995,5.6142344,4.448175,4.0949273,4.554492,4.8837323,4.3692946,4.32471,4.2698364,4.214963,4.65395,5.703404,7.4044795,8.30646,8.131552,7.7680154,7.6445503,6.526505,6.310441,7.116394,7.2638664,4.5030484,3.841138,4.99005,6.385892,5.2026844,4.1429415,4.6436615,6.7871537,9.462232,10.39165,10.964391,14.887839,21.69557,31.644804,45.74384,51.481537,50.517822,48.23715,45.07507,36.528538,35.25959,26.665043,22.12427,28.818823,49.742737,53.697052,40.112453,26.953129,21.565247,20.659836,22.271742,21.712719,19.747564,17.267973,15.289101,10.63858,8.203573,6.7631464,5.662249,4.8082814,3.9268777,3.673088,4.280125,5.446185,6.3001523,2.836269,1.9857311,2.4315774,2.867135,1.9994495,1.3512574,1.3546871,1.5433143,1.6359133,1.5261664,3.9303071,5.521636,6.831738,7.1061053,4.2869844,3.309552,4.6127954,5.871454,6.135532,5.844017,6.9654922,10.285333,10.8958,7.915488,4.4859004,5.377593,6.121814,6.451054,6.307011,5.844017,5.1100855,5.295283,5.6656785,5.442755,3.7691166,4.0366244,4.2046742,3.9474552,3.4913201,3.6010668,4.249259,6.0566516,7.2295704,7.2432885,6.852316,7.205563,7.191845,5.219832,2.4795918,2.9288676,4.835718,4.2115335,3.5153272,4.396731,7.706283,7.3255987,5.007198,3.8720043,4.73969,6.118384,7.4627824,7.7611566,7.9875093,8.361334,8.361334,7.7268605,6.2864337,5.346727,4.931747,3.782835,3.8685746,4.496189,5.3673043,6.691125,9.170717,9.853205,9.712592,9.547972,9.424506,8.666568,8.64256,9.441654,11.008976,12.891819,14.2362175,11.979549,10.690024,9.678296,8.745448,8.210432,7.8674736,5.9880595,4.7602673,4.705394,4.6676683,9.002667,11.249047,9.668007,6.327589,7.0958166,6.608815,6.2384195,6.138962,6.3001523,6.5299344,7.0203657,6.3001523,4.400161,2.2600982,1.7250825,2.1023371,1.7765263,1.6667795,1.8416885,1.5090185,1.6084765,1.7147937,1.6736387,1.5090185,1.4335675,1.4472859,1.2380811,1.097468,1.1489118,1.3443983,1.0734608,0.8711152,0.6859175,0.53501564,0.47328308,0.65505123,0.8025235,0.88826317,0.91912943,0.9294182,0.980862,1.1008976,1.1077567,0.9431366,0.6859175,0.61389613,0.58645946,0.4938606,0.33952916,0.22978236,0.16804978,0.19891608,0.34981793,0.5761707,0.7476501,0.5041494,0.34981793,0.28465575,0.28122616,0.30523327,0.65848076,0.8676856,0.85396725,0.6790583,0.5178677,0.5555932,0.7305021,0.8093826,0.8162418,1.0220171,0.91227025,1.0494537,1.1180456,1.039165,0.9774324,1.0871792,1.0117283,0.7990939,0.5418748,0.3806842,0.5144381,0.7682276,0.94656616,0.9842916,0.94656616,0.7373613,0.6859175,0.7305021,0.77508676,0.70306545,0.7510797,0.71678376,0.77851635,0.90884066,0.8848336,0.8471081,1.0940384,1.4987297,1.7730967,1.4815818,1.5638919,1.4575747,1.2209331,1.1489118,1.786815,1.5913286,1.4507155,1.3101025,1.1489118,0.9774324,1.0631721,1.4404267,1.7936742,1.8176813,1.2209331,0.90198153,0.84367853,1.0323058,1.1763484,0.6859175,0.61389613,2.5619018,5.23698,6.3001523,2.3972816,1.0666018,2.8465576,3.5016088,2.0508933,0.7922347,2.1469216,3.8617156,3.8479972,2.4487255,2.411,4.0091877,4.3452873,3.2409601,1.3992717,0.4115505,0.38754338,0.29837412,0.4938606,1.0700313,1.8759843,4.0023284,6.444195,7.610255,7.0923867,5.675967,3.4192986,1.6633499,0.7956643,0.9294182,1.8931323,4.4550343,9.373062,14.887839,22.237446,35.626556,35.945507,22.504953,12.312219,10.88894,12.267634,14.441993,17.933313,20.845032,22.230585,22.11055,24.905664,26.445549,25.787067,23.022821,19.288,19.178253,20.155685,21.431492,22.902784,25.162884,27.724785,30.334702,34.3336,39.100727,42.067318,40.46913,37.214455,33.25671,30.60221,32.286137,29.419,26.02028,22.210009,17.947031,13.015285,10.525404,10.131001,10.731179,12.507706,16.938732,13.958421,12.655178,12.555719,11.7257595,6.742569,7.939495,7.764586,6.334448,4.3692946,3.1723683,2.843128,2.194936,2.7916842,4.389872,4.928317,4.245829,8.457363,14.79524,18.410025,12.404818,4.9831905,5.90232,10.021255,12.744347,10.010965,9.191295,9.115844,8.491658,6.6876955,3.724532,4.4550343,4.6745276,6.262427,8.378482,7.4765005,4.938606,2.8122618,2.201795,3.0317552,4.0434837,2.6167753,1.762808,1.1763484,0.7613684,0.6241849,0.5144381,0.48014224,0.6927767,0.9328478,0.5796003,1.2895249,1.786815,1.5227368,0.8196714,0.8711152,0.9294182,1.2929544,1.471293,1.2895249,0.90198153,0.97400284,2.0440342,3.350707,4.3521466,4.729401,3.6936657,5.055212,6.341307,6.6396813,6.591667,7.740579,9.911508,10.47396,8.652849,5.5559316,4.0880685,4.537344,5.5387836,5.98463,5.020916,4.506478,3.57363,2.760818,2.534465,3.2649672,1.5193073,1.313532,1.1420527,0.5693115,0.22978236,0.37382504,1.1180456,2.0063086,2.452155,1.7079345,2.6236343,4.4447455,5.6656785,5.830299,5.5250654,4.413879,4.822,8.22758,12.977559,14.280802,12.377381,10.7757635,10.39165,11.375941,13.121602,10.168727,8.477941,8.31332,9.678296,12.329367,12.682614,12.075578,12.38767,13.557159,13.581166,16.667795,17.514904,13.697772,7.3221693,4.99005,1.903421,0.77165717,1.4507155,3.2649672,5.0346346,4.547633,4.7259717,4.4413157,3.8548563,4.4413157,3.5976372,2.8465576,1.4987297,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.010288762,0.010288762,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0274367,0.041155048,0.034295876,0.017147938,0.030866288,0.041155048,0.0274367,0.01371835,0.01371835,0.01371835,0.01371835,0.024007112,0.024007112,0.017147938,0.030866288,0.030866288,0.030866288,0.024007112,0.01371835,0.01371835,0.0034295875,0.010288762,0.01371835,0.0274367,0.07545093,0.07545093,0.15090185,0.17833854,0.15433143,0.16804978,0.14404267,0.15433143,0.16119061,0.14747226,0.12346515,0.12346515,0.15090185,0.15433143,0.13032432,0.106317215,0.09602845,0.1097468,0.26407823,0.490431,0.5658819,0.89512235,0.64819205,0.31209245,0.11317638,0.01371835,0.08916927,0.82996017,1.9891608,2.9117198,2.534465,3.3747141,4.3007026,3.9886103,2.843128,2.9906003,2.452155,1.4027013,0.53158605,0.1097468,0.0,0.0,0.28465575,0.59674823,0.7099246,0.4424168,0.6756287,1.3101025,1.7319417,1.6427724,1.0666018,0.89855194,0.89855194,1.1249046,1.4335675,1.4953002,1.4575747,2.0097382,2.5824795,2.8911421,2.9151495,3.9165888,3.9268777,4.105216,4.6916757,5.020916,5.06893,5.1169443,5.1238036,5.206114,5.645101,7.915488,9.2153015,9.314759,8.97523,9.962952,9.80519,10.690024,12.624311,14.55174,14.342535,14.476289,14.527733,15.830976,17.79613,17.929884,14.071597,12.044711,10.89237,9.595985,7.0786686,6.138962,4.722542,3.6936657,3.2375305,2.884283,1.9685832,1.529596,1.2723769,1.0940384,1.0837497,0.8745448,0.64133286,0.51100856,0.4664239,0.31895164,0.31895164,0.34638834,0.35324752,0.32581082,0.29151493,0.25378948,0.216064,0.16119061,0.09945804,0.07545093,0.07545093,0.08573969,0.09602845,0.116605975,0.15090185,0.16462019,0.15776102,0.13375391,0.13032432,0.22978236,8.663138,9.280463,8.124693,7.390761,7.4524937,6.8454566,6.1286726,5.6005163,5.0106273,4.530485,4.7602673,4.6436615,4.633373,4.7191124,5.7308407,9.318189,13.125031,12.936404,10.388221,7.366754,6.0052075,4.7842746,4.5510626,4.746549,4.870014,4.5167665,4.7842746,5.0003386,5.0346346,5.147811,5.994919,6.694555,8.158989,8.556821,7.9909387,8.522525,7.81603,7.2364297,7.239859,7.3564653,6.2144127,4.431027,5.06893,5.754848,5.4324665,4.3349986,4.3007026,5.703404,9.5205345,14.476289,17.055338,15.148488,17.662374,26.143745,40.177616,57.404434,56.159496,55.21293,54.660767,50.438942,34.35761,28.907993,42.427425,69.106186,94.60517,96.06618,61.35189,36.507957,26.157463,26.215767,23.907654,19.843594,16.726099,14.205351,12.253916,11.163307,7.8606143,6.1492505,5.305572,4.955754,5.086078,3.6799474,3.117495,3.3850029,4.7088237,7.548522,3.4947495,1.8416885,1.8656956,2.5756202,2.6956558,3.923448,5.579939,5.164959,3.7931237,6.200694,6.0566516,5.2301207,4.307562,7.3873315,22.096832,20.21056,11.773774,6.560801,6.334448,4.8322887,5.1340923,9.434795,11.945253,9.80862,3.1072063,4.2698364,5.1580997,5.7651367,5.9571934,5.453044,4.3007026,4.32128,5.6005163,7.051232,6.392751,6.1732574,5.9983487,5.0826488,3.758828,3.4776018,3.82399,4.5613513,4.9420357,5.0483527,5.7891436,6.708273,7.857185,7.2878733,5.545643,5.662249,4.3761535,3.666229,3.9886103,5.761707,9.352485,7.8023114,6.8969,7.4353456,9.054111,10.206452,8.961512,10.034973,10.906088,10.38479,8.604835,6.7802944,5.4599032,5.5113473,6.307011,5.7239814,5.878313,6.9037595,7.6342616,8.076678,9.403929,9.997248,9.301042,8.824328,8.707723,7.7268605,9.314759,10.861504,11.019264,10.374502,11.454823,10.436234,9.544542,8.549961,7.548522,6.9654922,6.728851,6.108095,4.9523244,3.7759757,3.7279615,5.5319247,6.8557453,6.4064693,5.1580997,6.327589,5.2438393,4.8837323,5.0757895,5.4016004,5.223262,4.8254294,5.3398676,4.6573796,3.069481,3.275256,3.5153272,2.5481834,2.0268862,2.2669573,2.2292318,1.879414,1.9480057,1.8999915,1.6016173,1.3238207,1.2380811,1.1111864,1.2929544,1.529596,0.96371406,0.91227025,0.90541106,0.8025235,0.7133542,1.0220171,1.0288762,1.1043272,1.1146159,1.0220171,0.8711152,0.8505377,0.9568549,1.0151579,0.9877212,0.96714365,1.1180456,0.91227025,0.58645946,0.30866286,0.18176813,0.17833854,0.15776102,0.17833854,0.24007112,0.28465575,0.24350071,0.26064864,0.29494452,0.33609957,0.39097297,0.490431,0.5453044,0.64133286,0.7373613,0.66533995,0.59331864,0.65505123,0.7373613,0.90884066,1.3889829,1.1626302,0.9774324,0.980862,1.1214751,1.1489118,0.85739684,0.8093826,0.77165717,0.65848076,0.52815646,0.7888051,1.0597426,1.0906088,0.8848336,0.70306545,0.805953,0.7305021,0.764798,0.9568549,1.1180456,0.94999576,0.75450927,0.71678376,0.8471081,0.97057325,1.0425946,1.5433143,1.9171394,1.8519772,1.2860953,1.4095604,1.2758065,1.5536032,2.311542,3.0043187,1.5398848,1.0906088,1.1934965,1.488441,1.7079345,1.5604624,1.3958421,1.2175035,1.0220171,0.7922347,0.7888051,0.7990939,1.0117283,1.3203912,1.3101025,0.7579388,1.0940384,1.6976458,1.879414,0.881404,2.277246,6.5642304,6.6636887,2.7985435,2.4898806,6.667118,7.795452,5.7377,2.2463799,0.97057325,1.6427724,2.061182,1.9137098,1.2517995,0.4972902,0.4046913,1.0528834,2.767677,4.389872,3.2821152,2.0646117,2.860276,3.882293,4.0709205,3.1243541,1.5124481,0.83338976,1.2106444,2.668219,5.127233,7.250148,12.504276,18.773561,25.708187,34.714283,34.875473,25.471546,16.53404,12.528283,12.3533745,13.138749,14.342535,15.635489,16.890718,18.20425,23.547548,25.564144,25.351511,24.007113,22.655855,23.122278,23.11199,23.087982,23.238884,23.465237,23.959099,26.246634,30.200947,34.728004,37.773476,38.593147,35.811752,30.732533,25.313786,22.155134,24.874798,25.51956,22.830763,17.641798,12.905538,17.895588,17.549198,15.182784,13.63261,15.241087,12.456262,10.456812,9.89093,10.319629,10.2236,8.471081,7.2638664,6.790583,7.205563,8.618553,9.499957,11.523414,10.573419,6.550512,3.3678548,7.281014,14.63062,17.95046,14.658057,7.0718093,3.340418,5.693115,10.021255,12.466551,9.448513,5.15467,3.4981792,3.0351849,3.1895163,4.249259,4.57164,5.857735,8.570539,11.105004,9.818909,6.677407,7.4524937,8.56025,8.31675,6.948344,5.079219,4.2595477,4.07435,3.8548563,2.6750782,1.1111864,0.65162164,0.64133286,0.72364295,0.8471081,1.5673214,1.8965619,1.6359133,1.1317638,1.2963841,1.5536032,1.1660597,0.9877212,1.3855534,2.2566686,1.879414,3.1963756,4.2698364,4.2526884,3.4124396,3.8685746,5.0312047,5.9400454,6.186976,5.9331865,7.500508,8.261876,8.80718,9.14328,8.680285,7.2432885,6.307011,5.360445,4.3109913,3.4947495,4.3795834,4.0366244,3.316411,2.7333813,2.4590142,1.9754424,2.0577524,1.6770682,1.0597426,1.704505,1.196926,1.3821237,1.2620882,0.97057325,1.7696671,3.8274195,6.2075534,6.831738,5.909179,5.926327,6.142391,7.2878733,10.131001,13.570878,14.623761,11.362224,8.834618,7.301592,7.0443726,8.351046,8.501947,6.2692857,4.979761,7.0306544,13.87954,12.610593,9.952662,10.491108,14.147048,16.143068,19.339443,18.842154,15.782962,11.530273,7.675417,4.7019644,3.100347,2.9082901,3.7451096,4.791134,4.3521466,4.6848164,4.4241676,3.4638834,2.9254382,1.2655178,0.64476246,0.31209245,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.006859175,0.01371835,0.017147938,0.0274367,0.0274367,0.017147938,0.030866288,0.034295876,0.024007112,0.01371835,0.01371835,0.01371835,0.024007112,0.020577524,0.017147938,0.017147938,0.017147938,0.006859175,0.006859175,0.0034295875,0.006859175,0.01371835,0.01371835,0.01371835,0.020577524,0.034295876,0.06516216,0.082310095,0.18519773,0.23321195,0.18862732,0.09602845,0.07888051,0.116605975,0.12346515,0.08916927,0.08573969,0.07545093,0.09945804,0.11317638,0.09602845,0.082310095,0.061732575,0.072021335,0.15090185,0.30523327,0.5144381,0.65848076,0.6824879,0.5418748,0.3018037,0.12346515,0.15090185,0.5212973,0.9328478,1.2449403,1.4815818,2.3629858,3.3266997,3.415869,2.8088322,2.8088322,2.750529,2.3904223,1.488441,0.3841138,0.0,0.0,0.26064864,0.7339317,1.0185875,0.37039545,0.58302987,1.0425946,1.2312219,1.0837497,1.0185875,0.9842916,1.0734608,1.2620882,1.3752645,1.1043272,1.2243627,1.5330256,2.1434922,2.7813954,2.8156912,2.7059445,2.5790498,2.6853669,3.234101,4.386442,4.149801,4.187526,4.400161,4.822,5.6210938,7.1884155,8.47451,9.239308,9.5205345,9.623423,10.878652,13.063298,15.055889,16.180794,16.187653,15.87213,16.13278,17.833855,20.550089,22.580404,19.356592,16.396858,13.745787,11.331357,8.971801,7.8674736,5.720552,3.9063,3.0146074,2.8465576,2.194936,1.6907866,1.3032433,1.0597426,1.0597426,1.0185875,0.85396725,0.71678376,0.6207553,0.45613512,0.3566771,0.32238123,0.32581082,0.32581082,0.29151493,0.23321195,0.1920569,0.15776102,0.12003556,0.07545093,0.08573969,0.082310095,0.07888051,0.08916927,0.116605975,0.1097468,0.09602845,0.07888051,0.058302987,0.058302987,8.361334,9.578837,10.264755,10.076128,9.006097,7.39762,6.8591747,6.1801167,5.501058,5.0655007,5.219832,5.1409516,4.5510626,3.9508848,4.3590055,7.3221693,10.449953,10.100135,7.9943686,5.8234396,5.212973,5.312431,5.394741,5.562791,5.7822843,5.8817425,6.7185616,7.596536,7.857185,7.7371492,8.375052,9.026674,9.595985,9.5033865,9.026674,9.270175,7.455923,6.9346256,7.332458,7.5210853,5.6039457,5.98463,7.8263187,8.251588,7.349606,8.155559,8.954653,8.742019,10.696883,15.470869,21.19485,29.419,32.443897,37.272755,47.019646,60.895756,57.93259,57.665085,58.217247,54.52701,38.34622,43.055042,64.20874,83.904854,89.09039,71.57206,44.677235,28.198069,23.022821,24.881657,24.3535,23.280039,17.04162,12.260776,10.64201,8.968371,6.0978065,4.4104495,4.6127954,5.844017,5.6793966,3.3952916,2.719663,3.0729103,4.214963,6.276145,3.8034124,2.1880767,1.704505,2.0508933,2.3389788,3.7279615,6.478491,7.716572,7.5759587,9.208443,6.8043017,5.576509,3.8034124,4.307562,14.455711,13.708061,10.127572,7.9429245,7.7542973,6.5642304,5.9228973,7.1198235,7.449064,5.751418,2.4041407,3.5118976,4.1189346,4.4584637,4.5819287,4.338428,3.9097297,4.149801,5.147811,6.310441,6.355026,6.142391,5.7754254,4.791134,3.649081,3.724532,3.799983,4.307562,4.787704,5.2026844,5.888602,7.0478024,7.740579,8.865483,9.465661,6.7048435,5.5902276,5.3707337,6.090947,7.682276,9.966381,8.539673,8.193284,8.484799,9.030104,9.489669,7.9292064,8.700864,8.453933,7.082098,7.723431,8.659708,7.431916,6.293293,6.0875177,6.245279,6.584808,6.992929,7.455923,7.953213,8.471081,7.64798,6.948344,7.5725293,8.611694,7.051232,8.9100685,10.120712,11.032983,11.790922,12.339656,11.537132,10.1481495,8.327039,6.5470824,5.5833683,5.336438,5.24041,4.5682106,3.8925817,5.0586414,6.715132,6.5127864,5.2644167,4.396731,5.960623,5.209543,4.537344,4.338428,4.4104495,3.9474552,3.2272418,3.7553983,3.6216443,2.7985435,3.1312134,3.450165,2.901431,2.4418662,2.4761622,2.8877127,2.1229146,2.1126258,2.0817597,1.7388009,1.2792361,1.3649758,1.2003556,1.1283343,1.1283343,0.823101,0.91912943,0.9602845,0.88826317,0.8162418,1.0597426,0.91227025,0.864256,0.86082643,0.8676856,0.864256,0.7613684,0.8505377,0.9602845,0.9877212,0.90198153,0.9842916,0.77851635,0.5007198,0.28808534,0.21263443,0.16804978,0.24007112,0.26407823,0.1920569,0.09602845,0.13032432,0.20234565,0.26750782,0.30866286,0.33952916,0.31552204,0.29837412,0.34638834,0.44584638,0.490431,0.5761707,0.61046654,0.66533995,0.7888051,0.9842916,0.83338976,0.7613684,0.881404,1.1043272,1.1454822,0.75450927,0.7339317,0.7990939,0.764798,0.5555932,0.7888051,0.9294182,0.9328478,0.89169276,1.0151579,1.0460242,0.8265306,0.84367853,1.2243627,1.7147937,1.3546871,1.1043272,1.0151579,1.0494537,1.0837497,0.8505377,1.1900668,1.6599203,1.8485477,1.371835,1.2963841,1.08032,1.4198492,2.1983654,2.4967396,1.313532,0.9328478,0.9911508,1.2243627,1.4541451,1.5810398,1.5536032,1.313532,0.9842916,0.88826317,0.9602845,0.8745448,0.99801,1.2620882,1.1454822,0.78194594,0.6310441,0.66533995,0.77851635,0.7888051,3.1483612,7.0443726,6.684266,2.5824795,1.587899,3.8685746,4.57507,3.4707425,1.4644338,0.61046654,0.61046654,0.7476501,0.7990939,0.65162164,0.29837412,0.3566771,1.2380811,2.74367,3.7759757,2.3595562,1.5913286,2.6853669,3.474172,3.216953,2.6167753,1.5364552,1.2037852,2.1915064,4.0023284,5.0757895,6.5333643,10.247607,14.79867,20.2037,27.930561,34.138115,27.656193,18.355152,12.116733,10.837497,12.579727,12.902108,12.843805,13.38911,15.443433,20.742146,25.207468,25.828222,23.93852,25.20061,23.986534,23.492674,23.36578,22.511812,19.102802,19.819586,24.6896,29.384705,32.296425,34.556522,36.363914,34.607967,30.797695,26.445549,23.057117,22.059107,22.350622,20.563807,16.695232,14.13333,20.231136,20.923914,18.416885,15.45715,15.319967,11.214751,10.175586,10.525404,10.590566,8.704293,10.155008,9.647429,10.155008,11.588576,10.792912,9.678296,11.626302,13.358243,12.250486,6.334448,12.1921835,17.785841,18.759844,14.606613,8.656279,6.018926,6.4716315,7.64798,7.8777623,6.2041235,4.98662,4.2698364,3.7965534,3.799983,4.9934793,7.8126,9.458802,10.906088,11.7086115,9.9869585,8.491658,10.734609,13.224489,13.848674,11.866373,9.098696,7.2535777,6.5710897,6.3618846,5.0106273,2.6133456,1.3341095,0.8711152,0.9911508,1.5193073,1.8965619,2.1091962,2.095478,2.0131679,2.2463799,1.99602,1.2003556,1.0871792,1.7730967,2.2463799,2.3732746,3.3747141,3.690236,3.1449318,2.935727,2.5653315,3.2889743,4.3041325,5.312431,6.5367937,7.8949103,7.613684,7.5690994,8.3922,9.4862385,7.9120584,6.2830043,5.0929375,4.465323,4.139512,4.338428,3.940596,4.1360826,4.6779575,3.8617156,3.7108135,3.2272418,2.8088322,2.6133456,2.5619018,2.0440342,2.5961976,2.9220085,2.8980014,3.5702004,6.111525,7.7714453,8.340756,8.330468,8.985519,12.212761,14.5243025,15.343974,14.623761,12.860953,8.460793,5.936616,4.6916757,4.9351764,7.6685576,7.082098,4.57507,3.117495,4.3281393,8.498518,8.820899,10.048691,11.718901,13.176475,13.581166,15.954441,15.906426,14.208781,11.626302,8.951223,4.616225,3.1620796,4.040054,5.7068334,5.5902276,4.773986,4.266407,3.765687,2.8945718,1.2106444,0.6241849,0.2777966,0.15090185,0.13032432,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.006859175,0.01371835,0.01371835,0.010288762,0.0,0.006859175,0.01371835,0.024007112,0.020577524,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.017147938,0.017147938,0.01371835,0.01371835,0.006859175,0.006859175,0.0034295875,0.0034295875,0.006859175,0.006859175,0.01371835,0.01371835,0.030866288,0.061732575,0.06859175,0.09602845,0.16804978,0.19548649,0.14747226,0.07545093,0.09259886,0.082310095,0.06516216,0.048014224,0.048014224,0.044584636,0.058302987,0.07545093,0.082310095,0.08573969,0.06859175,0.072021335,0.1097468,0.1920569,0.31895164,0.37382504,0.4115505,0.35324752,0.274367,0.40126175,0.764798,0.58645946,0.41840968,0.59331864,1.2106444,2.2498093,2.8534167,2.8019729,2.435007,2.6613598,2.1812177,2.3321195,1.99602,1.0220171,0.20920484,0.041155048,0.10288762,0.4389872,0.77508676,0.50757897,0.59674823,0.91569984,1.0768905,1.1111864,1.4747226,1.4610043,1.4232788,1.3272504,1.155771,0.88826317,1.1797781,1.4575747,1.9411465,2.5138876,2.7093742,2.627064,2.5241764,2.435007,2.6819375,3.9063,3.9954693,3.9303071,4.3109913,5.267846,6.468202,6.9654922,7.953213,9.283894,10.662587,11.633161,12.929544,14.3974085,15.854982,17.158226,18.231688,16.976458,17.151367,18.6158,20.505503,21.19828,18.608942,16.204802,14.222499,12.490558,10.443094,8.64942,6.3310184,4.413879,3.3232703,2.976882,2.4761622,2.1194851,1.7079345,1.313532,1.2998136,1.3375391,1.1111864,0.91912943,0.805953,0.5624523,0.38754338,0.31552204,0.29151493,0.274367,0.24350071,0.18176813,0.14747226,0.12689474,0.11317638,0.09602845,0.106317215,0.106317215,0.10288762,0.10288762,0.106317215,0.08573969,0.06859175,0.044584636,0.024007112,0.01371835,9.208443,9.925226,10.690024,10.388221,8.875772,6.989499,7.431916,7.39762,7.0546613,6.5196457,5.8405876,5.40503,4.5030484,3.6079261,3.2958336,4.232111,5.552502,5.2266912,4.420738,4.2869844,5.9640527,8.186425,8.844906,8.021805,6.7391396,6.941485,8.303031,11.122152,12.648318,12.325937,11.784062,12.30193,12.079007,11.22161,10.069269,9.1810055,7.0958166,7.1987042,8.042382,8.282454,6.6705475,8.652849,10.158438,9.547972,8.182996,10.439664,10.261326,9.578837,11.252477,17.391438,29.360699,67.823524,81.20577,77.72817,70.32026,76.62727,75.37891,82.694214,87.45791,80.56787,54.921413,56.69794,67.40854,69.61377,58.52591,42.00559,28.5959,19.05136,15.817257,17.556059,19.133669,22.673002,16.414005,11.036412,9.637141,7.723431,5.161529,3.3541365,3.5873485,5.0003386,4.5853586,2.901431,2.8499873,3.4124396,3.9783216,4.3521466,4.2046742,4.190956,3.2821152,2.1332035,3.0866287,4.770556,8.018375,9.091836,7.932636,8.1487,6.2247014,5.1992545,4.4413157,4.2218223,5.6965446,5.6073756,6.9209075,7.407909,6.5539417,5.576509,5.24041,4.633373,3.875434,3.2649672,3.2581081,4.0949273,4.0846386,4.2698364,5.0106273,5.994919,5.079219,5.003768,5.874883,6.9552035,6.6225333,5.9812007,5.411889,4.4756117,3.6696587,4.400161,5.528495,7.98065,9.1810055,8.152129,5.5113473,6.9860697,6.944915,7.8126,8.738589,5.610805,5.8817425,6.9654922,7.6857057,7.8846216,8.440215,7.599966,7.2295704,6.725421,6.1492505,6.2247014,6.660259,6.958633,6.416758,6.138962,9.012956,10.816919,9.369633,7.2947326,6.1046658,6.1904054,6.917478,7.414768,7.8331776,8.196714,8.385342,7.7885933,7.2467184,7.7131424,8.937505,9.438225,8.776315,8.525954,9.510246,11.375941,12.566009,12.617453,11.358793,8.707723,5.6828265,4.4104495,5.768566,5.9400454,5.1238036,4.290414,5.188966,7.116394,6.495639,5.751418,5.8165803,6.142391,5.2609873,4.588788,4.232111,4.0057583,3.433017,2.5996273,2.8705647,2.8054025,2.318401,2.6785078,3.5633414,3.4776018,2.935727,2.6476414,3.4913201,2.5893385,2.1160555,1.7971039,1.488441,1.1763484,1.2689474,1.2346514,1.0528834,0.83338976,0.82996017,0.9294182,0.97400284,0.94656616,0.89169276,0.9259886,0.77165717,0.64133286,0.66533995,0.8162418,0.89855194,0.72364295,0.7682276,0.86082643,0.8848336,0.77851635,0.7579388,0.64133286,0.53844523,0.45613512,0.32238123,0.19548649,0.22292319,0.23664154,0.16462019,0.058302987,0.09602845,0.14747226,0.1920569,0.22635277,0.25378948,0.2503599,0.23321195,0.216064,0.216064,0.25378948,0.4698535,0.53158605,0.58988905,0.6790583,0.7407909,0.52472687,0.6173257,0.7579388,0.7956643,0.7099246,0.5590228,0.6893471,0.8471081,0.84367853,0.5624523,0.7579388,0.77508676,0.7476501,0.8196714,1.1694894,1.0597426,0.83338976,0.8779744,1.313532,1.9720128,1.3889829,1.1077567,1.08032,1.1523414,1.0666018,0.8196714,0.96371406,1.2483698,1.4095604,1.196926,1.196926,1.1214751,1.3272504,1.7388009,1.862266,1.1934965,0.9568549,0.90198153,0.91227025,0.9877212,1.3341095,1.5124481,1.4369972,1.2415106,1.2895249,1.4267083,1.2277923,1.1797781,1.2620882,0.9568549,0.7442205,0.6379033,0.8745448,1.2586586,1.1660597,2.6579304,4.431027,3.9646032,1.6221949,0.64133286,0.96714365,1.4438564,1.4987297,1.0768905,0.65162164,0.48357183,0.45956472,0.42869842,0.36010668,0.33609957,0.37039545,1.3238207,2.0303159,2.0920484,1.8828435,3.7794054,5.429037,5.086078,3.2306714,2.5619018,1.8965619,2.287535,3.391862,4.3109913,3.5804894,4.1326528,6.1321025,9.078118,13.591455,21.417774,33.6614,30.159792,20.457489,12.079007,10.563129,12.809509,13.488567,12.373952,10.868362,12.000127,15.861842,20.61182,22.144846,21.568676,25.224615,23.671013,22.666143,22.26831,21.28402,17.254255,18.708399,24.53184,28.170631,28.537598,30.039757,31.950037,31.205816,29.75167,27.947708,24.562706,19.504065,18.807858,18.650097,17.350283,15.361122,18.656956,19.579515,18.187103,15.529172,13.629181,10.6317215,13.660047,16.678083,16.023033,10.412228,12.662037,12.926115,12.943263,13.066729,12.257345,8.663138,11.993267,17.226818,19.085653,12.065289,15.217079,17.909306,15.728088,9.753747,6.5710897,5.528495,5.302142,5.079219,4.8254294,5.271276,7.6033955,8.505377,7.881192,6.5813785,6.40304,11.790922,14.692352,15.172495,14.068168,12.987847,12.147599,14.0750265,16.352274,17.151367,15.22051,12.607163,10.823778,9.774324,8.882631,7.0923867,5.0449233,2.8911421,1.4815818,1.1934965,1.903421,2.784825,2.49331,2.8054025,3.4947495,2.3424082,1.937717,1.4095604,1.5193073,2.0508933,1.8005334,2.7299516,2.726522,2.3046827,1.9651536,2.201795,1.7147937,2.1812177,3.2032347,4.6608095,6.701414,6.835168,6.5024977,6.5470824,7.3598948,8.920357,7.795452,6.619104,5.895461,5.689686,5.6519604,5.586798,4.979761,5.1066556,5.7719955,5.31929,4.715683,3.9508848,3.2443898,2.9254382,3.426158,3.4227283,4.249259,4.979761,5.336438,5.6999745,7.3084507,8.694004,9.156999,8.958082,9.321619,13.629181,16.47231,16.266533,13.759505,12.041282,9.3764925,7.5519514,6.711703,7.082098,8.988949,7.363324,4.9008803,3.9200184,5.2026844,7.9875093,8.251588,9.849775,10.9198065,10.902658,10.521975,12.260776,13.029003,12.2093315,9.880642,6.8454566,3.74168,3.0248961,4.170378,5.90232,6.183546,5.802862,4.4859004,3.357566,2.4452958,0.69963586,1.0117283,0.6241849,0.2503599,0.12346515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.006859175,0.010288762,0.006859175,0.006859175,0.006859175,0.006859175,0.017147938,0.01371835,0.0,0.0,0.010288762,0.010288762,0.010288762,0.01371835,0.01371835,0.010288762,0.010288762,0.010288762,0.006859175,0.0,0.01371835,0.006859175,0.0034295875,0.006859175,0.006859175,0.01371835,0.01371835,0.030866288,0.0548734,0.06516216,0.12346515,0.15090185,0.13032432,0.082310095,0.06859175,0.09602845,0.06516216,0.037725464,0.041155048,0.037725464,0.0274367,0.044584636,0.07888051,0.11317638,0.14747226,0.12346515,0.106317215,0.12689474,0.18176813,0.23664154,0.216064,0.17833854,0.13032432,0.19548649,0.6207553,1.1111864,0.72364295,0.36696586,0.45270553,0.90198153,1.7971039,2.6064866,2.5996273,2.1194851,2.5824795,1.6770682,2.037175,2.3149714,1.8176813,0.51100856,0.106317215,0.0034295875,0.13032432,0.37039545,0.53844523,0.58988905,0.8196714,1.0734608,1.3375391,1.7353712,1.7079345,1.587899,1.3272504,1.0151579,0.8711152,1.0323058,1.2655178,1.6873571,2.2738166,2.8637056,3.0386145,3.0866287,3.000889,2.9871707,3.4776018,3.6044965,3.5221863,3.974892,5.1992545,6.9380555,7.5039372,8.865483,10.861504,12.71691,13.042721,14.105893,14.853543,15.861842,17.185663,18.334574,16.846134,16.973028,17.844143,18.77699,19.243416,17.243965,15.608052,14.555169,13.725209,12.188754,10.192734,8.186425,6.1766872,4.40702,3.391862,2.7711067,2.452155,2.0920484,1.7147937,1.7079345,1.4953002,1.1763484,0.939707,0.7922347,0.5418748,0.3806842,0.31209245,0.28122616,0.2469303,0.20234565,0.14404267,0.11317638,0.106317215,0.11317638,0.12003556,0.12003556,0.12003556,0.116605975,0.12003556,0.13032432,0.08573969,0.0548734,0.030866288,0.01371835,0.01371835,9.709162,9.31133,9.551401,9.328478,8.172707,6.262427,7.915488,9.321619,9.650859,8.707723,6.9346256,6.012067,5.1100855,4.383013,3.7451096,2.8637056,2.7059445,2.3218307,2.393852,3.7348208,7.281014,10.652299,11.866373,10.419086,8.141841,9.205012,13.361672,19.222837,21.4555,19.140528,15.745236,15.8138275,15.062748,13.200482,10.741467,9.016385,7.7885933,8.608265,9.472521,9.554831,9.218731,11.132441,10.768905,8.786603,7.2878733,9.860064,7.8126,8.152129,11.526843,19.915615,36.607418,111.2764,144.51596,137.35841,112.178375,112.7031,118.65687,136.04488,140.35243,119.73376,75.01194,61.173553,53.772503,44.838425,34.67656,31.860868,22.007662,12.778643,8.196714,8.707723,11.194174,16.45173,12.991278,9.1981535,7.932636,6.5196457,4.6402316,3.0043187,2.3424082,2.4658735,2.253239,2.301253,3.0351849,3.542764,3.4021509,2.6750782,6.2864337,7.3255987,5.3158607,2.5824795,4.256118,6.3653145,9.3079,8.628842,5.086078,4.647091,4.588788,3.724532,4.7534084,6.6533995,4.664239,4.273266,5.56965,5.312431,3.2683969,2.1915064,2.9288676,3.0043187,3.2649672,3.9268777,4.5647807,4.863155,4.48933,4.756838,6.0978065,8.06639,5.9331865,5.669108,7.6033955,9.822338,8.200144,6.557371,5.878313,5.7068334,5.778855,6.0223556,8.001227,12.271064,13.680624,10.556271,4.722542,6.1766872,5.8337283,5.1409516,4.712253,4.355576,5.288424,6.9552035,7.4284863,6.6465406,6.433906,6.166398,5.751418,5.0003386,4.197815,4.1017866,6.4373355,6.5196457,6.7185616,8.162418,10.72775,10.864933,9.465661,7.81603,6.691125,6.341307,7.4799304,8.639131,9.043822,8.81061,8.97523,9.609704,9.081548,8.501947,9.294182,13.210771,9.56512,7.517656,6.999788,7.8606143,9.89436,11.773774,11.626302,8.968371,5.3090014,4.1120753,7.3187394,7.7131424,6.5710897,5.0483527,4.173808,5.188966,5.23698,6.5299344,8.340756,6.992929,5.3501563,4.6848164,4.482471,4.314421,3.8205605,2.8259802,2.8122618,2.5619018,2.1194851,2.8156912,4.297273,4.1635194,3.2615378,2.6407824,3.5633414,2.877424,2.0028791,1.3512574,1.0768905,1.0666018,0.9842916,1.2072148,1.2072148,0.94999576,0.8848336,0.881404,0.9259886,0.9602845,0.9328478,0.7990939,0.7888051,0.64819205,0.65162164,0.8093826,0.8471081,0.6790583,0.6790583,0.7099246,0.7133542,0.72021335,0.6824879,0.6344737,0.64133286,0.6276145,0.36353627,0.20577525,0.09602845,0.06516216,0.08573969,0.06859175,0.09602845,0.08916927,0.09259886,0.12003556,0.15776102,0.274367,0.32238123,0.28122616,0.17490897,0.11317638,0.31209245,0.41840968,0.5041494,0.6207553,0.8265306,0.5590228,0.65162164,0.607037,0.34295875,0.19548649,0.36353627,0.6241849,0.8128122,0.823101,0.6207553,0.77508676,0.7476501,0.64476246,0.6379033,0.9362774,0.84024894,0.7579388,0.90198153,1.3101025,1.8348293,1.1454822,0.864256,0.94656616,1.1283343,0.9259886,0.9534253,1.0117283,0.90198153,0.69963586,0.7476501,1.0597426,1.255229,1.3203912,1.3615463,1.6221949,1.196926,1.1214751,1.0700313,0.9328478,0.7956643,1.0700313,1.2655178,1.3546871,1.4232788,1.6530612,1.821111,1.6907866,1.5707511,1.4918705,1.2312219,1.0734608,1.1146159,1.4987297,1.8897027,1.4507155,1.2758065,0.94656616,0.7407909,0.6927767,0.6001778,0.7510797,1.5227368,1.9342873,1.587899,0.6790583,0.7305021,1.0117283,0.94656616,0.58302987,0.5693115,0.4698535,1.4541451,1.5090185,0.91569984,2.2292318,6.5333643,8.110974,6.451054,3.210094,2.1880767,1.9308578,3.4055803,4.448175,3.9886103,2.0440342,1.7936742,2.7951138,5.254128,10.041832,18.677534,32.731983,30.626217,21.37319,12.912396,12.113303,13.498857,15.035312,13.845244,10.672876,9.860064,12.212761,14.692352,15.9921665,17.367432,22.624989,23.081123,21.4555,20.244854,19.672113,17.71039,19.929333,23.993395,24.998262,23.482386,25.444109,27.254932,27.121178,27.258362,27.138325,23.496103,17.96761,17.62122,18.996485,19.068506,15.254805,15.059319,15.700651,15.539461,13.869251,10.909517,10.930096,18.015623,22.77932,21.126259,14.256795,14.534592,14.990726,14.520873,13.87954,15.700651,9.098696,13.509145,20.62897,23.76361,17.851004,14.843254,14.373401,9.496528,1.862266,1.7250825,3.0386145,4.245829,5.4084597,6.711703,8.443645,11.043272,12.504276,12.425395,11.266195,10.357354,14.994157,18.595222,19.058218,17.497755,18.259123,17.29884,17.86815,18.722118,18.804428,17.237106,15.443433,14.606613,13.567448,11.780633,9.314759,8.038953,5.0757895,2.452155,1.3032433,1.8656956,3.450165,2.702515,3.216953,4.437886,1.6496316,1.5673214,1.6907866,1.8965619,1.9411465,1.4507155,2.603057,1.7422304,1.1626302,1.4198492,1.3443983,1.7250825,2.2566686,3.069481,4.190956,5.552502,4.4413157,4.9523244,5.7822843,6.8043017,9.0644,9.218731,8.371623,7.4010496,6.725421,6.3035817,6.557371,6.258997,6.077229,6.15268,6.135532,4.2046742,3.5976372,2.668219,1.8965619,3.8891523,4.3795834,4.945465,5.645101,6.3893213,6.9380555,6.948344,8.64599,8.779744,7.0923867,6.3001523,9.325048,11.869802,12.614022,12.161317,13.032433,13.577737,12.5145645,11.444533,10.916377,10.401938,8.632272,6.4373355,6.0326443,8.169277,12.168177,10.786053,9.201583,8.704293,9.033533,8.378482,10.082987,11.153018,10.388221,7.596536,3.6010668,4.2046742,4.530485,4.372724,4.3624353,5.9743414,6.5470824,5.0929375,3.234101,1.8382589,1.039165,1.3409687,0.77851635,0.21263443,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.01371835,0.0034295875,0.010288762,0.010288762,0.0,0.0034295875,0.024007112,0.010288762,0.006859175,0.017147938,0.024007112,0.006859175,0.0,0.0,0.0034295875,0.0034295875,0.010288762,0.006859175,0.0034295875,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.017147938,0.041155048,0.16804978,0.15776102,0.08916927,0.041155048,0.07545093,0.07545093,0.0548734,0.048014224,0.0548734,0.044584636,0.0274367,0.06859175,0.13375391,0.1920569,0.23664154,0.17490897,0.1371835,0.15090185,0.20920484,0.2469303,0.18519773,0.09259886,0.034295876,0.13032432,0.5727411,0.84367853,0.66191036,0.48700142,0.4629943,0.4424168,0.85739684,2.2052248,2.6304936,2.1572106,2.7230926,1.9171394,2.054323,2.369845,2.1434922,0.6893471,0.14747226,0.0034295875,0.0,0.072021335,0.36353627,0.5007198,0.71678376,1.0494537,1.3889829,1.5055889,1.5124481,1.4061309,1.1866373,0.96371406,0.9534253,0.8505377,1.0597426,1.5158776,2.1674993,2.9700227,3.2958336,3.6182148,3.7725463,3.649081,3.1860867,2.843128,3.1346428,3.7142432,4.715683,6.7357097,8.440215,10.463672,12.775213,14.311668,12.9809885,14.424845,15.289101,16.143068,16.86671,16.664366,15.642348,15.745236,16.348843,17.322845,19.020493,17.672665,16.232237,15.247946,14.613472,13.560589,12.370522,10.930096,8.594546,5.7925735,4.0434837,3.1826572,2.6819375,2.335549,2.085189,2.0406046,1.5021594,1.214074,0.96714365,0.69963586,0.48357183,0.37382504,0.33609957,0.30866286,0.25721905,0.18176813,0.13375391,0.1097468,0.116605975,0.1371835,0.14747226,0.13375391,0.12346515,0.12003556,0.1371835,0.17490897,0.116605975,0.07545093,0.044584636,0.017147938,0.01371835,7.1712675,7.3187394,11.008976,13.138749,11.4754,6.6533995,8.080108,10.405369,11.101575,9.692014,7.750868,7.48336,6.262427,5.103226,4.437886,4.1189346,4.2183924,3.6936657,3.2718265,3.6559403,5.5250654,6.2075534,6.526505,7.8846216,11.365653,17.700102,31.418451,40.194763,38.476543,28.294096,19.288,18.554068,17.089634,14.359683,11.47197,11.153018,11.118723,10.731179,10.38479,10.511685,11.612583,11.30735,9.016385,7.1952744,7.346176,9.993818,8.639131,8.491658,11.238758,17.429163,26.476416,107.49013,161.46155,173.1873,158.62527,164.91171,189.495,204.35883,184.24773,131.10284,74.03451,60.168682,51.419804,43.716953,34.82746,24.3535,17.761833,12.908967,9.1810055,7.2878733,9.277034,11.4033785,9.325048,6.9620624,5.7239814,4.5167665,3.9063,3.059192,2.2223728,1.6427724,1.5570327,1.9480057,1.9548649,1.6599203,1.2826657,1.1592005,12.778643,9.3764925,3.9165888,2.085189,2.3046827,3.1209247,4.6093655,5.120374,4.5613513,4.3795834,2.3767042,1.7593783,2.6853669,4.297273,4.698535,4.6127954,5.65539,4.9831905,2.8396983,2.534465,2.7539587,2.9906003,3.223812,3.357566,3.234101,2.527606,3.1106358,3.2992632,2.7299516,2.3664153,1.5604624,3.5187566,8.39563,12.864383,10.117283,7.56567,7.239859,10.192734,13.361672,9.551401,7.8674736,7.8674736,6.9963584,5.2747054,5.3090014,5.1512403,5.0277753,5.0483527,5.586798,7.3084507,6.5024977,4.7191124,4.7602673,6.800872,8.361334,8.543102,8.903209,9.266746,9.253027,8.237869,7.5210853,7.6033955,7.4044795,6.6876955,6.0875177,6.5882373,6.9346256,6.842027,6.6705475,7.414768,8.56368,8.988949,8.628842,7.936065,7.888051,6.4716315,5.6519604,6.5299344,9.098696,12.22305,11.22161,8.711152,6.135532,4.461893,4.180667,7.8674736,8.954653,7.9600725,6.1766872,5.675967,6.5196457,7.0032177,7.301592,7.1026754,5.6142344,3.2581081,3.3301294,5.429037,8.056101,8.604835,6.6396813,4.722542,4.2526884,4.9077396,4.6402316,3.3198407,2.4967396,2.0680413,2.3286898,3.9508848,4.866585,4.108646,2.8637056,2.0131679,2.136633,1.9171394,1.9445761,1.7662375,1.371835,1.1900668,1.1660597,1.3889829,1.4129901,1.1523414,0.8848336,0.823101,0.84367853,0.89512235,0.8848336,0.70306545,0.8471081,0.7373613,0.5178677,0.36010668,0.45613512,0.4938606,0.5693115,0.59331864,0.58645946,0.67219913,0.6824879,0.5590228,0.40126175,0.24007112,0.044584636,0.034295876,0.048014224,0.072021335,0.082310095,0.044584636,0.06859175,0.058302987,0.0274367,0.0,0.0,0.23321195,0.40126175,0.34981793,0.16119061,0.1371835,0.19891608,0.32238123,0.40126175,0.45956472,0.65505123,0.97400284,0.86082643,0.48700142,0.20920484,0.548734,0.5624523,0.52815646,0.5144381,0.58302987,0.77851635,0.77851635,0.7339317,0.59331864,0.45956472,0.59674823,0.7407909,0.7407909,1.0768905,1.6393428,1.7250825,1.4061309,1.255229,1.2792361,1.2792361,0.84024894,0.7407909,0.70649505,0.548734,0.37039545,0.5658819,0.8093826,0.9431366,0.96714365,0.9842916,1.2037852,1.0940384,1.3512574,1.5638919,1.4918705,1.0528834,1.1008976,1.196926,1.2380811,1.2758065,1.4953002,1.3992717,1.7662375,2.0097382,2.0268862,2.1983654,2.5756202,2.5893385,2.1469216,1.546744,1.4507155,0.97400284,0.91912943,1.0597426,1.1249046,0.8093826,1.6016173,3.82399,4.5613513,3.0248961,0.53501564,0.7407909,1.9754424,2.1023371,0.97057325,0.39783216,0.59331864,1.4267083,1.3238207,0.5796003,1.371835,4.437886,5.2575574,4.341858,2.6407824,1.5398848,1.9068506,3.6936657,4.955754,4.413879,1.4335675,1.1523414,1.9720128,4.4859004,10.010965,20.567236,29.995173,23.232025,15.498305,13.173045,13.807519,13.954991,15.501736,16.595774,16.341984,14.815818,17.04848,18.02934,15.844694,13.495427,18.890167,22.137987,20.155685,18.173384,17.367432,14.87755,18.69811,20.652975,20.467777,20.478067,25.6053,27.909983,27.793377,26.35295,24.69303,23.911083,20.443771,21.966507,22.148275,18.526632,12.4974165,12.106443,14.352823,14.815818,12.97413,12.1921835,12.144169,15.601193,15.46744,11.4033785,9.825768,13.1593275,13.588025,17.069057,22.94051,23.94195,11.002116,8.443645,14.390549,22.11055,20.03565,11.784062,5.9400454,2.8637056,2.9322972,6.5470824,8.388771,10.377932,12.655178,14.496866,14.328816,12.483699,11.787492,14.586036,19.257133,20.172834,16.79126,15.999025,16.04361,16.770683,19.637817,21.479506,21.476076,21.726437,22.450079,21.973368,19.360022,17.7927,16.595774,15.172495,13.001566,10.827208,7.016936,3.6147852,1.7902447,1.8142518,1.8416885,1.9754424,2.352697,2.5653315,1.6633499,1.5913286,1.8108221,1.7010754,1.3032433,1.3272504,1.0357354,1.2277923,1.6736387,2.0028791,1.7079345,1.4644338,2.2738166,2.9940298,3.1723683,3.0351849,3.0489032,4.4721823,5.576509,7.281014,13.152468,15.155347,11.482259,7.720001,5.7925735,3.9371665,2.8980014,4.2869844,6.883182,8.711152,7.0478024,2.6304936,1.7730967,1.7422304,1.6530612,2.4727325,2.4967396,2.4007113,3.3541365,5.1580997,6.2555676,6.2555676,7.438775,7.2604365,5.456474,4.029765,6.1766872,8.251588,11.413667,14.596324,14.510585,14.30481,13.004995,10.912948,9.256456,10.206452,7.9875093,6.077229,5.5319247,6.636252,8.89635,9.211872,10.316199,11.447963,10.7586155,5.3261495,7.301592,7.8434668,6.708273,5.103226,5.675967,8.155559,9.294182,7.4765005,4.389872,5.0346346,5.254128,4.5784993,2.551613,0.22292319,0.1371835,0.12689474,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.017147938,0.030866288,0.024007112,0.0,0.0,0.017147938,0.017147938,0.0034295875,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.0,0.01371835,0.006859175,0.006859175,0.01371835,0.01371835,0.0034295875,0.010288762,0.010288762,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.20920484,0.19548649,0.1097468,0.06516216,0.1371835,0.08916927,0.048014224,0.037725464,0.044584636,0.044584636,0.044584636,0.1371835,0.23664154,0.28465575,0.26064864,0.11317638,0.06859175,0.09259886,0.12346515,0.07545093,0.11317638,0.06859175,0.030866288,0.037725464,0.061732575,0.09602845,0.18176813,0.29494452,0.4046913,0.4424168,0.37039545,1.155771,2.0474637,2.7333813,3.357566,3.3438478,2.6819375,1.7730967,0.94656616,0.45613512,0.09259886,0.0,0.0,0.020577524,0.106317215,0.36353627,0.6379033,0.84367853,0.9294182,0.8711152,1.0528834,0.9259886,0.78537554,0.78194594,0.91569984,1.0494537,1.5501735,1.99602,2.1880767,2.1503513,2.760818,3.5290456,3.8891523,3.7108135,3.2958336,2.4658735,3.9508848,5.0757895,5.3570156,6.5162163,8.796892,10.017825,11.197603,12.38424,12.665466,15.776102,17.278261,17.95732,17.737827,15.6869335,14.637479,14.373401,16.12592,18.934752,19.668684,19.325726,17.19938,15.086755,13.684054,12.572867,13.255356,12.22648,9.530824,6.2898636,4.715683,3.981751,3.175798,2.5790498,2.2258022,1.9068506,1.7010754,1.7936742,1.5673214,0.99801,0.65505123,0.48357183,0.432128,0.37382504,0.26407823,0.16804978,0.13032432,0.14061308,0.16462019,0.18176813,0.18176813,0.17147937,0.15776102,0.17833854,0.20920484,0.19891608,0.19891608,0.18862732,0.12346515,0.0274367,0.01371835,4.290414,4.681387,8.330468,10.487679,10.024684,9.410788,10.751757,11.633161,11.032983,9.582268,9.595985,11.581717,10.734609,9.736599,9.211872,7.73372,6.2967224,5.1100855,4.911169,5.7891436,7.208993,8.049242,7.846896,9.115844,13.478279,21.678423,30.694807,33.363026,28.883986,20.159115,13.807519,12.936404,12.281353,11.396519,10.744898,11.667457,10.9369545,10.621432,13.176475,16.986746,16.335125,11.166737,8.700864,8.076678,8.573969,9.592556,7.5931067,6.9689217,7.9189177,10.909517,16.684942,47.510075,74.850746,89.67342,97.75353,119.70289,160.92996,190.8634,181.0445,132.41295,75.31717,55.79596,44.152508,37.204166,31.487043,23.280039,17.799559,14.983868,13.169616,11.629731,10.583707,10.079557,8.237869,6.2418494,4.756838,3.9303071,3.309552,2.8259802,2.3595562,1.9274281,1.6667795,1.6873571,1.7593783,1.6153357,1.7319417,3.3678548,9.383351,8.827758,6.334448,4.0366244,1.5707511,2.4761622,4.2938433,4.3658648,2.942586,3.1586502,4.945465,4.98662,4.5956473,4.705394,5.857735,5.079219,4.695105,3.858286,2.6956558,2.311542,2.2978237,3.3712845,4.184097,4.108646,3.234101,3.2203827,4.664239,5.885172,6.0497923,5.195825,6.56766,8.340756,9.554831,9.187865,6.138962,6.358455,6.7048435,7.2021337,7.3221693,5.9743414,6.3035817,5.254128,4.3349986,4.5819287,6.543653,4.9008803,4.756838,4.976331,5.0003386,4.856296,5.9640527,5.9469047,6.5710897,8.124693,9.424506,9.959522,10.14129,9.338767,7.81603,6.715132,6.6293926,6.279575,6.118384,5.9160385,4.770556,5.5730796,6.492209,6.694555,6.001778,4.9008803,5.610805,5.844017,5.9126086,6.327589,7.7920227,7.164408,6.1458206,5.2747054,5.703404,9.218731,10.590566,9.692014,8.076678,6.5813785,5.305572,5.9331865,7.2432885,8.213862,8.399059,7.9463544,7.3530354,5.8817425,6.0052075,8.114404,10.511685,6.464772,4.962613,7.425057,11.341646,10.278474,7.0032177,5.0140567,4.5819287,4.90431,4.0880685,4.166949,3.9783216,3.9954693,4.5647807,5.90575,4.2423997,3.3061223,2.726522,2.3218307,2.1126258,1.6976458,1.6770682,1.6359133,1.4644338,1.3615463,1.1111864,1.3306799,1.6324836,1.6530612,1.0323058,0.939707,0.85396725,0.7510797,0.6310441,0.50757897,0.47671264,0.47671264,0.45613512,0.42526886,0.44584638,0.48357183,0.490431,0.4664239,0.44584638,0.51100856,0.5727411,0.5178677,0.37039545,0.19548649,0.106317215,0.06516216,0.05144381,0.061732575,0.06859175,0.034295876,0.08573969,0.10288762,0.06516216,0.0,0.0,0.06516216,0.14747226,0.21263443,0.23664154,0.20920484,0.2503599,0.22635277,0.25721905,0.3841138,0.5693115,0.6344737,0.4664239,0.41840968,0.5453044,0.5727411,0.45956472,0.40126175,0.51100856,0.6927767,0.64476246,0.65505123,0.9602845,1.138623,1.0220171,0.71678376,0.6207553,0.6379033,0.83681935,1.1008976,1.138623,1.0837497,0.939707,0.83338976,0.77165717,0.64476246,0.7510797,0.9877212,1.1283343,1.2003556,1.4918705,1.1592005,1.1729189,1.1317638,0.97400284,0.94999576,1.0357354,1.2517995,1.3032433,1.1420527,0.9568549,1.0425946,1.1317638,1.1660597,1.1694894,1.2620882,1.2723769,1.3478279,1.4918705,1.6736387,1.7936742,2.1812177,2.1812177,1.8656956,1.5604624,1.8656956,1.7799559,1.6256244,1.4507155,1.1763484,0.5761707,1.0082988,1.9308578,2.061182,1.2106444,0.3018037,0.8128122,1.5433143,1.5055889,0.7442205,0.34638834,0.5521636,0.922559,0.9259886,0.7305021,1.2037852,1.845118,2.3458378,2.294394,1.8039631,1.5158776,1.8245405,2.6133456,3.5153272,3.4844608,0.7990939,0.939707,2.4315774,5.7136927,11.561139,21.10568,20.7833,14.932424,11.832077,12.830087,12.332796,11.091286,11.135871,11.705182,12.229909,12.325937,16.221949,19.86417,20.025362,17.45317,16.852993,19.514353,18.512913,16.11906,13.533153,10.88551,12.548861,13.903547,12.339656,9.187865,9.72288,13.214201,16.407146,19.171394,20.61868,19.12681,14.651197,14.846684,15.357693,14.38026,12.668896,13.166186,11.05699,9.283894,9.493098,12.034423,14.572317,13.841815,11.262765,9.1810055,10.875222,9.043822,10.216741,12.847235,15.46744,16.702091,15.343974,18.115082,22.52553,25.385807,22.793037,11.787492,7.040943,6.680836,8.268735,8.81747,11.002116,13.594885,16.616352,18.999914,18.62609,16.558048,16.835844,18.756414,20.488356,19.061647,15.182784,13.05301,12.740917,14.411126,18.296848,22.19972,25.756203,26.551867,24.655304,22.607841,21.506943,21.057667,19.384027,16.914726,16.383139,13.474849,9.355915,5.6142344,2.942586,1.1317638,1.1866373,1.1214751,1.3169615,1.7696671,2.1160555,2.6579304,2.935727,2.8877127,2.5619018,2.095478,1.0700313,1.1900668,1.8416885,2.2738166,1.5981878,2.1160555,2.5001693,3.210094,4.1463714,4.647091,4.9831905,5.4016004,5.3913116,6.667118,13.152468,14.177915,9.952662,5.9812007,4.3178506,3.5461934,3.923448,5.271276,5.3673043,4.249259,4.2286816,3.0146074,2.4898806,2.4967396,2.74367,2.8019729,2.2600982,2.177788,2.935727,4.482471,6.341307,5.0826488,5.5833683,6.001778,5.7925735,5.7136927,5.206114,5.7308407,7.051232,8.594546,9.445084,8.447074,7.9257765,9.335337,11.050131,8.388771,7.0478024,4.9831905,3.7553983,3.5016088,2.9391565,4.7019644,8.268735,10.508256,9.9801,6.948344,8.632272,8.375052,7.641121,7.3050213,7.654839,7.641121,7.040943,5.40503,3.2443898,2.0097382,1.8554068,1.255229,0.66533995,0.29151493,0.08916927,0.037725464,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.010288762,0.0034295875,0.006859175,0.01371835,0.01371835,0.01371835,0.024007112,0.020577524,0.006859175,0.01371835,0.01371835,0.017147938,0.010288762,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.0,0.01371835,0.006859175,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0034295875,0.01371835,0.0548734,0.058302987,0.05144381,0.06516216,0.1371835,0.106317215,0.116605975,0.13375391,0.12689474,0.058302987,0.106317215,0.30523327,0.37382504,0.26407823,0.16119061,0.07545093,0.041155048,0.048014224,0.061732575,0.05144381,0.048014224,0.09602845,0.20577525,0.28122616,0.1097468,0.36010668,0.70306545,0.66876954,0.31552204,0.23664154,0.5624523,0.83338976,1.3341095,2.1332035,3.0900583,2.2086544,2.3149714,2.5893385,2.4658735,1.6530612,1.0425946,0.3841138,0.030866288,0.017147938,0.082310095,0.30866286,0.71678376,0.99801,0.96371406,0.5418748,0.5658819,0.53158605,0.5041494,0.5007198,0.48700142,0.61389613,0.86082643,1.2449403,1.6599203,1.9068506,2.4384367,2.9940298,3.5118976,3.875434,3.9303071,3.6868064,5.429037,7.2638664,8.333898,8.81061,11.015835,13.029003,14.1299,14.538021,15.436573,16.331696,17.103354,17.864721,18.45461,18.44432,17.110212,16.756964,19.329155,23.321196,23.770472,19.150816,16.863281,16.61292,17.171944,16.393429,16.239098,15.151917,12.346515,8.663138,6.5710897,5.936616,4.9694724,3.99204,3.1483612,2.4315774,1.978872,1.903421,1.5844694,1.0288762,0.864256,0.7510797,0.6927767,0.5624523,0.37039545,0.25378948,0.15776102,0.13032432,0.14404267,0.17147937,0.17147937,0.14747226,0.14061308,0.15433143,0.16804978,0.1371835,0.12689474,0.15090185,0.13375391,0.08573969,0.11317638,5.0895076,5.7754254,7.3564653,8.128122,8.117833,9.084977,11.019264,12.761495,17.031332,25.039417,36.473663,34.07638,25.711617,18.62266,15.3302555,13.670336,10.995257,8.2481575,6.8557453,6.6705475,5.953764,6.327589,7.4113383,8.447074,9.8429165,13.173045,17.844143,19.03421,16.935303,13.419975,12.0138445,12.408247,11.592006,10.799771,10.906088,12.408247,12.6757555,14.006435,16.252815,17.480608,13.954991,8.546532,6.7871537,6.725421,7.006647,6.8900414,6.7528577,7.1095347,7.7680154,9.112414,12.120162,18.348293,27.553307,41.628334,64.35621,101.4129,138.58963,159.9251,154.66411,124.27453,82.44728,51.406086,35.681427,29.08633,25.67732,19.740705,16.167076,13.738928,11.845795,10.233889,9.006097,8.491658,7.0958166,5.4736214,4.1017866,3.2889743,2.843128,2.6407824,2.527606,2.411,2.2600982,2.0989075,2.1091962,2.3046827,3.1072063,5.360445,6.375603,7.373613,6.944915,5.1238036,3.3850029,2.9631636,4.0091877,4.2698364,3.6970954,4.4447455,5.717122,5.7719955,5.658819,6.427047,9.132992,5.5662203,3.649081,2.7402403,2.5481834,3.1277838,3.508468,5.3090014,6.3447366,5.8645945,4.5613513,4.729401,8.755736,10.161868,7.4627824,4.1943855,7.3187394,7.5382333,5.9812007,4.1772375,4.0709205,4.8185706,5.442755,6.046363,6.601956,6.9380555,9.760606,9.294182,7.291303,5.638242,6.3310184,5.48734,5.6656785,6.4819202,7.0752387,6.135532,6.677407,7.2295704,8.22758,9.23245,8.920357,8.848335,8.855195,8.052671,6.691125,6.1766872,5.377593,4.852866,4.9351764,5.3981705,5.429037,5.977771,7.0135064,7.507367,7.133542,6.2692857,6.2144127,6.4236174,6.2555676,6.018926,6.9689217,6.7048435,6.5162163,5.8817425,5.7068334,8.330468,9.22902,8.858624,8.529384,8.399059,7.490219,5.9640527,6.3001523,7.2295704,8.1041155,8.906639,9.033533,6.677407,5.5833683,7.5279446,12.339656,9.541112,7.5519514,8.683716,11.341646,10.045261,7.1061053,5.6348124,5.329579,5.439326,4.756838,4.619654,4.307562,4.3281393,4.856296,5.7068334,4.6093655,3.292404,2.393852,2.020027,1.7490896,1.6667795,1.6839274,1.7079345,1.6153357,1.2655178,0.9534253,1.08032,1.4095604,1.5741806,1.0871792,1.1489118,1.1351935,0.91227025,0.5693115,0.39440256,0.4972902,0.5178677,0.44927597,0.37382504,0.45956472,0.47671264,0.48357183,0.44927597,0.39440256,0.39097297,0.4355576,0.42526886,0.31895164,0.16119061,0.08573969,0.06516216,0.034295876,0.024007112,0.0274367,0.01371835,0.037725464,0.048014224,0.030866288,0.0,0.0,0.010288762,0.06859175,0.12689474,0.15776102,0.15433143,0.2503599,0.24007112,0.25721905,0.33952916,0.42183927,0.37039545,0.274367,0.39440256,0.6276145,0.4972902,0.4081209,0.36010668,0.45956472,0.61389613,0.51100856,0.5144381,0.86082643,1.0151579,0.85739684,0.6927767,0.71678376,0.8025235,0.90541106,0.96371406,0.90198153,0.83338976,0.6962063,0.58988905,0.5624523,0.6241849,0.8471081,1.0048691,1.0220171,1.0220171,1.2929544,1.3958421,1.2209331,0.922559,0.6893471,0.72021335,0.89855194,1.0631721,1.0734608,0.9431366,0.8196714,0.9911508,1.0837497,1.1420527,1.1592005,1.0597426,1.0597426,1.0940384,1.1832076,1.2483698,1.1077567,1.4918705,1.6839274,1.7799559,1.7936742,1.6496316,1.3889829,1.2723769,1.1077567,0.83338976,0.53844523,1.1043272,2.5070283,3.1895163,2.527606,0.8196714,1.1008976,1.2689474,1.0117283,0.52472687,0.52815646,1.196926,1.6804979,1.6942163,1.3409687,1.1317638,1.3512574,1.5776103,1.7456601,1.8348293,1.8588364,2.0714707,2.8054025,3.6559403,3.6216443,1.097468,1.0494537,2.2326615,5.3501563,10.007536,14.712931,13.104454,9.277034,7.2707253,7.582818,7.174697,5.953764,6.0875177,7.010077,8.189855,9.122703,12.72034,17.075916,19.21255,19.027351,19.308577,21.795029,19.576086,15.097044,10.823778,9.266746,8.995808,9.273604,8.450503,7.164408,8.333898,9.373062,10.072699,11.063849,11.760056,10.367643,9.774324,10.343636,9.791472,7.970361,6.8969,7.888051,7.0375133,6.427047,7.1987042,9.55826,12.860953,12.185325,9.609704,8.1487,11.760056,11.2593355,13.5503,17.333136,20.649546,20.896477,24.758192,28.544456,29.419,26.496992,20.848463,11.825217,7.7885933,7.81603,10.600855,14.438563,19.013634,21.723007,22.624989,21.846472,19.589804,16.753534,15.450292,15.827546,17.147938,17.785841,14.095605,13.070158,13.516005,15.289101,19.294859,23.869928,27.892836,29.079472,27.594461,26.051146,24.981115,22.542679,20.337454,18.95533,17.977898,16.420864,14.452282,11.132441,6.848886,3.3061223,2.2223728,1.5501735,1.214074,1.3169615,2.136633,3.0900583,3.192946,2.7882545,2.2292318,1.8759843,1.0288762,1.2072148,1.7388009,2.0234566,1.5158776,3.4124396,3.758828,4.5956473,6.200694,7.1026754,6.667118,7.2192817,7.81603,8.47451,10.179015,11.814929,9.688584,6.9826403,5.144381,3.8617156,4.513337,5.003768,4.5510626,3.5187566,3.433017,3.2306714,2.702515,2.7333813,3.3369887,3.6696587,3.1415021,2.9974594,3.1655092,4.1943855,7.2432885,6.81802,6.6636887,6.135532,5.4736214,5.8405876,5.1169443,5.48734,5.936616,6.15268,6.5230756,6.944915,7.0443726,8.40249,9.417647,5.2987127,4.928317,3.7279615,2.6750782,2.386993,3.1140654,3.7691166,4.90431,6.138962,7.0032177,6.924337,8.762596,9.016385,8.659708,8.056101,6.948344,7.2947326,6.8111606,4.513337,1.4267083,0.5727411,0.432128,0.274367,0.26750782,0.32924038,0.14061308,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.0,0.0034295875,0.0034295875,0.006859175,0.01371835,0.006859175,0.01371835,0.020577524,0.01371835,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.01371835,0.020577524,0.017147938,0.010288762,0.01371835,0.024007112,0.034295876,0.048014224,0.07545093,0.12003556,0.1097468,0.13375391,0.19891608,0.24007112,0.12346515,0.16462019,0.6310441,0.65162164,0.19548649,0.082310095,0.061732575,0.044584636,0.041155048,0.044584636,0.044584636,0.0274367,0.082310095,0.28808534,0.47671264,0.2503599,0.32924038,0.6790583,0.6001778,0.15090185,0.12689474,0.31209245,0.41840968,0.77165717,1.5021594,2.5550427,1.5158776,1.4232788,1.6084765,1.5981878,1.138623,0.97400284,0.5727411,0.20234565,0.006859175,0.030866288,0.18519773,0.490431,0.7407909,0.7442205,0.34638834,0.29837412,0.36010668,0.4629943,0.52815646,0.4629943,0.7339317,0.89855194,1.1111864,1.3615463,1.4815818,2.1983654,2.3629858,2.4555845,2.7813954,3.457024,4.1155047,5.4839106,7.3050213,8.940934,9.383351,11.2250395,12.864383,13.663476,14.171056,16.091625,17.408587,18.03277,18.917604,19.994495,20.159115,18.77699,18.392878,20.982216,25.10458,25.93111,21.53781,19.648108,19.991066,20.94792,19.565796,17.923023,16.595774,14.5414505,11.7086115,9.002667,7.373613,6.0497923,4.9831905,4.1292233,3.450165,2.7128036,2.294394,1.8588364,1.3649758,1.08032,0.89512235,0.8711152,0.7510797,0.5041494,0.32924038,0.20577525,0.16462019,0.18176813,0.21263443,0.21263443,0.17490897,0.14747226,0.1371835,0.13032432,0.08573969,0.06516216,0.082310095,0.08573969,0.07888051,0.09945804,7.610255,7.7680154,8.203573,9.246168,10.041832,8.543102,11.578287,19.099373,35.33847,59.547928,85.9969,66.86667,42.351974,26.116308,20.96164,18.821575,15.337115,11.849225,9.249598,7.5107965,5.6656785,5.895461,7.3564653,8.052671,7.6616983,7.5382333,8.944365,9.9801,11.029553,12.233338,13.461131,13.96185,12.9638405,12.082437,12.312219,13.996146,15.165636,17.04162,17.432592,15.419425,11.345076,8.327039,6.307011,5.5559316,5.645101,5.439326,6.495639,7.0306544,7.442205,8.40249,10.851214,9.630281,12.195613,26.946268,54.513294,87.74943,102.58925,106.71162,102.304596,91.03497,74.06537,43.260815,26.942839,20.515793,18.581505,14.925565,13.066729,11.46854,9.928656,8.484799,7.4181976,7.0272245,5.703404,4.266407,3.1723683,2.5138876,2.253239,2.4315774,2.9322972,3.5221863,3.8548563,3.7313912,3.5050385,3.4981792,3.9474552,4.9934793,4.0777793,4.945465,5.98463,6.135532,4.9180284,3.6627994,3.6010668,3.6868064,3.7039545,4.262977,4.0846386,4.3933015,4.9934793,6.0978065,8.354475,4.7362604,2.8499873,3.6285036,5.9400454,6.5882373,5.284994,6.728851,7.747438,7.239859,6.1629686,6.5950966,9.530824,9.31133,5.470192,2.7573884,7.06495,6.5230756,4.098357,2.5207467,4.2595477,4.8425775,5.2266912,5.8474464,6.6533995,7.116394,9.856634,9.962952,8.337327,6.416758,6.1904054,6.478491,6.444195,7.3839016,8.700864,7.881192,7.720001,7.857185,8.940934,10.196163,9.445084,8.093826,7.239859,6.3173003,5.5422134,5.895461,4.839148,4.664239,5.0449233,5.586798,5.826869,6.2487082,7.239859,7.5382333,7.1266828,7.250148,7.4696417,8.018375,7.486789,6.2830043,6.6396813,6.81802,6.6636887,6.39961,6.7940125,9.15014,9.863494,8.776315,8.742019,10.134431,10.834066,8.711152,7.39762,6.701414,6.6876955,7.6616983,9.22216,7.3084507,5.610805,6.3481665,10.257896,9.753747,8.436785,8.8929205,10.686595,10.374502,7.6033955,6.4819202,6.090947,5.754848,5.0449233,4.996909,4.6093655,4.4447455,4.6779575,5.0895076,5.0174866,3.6353626,2.4898806,2.1263442,2.0920484,1.9342873,1.8759843,1.786815,1.5776103,1.1763484,0.9568549,0.9568549,1.1934965,1.430138,1.1729189,1.3478279,1.4267083,1.1900668,0.72021335,0.39440256,0.61389613,0.70649505,0.58302987,0.38754338,0.48014224,0.50757897,0.5144381,0.47671264,0.39440256,0.31209245,0.29151493,0.26407823,0.1920569,0.08916927,0.037725464,0.037725464,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.08573969,0.09259886,0.09945804,0.19548649,0.24007112,0.25721905,0.26750782,0.29837412,0.2194936,0.18862732,0.31209245,0.48700142,0.38754338,0.31895164,0.32238123,0.37382504,0.41498008,0.34981793,0.3566771,0.58302987,0.66533995,0.548734,0.51100856,0.7682276,0.85739684,0.89169276,0.8779744,0.7476501,0.6927767,0.58645946,0.5007198,0.4972902,0.61046654,0.89855194,0.90884066,0.764798,0.65848076,0.8779744,1.2072148,1.0528834,0.71678376,0.48014224,0.6036074,0.7476501,0.823101,0.8162418,0.7442205,0.65505123,0.90541106,1.0185875,1.097468,1.1111864,0.89512235,0.8848336,0.9534253,1.0151579,1.0014396,0.864256,1.0117283,1.3272504,1.6907866,1.8348293,1.3375391,1.0597426,0.90884066,0.823101,0.8093826,0.9534253,1.1832076,4.187526,6.358455,5.638242,1.5158776,1.1489118,0.88826317,0.6310441,0.45270553,0.6207553,1.4610043,1.862266,2.037175,1.920569,1.1763484,1.3272504,1.4129901,1.704505,2.0577524,1.9239986,2.4315774,3.223812,3.8308492,3.5839188,1.6290541,1.2586586,2.2909644,4.6745276,7.3839016,8.4264965,7.3701835,5.0243454,3.4192986,3.3061223,4.170378,4.32128,5.24041,5.994919,6.375603,6.910619,10.257896,14.942713,18.512913,20.742146,23.629858,26.232914,22.830763,16.016174,10.048691,10.868362,9.523964,8.045813,6.7802944,6.358455,7.6925645,7.2947326,7.3118806,8.158989,9.729739,11.4205265,12.322508,11.694893,11.4205265,11.7086115,11.087856,14.239647,9.9801,6.680836,7.2192817,8.988949,12.610593,12.277924,10.082987,8.831187,12.024134,14.483148,19.215979,24.912523,28.359259,24.425522,27.323523,29.871706,29.43615,25.629307,20.28944,13.392539,9.674867,9.510246,12.425395,17.093063,22.690151,25.406384,24.576424,21.10568,17.436022,15.865272,14.3974085,15.049029,17.511473,19.140528,16.753534,16.352274,16.540901,17.141079,19.20569,22.95423,26.19176,27.484715,27.323523,28.115759,29.68994,26.112879,23.180582,22.415783,21.095392,20.598103,20.265432,18.077356,13.704632,8.505377,6.7494283,4.125794,1.9925903,1.2072148,2.1057668,3.1106358,2.9940298,2.7745364,2.5550427,1.5364552,0.99801,1.3889829,1.8759843,2.085189,2.095478,4.846007,6.077229,7.3221693,8.56368,8.2481575,8.8929205,10.364213,11.777204,12.240198,10.854645,11.105004,9.990388,8.584257,7.257007,5.662249,5.672538,5.5147767,4.98662,4.173808,3.4467354,3.309552,2.6407824,2.534465,3.1792276,3.865145,3.8891523,3.9954693,3.7348208,3.782835,5.9434752,6.848886,7.1369715,6.3378778,4.9591837,4.479041,4.6882463,5.144381,5.5593615,5.720552,5.4770513,7.034084,6.447624,6.5470824,6.7665763,3.1380725,3.1792276,2.784825,2.1572106,2.0989075,4.0263357,4.9248877,4.7328305,4.8082814,5.501058,6.125243,7.9600725,8.772884,8.570539,7.4353456,5.5387836,7.3118806,7.1712675,4.57164,1.0288762,0.13375391,0.12346515,0.52815646,0.70649505,0.48357183,0.13375391,0.06516216,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.01371835,0.0,0.0,0.0,0.006859175,0.01371835,0.006859175,0.006859175,0.01371835,0.010288762,0.010288762,0.020577524,0.017147938,0.01371835,0.010288762,0.006859175,0.010288762,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.006859175,0.01371835,0.010288762,0.010288762,0.010288762,0.010288762,0.01371835,0.017147938,0.01371835,0.010288762,0.01371835,0.0274367,0.037725464,0.048014224,0.06859175,0.09602845,0.10288762,0.12003556,0.17833854,0.23664154,0.15433143,0.16119061,0.53501564,0.52815646,0.13375391,0.07545093,0.058302987,0.06516216,0.058302987,0.041155048,0.041155048,0.024007112,0.12689474,0.28465575,0.45956472,0.6276145,0.5555932,0.50757897,0.30523327,0.041155048,0.09259886,0.16462019,0.18519773,0.5453044,1.3649758,2.5070283,1.1832076,0.71678376,0.59674823,0.5178677,0.38754338,0.5007198,0.45270553,0.2503599,0.01371835,0.0,0.06516216,0.2469303,0.39097297,0.39097297,0.16462019,0.25721905,0.4972902,0.66876954,0.64476246,0.39783216,0.66876954,0.78537554,0.90541106,1.0597426,1.1317638,1.9239986,2.1194851,2.1160555,2.2635276,2.877424,4.0674906,5.6142344,7.534804,9.325048,9.938945,11.1393,12.600305,13.073587,13.193623,15.45715,17.902447,18.554068,19.312008,20.61182,21.434921,21.500084,22.415783,24.0174,25.625877,26.064865,23.928232,23.146286,23.098272,22.964518,21.705858,19.363451,18.320856,17.062197,14.898128,11.938394,9.002667,7.421627,6.2727156,5.195825,4.417309,3.5359046,2.7093742,2.1160555,1.7490896,1.4232788,1.1008976,0.9431366,0.78537554,0.5796003,0.40126175,0.25378948,0.19891608,0.20577525,0.23321195,0.23664154,0.18862732,0.15090185,0.12346515,0.09602845,0.048014224,0.024007112,0.024007112,0.030866288,0.044584636,0.07545093,8.985519,8.035523,9.6645775,13.893259,17.233677,12.6929035,15.505165,31.147512,60.25785,99.02248,139.18637,98.77212,56.330975,30.866287,24.281479,21.342323,18.012194,15.2033615,12.339656,9.56512,7.7131424,7.689135,7.9086285,8.361334,8.934075,9.403929,9.012956,9.592556,11.893809,14.815818,15.426285,16.616352,16.259674,15.134769,14.373401,15.470869,16.983316,17.511473,15.824117,12.603734,10.429376,10.113853,7.531374,5.926327,6.0737996,6.2487082,7.0889573,7.0889573,7.2878733,8.505377,11.365653,10.573419,14.2190695,29.803116,53.138027,68.34482,60.18583,53.172325,48.940212,48.110252,50.274323,32.474762,19.871029,13.660047,12.099585,10.508256,10.069269,9.959522,9.424506,8.237869,6.7219915,5.8817425,4.417309,3.0866287,2.2463799,1.8485477,1.7113642,2.510458,3.666229,4.671098,5.099797,5.147811,4.588788,3.9886103,3.542764,3.07634,2.8808534,2.5927682,4.307562,6.7974424,5.528495,4.4756117,3.590778,2.9494452,2.534465,2.2669573,1.7422304,2.3286898,3.2786856,3.981751,3.957744,2.9151495,2.7299516,5.545643,9.582268,9.136421,5.5902276,5.926327,6.773435,6.701414,6.2418494,6.835168,5.892031,3.8308492,1.9891608,2.6133456,6.368744,6.262427,4.8768735,4.180667,5.5319247,6.042933,5.8817425,5.6176643,5.453044,5.23698,5.9743414,6.416758,6.7357097,6.8969,6.6876955,6.8283086,6.183546,6.7700057,8.289313,8.14527,8.080108,7.610255,8.399059,10.028113,10.000677,7.6616983,6.166398,5.206114,4.880303,5.6999745,5.2301207,5.593657,6.094377,6.2041235,5.56965,5.919468,6.632822,6.39961,5.658819,6.5985265,7.963502,9.0644,8.405919,6.7185616,6.9552035,7.7028537,6.9209075,6.4304767,7.281014,9.740028,11.502836,9.729739,9.030104,10.950673,13.96185,12.55915,10.398509,7.9120584,5.919468,5.5902276,8.1487,7.4696417,6.23156,5.9126086,6.8111606,8.282454,7.956643,8.196714,9.554831,10.7586155,8.2481575,7.4181976,6.8557453,6.025785,5.2781353,5.658819,5.453044,4.9488945,4.547633,4.763697,5.113515,4.07435,3.275256,3.223812,3.2958336,2.335549,2.0303159,1.8142518,1.471293,1.1351935,1.0528834,1.0014396,1.1351935,1.3306799,1.1832076,1.3306799,1.471293,1.3341095,0.91569984,0.490431,0.7956643,0.91569984,0.7510797,0.45956472,0.48357183,0.5521636,0.52815646,0.45613512,0.36010668,0.23664154,0.17147937,0.12346515,0.06516216,0.01371835,0.0,0.0,0.030866288,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.05144381,0.07888051,0.09602845,0.106317215,0.12003556,0.16804978,0.19548649,0.20920484,0.28465575,0.18519773,0.16119061,0.20577525,0.274367,0.29151493,0.1920569,0.274367,0.32238123,0.2777966,0.26407823,0.22978236,0.31895164,0.39440256,0.39097297,0.33266997,0.6927767,0.7099246,0.69963586,0.7133542,0.5418748,0.5727411,0.5144381,0.45613512,0.45956472,0.5761707,0.86082643,0.805953,0.6344737,0.53501564,0.65848076,0.72707254,0.7476501,0.6276145,0.47671264,0.58988905,0.6824879,0.6790583,0.64819205,0.6241849,0.6001778,0.8779744,1.0117283,1.039165,0.96371406,0.7339317,0.8025235,0.90198153,0.9602845,0.97400284,1.0151579,0.8848336,1.1454822,1.4850113,1.6084765,1.2277923,1.1180456,0.8779744,0.8676856,1.1694894,1.5673214,1.1317638,4.866585,7.8023114,7.0306544,1.7182233,0.90884066,0.61046654,0.59331864,0.65162164,0.6241849,1.0734608,1.471293,2.5653315,3.391862,1.2655178,1.138623,1.4678634,2.1503513,2.6064866,1.7593783,2.411,3.000889,3.2375305,2.9665933,2.170929,1.646202,2.7128036,4.201245,5.2026844,5.055212,3.542764,2.218943,2.2155135,3.5187566,4.979761,5.8508763,7.222711,7.4010496,6.40304,5.994919,9.23245,13.941273,17.977898,21.157125,25.258911,27.93399,24.6896,17.36057,10.823778,12.987847,12.627741,10.079557,7.2947326,5.5730796,5.5319247,5.4187484,7.3393173,10.261326,13.824667,18.348293,17.134218,14.592895,15.830976,19.78529,19.21255,23.94195,14.544881,7.442205,8.032094,10.696883,13.540011,12.288212,10.878652,11.393089,14.057879,16.338554,22.573545,29.196077,31.565924,23.976246,23.211449,23.965958,24.10314,22.971376,21.410915,15.971589,13.207341,13.677195,15.937293,16.530611,21.071384,23.516682,22.659285,19.390888,16.726099,17.580065,16.96617,18.392878,21.45207,21.812176,20.474638,19.665255,19.099373,18.670673,18.46147,21.3629,23.965958,25.173172,25.780209,28.465576,32.74913,30.389574,27.741934,26.836521,25.375517,24.535269,24.120289,23.372639,20.886189,14.592895,12.836946,8.011517,3.865145,2.1160555,2.4795918,3.0283258,2.7951138,3.069481,3.426158,1.7593783,1.3821237,1.9137098,2.4761622,2.942586,3.9337368,6.8626046,8.848335,10.244178,10.7757635,9.541112,11.989838,13.564018,14.850114,15.638919,14.904987,12.168177,10.041832,9.146709,9.102125,8.519095,8.008087,7.671987,6.7631464,5.3330083,4.2218223,4.6882463,3.7931237,3.0489032,3.0557625,3.5050385,4.081209,4.3452873,3.8891523,3.0523329,2.9151495,4.232111,5.4324665,5.48734,4.331569,2.8637056,3.6559403,4.033195,4.8905916,5.768566,4.8494368,6.7528577,5.2987127,4.4241676,4.5510626,2.5996273,2.8739944,2.8088322,2.4144297,2.3561265,3.957744,6.790583,7.39762,6.9620624,6.2075534,5.3981705,7.7714453,8.553391,7.864044,6.2487082,4.6779575,7.0615206,6.958633,4.914599,2.0749004,0.20234565,0.47671264,1.2346514,1.3889829,0.7579388,0.06859175,0.07545093,0.0548734,0.024007112,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.006859175,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.017147938,0.030866288,0.017147938,0.01371835,0.01371835,0.01371835,0.0,0.01371835,0.010288762,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.006859175,0.010288762,0.01371835,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.006859175,0.020577524,0.030866288,0.034295876,0.048014224,0.061732575,0.06859175,0.08573969,0.08573969,0.09259886,0.11317638,0.116605975,0.106317215,0.1097468,0.1097468,0.11317638,0.13032432,0.06859175,0.07545093,0.06516216,0.0274367,0.024007112,0.06516216,0.2503599,0.28808534,0.36010668,1.1351935,1.0014396,0.4115505,0.024007112,0.020577524,0.1097468,0.2194936,0.17833854,0.5590228,1.4472859,2.469303,1.0117283,0.5212973,0.34638834,0.18176813,0.072021335,0.082310095,0.14747226,0.12689474,0.030866288,0.0,0.0,0.09602845,0.13032432,0.07545093,0.037725464,0.90198153,1.2072148,1.0940384,0.70649505,0.18176813,0.29494452,0.5007198,0.764798,0.9911508,0.99801,1.5776103,2.0920484,2.3424082,2.352697,2.3732746,3.4227283,5.40503,7.641121,9.47938,10.30934,10.847785,13.55373,14.393978,13.37882,14.586036,17.278261,18.362011,19.54522,21.37319,23.249174,25.639595,28.489584,29.00745,27.289227,26.318655,25.76649,25.913963,25.365229,24.055126,23.262892,21.428062,20.827885,19.761284,17.573206,14.640909,10.89237,9.129561,7.7920227,6.3378778,5.2472687,4.461893,3.3815732,2.5001693,2.0097382,1.762808,1.4164196,1.0494537,0.78537554,0.6379033,0.50757897,0.3566771,0.274367,0.25721905,0.2709374,0.2777966,0.21263443,0.15433143,0.11317638,0.07888051,0.030866288,0.006859175,0.0,0.0,0.01371835,0.061732575,5.4324665,4.149801,9.211872,18.986197,28.304386,28.486153,26.253492,44.581207,74.15454,111.794266,160.47383,115.52908,67.83724,35.794605,23.475527,20.646116,19.387459,18.149376,16.489456,14.119612,10.909517,8.748878,7.349606,8.025234,10.456812,12.665466,12.017275,11.88352,12.566009,13.437123,12.922686,21.407484,23.262892,20.20027,15.553179,14.29795,16.444872,14.832966,11.821788,9.208443,8.193284,8.241299,7.9909387,8.128122,8.447074,7.8126,8.680285,9.873782,11.327928,12.535142,12.572867,9.9869585,11.88352,20.659836,33.983784,44.786983,45.836437,48.06567,47.37632,42.033024,32.67025,25.029129,17.394867,11.705182,8.848335,8.652849,10.127572,10.497967,9.619993,7.8091707,5.844017,5.051782,4.1189346,3.234101,2.4830213,1.862266,1.8005334,3.5804894,4.715683,4.256118,2.7916842,2.9391565,2.1332035,1.5707511,1.9274281,3.357566,3.2581081,2.4830213,3.3815732,5.7377,6.773435,6.138962,5.192395,3.858286,2.4624438,1.7559488,2.6956558,2.2326615,2.7642474,4.0057583,3.0077481,2.0920484,3.8102717,4.530485,3.340418,2.0440342,1.4472859,1.5913286,2.1332035,2.5790498,2.2738166,1.9308578,1.5090185,1.5570327,2.3321195,3.782835,3.0900583,3.2889743,3.8034124,4.396731,5.2026844,5.751418,5.295283,4.280125,3.5050385,4.0880685,5.284994,6.992929,8.549961,9.071259,7.4456344,4.870014,4.383013,4.962613,5.802862,6.3035817,6.667118,6.7494283,6.7802944,6.667118,5.9983487,4.605936,5.1992545,5.9400454,6.0806584,5.9812007,5.919468,6.0532217,6.210983,6.2658563,6.118384,5.6176643,5.363875,5.079219,5.0346346,6.0737996,7.781734,9.14328,8.800322,7.284444,7.0032177,8.004657,8.06296,7.1541195,6.111525,6.636252,9.407358,9.716022,8.766026,8.98209,14.023583,13.509145,13.766364,11.746337,7.936065,6.3481665,8.594546,8.64256,8.128122,7.8846216,7.936065,10.216741,9.431366,7.191845,5.693115,7.706283,7.8537555,8.2653055,8.014946,7.3530354,7.720001,7.0375133,6.8557453,5.672538,4.0057583,4.4104495,5.130663,4.513337,4.647091,5.442755,4.6402316,2.417859,1.7971039,1.845118,1.7833855,0.9774324,0.85396725,1.0082988,1.0940384,0.9877212,0.7922347,0.7922347,1.0220171,1.039165,0.7956643,0.6241849,1.2586586,1.0700313,0.65505123,0.39783216,0.45613512,0.5178677,0.42526886,0.28465575,0.16119061,0.07545093,0.09945804,0.16119061,0.15090185,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.09602845,0.116605975,0.1097468,0.106317215,0.16804978,0.082310095,0.041155048,0.12689474,0.30866286,0.4424168,0.23664154,0.20234565,0.22635277,0.24350071,0.24350071,0.12346515,0.274367,0.432128,0.48357183,0.47328308,0.25378948,0.28122616,0.35324752,0.4046913,0.5041494,0.6001778,0.5418748,0.53844523,0.5418748,0.26064864,0.22292319,0.22292319,0.26407823,0.3806842,0.6241849,0.77165717,0.7339317,0.6859175,0.65848076,0.548734,0.548734,0.48357183,0.5041494,0.58988905,0.5658819,0.84367853,0.88826317,0.8745448,0.89512235,0.9294182,1.138623,1.2175035,1.0460242,0.7099246,0.5041494,0.7956643,0.9534253,1.0117283,0.96714365,0.7476501,0.8711152,0.97400284,1.1694894,1.3855534,1.371835,0.9842916,0.84024894,0.9842916,1.3238207,1.6187652,1.4335675,1.7079345,1.587899,0.99801,0.65505123,0.70649505,1.1283343,1.3478279,1.1866373,0.8711152,0.5761707,2.3629858,6.0737996,8.076678,1.2655178,1.1694894,2.5070283,4.046913,4.40702,2.0749004,1.2346514,1.4335675,1.8416885,2.2292318,2.976882,2.609916,2.784825,3.6868064,4.4584637,3.1895163,1.138623,2.1915064,5.9331865,9.400499,7.0786686,4.0537724,4.3933015,5.223262,5.346727,5.2506986,6.7391396,9.767465,12.593445,14.88441,17.717249,19.853882,18.471758,15.158776,11.547421,9.338767,13.841815,13.797231,11.948683,10.487679,11.063849,9.719451,10.034973,10.844356,11.022695,9.462232,7.349606,7.205563,8.224151,8.152129,3.2821152,2.4658735,2.3595562,3.0729103,5.4736214,11.183885,9.47595,6.8969,8.790032,15.645778,23.11542,17.37772,18.71183,23.009102,26.35981,25.039417,24.672453,24.4461,22.100262,18.71526,18.677534,17.017612,17.892159,20.906765,23.02625,18.571217,21.976797,23.166862,23.338343,23.880217,26.380386,26.503853,22.974806,20.539799,20.430052,20.37175,16.671225,16.259674,17.597214,19.548649,21.393766,26.469557,29.542467,30.770258,30.77369,30.639935,28.465576,28.719366,29.964306,30.1838,26.77822,24.336353,22.69358,22.961088,22.94394,17.1205,14.826107,10.679735,7.298162,5.394741,3.782835,3.210094,3.093488,2.7470996,2.369845,3.0523329,2.8808534,3.0317552,3.5016088,4.7259717,7.582818,10.844356,10.823778,10.902658,12.689473,16.019604,15.8138275,13.838386,13.248496,14.452282,15.138199,12.195613,8.906639,7.531374,8.580828,10.803201,11.705182,11.190743,9.506817,7.5553813,6.8969,10.206452,8.927217,6.495639,4.7774153,4.0434837,4.1292233,3.2546785,2.4487255,2.1332035,2.1194851,1.6804979,1.9754424,2.6579304,3.3026927,3.3884325,2.7162333,3.1895163,4.372724,4.8014226,1.9685832,4.9351764,5.857735,4.9488945,3.2958336,2.867135,4.6265135,4.664239,4.033195,3.7759757,4.897451,8.073249,7.6651278,7.0306544,6.9380555,5.56965,11.039842,11.149589,8.704293,6.0086374,4.897451,5.0929375,5.2781353,4.4241676,2.4830213,0.39783216,1.4335675,1.9514352,1.7662375,1.0082988,0.09259886,0.09259886,0.072021335,0.041155048,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.006859175,0.017147938,0.030866288,0.017147938,0.01371835,0.01371835,0.01371835,0.0,0.01371835,0.024007112,0.024007112,0.01371835,0.01371835,0.041155048,0.037725464,0.024007112,0.01371835,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.044584636,0.044584636,0.0548734,0.08573969,0.106317215,0.044584636,0.034295876,0.030866288,0.024007112,0.017147938,0.030866288,0.07888051,0.12003556,0.15090185,0.16804978,0.16804978,0.106317215,0.0548734,0.024007112,0.01371835,0.0,0.19548649,0.40126175,0.45956472,0.59674823,1.4027013,1.0254467,0.41840968,0.044584636,0.037725464,0.18176813,0.14747226,0.20234565,0.4081209,0.6756287,0.7476501,0.6859175,0.78194594,0.65848076,0.30523327,0.061732575,0.01371835,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.037725464,0.18176813,3.1483612,2.9391565,1.6942163,0.6310441,0.044584636,0.082310095,0.89855194,1.6667795,1.8279701,1.0837497,1.1934965,1.4232788,1.4267083,1.2517995,1.313532,1.6290541,2.5413244,4.629943,7.233,8.453933,8.796892,15.271953,18.420315,16.355703,14.754086,15.584045,18.355152,22.426073,26.164322,26.946268,30.060333,32.807434,34.155262,33.58252,31.065203,28.503302,27.495003,27.76937,27.93742,25.495554,24.826784,23.34863,21.390337,18.948471,15.700651,12.490558,10.233889,8.669997,7.4936485,6.3310184,5.8817425,5.0346346,3.5702004,2.0337453,1.7388009,1.762808,1.5055889,1.138623,0.823101,0.70306545,0.6276145,0.51100856,0.45956472,0.48357183,0.47328308,0.33952916,0.20577525,0.12003556,0.07888051,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,6.543653,8.06296,11.255906,14.13333,15.230798,13.594885,16.770683,24.624437,34.614826,48.079388,70.25853,59.54107,40.801804,32.93433,39.99585,51.186592,33.788296,27.714497,24.374079,20.080235,16.050468,12.483699,11.331357,11.2593355,10.912948,8.8929205,8.460793,8.848335,11.989838,19.579515,33.08866,41.474003,36.473663,27.045727,19.325726,16.592344,14.5414505,11.746337,9.743458,8.827758,8.05953,8.255017,12.5145645,13.227919,9.23245,5.785714,10.734609,11.633161,11.780633,12.428825,12.768354,15.484588,18.495766,21.626978,25.097721,29.51503,34.196415,40.434837,43.42201,41.30595,35.18414,25.725336,17.141079,11.080997,8.052671,7.4181976,8.203573,8.114404,7.267296,5.967482,4.695105,4.0880685,3.532475,3.1483612,2.8259802,2.253239,1.7799559,2.4384367,2.9734523,2.7916842,1.961724,2.1674993,1.8073926,1.6359133,2.1434922,3.5530527,1.961724,1.6839274,1.8416885,2.1194851,2.7470996,2.7368107,2.4658735,1.8691251,1.6873571,3.5016088,2.369845,2.527606,2.8637056,3.07634,3.6765177,3.2992632,3.1689389,2.6853669,2.0097382,2.0817597,2.07833,2.4212887,2.8225505,3.100347,3.1655092,3.117495,3.093488,2.9048605,2.5893385,2.4418662,1.920569,2.16064,2.9048605,4.029765,5.521636,4.3109913,3.642222,3.4055803,3.6387923,4.5167665,5.3501563,6.046363,6.279575,5.672538,3.782835,3.2409601,5.3398676,6.5162163,6.0978065,6.3138704,5.099797,4.1635194,3.5393343,3.210094,3.1037767,3.683377,4.846007,6.5367937,7.891481,7.226141,6.217842,5.453044,4.722542,4.3658648,5.2644167,7.654839,8.014946,7.2535777,6.245279,5.8165803,5.456474,6.0223556,6.392751,6.0326443,4.99005,5.8234396,5.878313,5.360445,5.188966,7.0032177,11.249047,14.225929,12.315649,7.822889,8.958082,12.583157,13.282792,11.413667,8.3922,6.677407,8.2310095,10.113853,10.045261,8.577398,9.105555,12.0138445,11.129011,8.748878,6.7974424,6.8385973,6.684266,6.944915,7.085528,7.0135064,7.085528,7.5931067,7.7714453,6.8043017,5.31929,5.360445,5.0174866,4.0537724,4.033195,4.8494368,4.7499785,3.0248961,2.6853669,2.784825,2.5413244,1.3066728,0.94999576,0.939707,0.96371406,0.91912943,0.939707,0.86082643,1.0048691,1.1592005,1.1763484,0.96714365,1.2106444,1.1077567,0.94999576,0.90541106,0.9945804,0.607037,0.40126175,0.26750782,0.16462019,0.08916927,0.044584636,0.037725464,0.030866288,0.01371835,0.0,0.0,0.0,0.01371835,0.030866288,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.041155048,0.034295876,0.07545093,0.17147937,0.25378948,0.17833854,0.16804978,0.18176813,0.1920569,0.20920484,0.09945804,0.09259886,0.16119061,0.2503599,0.26750782,0.06859175,0.06859175,0.1371835,0.20920484,0.31552204,0.15433143,0.15090185,0.18519773,0.20920484,0.2469303,0.3841138,0.490431,0.5418748,0.5178677,0.39440256,0.31895164,0.30866286,0.37039545,0.490431,0.6379033,0.64819205,0.5624523,0.490431,0.4355576,0.31895164,0.30866286,0.32238123,0.38754338,0.48014224,0.5041494,0.5796003,0.5796003,0.6241849,0.72707254,0.77165717,0.7442205,0.72364295,0.6962063,0.6790583,0.6859175,0.85396725,0.78537554,0.764798,0.83681935,0.8196714,0.84367853,0.88826317,0.980862,1.0597426,0.9568549,1.0254467,0.9774324,1.0460242,1.2895249,1.5913286,1.7422304,1.821111,1.6839274,1.5227368,1.8656956,1.5913286,1.4747226,1.4232788,1.2209331,0.5041494,0.8162418,4.5167665,8.258447,8.625413,2.1469216,1.3546871,1.8313997,2.568761,2.6236343,1.1111864,0.9328478,2.170929,3.625074,4.602506,4.928317,5.0586414,4.4516044,4.122364,4.040054,3.0900583,3.7348208,5.439326,5.9297566,4.880303,3.9200184,4.9248877,6.800872,7.3873315,6.1629686,4.249259,4.6745276,5.778855,7.0615206,8.477941,10.439664,12.068718,11.910957,11.447963,11.461681,12.034423,16.023033,15.4742985,13.255356,12.274493,15.494876,18.416885,19.404606,20.443771,21.795029,21.959648,18.842154,20.433481,21.884197,20.443771,15.436573,11.770344,9.414218,8.453933,8.827758,10.343636,7.1884155,6.0875177,7.4799304,10.477389,12.850664,13.197053,19.006773,25.337791,28.479294,25.979126,22.264881,18.708399,17.549198,17.700102,14.733508,19.500635,21.592682,22.587263,22.8582,21.596113,23.098272,23.770472,23.060547,21.170843,19.03421,21.273731,21.849901,22.011093,21.098822,16.53747,15.642348,17.748116,21.386908,24.957108,26.702768,28.060884,28.153484,29.189219,31.150944,31.785418,27.865398,27.309805,26.675331,24.675882,22.18943,22.474087,21.246294,19.678972,18.44775,17.741257,18.818146,14.592895,9.993818,7.442205,6.848886,6.0978065,6.632822,6.852316,6.715132,7.750868,5.8337283,4.3521466,3.8925817,5.0655007,8.498518,11.38623,12.579727,12.8197975,12.878101,13.543441,13.540011,12.535142,10.988399,9.8429165,10.487679,10.912948,9.914937,9.6988735,10.72089,11.681175,12.274493,13.121602,12.79922,11.832077,12.696333,13.766364,12.185325,10.103564,7.936065,4.3624353,3.5187566,3.2032347,3.3198407,3.508468,3.1449318,2.0920484,2.2155135,2.4555845,2.6167753,3.3884325,4.180667,4.434457,5.3090014,6.276145,5.0929375,5.4633327,5.885172,5.641671,5.271276,6.543653,6.893471,6.543653,5.5593615,4.671098,5.2781353,7.191845,6.924337,6.2144127,6.0635104,6.7185616,9.283894,9.770895,8.378482,6.138962,4.911169,6.169828,5.2747054,3.0146074,0.82996017,0.8128122,1.371835,1.8039631,1.7490896,1.1866373,0.45613512,0.22292319,0.072021335,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.006859175,0.006859175,0.0,0.0034295875,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.020577524,0.024007112,0.024007112,0.017147938,0.017147938,0.024007112,0.0274367,0.024007112,0.01371835,0.01371835,0.024007112,0.030866288,0.024007112,0.01371835,0.030866288,0.024007112,0.017147938,0.01371835,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.024007112,0.0034295875,0.0,0.006859175,0.017147938,0.020577524,0.020577524,0.017147938,0.020577524,0.030866288,0.010288762,0.006859175,0.006859175,0.010288762,0.017147938,0.017147938,0.0274367,0.044584636,0.048014224,0.044584636,0.044584636,0.034295876,0.05144381,0.048014224,0.01371835,0.0,0.06859175,0.38754338,0.5212973,0.42869842,0.4629943,0.28122616,0.1097468,0.037725464,0.072021335,0.15776102,0.14061308,0.45613512,0.78194594,0.86082643,0.5144381,0.38754338,0.48014224,0.53158605,0.4115505,0.1097468,0.020577524,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.09945804,0.5007198,1.903421,1.8656956,1.2758065,0.6893471,0.33952916,0.15090185,0.432128,0.7956643,0.99801,0.9362774,1.3203912,1.4644338,1.4267083,1.4610043,2.020027,2.8054025,2.877424,3.5530527,5.346727,7.963502,9.829198,12.644889,14.143619,14.671775,17.185663,20.817596,22.85477,25.728765,29.645353,32.574223,35.25616,36.950375,37.207596,36.24388,34.961216,31.528198,29.401854,29.583622,30.705097,29.0246,26.555296,24.902235,23.163433,20.7833,17.545769,14.225929,12.154458,10.844356,9.884071,8.920357,6.9552035,5.576509,4.2286816,2.9151495,2.201795,1.6530612,1.3581166,1.1249046,0.8711152,0.65162164,0.6173257,0.59674823,0.59331864,0.59331864,0.5693115,0.4355576,0.29494452,0.17490897,0.09259886,0.0548734,0.034295876,0.010288762,0.0,0.0,0.0,5.329579,7.870903,9.301042,8.889491,7.5690994,7.905199,11.760056,15.885849,19.46291,22.834194,27.505291,25.481834,26.977135,43.5832,69.96701,83.84998,48.55953,35.58883,29.857988,23.873358,17.717249,12.826657,11.170166,10.525404,9.3936405,7.006647,8.1384115,10.220171,17.315987,33.32873,61.98979,60.25099,44.31027,28.753662,20.488356,18.71183,14.164196,11.190743,10.31277,10.412228,8.759167,8.889491,11.273054,11.365653,9.386781,10.30591,16.0539,14.582606,13.509145,15.515453,18.355152,16.187653,14.911846,15.4914465,17.37772,18.526632,21.386908,29.662502,36.398212,38.22275,35.34533,28.626766,20.673553,14.201921,10.316199,8.501947,7.997798,7.010077,5.7891436,4.6402316,3.9165888,3.806842,3.4604537,3.1586502,2.9391565,2.5961976,2.1983654,2.318401,2.4555845,2.4624438,2.551613,2.369845,1.6804979,1.2895249,1.4781522,2.0268862,1.3924125,1.5433143,1.5536032,1.2998136,1.4369972,1.9925903,1.5844694,1.1832076,1.5330256,3.1312134,6.193835,9.873782,9.458802,5.6313825,4.448175,3.9337368,3.018037,2.9803114,4.0880685,5.579939,5.1169443,4.5030484,3.7108135,3.1209247,3.5050385,3.5804894,3.5153272,3.234101,2.7951138,2.369845,2.0337453,2.2841053,2.9665933,3.7691166,4.190956,3.8308492,3.9131594,3.724532,3.532475,4.5853586,4.773986,4.5613513,4.245829,3.9611735,3.6936657,2.952875,4.8322887,5.960623,5.597087,5.6039457,4.372724,3.9851806,4.3658648,5.3158607,6.509357,5.8165803,5.4496145,6.543653,8.210432,7.5279446,6.636252,5.8543057,5.0483527,4.3590055,4.2081037,6.9689217,8.766026,9.259886,8.385342,6.385892,5.586798,6.9723516,8.279024,8.323608,6.992929,7.4353456,7.8949103,7.3050213,6.293293,7.1678376,12.46998,16.29397,14.500296,9.047252,7.98408,12.864383,14.493437,13.323947,10.487679,7.7748747,9.287323,11.094715,10.696883,8.447074,7.548522,8.995808,8.923786,8.303031,7.610255,6.8043017,6.5059276,6.893471,6.9037595,6.475061,6.5333643,7.582818,8.028665,7.4284863,6.2144127,5.6828265,5.5319247,4.6916757,4.266407,4.5956473,5.2609873,4.057202,3.5976372,3.5187566,3.2443898,2.020027,1.3786942,1.4369972,1.6221949,1.5364552,0.9568549,1.1523414,1.2483698,1.4095604,1.611906,1.6564908,1.4610043,1.2517995,1.2963841,1.4575747,1.2106444,0.6173257,0.3841138,0.25378948,0.12346515,0.072021335,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.006859175,0.044584636,0.12346515,0.17490897,0.13032432,0.12689474,0.12689474,0.1097468,0.061732575,0.048014224,0.05144381,0.106317215,0.18862732,0.22978236,0.07545093,0.020577524,0.048014224,0.1371835,0.29151493,0.2194936,0.20577525,0.18862732,0.16462019,0.20920484,0.33609957,0.38754338,0.4664239,0.5212973,0.36353627,0.30866286,0.36353627,0.44927597,0.5178677,0.5590228,0.5693115,0.45613512,0.32924038,0.25378948,0.2503599,0.274367,0.31895164,0.36353627,0.39440256,0.38754338,0.4115505,0.4698535,0.5178677,0.52472687,0.48357183,0.47328308,0.4629943,0.47671264,0.5041494,0.5212973,0.6207553,0.59674823,0.6207553,0.7305021,0.8471081,0.84024894,0.83338976,0.864256,0.8745448,0.71678376,0.7682276,0.82996017,0.9534253,1.1729189,1.4850113,1.8931323,1.8416885,1.6359133,1.6530612,2.3492675,1.7696671,1.3546871,1.039165,0.7476501,0.3841138,0.8471081,3.6010668,5.5250654,4.880303,1.313532,0.764798,0.94999576,1.313532,1.3958421,0.8505377,0.85396725,1.5604624,2.5790498,3.673088,4.756838,4.9351764,3.9611735,3.0077481,2.5824795,2.534465,4.791134,6.1801167,5.2747054,2.9974594,2.6167753,4.2046742,6.392751,7.222711,6.121814,3.9063,3.5016088,3.7279615,4.2286816,4.8837323,5.802862,6.8557453,7.373613,7.891481,8.663138,9.661148,12.356804,12.860953,12.6929035,12.713481,13.13189,13.951562,14.373401,16.304258,19.654966,22.347193,20.663265,19.239986,18.317427,17.604073,16.29054,12.397959,9.325048,8.591117,9.47595,8.995808,7.208993,7.7542973,8.827758,9.853205,11.502836,11.921246,16.235666,22.11398,26.054577,23.403505,20.930773,16.815268,15.223939,16.077906,15.066177,18.883308,21.290878,22.11055,21.77788,21.318316,21.987085,20.985645,19.013634,16.839275,15.29253,17.2131,19.819586,21.486366,21.211998,18.62609,20.03565,23.478956,26.836521,29.062325,30.18037,32.615376,33.726562,33.781437,32.526207,29.189219,26.781649,27.056015,27.237783,26.380386,25.382378,24.94682,23.238884,21.61326,20.567236,19.720127,20.412905,17.19938,13.262215,10.357354,8.776315,8.364764,8.525954,8.666568,8.690575,9.009526,6.9517736,5.453044,5.9126086,8.433355,11.80464,12.651748,12.730629,12.415107,12.22305,12.823228,13.810948,11.543991,9.925226,10.443094,12.161317,12.061859,11.146159,10.744898,11.207891,11.928105,13.423406,14.956431,15.316538,14.520873,13.824667,13.149038,12.312219,11.653738,10.600855,7.671987,6.444195,6.0806584,6.7357097,7.699424,7.394191,5.645101,4.5510626,3.57363,2.9803114,3.8548563,4.1943855,4.479041,4.547633,4.7842746,6.094377,4.3178506,4.280125,5.638242,7.531374,8.570539,7.486789,7.4799304,7.4456344,7.034084,6.6533995,8.443645,10.933525,12.199042,11.907528,11.324498,10.714031,10.240748,9.259886,7.7714453,6.4407654,6.8626046,5.4599032,3.1209247,1.2586586,1.8039631,1.5776103,1.5261664,1.3203912,0.89855194,0.44927597,0.19891608,0.061732575,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.006859175,0.017147938,0.024007112,0.020577524,0.010288762,0.010288762,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.010288762,0.010288762,0.01371835,0.006859175,0.01371835,0.030866288,0.034295876,0.0274367,0.01371835,0.01371835,0.024007112,0.030866288,0.030866288,0.034295876,0.0274367,0.037725464,0.044584636,0.034295876,0.01371835,0.020577524,0.017147938,0.010288762,0.082310095,0.39440256,0.89169276,0.42869842,0.024007112,0.010288762,0.020577524,0.010288762,0.0034295875,0.006859175,0.01371835,0.01371835,0.01371835,0.010288762,0.010288762,0.01371835,0.010288762,0.0034295875,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.010288762,0.010288762,0.006859175,0.01371835,0.01371835,0.024007112,0.020577524,0.006859175,0.010288762,0.05144381,0.24350071,0.32581082,0.24350071,0.1371835,0.0548734,0.85739684,1.1111864,0.5693115,0.17833854,0.08573969,0.31552204,0.59331864,0.6859175,0.39440256,0.24007112,0.32581082,0.42526886,0.4081209,0.22292319,0.05144381,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.19548649,0.97400284,1.3649758,1.313532,1.2449403,1.2483698,1.08032,0.4629943,0.25378948,0.31895164,0.4938606,0.58988905,0.980862,1.6496316,2.0406046,2.0646117,2.0886188,2.411,2.4418662,2.952875,4.695105,8.354475,8.879202,9.122703,11.266195,15.820687,21.644127,24.075705,24.329493,26.301506,30.59878,34.556522,39.608307,42.07075,42.122192,40.753788,39.769497,38.281055,36.42222,35.386482,34.628544,31.867727,28.67135,26.610168,24.998262,23.005672,19.661825,16.86671,14.712931,13.2862215,12.517994,12.195613,10.017825,7.699424,5.5593615,3.8960114,2.9700227,2.2360911,1.6770682,1.2895249,1.0460242,0.89855194,0.7990939,0.7442205,0.7339317,0.7339317,0.6859175,0.52472687,0.34981793,0.20920484,0.116605975,0.08916927,0.048014224,0.0274367,0.01371835,0.010288762,0.010288762,5.5730796,7.7268605,7.291303,5.7136927,4.629943,5.861165,8.152129,10.847785,12.984418,13.72178,12.360233,13.742357,30.739393,65.25476,99.746124,97.24595,51.131718,33.92891,27.296087,21.500084,15.419425,11.670886,10.13786,9.410788,8.567109,7.14726,8.498518,11.348505,25.19718,55.967438,106.02913,81.655045,51.995975,30.818274,22.148275,20.244854,14.760944,13.433694,13.481709,12.538571,8.64942,9.177576,10.034973,10.652299,12.082437,16.993607,18.639809,14.112752,12.161317,15.940722,23.005672,16.383139,11.080997,11.749766,16.914726,18.972477,15.824117,21.407484,28.722795,33.513927,34.24786,31.116648,25.783638,20.152256,15.354263,11.7257595,9.424506,7.191845,5.3227196,4.0229063,3.415869,3.426158,3.192946,2.952875,2.7813954,2.6167753,2.2909644,2.1194851,2.0508933,2.1057668,2.369845,2.1812177,1.5090185,0.9877212,0.8265306,0.805953,0.97400284,1.3341095,1.8656956,2.16064,1.4198492,2.1846473,1.8862731,1.5707511,1.7388009,2.3389788,7.1712675,10.628291,9.832627,6.0154963,4.5167665,4.1326528,3.426158,3.590778,4.7191124,5.8062916,5.0243454,4.434457,4.0846386,3.8685746,3.5187566,3.590778,3.666229,3.5461934,3.234101,2.9563043,2.8122618,3.059192,3.4021509,3.4398763,2.6750782,2.8808534,3.2066643,3.450165,3.7622573,4.6608095,4.5099077,4.1189346,3.6147852,3.3198407,3.7348208,3.210094,4.1772375,4.636802,4.32128,4.698535,4.201245,4.1600895,4.880303,6.125243,7.1198235,6.385892,5.7239814,6.090947,6.9654922,6.3378778,6.200694,6.4887795,6.550512,5.960623,4.5270553,6.756287,9.112414,10.425946,10.175586,8.501947,7.174697,8.189855,9.537683,10.124143,9.760606,9.541112,10.213311,9.921797,8.615124,8.011517,12.435684,15.951012,15.004445,10.64201,8.532814,13.2690735,15.0250225,14.651197,12.734058,9.599416,9.949233,10.357354,9.740028,8.001227,6.0532217,6.324159,6.711703,7.421627,7.8434668,6.560801,6.169828,6.8214493,7.006647,6.3790326,5.751418,6.691125,7.459353,7.226141,6.138962,5.3330083,5.2918534,4.647091,3.981751,3.8445675,4.7602673,4.554492,4.461893,4.3624353,3.998899,2.983741,1.8382589,1.8142518,2.277246,2.4247184,1.2758065,1.3203912,1.3238207,1.5227368,1.9171394,2.2806756,1.7490896,1.3649758,1.2483698,1.2346514,0.881404,0.47328308,0.33952916,0.2777966,0.20234565,0.14747226,0.10288762,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.030866288,0.037725464,0.05144381,0.07545093,0.06516216,0.048014224,0.044584636,0.06859175,0.08916927,0.037725464,0.044584636,0.058302987,0.08916927,0.13375391,0.16804978,0.08573969,0.037725464,0.044584636,0.1097468,0.20920484,0.22292319,0.22978236,0.20577525,0.16462019,0.18519773,0.25721905,0.31895164,0.4081209,0.4424168,0.20920484,0.1920569,0.32924038,0.4389872,0.4424168,0.34981793,0.38754338,0.32924038,0.2503599,0.20577525,0.22635277,0.22978236,0.28122616,0.31895164,0.31552204,0.26407823,0.30866286,0.3806842,0.4046913,0.37039545,0.32581082,0.36696586,0.4046913,0.40126175,0.3566771,0.31895164,0.38754338,0.42869842,0.47671264,0.5590228,0.6893471,0.6859175,0.7133542,0.7922347,0.83338976,0.65162164,0.65162164,0.83681935,1.0117283,1.1249046,1.2346514,1.7250825,1.6221949,1.3581166,1.3169615,1.8382589,1.5055889,1.1660597,0.7990939,0.4938606,0.45270553,0.6824879,1.7525192,2.1812177,1.5673214,0.58645946,0.5555932,0.6276145,0.72364295,0.77165717,0.6927767,0.8505377,0.97400284,1.3684053,2.1503513,3.2443898,3.3850029,2.8534167,2.1915064,1.920569,2.5241764,4.3795834,5.2266912,4.2766957,2.318401,1.7490896,2.5173173,3.865145,4.705394,4.48933,3.192946,2.5961976,2.633923,2.7470996,2.8156912,3.1209247,3.9337368,4.5922174,5.0655007,5.6485305,6.9654922,8.2310095,9.80519,10.748327,10.4533825,8.632272,8.4093485,9.537683,12.452832,16.647217,20.687271,21.997374,18.427174,15.028452,14.030442,14.850114,12.247057,10.319629,10.714031,12.257345,10.943813,10.117283,9.585697,8.851766,8.666568,11.032983,12.459691,14.654627,19.21255,23.989964,23.091412,22.402065,18.78042,16.221949,15.563468,14.476289,16.016174,19.068506,20.841602,20.742146,20.399187,20.683842,19.315437,17.53891,15.806969,13.783512,14.832966,18.224829,20.824455,21.647556,21.839613,24.233465,27.227495,29.419,30.50961,31.298416,33.5688,34.32331,32.924038,29.110338,23.019392,23.44809,25.228045,27.035439,27.982004,27.628757,25.670462,23.866499,23.10856,23.170294,22.703869,22.450079,19.973917,16.897577,14.291091,12.665466,10.518545,9.163857,9.517105,10.789482,10.484249,7.9017696,6.101236,7.2947326,10.964391,13.872682,13.310229,12.240198,11.063849,10.494537,11.585147,12.620882,11.681175,11.873232,13.629181,14.743796,13.104454,11.543991,10.882081,11.451392,13.118172,15.892709,16.750105,16.530611,15.971589,15.717799,14.579176,13.210771,12.466551,12.0138445,10.319629,10.864933,9.6988735,9.547972,10.731179,11.173596,9.373062,7.380472,7.0958166,8.028665,7.267296,5.7582774,5.4496145,5.6999745,6.2692857,7.3255987,4.40359,3.7142432,5.586798,8.601405,9.575408,8.995808,10.182446,10.964391,10.425946,8.886061,11.05356,14.987297,17.785841,18.235117,16.835844,13.368532,11.900668,10.988399,9.956093,8.89635,8.244728,5.5662203,3.1380725,2.085189,2.369845,1.5330256,1.0666018,0.7956643,0.5796003,0.32581082,0.1371835,0.041155048,0.006859175,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.010288762,0.017147938,0.030866288,0.030866288,0.024007112,0.020577524,0.017147938,0.006859175,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.006859175,0.01371835,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.017147938,0.030866288,0.037725464,0.0274367,0.01371835,0.024007112,0.037725464,0.041155048,0.037725464,0.044584636,0.037725464,0.041155048,0.041155048,0.034295876,0.01371835,0.020577524,0.024007112,0.06516216,0.3018037,1.0220171,2.4624438,1.8142518,0.7373613,0.1097468,0.020577524,0.010288762,0.010288762,0.017147938,0.024007112,0.0274367,0.024007112,0.017147938,0.01371835,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0034295875,0.010288762,0.048014224,0.10288762,0.12003556,0.09602845,0.044584636,0.020577524,0.85739684,1.1214751,0.5693115,0.16119061,0.0548734,0.14061308,0.34295875,0.5144381,0.45613512,0.34981793,0.30866286,0.28122616,0.24350071,0.17490897,0.041155048,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.21263443,0.9602845,0.9842916,0.97400284,1.2483698,1.7730967,2.1674993,1.0563129,0.5007198,0.34981793,0.40126175,0.39440256,0.83681935,1.7353712,2.301253,2.469303,2.9048605,2.2395205,2.2052248,2.9494452,4.681387,7.689135,7.346176,8.23444,12.041282,18.056778,23.177153,22.474087,23.712168,27.92027,34.227283,39.896393,43.349987,45.22254,45.418026,44.608643,44.24511,44.73211,43.66551,41.48086,38.438816,34.60111,31.517908,28.904564,26.743923,24.754763,22.395206,19.552078,17.29198,15.858413,15.498305,16.45516,15.230798,12.061859,8.440215,5.501058,4.0263357,3.234101,2.4212887,1.821111,1.4850113,1.2860953,1.1934965,1.08032,0.9842916,0.90884066,0.84024894,0.6790583,0.4938606,0.32581082,0.20577525,0.16119061,0.106317215,0.072021335,0.041155048,0.020577524,0.01371835,6.217842,7.3084507,5.919468,4.650521,4.5682106,5.192395,5.4633327,6.8797526,8.357904,9.22902,9.235879,14.997586,38.936108,75.944786,102.877335,78.589,37.608856,22.95423,17.995045,14.195063,11.091286,10.947243,10.532263,9.908078,9.2153015,8.656279,9.030104,15.385129,43.63807,95.308235,157.52782,102.41777,58.474464,32.776566,23.68473,20.800447,16.21166,18.12537,18.598652,14.654627,8.2653055,9.6645775,10.799771,12.504276,15.837835,22.100262,18.979338,11.869802,9.31133,15.021593,27.92027,20.11453,11.97269,13.88983,23.427511,25.306927,16.091625,15.741806,20.382038,26.373528,30.296976,30.252392,28.791388,25.488693,20.78673,15.9921665,12.21619,8.930646,6.3824625,4.6127954,3.4707425,3.1072063,2.976882,2.8945718,2.7470996,2.5001693,2.0886188,1.7216529,1.605047,1.6839274,1.6324836,1.5741806,1.3581166,0.9842916,0.6036074,0.50757897,0.5693115,0.980862,2.0131679,2.8568463,1.6221949,2.194936,2.253239,2.0886188,2.318401,3.8685746,5.2918534,4.170378,3.2135234,3.3061223,3.532475,3.6936657,3.6387923,3.2992632,2.784825,2.3767042,2.3904223,2.8499873,4.0606318,5.038064,3.5016088,3.5530527,3.9337368,3.9508848,3.566771,3.3815732,3.4535947,3.5770597,3.4638834,2.901431,1.7559488,1.4404267,1.3546871,2.3046827,3.9131594,4.619654,4.6265135,4.705394,4.2835546,3.4981792,3.1860867,3.542764,3.8308492,3.4981792,3.0420442,3.974892,4.3041325,3.9131594,3.8548563,4.170378,3.8891523,4.787704,5.188966,5.3913116,5.5490727,5.6999745,5.8543057,6.6396813,7.4044795,7.531374,6.420188,8.207003,9.462232,10.199594,10.645439,11.279913,9.554831,8.704293,8.748878,9.619993,11.153018,10.13786,10.587136,11.502836,11.955542,11.101575,13.327377,15.920145,15.134769,11.314209,8.903209,12.0138445,13.197053,13.694343,13.416546,10.978109,9.609704,9.119273,9.019815,8.570539,6.7700057,6.3447366,6.1732574,6.90033,7.6857057,6.23156,5.7754254,6.615674,7.3873315,7.099246,5.15467,5.7582774,6.632822,6.625963,5.778855,5.3398676,4.729401,4.1120753,3.5359046,3.216953,3.5187566,4.033195,4.6848164,4.9591837,4.605936,3.642222,2.1503513,1.9411465,2.5173173,2.9631636,1.9685832,1.3546871,1.1454822,1.3649758,1.8862731,2.4075704,1.8656956,1.4369972,1.0357354,0.65848076,0.4046913,0.28465575,0.274367,0.31209245,0.33609957,0.24350071,0.18862732,0.116605975,0.048014224,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.048014224,0.06859175,0.06859175,0.048014224,0.0,0.0,0.006859175,0.048014224,0.09259886,0.072021335,0.0548734,0.06516216,0.082310095,0.09602845,0.09602845,0.072021335,0.058302987,0.061732575,0.06516216,0.048014224,0.106317215,0.15433143,0.17833854,0.16804978,0.116605975,0.13375391,0.274367,0.36353627,0.30523327,0.08916927,0.06516216,0.20920484,0.32238123,0.30866286,0.15776102,0.17490897,0.20234565,0.22978236,0.22978236,0.18176813,0.14061308,0.23321195,0.30523327,0.28808534,0.20234565,0.23664154,0.25378948,0.26064864,0.2777966,0.32581082,0.39097297,0.45613512,0.41498008,0.29151493,0.26064864,0.30866286,0.32924038,0.33266997,0.33952916,0.40126175,0.41840968,0.5178677,0.6859175,0.805953,0.6790583,0.77165717,1.0460242,1.1832076,1.0837497,0.8848336,1.2620882,1.1934965,0.9534253,0.78194594,0.89512235,1.1694894,1.1180456,0.88826317,0.65162164,0.6001778,0.45613512,0.42183927,0.4355576,0.47328308,0.5418748,0.8025235,0.75450927,0.64476246,0.5693115,0.47328308,0.8265306,0.922559,1.1111864,1.430138,1.5913286,1.786815,2.0680413,2.1194851,2.1126258,2.7162333,3.0351849,3.5633414,3.1106358,1.8073926,1.0940384,1.5673214,1.4575747,1.6564908,2.177788,2.177788,1.99602,2.1263442,2.0097382,1.7353712,2.0234566,2.8054025,3.2546785,3.6799474,4.513337,6.327589,6.1492505,7.8674736,8.275595,6.8111606,5.552502,6.574519,9.115844,12.188754,15.505165,19.473198,22.799898,20.29287,16.756964,14.692352,14.291091,13.203912,13.279363,14.38369,15.319967,13.828096,13.275933,10.419086,7.7131424,6.8043017,8.519095,11.7257595,13.738928,17.487467,22.240875,23.623,24.185452,22.072824,19.435472,16.80498,13.104454,14.249936,17.346853,19.099373,18.890167,18.763273,19.648108,19.270851,18.4649,17.20281,14.572317,14.195063,16.750105,19.572655,21.462358,22.676432,24.487255,26.147175,28.081463,30.067194,31.226395,30.022608,28.290667,26.082012,23.19773,19.185112,21.983656,23.845922,25.571005,26.719915,25.636166,25.550426,25.046278,24.583282,24.658733,25.800787,25.18346,23.057117,20.773012,19.11652,18.296848,12.576297,9.3079,10.038403,12.922686,12.754636,9.695444,7.085528,7.7028537,11.005547,13.13189,12.586586,11.540562,9.956093,8.766026,9.89436,10.902658,13.670336,15.999025,16.736387,15.803539,13.313659,11.674315,11.111863,11.893809,14.335675,17.693241,17.909306,17.29198,17.569777,19.901896,19.483486,16.918156,14.757515,13.491997,11.585147,13.639469,11.794352,10.39508,11.063849,12.699762,12.034423,10.055551,11.231899,14.287662,12.202472,9.709162,8.611694,9.788043,11.5645685,9.72288,6.118384,5.120374,6.4819202,9.016385,10.593996,12.0138445,14.335675,15.049029,13.495427,10.854645,12.72034,15.937293,18.835295,20.083664,18.694681,14.352823,12.953552,12.336226,11.547421,10.847785,9.846346,5.6485305,2.8808534,2.6853669,2.6922262,1.4472859,0.6927767,0.41840968,0.40126175,0.20577525,0.07888051,0.020577524,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0,0.030866288,0.037725464,0.030866288,0.020577524,0.034295876,0.020577524,0.006859175,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.0034295875,0.0,0.010288762,0.01371835,0.01371835,0.017147938,0.024007112,0.0274367,0.030866288,0.030866288,0.020577524,0.044584636,0.061732575,0.06516216,0.058302987,0.061732575,0.05144381,0.0274367,0.024007112,0.030866288,0.017147938,0.024007112,0.034295876,0.12689474,0.51100856,1.5261664,3.5976372,3.223812,1.7730967,0.4046913,0.041155048,0.01371835,0.0274367,0.044584636,0.048014224,0.05144381,0.037725464,0.024007112,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.024007112,0.020577524,0.010288762,0.0,0.010288762,0.0274367,0.048014224,0.06516216,0.08573969,0.048014224,0.072021335,0.22292319,0.48700142,0.7579388,0.72021335,0.432128,0.15776102,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.13032432,0.45270553,0.5521636,0.70649505,1.1180456,1.8999915,3.0660512,1.7765263,1.0768905,0.9945804,1.1900668,0.939707,1.3272504,1.7902447,2.020027,2.435007,4.187526,3.2409601,2.760818,3.2478194,4.547633,5.861165,6.6396813,10.045261,14.387119,18.338005,20.920483,18.95533,23.153145,32.094078,44.118214,57.335842,53.44669,49.008804,46.70069,47.13282,48.857903,50.065117,49.61241,47.071087,42.8767,38.32907,35.112118,31.895163,28.825684,26.339231,25.169743,21.572105,19.065077,18.070496,18.866161,21.596113,21.740154,18.279701,13.173045,8.361334,5.7582774,4.705394,3.532475,2.620205,2.0714707,1.7422304,1.7147937,1.5810398,1.3786942,1.1660597,1.039165,0.91227025,0.7442205,0.5521636,0.3841138,0.3018037,0.22978236,0.16804978,0.1097468,0.0548734,0.024007112,1.3581166,1.8348293,2.6133456,3.333559,4.386442,6.910619,5.7754254,6.245279,7.7028537,8.673427,6.8043017,10.2236,20.855322,34.09696,40.088448,23.732746,12.778643,10.957532,10.240748,8.429926,9.126132,12.617453,13.670336,12.3911,10.244178,10.086417,11.2593355,33.273857,92.02612,165.67651,194.68396,112.044624,56.38585,28.211786,20.762722,20.018501,18.79757,24.315775,24.418663,17.065628,10.316199,12.3911,11.773774,11.622872,14.520873,22.491234,24.065414,15.789821,12.46312,21.28059,41.82382,31.16809,17.573206,19.37374,30.25925,19.288,10.912948,7.164408,8.958082,14.490007,19.226267,22.755312,24.552416,24.233465,22.131128,19.288,15.940722,12.771784,9.860064,7.205563,4.715683,3.9714622,3.9954693,4.0263357,3.6696587,2.9151495,2.4247184,2.0028791,1.9102802,2.2566686,2.976882,1.8519772,1.5913286,1.3169615,0.77508676,0.33609957,0.4938606,1.0563129,1.1214751,0.8265306,1.3272504,1.5090185,1.0906088,1.0837497,3.5393343,11.533703,7.507367,2.8945718,0.7888051,1.313532,1.6187652,2.0817597,2.0406046,1.4918705,0.91227025,1.2655178,3.9268777,4.4104495,4.5819287,4.7808447,3.8308492,4.0366244,4.170378,3.683377,2.819121,2.6236343,2.976882,2.620205,2.2463799,2.0097382,1.5090185,0.91227025,0.90884066,1.5090185,2.5824795,3.875434,4.3041325,4.712253,4.852866,4.6127954,4.029765,3.8102717,3.3884325,3.1552205,3.2649672,3.6319332,4.400161,3.7691166,3.2306714,3.3644254,3.8137012,4.448175,4.187526,4.722542,6.8111606,10.254466,8.433355,5.627953,4.602506,6.0806584,8.7283,10.521975,9.167287,8.131552,9.14328,12.205902,12.377381,10.388221,8.001227,7.1987042,10.179015,8.505377,8.436785,11.688034,16.715809,18.708399,20.172834,21.599543,17.809847,10.501397,8.255017,6.619104,8.032094,9.89436,10.611144,9.599416,8.865483,11.05356,12.610593,12.30193,11.214751,8.591117,6.773435,6.783724,7.795452,7.1095347,6.684266,7.3255987,8.491658,8.766026,5.874883,6.742569,6.848886,6.8111606,7.0478024,7.781734,6.0978065,5.2472687,5.0140567,4.7774153,3.4947495,2.5070283,3.1826572,4.262977,4.5682106,3.0043187,2.2360911,2.2566686,2.3218307,2.3218307,2.760818,1.6016173,0.9842916,0.94656616,1.2963841,1.6016173,1.6256244,1.5947582,1.5604624,1.3958421,0.8093826,0.3566771,0.25378948,0.26064864,0.23321195,0.12346515,0.13375391,0.1371835,0.08916927,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.037725464,0.0,0.0,0.048014224,0.024007112,0.017147938,0.037725464,0.0,0.01371835,0.061732575,0.072021335,0.037725464,0.0,0.0,0.0548734,0.14747226,0.20234565,0.09259886,0.12689474,0.16462019,0.2194936,0.2709374,0.26064864,0.08916927,0.06516216,0.12346515,0.2194936,0.30523327,0.23321195,0.19548649,0.15776102,0.12003556,0.106317215,0.15433143,0.41498008,0.53158605,0.42183927,0.274367,0.15090185,0.16804978,0.18519773,0.1920569,0.29151493,0.4115505,0.48014224,0.38754338,0.2469303,0.3806842,0.3806842,0.35324752,0.29151493,0.22978236,0.22978236,0.26407823,0.31895164,0.41840968,0.5453044,0.65505123,0.8745448,1.1214751,1.0940384,0.7990939,0.5796003,0.7133542,0.77508676,0.7133542,0.66191036,0.9294182,1.2346514,1.2209331,1.0666018,0.881404,0.6859175,0.4424168,0.36353627,0.38754338,0.45613512,0.5178677,0.4938606,0.37039545,0.30866286,0.36353627,0.47328308,0.7305021,1.039165,1.3752645,1.5913286,1.4198492,1.7250825,1.937717,1.7971039,1.4472859,1.4335675,1.762808,2.3218307,1.821111,0.8025235,1.6324836,4.1360826,2.976882,1.7353712,1.7388009,2.0440342,2.3972816,2.452155,2.1469216,1.8656956,2.4247184,2.767677,3.0351849,4.5990767,6.9620624,7.7680154,5.717122,6.310441,6.495639,5.7994323,6.3481665,5.9331865,6.927767,8.06296,9.657719,13.625751,13.797231,14.627191,15.45715,15.121051,11.948683,11.14273,11.729189,11.489118,10.103564,9.139851,10.823778,10.247607,9.709162,9.153569,6.166398,4.616225,8.155559,12.734058,15.810398,16.37285,19.572655,21.633839,21.53095,19.377169,16.448301,19.438902,18.8593,16.180794,13.512574,13.612033,17.748116,17.391438,15.134769,14.339106,19.150816,14.925565,13.450842,14.939283,17.864721,18.9519,18.927893,20.779871,25.234905,30.615927,32.8383,26.77136,24.291767,23.845922,25.18003,29.34355,32.392452,29.707087,26.483274,24.391226,21.544668,32.50906,35.42078,32.546783,27.961426,27.556736,26.287788,25.26577,24.85765,24.387796,22.155134,14.05102,10.093276,10.172156,12.435684,13.289652,12.703192,10.213311,8.7317295,9.091836,10.055551,10.251037,10.528833,10.096705,9.403929,10.161868,14.520873,18.12537,18.821575,17.062197,15.913286,13.7526455,13.708061,13.22106,12.027563,12.161317,14.116182,17.20281,19.819586,21.723007,24.0174,24.504402,23.60928,21.60983,18.430603,13.670336,10.521975,10.028113,9.72288,9.599416,12.099585,14.102464,12.898679,11.30735,11.166737,13.351384,14.706071,14.349394,15.247946,16.386568,12.785502,7.366754,7.7131424,9.661148,11.314209,13.059869,15.12448,16.609491,16.300829,13.978998,10.4533825,9.623423,12.178465,14.267084,13.776653,10.347065,9.822338,10.477389,11.197603,11.204462,10.055551,9.640571,6.0840883,3.6079261,3.4981792,4.1189346,2.253239,0.9877212,0.39097297,0.24007112,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.020577524,0.044584636,0.020577524,0.01371835,0.01371835,0.01371835,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0034295875,0.010288762,0.010288762,0.006859175,0.030866288,0.017147938,0.01371835,0.0274367,0.044584636,0.044584636,0.058302987,0.08916927,0.106317215,0.1097468,0.12346515,0.072021335,0.034295876,0.0274367,0.041155048,0.030866288,0.006859175,0.017147938,0.041155048,0.31895164,1.3443983,2.2841053,2.2600982,1.7559488,1.0151579,0.07545093,0.05144381,0.06516216,0.09602845,0.11317638,0.07545093,0.05144381,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.01371835,0.024007112,0.12689474,0.48700142,1.3443983,1.2586586,0.7133542,0.2194936,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.17147937,0.5178677,0.8745448,1.430138,2.8225505,2.2738166,1.6427724,2.3424082,3.724532,3.0523329,2.6853669,2.2086544,1.7936742,2.037175,3.9680326,5.5422134,4.314421,3.1552205,3.3438478,4.5784993,8.189855,11.153018,11.869802,12.325937,18.11165,22.299177,26.02714,38.088997,62.26759,97.36256,83.63049,61.574814,48.655556,49.482086,55.816536,56.6705,56.1252,54.256073,50.70645,44.677235,39.13502,35.35219,32.231262,29.26124,26.490133,22.36434,19.006773,19.061647,22.597551,27.114319,27.68706,24.919382,19.507494,13.227919,8.958082,7.051232,4.938606,3.2958336,2.4247184,2.2429502,2.1469216,2.085189,1.8965619,1.5776103,1.2963841,1.138623,1.0082988,0.83681935,0.64476246,0.53501564,0.42526886,0.36010668,0.28122616,0.17147937,0.061732575,5.4599032,8.512236,6.2830043,3.8479972,3.5118976,4.787704,4.5819287,4.4516044,4.791134,5.446185,5.7068334,8.899779,11.015835,13.742357,16.331696,15.597764,14.335675,14.699212,14.009865,12.065289,11.149589,12.1921835,12.932974,12.833516,12.048141,11.441104,18.921034,64.51397,136.81653,194.05635,164.15721,92.09471,50.178295,30.845709,25.217756,23.094843,21.397196,20.392326,18.067066,15.073037,14.757515,12.459691,11.303921,10.323058,10.22703,13.433694,20.594673,22.714157,22.048819,23.413794,34.182697,24.367218,17.586924,19.925903,25.324074,15.601193,11.338216,8.659708,8.134981,9.630281,12.30536,15.206791,18.070496,19.86074,20.080235,18.79757,16.156786,13.419975,11.015835,8.868914,6.385892,4.7534084,4.0366244,3.6765177,3.3438478,2.9391565,2.6373527,2.551613,3.175798,4.0709205,3.8548563,2.9940298,2.4041407,1.7490896,1.0014396,0.44584638,0.32238123,0.5418748,0.58988905,0.5693115,1.2037852,1.3992717,1.4404267,1.4644338,2.7230926,7.5931067,4.3658648,2.1263442,1.0597426,0.89855194,0.90884066,1.9411465,3.000889,3.5393343,3.5153272,3.391862,4.4687524,4.32128,3.9268777,3.799983,3.9886103,4.372724,4.763697,4.804852,4.40359,3.7108135,3.957744,3.1895163,2.1400626,1.3443983,1.155771,0.8025235,0.8745448,1.2895249,1.9308578,2.668219,3.4467354,3.899441,3.9268777,3.6353626,3.333559,3.4638834,3.4604537,3.3644254,3.6182148,5.0586414,4.139512,4.1772375,5.3501563,7.2947326,9.112414,7.870903,7.023795,7.4936485,9.369633,11.914387,9.585697,8.31675,9.277034,11.4205265,11.461681,8.06296,5.994919,5.360445,6.23156,8.632272,8.615124,8.2653055,7.905199,8.344186,10.871792,9.122703,8.169277,10.30934,14.280802,15.265094,15.138199,13.347955,10.707172,8.56368,8.827758,10.257896,12.027563,13.474849,13.670336,11.417097,8.515666,7.6925645,6.9654922,6.5950966,9.091836,8.879202,7.8983397,7.6514096,8.244728,8.378482,8.97866,8.06296,7.0786686,6.632822,6.4716315,7.630832,7.9737906,7.750868,7.140401,6.23156,6.0223556,5.874883,5.1409516,3.865145,2.7985435,3.0111778,2.8739944,2.9974594,3.1723683,2.369845,2.452155,2.8054025,3.093488,3.275256,3.6285036,1.8245405,1.3066728,1.471293,1.7010754,1.3821237,1.2106444,1.2277923,1.1797781,0.9294182,0.42869842,0.32924038,0.2194936,0.14747226,0.11317638,0.072021335,0.15433143,0.17490897,0.12003556,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.037725464,0.034295876,0.024007112,0.024007112,0.037725464,0.020577524,0.030866288,0.09602845,0.15776102,0.061732575,0.01371835,0.0548734,0.14061308,0.2194936,0.22635277,0.22292319,0.16804978,0.2777966,0.5212973,0.6241849,0.28808534,0.09259886,0.12689474,0.34295875,0.53844523,0.4355576,0.30866286,0.19891608,0.12689474,0.09602845,0.12346515,0.24007112,0.29151493,0.25721905,0.23664154,0.22292319,0.22292319,0.19548649,0.17490897,0.25378948,0.39440256,0.39440256,0.26407823,0.13375391,0.26064864,0.29837412,0.26750782,0.216064,0.17147937,0.13032432,0.1097468,0.15090185,0.22635277,0.34638834,0.53501564,0.64476246,0.7339317,0.72021335,0.6173257,0.5418748,0.66876954,0.6893471,0.7133542,0.7956643,0.96714365,1.0185875,0.91227025,0.8505377,0.8196714,0.5658819,0.37039545,0.37382504,0.4081209,0.41498008,0.45613512,0.5418748,0.7339317,0.6790583,0.44927597,0.5590228,0.64819205,0.6344737,0.70649505,0.939707,1.2860953,1.786815,1.5364552,1.2860953,1.3306799,1.4815818,1.313532,1.7422304,2.1880767,2.194936,1.4129901,1.4644338,1.4781522,1.8313997,2.2978237,2.0577524,1.9411465,1.8828435,2.0234566,2.4315774,3.1106358,4.046913,4.0846386,4.5956473,5.5593615,5.545643,4.091498,4.2115335,4.537344,4.3487167,3.5873485,3.3781435,3.8479972,7.0032177,10.943813,9.853205,10.964391,13.001566,12.590015,9.914937,8.7145815,9.585697,10.923236,11.015835,10.203023,10.847785,8.899779,7.8983397,8.337327,10.847785,16.187653,16.901007,13.975569,14.085316,17.902447,20.083664,18.104792,17.748116,18.067066,17.95389,16.11906,15.46744,15.786391,15.391989,14.445422,14.953001,19.970488,20.124819,18.272842,16.115631,14.205351,12.432255,11.4754,13.334236,17.408587,20.478067,19.250275,20.378609,23.046827,25.26234,23.852781,18.410025,16.266533,16.743246,19.147387,22.762173,23.238884,22.227156,23.242313,26.164322,27.244642,29.840841,30.969175,29.477304,26.061436,23.28347,21.839613,22.648996,23.715597,23.712168,21.983656,20.69413,18.87302,18.132229,17.61779,13.999576,12.905538,13.179905,12.833516,11.533703,10.604284,10.439664,10.539123,9.685155,8.361334,8.745448,14.373401,18.392878,20.663265,21.050808,19.456049,17.195951,15.662926,14.815818,14.925565,16.554619,18.224829,20.738716,22.295748,22.515242,22.419212,22.223726,20.910194,19.301718,17.29198,13.831526,13.042721,12.092726,11.499407,11.835506,13.711491,14.46257,14.112752,13.646329,13.234778,12.21619,11.276484,10.755186,11.893809,12.490558,6.927767,6.2830043,9.537683,12.548861,13.684054,13.817808,14.037301,15.6697855,14.411126,10.789482,10.172156,10.182446,9.410788,8.988949,8.81061,7.5382333,7.7268605,8.237869,8.553391,8.611694,8.824328,8.272165,5.5319247,3.4295874,2.9048605,3.0214665,2.0131679,0.9945804,0.44584638,0.32238123,0.058302987,0.12003556,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.020577524,0.034295876,0.020577524,0.006859175,0.0034295875,0.0034295875,0.0,0.010288762,0.01371835,0.006859175,0.0034295875,0.0034295875,0.0,0.0034295875,0.006859175,0.01371835,0.017147938,0.017147938,0.01371835,0.024007112,0.034295876,0.034295876,0.0548734,0.06516216,0.06516216,0.061732575,0.072021335,0.09259886,0.0548734,0.048014224,0.082310095,0.07888051,0.024007112,0.017147938,0.024007112,0.08916927,0.30523327,0.5418748,0.5658819,0.48700142,0.34638834,0.08916927,0.11317638,0.15090185,0.15776102,0.12689474,0.09945804,0.08573969,0.048014224,0.020577524,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.0034295875,0.041155048,0.14747226,0.37725464,0.35324752,0.18862732,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.082310095,0.4355576,0.70306545,0.94656616,1.6633499,2.8705647,3.5873485,3.9097297,3.957744,3.882293,3.8171308,3.5633414,5.223262,7.1198235,3.7965534,4.0537724,3.175798,2.5584722,2.6716487,3.07634,4.2286816,5.8062916,7.06495,8.584257,12.288212,20.941061,25.59501,34.817173,65.29935,141.87175,151.0459,119.89838,84.292404,64.26704,64.08184,68.176765,64.661446,60.216698,56.639637,50.843636,44.64637,41.189346,38.2399,34.51537,29.67622,22.923363,19.507494,19.188541,22.079683,28.678211,32.807434,31.833431,26.953129,20.04251,13.680624,10.192734,7.2295704,5.0757895,3.7965534,3.2306714,2.8396983,2.6407824,2.5447538,2.4384367,2.1743584,1.8519772,1.6187652,1.4815818,1.3821237,1.1934965,0.89855194,0.7579388,0.65505123,0.5144381,0.31895164,4.479041,7.56224,8.429926,9.983529,12.593445,14.105893,10.031544,5.8371577,3.6319332,3.6525106,4.280125,6.999788,7.2158523,7.2707253,8.666568,12.082437,14.033872,16.283682,16.060759,12.919256,8.772884,9.407358,12.408247,15.731518,18.800999,22.518671,37.852356,97.57862,158.16571,178.64035,120.64946,72.25455,46.38174,33.83974,28.105469,25.337791,23.410364,20.913624,18.468328,16.499744,15.237658,12.459691,11.30735,10.532263,9.613133,8.769455,14.743796,17.401728,16.407146,14.654627,18.255693,15.086755,13.258785,15.999025,20.004784,15.45715,11.760056,9.1810055,8.2481575,8.597976,8.971801,10.100135,12.360233,14.534592,15.848124,15.9750185,14.726648,13.059869,11.327928,9.527394,7.291303,5.4496145,4.616225,4.0606318,3.4535947,2.8808534,4.887162,5.8200097,5.096367,3.525616,3.3232703,3.1586502,2.5619018,1.7799559,1.097468,0.8128122,0.6824879,0.58645946,0.5521636,0.6790583,1.138623,1.3409687,1.5398848,1.4507155,1.5707511,3.192946,2.2600982,1.9857311,1.9857311,2.2360911,3.0660512,2.9288676,3.3609958,3.8342788,3.9611735,3.4810312,4.15666,4.2252517,3.9337368,3.6868064,4.0366244,4.0709205,4.3590055,4.2869844,3.7965534,3.3884325,3.4398763,3.1963756,2.4384367,1.5433143,1.4987297,1.3821237,1.4438564,1.7422304,2.2395205,2.8328393,3.1346428,3.117495,2.9665933,2.8122618,2.719663,3.0043187,3.4467354,3.8342788,4.2835546,5.2164025,5.6142344,6.1561093,7.1781263,8.594546,9.904649,8.872343,7.7371492,6.9620624,7.085528,8.721441,8.889491,9.705732,10.988399,12.710052,14.994157,9.259886,6.245279,5.8165803,6.776865,6.866034,5.874883,5.5147767,5.5422134,6.135532,7.881192,8.988949,10.1652975,12.662037,15.138199,13.63604,11.866373,11.108434,10.700313,10.161868,9.191295,10.079557,11.849225,13.37882,13.862392,12.812939,9.798331,7.548522,5.9331865,5.593657,7.9463544,9.06097,9.966381,10.731179,11.105004,10.511685,9.205012,8.251588,7.222711,6.252138,6.046363,6.509357,7.613684,8.447074,8.196714,6.1458206,5.346727,5.717122,5.254128,3.707384,2.6167753,2.9906003,2.877424,2.7745364,2.767677,2.5619018,3.1826572,3.7691166,4.448175,5.1580997,5.658819,3.1723683,1.7388009,1.3889829,1.6256244,1.4267083,1.1934965,1.0528834,0.83338976,0.50757897,0.20920484,0.216064,0.12689474,0.05144381,0.041155048,0.05144381,0.12689474,0.10288762,0.05144381,0.017147938,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.010288762,0.006859175,0.017147938,0.017147938,0.041155048,0.106317215,0.15776102,0.07545093,0.01371835,0.0274367,0.09259886,0.16804978,0.21263443,0.2469303,0.15090185,0.19548649,0.3841138,0.4972902,0.274367,0.09259886,0.12003556,0.30523327,0.3841138,0.274367,0.25378948,0.18519773,0.06516216,0.037725464,0.061732575,0.11317638,0.14061308,0.14404267,0.15433143,0.21263443,0.25378948,0.22978236,0.15776102,0.13375391,0.2503599,0.23664154,0.14404267,0.06516216,0.12689474,0.15433143,0.14404267,0.13032432,0.12689474,0.106317215,0.0548734,0.061732575,0.12003556,0.2194936,0.34638834,0.39783216,0.39783216,0.39783216,0.4046913,0.4046913,0.490431,0.5590228,0.64476246,0.7373613,0.8128122,0.70306545,0.6207553,0.6756287,0.78194594,0.64476246,0.39440256,0.33609957,0.32924038,0.33952916,0.39783216,0.5418748,0.6790583,0.5727411,0.36696586,0.5693115,0.764798,0.65162164,0.5658819,0.7339317,1.2689474,1.9857311,1.6907866,1.4198492,1.4644338,1.3684053,1.6976458,1.9891608,2.1297739,1.9102802,1.0185875,0.6927767,0.82996017,1.1729189,1.4610043,1.4267083,1.4369972,1.9445761,2.8568463,3.981751,5.0483527,5.446185,4.671098,3.9543142,3.7039545,3.4981792,2.609916,2.7333813,3.018037,2.935727,2.2566686,2.510458,4.7499785,7.06838,8.042382,6.742569,8.779744,10.021255,9.325048,7.473071,7.143831,8.351046,8.405919,7.599966,6.691125,6.9380555,5.113515,4.4927597,5.5593615,8.56025,13.529722,15.419425,13.145609,12.926115,16.139639,19.336014,17.398296,16.660936,17.329706,18.176813,16.540901,13.87954,13.399398,13.965281,14.96672,16.331696,16.434584,15.265094,14.476289,13.862392,11.348505,9.904649,9.9801,11.499407,13.924125,16.280252,15.093615,14.654627,15.45715,16.684942,16.232237,13.077017,11.30735,10.827208,11.561139,13.426835,13.865822,14.754086,16.503176,19.795578,25.584723,29.902573,30.324413,28.551315,25.955118,23.588703,23.660725,24.950249,26.095732,26.226055,24.970827,25.76649,25.77678,25.468117,24.096281,19.70641,16.952452,16.37971,16.47231,16.29054,15.46744,16.191082,14.328816,11.938394,10.978109,13.29994,16.70895,19.1954,20.94449,21.52066,19.853882,18.327715,16.37628,17.072487,19.589804,19.20912,19.425184,19.843594,20.11453,20.162544,20.169403,18.821575,16.70552,14.88098,13.63261,12.4802685,13.29994,12.634601,11.914387,12.127021,13.810948,14.846684,15.059319,14.887839,14.263655,12.627741,10.864933,9.592556,9.0644,8.824328,7.7131424,8.035523,11.077567,13.903547,15.731518,17.95389,18.097933,17.19938,14.898128,12.281353,11.8869505,11.043272,9.781183,9.2153015,9.129561,7.98065,7.8777623,8.320179,8.742019,8.587687,7.31531,7.3084507,5.329579,3.7039545,3.2306714,3.1586502,1.8897027,1.1900668,0.6824879,0.25721905,0.07888051,0.12689474,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.017147938,0.0274367,0.0274367,0.024007112,0.020577524,0.01371835,0.006859175,0.0,0.006859175,0.010288762,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.020577524,0.030866288,0.041155048,0.058302987,0.072021335,0.06516216,0.0548734,0.08916927,0.13375391,0.11317638,0.10288762,0.116605975,0.1097468,0.106317215,0.08916927,0.082310095,0.09259886,0.12003556,0.16462019,0.20577525,0.26750782,0.34295875,0.40126175,0.34295875,0.31552204,0.26750782,0.18862732,0.09602845,0.06516216,0.034295876,0.020577524,0.01371835,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.017147938,0.034295876,0.0548734,0.05144381,0.024007112,0.0034295875,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.26064864,0.4698535,0.5796003,0.66876954,1.4678634,2.428148,3.234101,3.7313912,3.9508848,4.1635194,4.695105,5.5147767,5.6142344,3.0043187,3.3472774,3.3884325,4.105216,5.40503,6.142391,4.2183924,3.865145,4.8185706,6.6053853,8.553391,15.484588,21.139977,28.805105,48.295452,95.977005,119.94296,119.46282,110.53217,104.66072,108.90655,107.28779,94.92755,78.40723,63.25188,53.94741,48.751587,45.82958,41.871834,35.921497,29.34698,23.832203,20.488356,20.025362,22.758743,28.647345,34.01465,35.02638,32.070072,26.047716,18.341434,13.241637,9.410788,6.601956,4.6916757,3.6799474,3.2306714,3.093488,3.0454736,2.901431,2.5070283,2.1469216,2.0680413,2.0303159,1.8999915,1.6324836,1.2037852,0.96714365,0.8848336,0.86082643,0.7579388,3.9474552,7.905199,12.854094,16.527182,17.943602,17.391438,11.38623,6.138962,3.4227283,3.1620796,3.4604537,4.8082814,5.2987127,6.0497923,7.507367,9.438225,10.916377,13.022143,13.203912,10.7757635,6.910619,8.549961,13.670336,19.651537,27.066305,39.711193,67.2062,120.087006,154.90761,146.08328,85.91802,56.907146,42.83555,35.451645,30.60221,28.211786,25.430391,22.69701,20.61525,18.9519,16.640358,13.461131,12.456262,12.240198,11.2250395,7.630832,12.751206,11.897239,9.304471,8.196714,10.765475,11.197603,10.882081,12.120162,14.188204,13.344524,10.367643,8.275595,7.5690994,7.73029,7.239859,6.7219915,7.781734,9.462232,11.026124,11.982979,12.000127,11.441104,10.491108,9.225591,7.6205435,6.0566516,5.3227196,4.6265135,3.7965534,3.2786856,7.9875093,8.834618,6.4373355,3.175798,3.175798,2.9048605,2.3732746,1.8554068,1.488441,1.2758065,1.0631721,0.881404,1.0357354,1.3958421,1.371835,1.4027013,1.7456601,1.762808,1.5090185,1.7147937,2.0680413,2.1229146,2.3801336,3.069481,4.1600895,3.2443898,3.2306714,3.6868064,3.957744,3.1449318,3.8925817,4.32471,4.1635194,3.6353626,3.4947495,3.2958336,3.566771,3.542764,3.117495,2.8328393,3.0283258,3.2992632,3.0420442,2.4007113,2.2806756,2.0646117,2.085189,2.3732746,2.8396983,3.2821152,3.1826572,2.9117198,2.702515,2.6064866,2.5001693,2.603057,3.2649672,3.8137012,4.07435,4.3487167,5.442755,5.977771,6.4304767,7.0375133,7.7885933,7.881192,7.421627,6.293293,5.3501563,6.3961806,7.9257765,8.985519,9.650859,10.926665,14.7369375,10.446524,7.48336,7.654839,10.340206,12.4974165,10.302481,8.666568,7.8194594,7.81603,8.512236,10.504827,12.459691,14.520873,15.505165,12.88496,10.347065,10.14129,10.360784,9.997248,8.961512,9.0644,10.30591,11.506266,12.30536,13.169616,11.736049,9.9801,8.155559,6.927767,7.366754,8.790032,10.532263,12.096155,12.864383,12.103014,9.431366,8.309891,7.56224,6.684266,5.8508763,6.3173003,6.9209075,7.750868,8.018375,6.0532217,4.9523244,5.552502,5.429037,4.1326528,3.1963756,3.2135234,3.1963756,3.0660512,2.836269,2.627064,3.333559,3.998899,4.8254294,5.645101,5.9331865,3.216953,1.7730967,1.471293,1.6873571,1.313532,1.1866373,0.922559,0.59674823,0.3018037,0.13375391,0.1097468,0.06516216,0.024007112,0.010288762,0.044584636,0.09259886,0.041155048,0.010288762,0.034295876,0.07888051,0.058302987,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.030866288,0.01371835,0.030866288,0.07545093,0.106317215,0.06859175,0.024007112,0.024007112,0.058302987,0.106317215,0.17147937,0.23321195,0.12689474,0.09259886,0.18519773,0.28465575,0.17490897,0.06859175,0.09259886,0.20234565,0.20234565,0.12003556,0.18176813,0.19548649,0.116605975,0.024007112,0.030866288,0.05144381,0.072021335,0.08916927,0.106317215,0.16462019,0.22978236,0.22635277,0.14747226,0.048014224,0.12346515,0.13032432,0.09602845,0.058302987,0.0548734,0.058302987,0.0548734,0.06516216,0.082310095,0.07545093,0.044584636,0.06859175,0.16119061,0.28122616,0.35324752,0.30523327,0.23664154,0.2469303,0.31209245,0.3018037,0.36353627,0.48014224,0.607037,0.70649505,0.7442205,0.5453044,0.50757897,0.66191036,0.8505377,0.7305021,0.36696586,0.24007112,0.22635277,0.25721905,0.31895164,0.44584638,0.51100856,0.45613512,0.40126175,0.65505123,1.3238207,1.2758065,1.0185875,0.9259886,1.2517995,2.1194851,2.1126258,1.8348293,1.5913286,1.4164196,1.5055889,1.6256244,1.5673214,1.2792361,0.83681935,0.6756287,0.72364295,0.8471081,0.980862,1.1420527,1.3855534,2.4487255,3.8891523,5.4736214,7.1952744,7.579388,6.2967224,4.681387,3.5530527,3.2478194,2.5378947,2.3321195,3.059192,3.7313912,1.9171394,2.393852,4.7328305,5.844017,5.528495,6.4716315,7.191845,6.9860697,6.4990683,6.1904054,6.351596,7.4627824,6.2692857,4.897451,4.1189346,3.3541365,2.5173173,2.287535,3.2649672,5.353586,7.7783046,9.31133,8.899779,9.187865,11.074138,13.704632,13.512574,13.831526,14.4145565,14.441993,12.538571,12.349944,12.195613,12.627741,13.756075,15.223939,12.689473,10.967821,10.377932,10.299051,9.184435,7.9463544,7.5279446,7.932636,8.844906,9.630281,9.3764925,8.64942,8.580828,9.541112,11.129011,10.319629,8.868914,7.226141,6.135532,6.6465406,7.747438,9.383351,11.149589,14.201921,21.246294,26.798796,27.652763,26.136887,24.398085,24.391226,25.560715,26.490133,27.560165,28.338682,27.567024,28.791388,29.861418,30.307264,29.638494,27.35096,23.647005,21.232576,20.61868,21.297739,21.753874,20.841602,17.724108,15.175924,15.059319,18.303709,20.138538,21.44178,21.640697,20.749004,19.342873,19.895037,18.818146,19.579515,21.308027,18.814716,18.097933,17.569777,16.890718,16.170506,15.988737,14.88098,13.1421795,11.780633,11.262765,11.533703,13.039291,12.679185,12.144169,12.373952,13.560589,14.263655,14.088745,13.543441,12.984418,12.627741,11.4376745,10.189304,8.357904,6.9792104,8.656279,9.201583,11.2421875,13.670336,16.105343,18.886738,19.435472,17.748116,15.854982,14.507155,13.145609,12.524854,11.276484,10.082987,9.184435,8.347616,7.8194594,8.333898,9.033533,9.043822,7.486789,6.5127864,4.616225,3.5393343,3.5050385,3.2443898,1.8382589,1.2723769,0.77165717,0.19891608,0.061732575,0.072021335,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.01371835,0.006859175,0.006859175,0.017147938,0.024007112,0.041155048,0.058302987,0.058302987,0.044584636,0.037725464,0.034295876,0.030866288,0.01371835,0.01371835,0.020577524,0.020577524,0.017147938,0.020577524,0.017147938,0.020577524,0.0274367,0.037725464,0.044584636,0.048014224,0.07545093,0.082310095,0.082310095,0.13032432,0.19891608,0.2469303,0.25378948,0.22292319,0.18176813,0.22978236,0.3018037,0.32581082,0.3018037,0.28465575,0.2503599,0.25378948,0.3018037,0.39097297,0.5007198,0.4355576,0.35324752,0.26750782,0.18176813,0.08573969,0.048014224,0.020577524,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09259886,0.29151493,0.4424168,0.216064,0.28808534,0.805953,1.5364552,2.1812177,2.4007113,2.8499873,3.882293,4.139512,3.350707,2.3424082,2.5550427,2.9494452,3.99204,5.4496145,6.392751,4.0434837,3.0729103,3.6216443,5.0929375,6.111525,10.511685,16.184223,22.751883,31.565924,45.7164,67.16161,85.99004,102.97679,120.88267,144.46794,160.13773,153.40544,124.171646,84.57706,59.03692,51.759335,49.015663,44.437164,36.6863,29.467016,24.45296,21.057667,20.62897,23.478956,28.897703,34.213566,36.593697,34.604538,28.678211,21.095392,15.4914465,10.998687,7.6274023,5.3158607,3.923448,3.5770597,3.649081,3.6353626,3.3266997,2.7985435,2.4384367,2.417859,2.4007113,2.218943,1.8897027,1.4781522,1.214074,1.1111864,1.097468,1.0254467,4.5853586,10.64201,18.145947,20.248285,16.37971,12.250486,7.2158523,4.297273,3.1792276,3.1826572,3.2581081,3.0557625,4.016047,6.0326443,7.7371492,6.475061,6.3001523,6.7494283,7.164408,7.3118806,7.380472,10.017825,15.426285,22.967947,35.475655,59.242695,98.16165,130.34148,139.0149,117.56283,69.5246,47.98679,38.366795,33.97349,31.387585,30.489033,26.064865,22.796469,20.776442,19.696121,18.825006,15.577187,14.812388,14.634049,13.317088,9.297611,13.704632,10.100135,6.9792104,7.9600725,11.784062,11.05699,10.151579,9.455373,9.23245,9.599416,7.939495,6.728851,6.0875177,5.8165803,5.4016004,4.297273,4.4413157,5.4016004,6.691125,7.764586,8.549961,8.81061,8.594546,8.014946,7.2535777,6.228131,5.6348124,4.976331,4.3590055,4.5167665,9.626852,9.091836,6.108095,3.4707425,3.590778,2.5824795,2.0989075,2.020027,2.0268862,1.6084765,1.1729189,1.0460242,1.4232788,1.9823016,1.8519772,1.6221949,1.9925903,2.201795,2.218943,2.7128036,2.9322972,2.2738166,2.0097382,2.4418662,2.8877127,2.4727325,2.7128036,3.3884325,3.8274195,2.8945718,3.5839188,4.341858,4.372724,3.6970954,3.192946,3.3952916,3.6868064,3.875434,3.765687,3.1655092,3.5839188,3.9508848,4.033195,3.765687,3.2581081,2.6236343,2.568761,2.8637056,3.2512488,3.4467354,3.340418,3.2066643,3.07634,2.9220085,2.6785078,2.4795918,3.0900583,3.5359046,3.5359046,3.5050385,3.789694,3.7691166,3.8342788,4.2286816,5.055212,6.217842,6.9552035,6.495639,5.48734,5.994919,7.4113383,6.9723516,6.557371,7.466212,10.422516,10.052121,8.419638,9.767465,15.309678,23.238884,19.723558,16.39,14.445422,13.780083,12.9809885,13.241637,13.505715,13.834956,13.666906,11.814929,10.103564,8.97866,8.114404,7.750868,8.656279,8.988949,9.355915,9.671436,10.323058,12.205902,12.847235,12.682614,10.786053,7.963502,6.7665763,8.073249,9.417647,10.971251,12.329367,12.521424,9.942374,8.042382,7.15069,6.931196,6.3790326,7.2192817,6.725421,6.584808,6.852316,5.9469047,5.3878818,5.662249,5.5113473,4.729401,4.180667,3.8960114,3.981751,3.8377085,3.2581081,2.4555845,2.8088322,3.5050385,4.245829,4.664239,4.32471,2.0440342,1.4267083,1.6667795,1.8965619,1.214074,1.0460242,0.7373613,0.48357183,0.33266997,0.17833854,0.06859175,0.0548734,0.041155048,0.01371835,0.041155048,0.06516216,0.030866288,0.020577524,0.06516216,0.1371835,0.116605975,0.048014224,0.0034295875,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.01371835,0.044584636,0.09602845,0.0274367,0.0034295875,0.020577524,0.058302987,0.06859175,0.041155048,0.048014224,0.05144381,0.06516216,0.1371835,0.20577525,0.12003556,0.05144381,0.07888051,0.17147937,0.09602845,0.041155048,0.05144381,0.1097468,0.12346515,0.08916927,0.13032432,0.19891608,0.216064,0.058302987,0.034295876,0.034295876,0.048014224,0.06859175,0.09259886,0.11317638,0.16462019,0.17833854,0.12689474,0.030866288,0.058302987,0.106317215,0.14061308,0.1371835,0.072021335,0.044584636,0.0274367,0.034295876,0.048014224,0.0274367,0.041155048,0.13032432,0.28465575,0.44584638,0.5144381,0.36696586,0.2469303,0.25721905,0.34638834,0.29837412,0.37382504,0.4972902,0.6379033,0.7579388,0.8093826,0.6173257,0.5555932,0.6927767,0.864256,0.66191036,0.26407823,0.1371835,0.14747226,0.20577525,0.26064864,0.29837412,0.42183927,0.5555932,0.69963586,0.91227025,1.862266,1.937717,1.5330256,1.0734608,1.0117283,1.786815,2.1057668,1.8828435,1.430138,1.4610043,0.805953,0.78537554,0.94999576,1.0425946,1.0117283,0.8093826,0.9294182,1.1832076,1.3992717,1.4369972,1.6359133,2.6613598,4.0229063,5.6999745,8.131552,9.925226,9.156999,7.438775,5.8508763,4.9180284,3.724532,2.8980014,4.108646,5.641671,2.4075704,2.585909,2.983741,3.673088,5.1340923,8.2310095,6.159539,4.671098,4.2389703,4.6608095,5.0757895,5.874883,4.616225,3.799983,3.7005248,2.3629858,1.7559488,1.5913286,2.0234566,2.860276,3.566771,3.8274195,3.9028704,4.105216,4.664239,5.6965446,6.5470824,7.963502,8.162418,6.944915,5.6999745,11.101575,13.13189,12.730629,11.495977,11.653738,11.05699,9.873782,8.357904,7.0889573,6.9963584,6.756287,5.435896,5.06893,5.562791,4.698535,5.31929,5.501058,5.7308407,6.560801,8.628842,9.6988735,8.899779,7.0135064,5.113515,4.554492,5.302142,6.2830043,8.388771,12.003556,17.021042,21.146837,22.916504,22.234016,21.016512,23.204588,24.734184,25.862518,27.807095,29.906002,29.614489,30.255821,31.641375,32.94119,33.788296,34.271866,30.454737,26.411253,24.27462,24.470106,25.718477,21.582394,19.082224,18.118511,18.691252,20.899906,22.552967,23.393215,22.374628,20.237995,19.514353,21.146837,21.150267,20.827885,20.179693,17.885298,16.578627,15.803539,14.459141,12.79922,12.415107,12.452832,11.369082,10.645439,10.899229,11.880091,12.912396,12.648318,12.545431,12.960411,13.145609,12.349944,11.115293,10.000677,9.736599,11.2421875,11.314209,10.9198065,9.256456,7.298162,7.781734,8.831187,10.251037,12.428825,14.760944,15.638919,16.393429,16.438013,16.194511,15.446862,13.341095,13.708061,12.205902,9.925226,8.014946,7.6959944,7.473071,8.097256,8.683716,8.875772,8.844906,6.276145,4.0023284,3.1655092,3.450165,3.0969174,2.1229146,1.4335675,0.881404,0.4081209,0.037725464,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.006859175,0.006859175,0.017147938,0.034295876,0.048014224,0.06516216,0.07888051,0.08573969,0.07545093,0.072021335,0.06859175,0.0548734,0.030866288,0.017147938,0.024007112,0.024007112,0.017147938,0.030866288,0.017147938,0.024007112,0.034295876,0.041155048,0.041155048,0.030866288,0.061732575,0.09602845,0.12003556,0.15776102,0.23664154,0.3566771,0.39783216,0.34295875,0.2709374,0.31895164,0.490431,0.5658819,0.5007198,0.42869842,0.32581082,0.2777966,0.2709374,0.29151493,0.31552204,0.32238123,0.22978236,0.14061308,0.09259886,0.061732575,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.01371835,0.05144381,0.024007112,0.006859175,0.0,0.01371835,0.072021335,0.044584636,0.01371835,0.0,0.0,0.0,0.0,0.0,0.1920569,0.42869842,0.23664154,0.18176813,0.11317638,0.10288762,0.15776102,0.23664154,0.78194594,1.7559488,2.4555845,2.5413244,2.0303159,1.6633499,1.6942163,1.961724,2.3904223,2.9803114,2.4624438,2.3424082,2.8396983,3.799983,4.6676683,7.599966,12.106443,17.734396,23.338343,27.1006,34.114105,46.57037,67.09988,98.44288,143.43907,191.44643,212.84706,184.54953,120.15217,69.91214,55.909134,51.522694,46.78643,38.80921,31.74426,25.392666,21.61326,21.20171,24.346642,30.615927,35.465363,38.555424,36.2576,29.151493,22.017952,16.304258,11.393089,8.004657,5.9914894,4.338428,4.033195,4.273266,4.2595477,3.7553983,3.1037767,2.6579304,2.5447538,2.4727325,2.2600982,1.8348293,1.5707511,1.3786942,1.2723769,1.196926,1.0597426,2.287535,9.040393,17.686382,19.871029,15.227368,11.382801,5.4016004,2.4590142,1.7525192,2.2566686,2.7470996,2.9048605,5.0243454,7.740579,8.697433,4.547633,3.765687,3.8445675,4.5784993,6.101236,8.89635,10.299051,13.488567,23.866499,44.704674,77.162285,113.90346,137.33783,135.62303,108.80709,68.8181,44.96532,32.804005,27.693918,26.634176,28.242653,21.93221,18.478617,16.496315,15.638919,16.602633,17.95732,17.826996,16.105343,13.838386,13.227919,9.530824,7.7440085,8.131552,8.597976,4.715683,3.5187566,4.1463714,5.8062916,7.9772205,10.405369,7.8674736,6.5470824,5.5079174,4.1189346,2.0440342,1.99602,2.1743584,2.6750782,3.3952916,4.029765,5.1752477,5.892031,6.108095,5.9469047,5.751418,5.2644167,4.9214582,4.8425775,5.3227196,6.835168,6.358455,4.57507,3.1517909,2.7745364,3.1277838,2.3218307,1.920569,1.920569,1.9994495,1.5090185,0.94999576,0.6344737,0.45613512,0.7407909,2.2429502,2.0234566,1.7936742,1.6290541,1.6256244,1.9068506,2.2738166,2.2360911,1.5776103,0.6893471,0.5796003,1.5947582,1.8999915,2.201795,2.5070283,2.1503513,2.1640697,3.5050385,4.4996185,4.7774153,5.2781353,6.8797526,6.728851,6.4716315,6.39961,5.446185,5.2026844,5.3878818,5.675967,5.528495,4.2115335,3.1860867,2.976882,3.0797696,3.199805,3.2512488,3.309552,3.309552,3.234101,3.1072063,2.959734,2.8877127,3.3541365,4.2218223,4.931747,4.5167665,4.383013,3.532475,3.1243541,3.6044965,4.715683,6.0806584,6.999788,6.4133286,4.7499785,3.9063,7.1884155,6.125243,4.386442,4.1463714,6.0875177,8.639131,8.937505,11.787492,18.903887,28.914852,23.640146,19.504065,17.929884,17.583494,14.373401,13.910407,12.154458,10.72775,9.9698105,8.958082,10.179015,9.403929,8.268735,8.05953,9.719451,10.39165,10.127572,9.616563,9.424506,10.010965,11.108434,11.667457,9.482809,5.813151,5.3878818,7.2775846,8.711152,9.743458,10.64201,11.8869505,9.239308,6.6636887,5.4839106,5.9743414,7.3530354,6.574519,7.514226,7.936065,7.4010496,7.2775846,6.8763227,5.8405876,5.103226,4.863155,4.6093655,4.695105,5.5490727,5.552502,4.3349986,2.760818,2.5173173,3.4467354,4.3178506,4.4104495,3.4947495,2.2498093,1.2346514,1.1043272,1.6770682,1.9239986,0.8848336,0.4698535,0.42183927,0.45956472,0.29151493,0.12003556,0.048014224,0.030866288,0.0274367,0.01371835,0.05144381,0.024007112,0.0,0.01371835,0.07545093,0.0274367,0.024007112,0.017147938,0.006859175,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.020577524,0.058302987,0.16804978,0.082310095,0.024007112,0.01371835,0.041155048,0.09259886,0.0548734,0.037725464,0.041155048,0.06516216,0.07545093,0.17490897,0.16119061,0.09602845,0.048014224,0.12346515,0.09602845,0.044584636,0.0274367,0.048014224,0.061732575,0.037725464,0.020577524,0.034295876,0.058302987,0.044584636,0.020577524,0.006859175,0.0,0.006859175,0.030866288,0.09259886,0.15090185,0.12346515,0.030866288,0.030866288,0.030866288,0.11317638,0.23664154,0.30523327,0.18176813,0.08573969,0.05144381,0.06516216,0.07545093,0.01371835,0.0274367,0.13032432,0.29494452,0.45613512,0.5041494,0.39440256,0.274367,0.28808534,0.39783216,0.39783216,0.53158605,0.6001778,0.6927767,0.7956643,0.8093826,0.8196714,0.5761707,0.41840968,0.4046913,0.31895164,0.18519773,0.116605975,0.12346515,0.19891608,0.31895164,0.2709374,0.45956472,0.84367853,1.255229,1.3889829,1.2037852,1.2963841,0.9842916,0.34981793,0.22978236,0.40126175,0.5624523,0.64133286,0.6790583,0.84024894,1.1214751,1.1797781,1.2415106,1.3684053,1.4644338,1.039165,1.2689474,1.7456601,2.061182,1.8142518,1.3992717,1.2963841,1.8039631,3.2581081,6.042933,10.827208,12.116733,11.533703,9.887501,7.140401,4.5784993,3.7519686,3.9474552,4.3109913,3.8617156,3.1415021,2.7779658,3.649081,5.751418,8.193284,5.65539,3.316411,1.9754424,1.670209,1.6942163,1.4369972,1.5570327,2.411,3.3129816,2.534465,1.0666018,0.78537554,1.0837497,1.2723769,0.5658819,0.30866286,0.20920484,0.17833854,0.29151493,0.77851635,0.6310441,1.0082988,1.1660597,1.6736387,4.3933015,12.891819,17.641798,16.263103,10.899229,8.224151,10.652299,9.102125,6.543653,4.8494368,4.7774153,6.108095,7.8023114,9.287323,9.434795,6.591667,6.420188,6.478491,7.4181976,8.529384,7.7371492,10.799771,11.832077,11.214751,9.242738,6.118384,3.8857226,3.7108135,5.768566,9.537683,13.810948,20.083664,21.908205,20.491785,18.324286,19.164536,21.77788,25.94483,30.663942,34.25129,34.36104,31.617367,33.09895,35.839188,37.859215,38.17817,33.50021,27.827673,24.466677,23.69159,22.751883,19.456049,19.29143,19.871029,20.237995,20.872469,21.143406,20.670124,20.406046,20.711279,21.345753,17.830425,16.722668,18.217968,21.109112,22.77932,19.178253,15.258235,12.88496,13.035862,15.806969,15.076467,11.550851,9.321619,10.134431,13.38225,12.490558,12.360233,12.651748,12.754636,11.763485,9.3593445,7.606825,6.4887795,6.4716315,8.484799,9.1810055,9.1981535,9.14328,8.903209,7.658269,8.464222,9.647429,11.38623,12.977559,12.816368,13.526293,14.994157,15.6526375,15.028452,13.732068,12.439114,11.218181,10.261326,9.270175,7.4765005,9.15014,9.623423,8.937505,7.9772205,8.453933,7.623973,5.5662203,3.9680326,3.4638834,3.6456516,3.316411,2.3561265,1.6736387,1.2449403,0.12346515,0.048014224,0.020577524,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.017147938,0.030866288,0.0548734,0.07888051,0.09259886,0.09602845,0.12346515,0.12346515,0.12346515,0.09602845,0.0548734,0.030866288,0.017147938,0.024007112,0.024007112,0.017147938,0.030866288,0.017147938,0.01371835,0.020577524,0.030866288,0.030866288,0.017147938,0.041155048,0.08573969,0.12346515,0.12346515,0.12346515,0.21263443,0.274367,0.2709374,0.26064864,0.26064864,0.2777966,0.28465575,0.28465575,0.31895164,0.33266997,0.33609957,0.30523327,0.25378948,0.22978236,0.16804978,0.08916927,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.06516216,0.030866288,0.0,0.072021335,0.36696586,0.2194936,0.072021335,0.0,0.0,0.0,0.0,0.0,0.09602845,0.23664154,0.21263443,0.6173257,0.48700142,0.28808534,0.23664154,0.31895164,0.61389613,1.2826657,1.7079345,1.7490896,1.7250825,1.5055889,1.2860953,1.2860953,1.4781522,1.587899,1.097468,1.7559488,2.6956558,3.542764,4.4104495,5.3501563,8.165848,13.207341,19.764713,26.061436,26.75764,29.669361,38.284485,58.16923,97.00245,144.50566,212.22974,218.26237,155.02078,89.12469,65.40566,55.147766,49.317467,43.048183,35.612835,28.520449,23.835632,23.081123,26.743923,34.302734,39.014988,42.845837,40.685196,32.454185,23.11542,15.107333,9.866923,7.6685576,7.160979,5.3398676,4.6436615,4.698535,4.57164,3.9200184,3.0043187,2.2498093,2.1160555,2.0920484,1.8348293,1.1763484,1.0288762,0.9911508,1.0837497,1.1934965,1.0837497,7.023795,28.17749,32.282707,22.786179,8.567109,3.899441,2.4898806,2.702515,2.8225505,2.503599,2.7951138,3.9097297,5.6519604,6.824879,6.7322803,5.1683884,5.8817425,5.9469047,5.2472687,4.7945633,6.711703,6.893471,12.867812,30.955456,61.6777,99.77013,128.81874,139.41959,123.736084,88.03408,52.69218,37.735752,29.35727,25.471546,24.94682,27.632187,23.44123,25.145735,30.958885,34.052376,22.559826,18.132229,18.931322,19.901896,18.509483,14.754086,9.386781,12.133881,14.493437,12.315649,5.8371577,8.673427,9.993818,8.690575,5.8405876,4.705394,4.197815,3.3541365,2.4898806,1.7662375,1.214074,1.3512574,1.2346514,1.2792361,1.6667795,2.318401,3.4364467,5.288424,6.5985265,7.1712675,7.9120584,11.410237,10.861504,9.191295,8.351046,9.325048,7.250148,5.576509,4.496189,3.9200184,3.4810312,3.234101,2.6922262,2.1160555,1.646202,1.3169615,1.1454822,0.8162418,0.5521636,0.6276145,1.3889829,2.0680413,2.2395205,2.0920484,1.762808,1.3203912,3.1140654,1.9102802,0.72707254,0.66533995,0.89855194,1.7147937,1.9891608,1.9548649,2.0817597,3.0557625,4.0434837,4.770556,4.245829,3.2443898,4.3041325,5.627953,6.677407,7.085528,6.927767,6.728851,6.708273,6.7459984,6.121814,4.880303,3.8445675,3.7176728,3.4913201,3.4055803,3.532475,3.7862647,3.5050385,3.0454736,2.7402403,2.719663,2.8739944,3.2786856,3.7553983,4.180667,4.5339146,4.9180284,4.9694724,4.2115335,3.4707425,3.0797696,2.8705647,3.40901,5.504488,6.543653,5.638242,3.6147852,4.914599,6.307011,6.444195,5.586798,5.576509,5.501058,6.210983,8.793462,13.358243,19.05136,20.399187,21.345753,20.19341,16.88386,12.9707,10.182446,8.930646,8.31675,7.864044,7.517656,8.279024,8.611694,8.656279,8.505377,8.193284,8.193284,8.076678,7.723431,7.486789,8.179566,8.89635,9.074688,8.886061,8.296172,7.058091,8.1212635,8.879202,9.407358,10.05898,11.458252,10.645439,9.3936405,8.56368,8.40249,8.549961,7.4970784,7.48336,8.2653055,8.937505,7.9257765,7.1712675,6.56766,5.761707,4.880303,4.547633,3.8137012,3.99204,4.6093655,5.0655007,4.6402316,4.0846386,3.5290456,3.40901,3.566771,3.2272418,2.0886188,1.0185875,0.7579388,1.2929544,1.8485477,0.9568549,0.4629943,0.28808534,0.29837412,0.3018037,0.30866286,0.23664154,0.19548649,0.16804978,0.041155048,0.058302987,0.030866288,0.006859175,0.006859175,0.0274367,0.037725464,0.0548734,0.0548734,0.044584636,0.07888051,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.0274367,0.05144381,0.13032432,0.2777966,0.09602845,0.020577524,0.0034295875,0.010288762,0.030866288,0.1097468,0.072021335,0.037725464,0.044584636,0.0274367,0.06516216,0.09259886,0.06859175,0.0274367,0.061732575,0.048014224,0.020577524,0.030866288,0.072021335,0.072021335,0.037725464,0.05144381,0.044584636,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.006859175,0.041155048,0.14404267,0.15433143,0.09945804,0.0274367,0.017147938,0.017147938,0.06516216,0.16804978,0.24350071,0.12346515,0.044584636,0.037725464,0.048014224,0.048014224,0.01371835,0.017147938,0.082310095,0.16462019,0.20920484,0.16119061,0.17833854,0.23664154,0.32238123,0.39097297,0.36010668,0.39783216,0.61046654,0.77165717,0.7407909,0.48014224,0.29494452,0.31209245,0.5144381,0.805953,1.0048691,0.89855194,0.6962063,0.4972902,0.42526886,0.6241849,0.64476246,0.59674823,0.7099246,0.922559,0.8505377,0.61046654,0.4972902,0.42869842,0.490431,0.9259886,1.3889829,1.1626302,0.8162418,0.72364295,1.0460242,1.4267083,1.5707511,1.4678634,1.1626302,0.7339317,1.2037852,1.9171394,2.428148,2.4007113,1.6221949,1.3821237,1.1763484,1.3546871,2.0268862,3.0523329,5.552502,7.514226,8.711152,9.009526,8.361334,5.8062916,4.7671266,4.6882463,4.870014,4.4447455,3.5118976,2.9254382,2.7779658,3.3987212,5.360445,4.07435,2.4007113,1.7662375,3.1209247,6.941485,6.7528577,9.9801,20.519222,28.187778,8.745448,1.9308578,0.65848076,0.85739684,0.59674823,0.11317638,0.12003556,0.11317638,0.12346515,0.15090185,0.18176813,0.2777966,0.66191036,0.6962063,0.6962063,1.9548649,6.8557453,13.111313,15.560039,13.296511,9.6645775,8.1384115,7.531374,6.691125,5.535354,5.0312047,6.2247014,9.983529,13.073587,13.646329,11.2421875,9.499957,6.944915,5.1100855,5.055212,7.3564653,10.744898,9.623423,8.014946,7.5382333,7.4010496,5.353586,4.098357,4.5270553,7.466212,13.663476,18.386019,19.147387,16.726099,14.037301,16.13621,21.153696,27.591032,33.66826,37.142433,35.33847,32.574223,32.317,32.02892,31.476753,32.721695,33.49335,33.452198,31.932888,28.647345,23.70188,21.352612,22.669573,23.252604,22.155134,21.911634,18.732407,19.630959,20.189981,18.828436,16.80498,15.693792,19.11995,21.424633,19.79901,14.284232,13.097594,13.776653,14.658057,15.234227,16.149927,15.45715,13.869251,13.423406,14.177915,14.212211,11.30049,10.590566,11.825217,13.498857,12.850664,10.933525,9.383351,8.021805,6.8866115,6.2247014,5.878313,5.5250654,6.478491,8.330468,8.930646,8.934075,10.7586155,12.140739,12.415107,12.500846,14.407697,15.724659,15.419425,13.858963,12.768354,11.523414,11.4205265,11.770344,12.034423,11.821788,11.718901,10.683165,9.47938,8.659708,8.587687,8.968371,7.4936485,5.9331865,4.9008803,3.841138,3.4433057,2.6785078,2.0440342,1.6290541,1.1111864,0.42183927,0.12346515,0.030866288,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0,0.006859175,0.024007112,0.048014224,0.07888051,0.08573969,0.09602845,0.14404267,0.19891608,0.19548649,0.216064,0.22635277,0.19891608,0.1371835,0.09259886,0.041155048,0.020577524,0.017147938,0.017147938,0.017147938,0.006859175,0.010288762,0.017147938,0.017147938,0.017147938,0.017147938,0.0274367,0.061732575,0.106317215,0.13375391,0.15433143,0.20577525,0.26407823,0.3018037,0.30866286,0.38754338,0.3806842,0.29494452,0.1920569,0.20920484,0.18519773,0.17833854,0.17147937,0.14404267,0.06859175,0.037725464,0.017147938,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.024007112,0.024007112,0.0034295875,0.0034295875,0.024007112,0.041155048,0.17490897,0.33609957,0.20920484,0.16804978,0.06516216,0.0,0.0,0.0,0.0,0.0,0.020577524,0.048014224,0.041155048,0.12346515,0.15776102,0.31209245,1.0323058,3.0420442,2.7402403,2.2120838,1.6221949,1.1729189,1.0906088,1.1729189,1.0666018,0.9877212,1.0700313,1.3546871,1.2860953,1.6530612,1.8416885,1.821111,2.1503513,2.877424,4.4756117,8.31675,14.634049,22.53582,24.52841,27.786518,33.778008,45.80557,69.02388,118.14586,169.29129,185.72588,159.83592,113.04949,83.489876,66.242485,56.749382,50.19887,41.535732,34.56681,28.544456,25.337791,26.606739,33.802013,40.82924,43.600346,41.48772,35.129265,26.42497,18.554068,11.924676,8.241299,7.346176,7.1952744,6.0806584,5.7136927,5.9571934,5.778855,3.2615378,2.1434922,2.3081124,2.369845,1.8245405,1.0288762,0.881404,0.78537554,0.823101,0.9774324,1.1214751,5.1340923,19.473198,19.963629,13.125031,5.4907694,3.5873485,3.3472774,3.1552205,2.5378947,1.7696671,1.8725548,2.767677,3.8342788,4.7499785,5.171818,4.73969,5.6348124,6.368744,5.977771,5.0449233,5.6793966,6.186976,15.261664,39.546574,77.23088,118.063545,137.9963,133.16402,104.11542,64.887794,42.976162,38.1473,39.820942,49.2283,61.715427,66.72605,39.72491,31.720255,34.529087,37.968964,29.85113,23.314335,21.551527,20.416334,17.744686,13.37882,12.082437,12.713481,11.924676,8.872343,5.2301207,8.388771,10.991828,10.093276,6.3618846,4.0846386,3.316411,2.3252604,1.5021594,1.0323058,0.89855194,1.1900668,1.2895249,1.4644338,1.9651536,3.018037,5.4016004,7.8263187,8.512236,7.671987,7.4936485,15.337115,13.05301,9.273604,7.8537555,7.8537555,6.5024977,5.453044,4.712253,4.245829,3.9543142,3.765687,3.3987212,2.6647894,1.9137098,2.0440342,1.5330256,1.2792361,1.3649758,1.5947582,1.4953002,2.0165975,2.1503513,2.0749004,1.8554068,1.430138,2.0646117,1.8656956,1.6187652,1.646202,1.8108221,1.7079345,2.0749004,2.4007113,2.7573884,3.782835,5.0826488,5.003768,4.3178506,4.1600895,5.9983487,5.593657,5.9228973,5.9228973,5.5902276,5.9983487,6.444195,6.8043017,6.4373355,5.3913116,4.40359,4.3487167,4.0777793,3.7965534,3.6970954,3.957744,3.525616,2.8499873,2.411,2.3252604,2.369845,2.5413244,2.867135,3.234101,3.6353626,4.1772375,4.3178506,4.0194764,3.590778,3.0454736,2.0989075,2.020027,4.170378,6.495639,7.1781263,4.6402316,4.184097,4.5853586,4.6676683,4.273266,4.256118,3.4947495,4.0606318,5.7994323,8.30646,10.9198065,15.752095,18.938183,18.44432,14.507155,9.633711,6.8145905,5.638242,5.079219,4.5922174,4.1155047,5.1752477,6.6396813,7.500508,7.4627824,6.941485,7.181556,7.2707253,7.1712675,7.0786686,7.4113383,7.613684,7.888051,8.423067,8.824328,8.107545,8.580828,8.862054,8.762596,8.786603,10.124143,12.487128,12.05843,11.30049,10.762046,9.088407,6.8214493,7.130112,8.47451,9.458802,8.81061,8.296172,7.936065,7.0272245,5.6176643,4.4859004,4.2115335,4.722542,5.4839106,5.826869,4.938606,4.5956473,4.0229063,3.9028704,4.1635194,3.9543142,3.0729103,2.253239,1.5673214,1.3478279,2.177788,0.805953,0.33609957,0.22978236,0.20577525,0.24007112,0.2469303,0.17490897,0.14061308,0.14061308,0.0548734,0.058302987,0.044584636,0.034295876,0.030866288,0.01371835,0.024007112,0.07888051,0.07545093,0.024007112,0.044584636,0.017147938,0.0034295875,0.0,0.006859175,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.07888051,0.106317215,0.116605975,0.15090185,0.044584636,0.006859175,0.0,0.030866288,0.16119061,0.12346515,0.058302987,0.024007112,0.024007112,0.01371835,0.030866288,0.06516216,0.07545093,0.058302987,0.044584636,0.034295876,0.01371835,0.024007112,0.058302987,0.06859175,0.037725464,0.037725464,0.034295876,0.024007112,0.017147938,0.0034295875,0.006859175,0.017147938,0.034295876,0.0548734,0.106317215,0.09602845,0.058302987,0.020577524,0.01371835,0.006859175,0.037725464,0.09259886,0.12689474,0.07888051,0.1371835,0.19891608,0.21263443,0.18519773,0.15090185,0.15090185,0.16462019,0.15776102,0.13032432,0.08573969,0.16462019,0.2469303,0.31895164,0.34638834,0.28808534,0.2469303,0.30866286,0.34981793,0.32238123,0.24007112,0.20577525,0.34638834,0.6001778,0.8745448,1.0460242,0.9945804,0.764798,0.5555932,0.5178677,0.7305021,0.72364295,0.5418748,0.51100856,0.64476246,0.6241849,0.4046913,0.39440256,0.4972902,0.71678376,1.1351935,1.6496316,1.7388009,1.3992717,0.8676856,0.6036074,0.96371406,1.2998136,1.1694894,0.65848076,0.36696586,0.7990939,1.5638919,2.4041407,2.9700227,2.843128,2.6064866,2.3561265,1.9239986,1.5501735,1.9102802,2.7642474,4.15666,5.6245236,6.835168,7.6033955,7.1712675,6.444195,5.3432975,4.098357,3.2649672,2.819121,2.7951138,2.5790498,2.2635276,2.6476414,2.3904223,1.546744,2.1160555,4.389872,6.9380555,4.040054,5.2266912,10.89237,14.918706,4.6882463,0.97057325,0.2503599,0.37725464,0.33266997,0.2194936,0.21263443,0.6173257,1.0117283,1.0048691,0.23321195,0.4424168,0.51100856,0.38754338,0.28808534,0.7099246,2.6064866,6.7494283,10.909517,13.557159,13.869251,11.838936,10.587136,9.465661,8.337327,7.596536,7.606825,8.718011,9.571979,9.602845,9.026674,8.3922,6.800872,6.6053853,8.128122,9.688584,9.078118,8.296172,8.224151,8.868914,9.369633,7.1026754,5.439326,5.8165803,8.779744,13.992717,16.098484,15.580616,13.896688,13.63604,18.485476,23.588703,26.630747,30.770258,35.31789,35.767166,31.42874,29.662502,28.225504,27.148615,28.719366,32.26213,33.994072,33.627106,30.811415,25.132017,24.953678,27.090311,27.237783,24.638157,22.089973,18.656956,18.879879,19.603521,18.752985,15.340545,15.920145,19.384027,20.097382,16.691803,12.061859,13.121602,14.0750265,15.004445,15.6526375,15.402277,15.354263,14.579176,13.2690735,11.910957,11.279913,10.161868,9.39707,9.6988735,10.823778,11.595435,11.30735,11.187314,10.220171,8.2653055,6.0635104,6.7631464,7.14726,8.303031,10.14472,11.38966,12.05843,12.850664,12.38424,10.916377,10.360784,12.620882,14.589465,14.791811,13.258785,11.547421,11.492548,11.592006,11.917816,12.343085,12.535142,11.478829,10.124143,9.595985,9.6988735,8.913498,9.006097,8.14527,7.116394,6.0669403,4.530485,3.6044965,2.6990852,2.0749004,1.6976458,1.2312219,0.59331864,0.25721905,0.08916927,0.01371835,0.006859175,0.0,0.0,0.0,0.0034295875,0.010288762,0.037725464,0.0274367,0.044584636,0.09945804,0.12689474,0.12003556,0.16119061,0.2194936,0.26064864,0.24007112,0.30866286,0.34638834,0.32581082,0.2503599,0.14404267,0.082310095,0.05144381,0.034295876,0.0274367,0.034295876,0.020577524,0.020577524,0.024007112,0.024007112,0.01371835,0.01371835,0.030866288,0.061732575,0.09602845,0.12003556,0.13032432,0.14061308,0.15776102,0.17833854,0.18176813,0.22978236,0.20920484,0.14404267,0.07888051,0.082310095,0.061732575,0.0548734,0.0548734,0.048014224,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.034295876,0.0548734,0.044584636,0.0,0.0034295875,0.017147938,0.16804978,0.36696586,0.29494452,0.116605975,0.044584636,0.017147938,0.0034295875,0.017147938,0.034295876,0.01371835,0.0,0.017147938,0.09259886,0.017147938,0.030866288,0.12689474,0.4938606,1.488441,1.4918705,1.196926,0.8128122,0.52472687,0.5007198,0.65162164,0.7133542,0.7339317,0.82996017,1.196926,1.2689474,1.3409687,1.214074,1.0048691,1.1489118,1.6153357,2.784825,5.435896,9.9869585,16.506605,19.442331,23.242313,28.372976,36.387924,49.941654,85.787704,121.650894,143.8952,147.90782,138.08548,122.642044,103.45693,84.364426,68.19392,56.78368,45.249977,34.49136,27.357819,25.492125,29.34698,35.3419,38.377083,38.363365,34.782875,26.68562,19.068506,12.459691,8.683716,8.025234,9.2153015,8.412778,8.035523,7.48336,6.228131,3.8308492,2.4007113,2.294394,2.1126258,1.4575747,0.9294182,0.78194594,0.69963586,0.6962063,0.7888051,0.97400284,2.7093742,7.191845,6.7048435,5.099797,4.2183924,3.865145,3.6456516,3.0146074,2.2326615,1.6599203,1.7525192,2.0234566,2.620205,3.6627994,4.6402316,4.396731,5.1512403,6.385892,6.4716315,5.4941993,5.2472687,5.9640527,16.067617,39.347656,74.50779,115.18613,132.95482,118.46824,84.63879,49.993095,38.672028,40.033573,48.027943,65.94754,86.86116,93.61402,51.39237,34.59425,32.371876,35.02638,34.021507,31.027477,29.563044,25.059996,17.923023,13.519434,14.2362175,11.746337,8.344186,5.778855,5.284994,6.7974424,8.419638,8.107545,5.970912,4.280125,3.2203827,2.2120838,1.7525192,1.8176813,1.879414,1.7490896,2.644212,3.3541365,3.4021509,3.0557625,5.0757895,7.6514096,8.416207,7.267296,6.368744,11.921246,9.537683,6.5950966,5.8988905,5.672538,6.111525,7.6685576,8.587687,7.936065,5.6073756,4.6608095,4.187526,3.4398763,2.5584722,2.5584722,1.6187652,1.5570327,1.8759843,2.061182,1.5741806,1.7319417,1.920569,1.9891608,1.9445761,1.9685832,1.8142518,2.6579304,3.0351849,2.5721905,1.9685832,1.529596,1.8828435,2.627064,3.5153272,4.4859004,5.144381,4.9351764,4.6573796,4.8837323,5.970912,4.8905916,4.7191124,4.355576,3.8857226,4.5682106,5.1992545,5.7308407,5.826869,5.4153185,4.7088237,4.7945633,4.629943,4.341858,4.1292233,4.256118,3.74168,2.884283,2.301253,2.1194851,1.9651536,1.8897027,2.0749004,2.4487255,2.9254382,3.4021509,3.450165,3.415869,3.4295874,3.2443898,2.2395205,1.8554068,3.2272418,5.171818,6.2247014,4.6265135,3.5050385,2.8054025,2.6647894,2.959734,3.3061223,2.5378947,2.7916842,4.461893,6.39961,5.919468,9.788043,13.001566,13.426835,10.738038,6.4304767,4.3933015,3.4535947,3.0420442,2.7128036,2.1640697,3.0454736,4.540774,5.638242,6.012067,6.0154963,6.8797526,7.3084507,7.425057,7.3427467,7.140401,7.140401,7.5931067,8.357904,9.019815,8.865483,8.220721,8.2653055,8.347616,8.467651,9.277034,12.932974,13.193623,12.38767,11.05699,7.9772205,6.3207297,6.9037595,8.207003,9.266746,9.6645775,9.448513,9.256456,8.484799,6.992929,5.127233,4.852866,5.518206,6.186976,6.108095,4.729401,4.506478,4.5613513,4.8185706,4.99005,4.57164,3.5359046,2.9048605,2.0886188,1.3786942,1.9239986,0.5761707,0.32238123,0.32924038,0.22978236,0.14404267,0.1371835,0.09602845,0.082310095,0.09945804,0.06859175,0.058302987,0.05144381,0.08573969,0.11317638,0.020577524,0.030866288,0.061732575,0.05144381,0.0274367,0.12003556,0.0548734,0.020577524,0.0034295875,0.006859175,0.0274367,0.044584636,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.12689474,0.14061308,0.09259886,0.034295876,0.017147938,0.024007112,0.020577524,0.037725464,0.15433143,0.07545093,0.0274367,0.010288762,0.01371835,0.010288762,0.0274367,0.048014224,0.061732575,0.06859175,0.082310095,0.037725464,0.01371835,0.037725464,0.08916927,0.1097468,0.07545093,0.06516216,0.08916927,0.12689474,0.13375391,0.08916927,0.06859175,0.058302987,0.048014224,0.048014224,0.05144381,0.037725464,0.024007112,0.01371835,0.01371835,0.037725464,0.061732575,0.07888051,0.07888051,0.07888051,0.18519773,0.2469303,0.2469303,0.20920484,0.19548649,0.20577525,0.1920569,0.15776102,0.12003556,0.1097468,0.20920484,0.26064864,0.2777966,0.26407823,0.2194936,0.16119061,0.12003556,0.10288762,0.13375391,0.25378948,0.3566771,0.48014224,0.6276145,0.77508676,0.84367853,0.7579388,0.6001778,0.53844523,0.6036074,0.69963586,0.58988905,0.41498008,0.37039545,0.4698535,0.5453044,0.34638834,0.48700142,0.7682276,1.0288762,1.1660597,1.4987297,1.7696671,1.529596,0.83338976,0.23321195,0.5041494,0.84367853,0.7339317,0.2777966,0.23321195,0.37039545,1.0254467,2.1332035,3.4227283,4.413879,4.7362604,4.633373,3.5873485,2.1091962,1.7456601,1.5536032,1.9925903,2.8019729,3.7759757,4.7602673,5.6348124,5.4736214,4.280125,2.6750782,1.9102802,1.8348293,2.0131679,2.0886188,2.1229146,2.5893385,2.1469216,1.3306799,1.7456601,3.216953,3.7759757,1.0734608,1.2072148,2.3801336,2.8225505,0.78194594,0.3018037,0.106317215,0.16119061,0.39783216,0.70306545,0.99801,1.8108221,2.2258022,1.7525192,0.32924038,0.44584638,0.34295875,0.2194936,0.17147937,0.20577525,0.47328308,2.136633,5.4941993,9.688584,12.706621,11.235329,9.630281,8.488229,8.320179,9.530824,10.31277,8.251588,5.8200097,4.5339146,4.962613,5.576509,5.686256,7.3530354,10.247607,11.653738,8.820899,7.7542973,8.2653055,9.685155,10.858074,10.377932,10.089847,10.034973,10.477389,11.880091,11.626302,10.717461,11.2250395,14.263655,20.015072,23.839062,25.43725,29.189219,34.690277,36.73088,31.888304,28.372976,25.896814,24.885086,26.469557,29.923151,31.58993,31.781986,30.286688,26.376957,27.85854,29.298965,28.654203,26.051146,23.76704,22.662714,21.829325,21.181131,20.19341,17.905876,19.12681,19.665255,17.55263,13.560589,11.194174,12.109874,12.106443,13.625751,16.47231,17.806417,17.734396,16.835844,14.143619,10.64201,9.266746,10.100135,8.97866,8.158989,8.539673,9.678296,9.585697,10.834066,11.105004,9.644,7.267296,8.285883,9.122703,9.801761,10.803201,13.066729,14.181344,14.466,13.440554,11.345076,9.132992,10.275044,12.185325,12.860953,11.80464,10.028113,11.091286,11.574858,11.897239,11.8869505,10.792912,9.499957,8.536243,8.505377,8.951223,8.357904,8.31332,8.388771,7.9292064,6.783724,5.3261495,4.4275975,3.2615378,2.4418662,1.9720128,1.2243627,0.7099246,0.34295875,0.116605975,0.030866288,0.09259886,0.048014224,0.06516216,0.072021335,0.044584636,0.0274367,0.061732575,0.058302987,0.10288762,0.18176813,0.20920484,0.20577525,0.24007112,0.274367,0.29494452,0.29151493,0.39783216,0.432128,0.4424168,0.432128,0.37039545,0.2503599,0.14747226,0.072021335,0.034295876,0.034295876,0.0274367,0.024007112,0.0274367,0.0274367,0.020577524,0.034295876,0.061732575,0.08916927,0.1097468,0.11317638,0.116605975,0.09602845,0.082310095,0.07888051,0.0548734,0.17833854,0.26064864,0.18176813,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.0034295875,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.044584636,0.044584636,0.0,0.0034295875,0.01371835,0.09259886,0.2194936,0.26064864,0.14747226,0.1371835,0.09602845,0.017147938,0.030866288,0.09945804,0.116605975,0.08573969,0.061732575,0.13375391,0.07545093,0.037725464,0.01371835,0.0,0.0,0.216064,0.28465575,0.28465575,0.26750782,0.26407823,0.36010668,0.53501564,0.6173257,0.71678376,1.2380811,1.0254467,0.89512235,0.8025235,0.7339317,0.6962063,0.980862,1.7765263,3.350707,6.351596,11.814929,16.647217,20.272291,23.550978,27.261791,32.0735,48.63155,69.17135,88.87433,105.75476,120.6666,131.16115,129.09311,117.5251,101.54665,88.274155,69.65492,50.991108,36.826912,29.295536,28.126047,31.32928,34.529087,36.4085,34.947495,27.405834,18.914175,12.082437,8.255017,7.64798,9.349055,10.2921915,10.329918,9.033533,6.680836,4.280125,2.633923,2.1229146,1.7216529,1.1454822,0.85396725,0.70306545,0.6241849,0.58645946,0.61389613,0.75450927,1.8862731,2.0577524,2.5001693,2.9974594,3.1312134,2.2841053,2.1057668,2.054323,2.0577524,2.1503513,2.4590142,2.2086544,2.5721905,3.532475,4.479041,4.2286816,4.955754,6.1046658,6.2864337,5.6313825,5.7891436,7.689135,17.463459,33.315014,56.653355,92.11872,113.38902,97.73638,69.07875,45.16081,37.526546,39.628883,47.36946,62.58997,79.47726,84.57706,49.73245,33.592808,29.405283,31.226395,33.92548,36.66229,37.852356,31.404732,20.141968,15.769243,14.767803,11.156448,7.949784,6.6396813,7.181556,6.1458206,4.955754,4.386442,4.355576,3.9063,3.0557625,2.3389788,2.3561265,2.9082901,3.0111778,2.74367,4.3795834,5.254128,4.5339146,3.223812,4.2835546,6.557371,7.1712675,5.892031,5.147811,4.0091877,3.309552,3.4398763,4.1463714,4.5442033,6.824879,10.357354,12.524854,11.694893,7.2192817,5.363875,4.623084,3.998899,3.1483612,2.3972816,1.3272504,1.4164196,1.6564908,1.5947582,1.3169615,1.3581166,1.7799559,2.0508933,2.218943,2.8945718,3.3952916,4.15323,4.0777793,3.0146074,1.7662375,1.5193073,1.6942163,2.5070283,3.758828,4.852866,4.7945633,4.938606,4.856296,4.400161,3.683377,3.426158,3.4192986,3.0660512,2.6476414,3.2992632,3.590778,4.0606318,4.40702,4.513337,4.417309,4.8837323,4.911169,4.7774153,4.647091,4.5819287,4.0263357,3.1140654,2.4452958,2.1503513,1.8588364,1.762808,1.8931323,2.2258022,2.668219,3.07634,2.9460156,2.9117198,3.2375305,3.5804894,3.0111778,2.6579304,3.1346428,3.5221863,3.4947495,3.2992632,2.4555845,1.8073926,1.8828435,2.551613,3.0248961,2.2498093,2.3046827,4.2595477,6.3310184,3.8891523,4.245829,6.0806584,7.0889573,6.293293,4.064061,2.8980014,2.6167753,2.627064,2.551613,2.2292318,2.534465,3.2409601,4.057202,4.756838,5.161529,6.355026,7.14726,7.5862474,7.641121,7.2192817,7.332458,7.7097125,8.39563,9.098696,9.184435,7.840037,8.021805,8.735159,9.39021,9.791472,12.13731,12.768354,11.749766,9.403929,6.3035817,6.5882373,6.8797526,7.6171136,8.796892,9.9801,9.424506,9.328478,9.273604,8.783174,7.3084507,6.159539,5.9469047,6.0978065,6.0566516,5.302142,4.962613,5.535354,5.802862,5.2987127,4.297273,3.0043187,2.6956558,2.4007113,1.8313997,1.3786942,0.48700142,0.45956472,0.5007198,0.31552204,0.08916927,0.15776102,0.16119061,0.13032432,0.09259886,0.06859175,0.061732575,0.061732575,0.12689474,0.18519773,0.041155048,0.058302987,0.048014224,0.041155048,0.08916927,0.26064864,0.13375391,0.061732575,0.020577524,0.0,0.0,0.07888051,0.041155048,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.07545093,0.12689474,0.12689474,0.07545093,0.01371835,0.024007112,0.048014224,0.041155048,0.010288762,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.020577524,0.024007112,0.0274367,0.048014224,0.12003556,0.037725464,0.01371835,0.061732575,0.14404267,0.16462019,0.13375391,0.16462019,0.2194936,0.26407823,0.26064864,0.18519773,0.13375391,0.08573969,0.041155048,0.034295876,0.020577524,0.006859175,0.006859175,0.01371835,0.01371835,0.08573969,0.12689474,0.14061308,0.1371835,0.12689474,0.14404267,0.1371835,0.11317638,0.08573969,0.10288762,0.12346515,0.12346515,0.12346515,0.13032432,0.14404267,0.22978236,0.2503599,0.2194936,0.17147937,0.16119061,0.13375391,0.14404267,0.17833854,0.2469303,0.39783216,0.4972902,0.53501564,0.5761707,0.6241849,0.6310441,0.432128,0.39783216,0.51100856,0.64133286,0.5453044,0.34981793,0.26750782,0.26750782,0.32581082,0.4389872,0.2777966,0.47328308,0.88826317,1.2346514,1.0666018,1.1934965,1.3375391,1.1626302,0.66533995,0.19548649,0.32581082,0.47328308,0.42526886,0.24350071,0.26750782,0.18176813,0.65162164,1.6839274,3.1792276,4.9248877,6.3310184,6.6293926,5.3501563,3.1415021,1.786815,1.097468,0.864256,0.8505377,0.97057325,1.2998136,1.9308578,2.277246,2.0474637,1.4815818,1.3615463,1.6256244,1.3615463,1.3478279,2.0474637,3.642222,2.4967396,1.3375391,0.65505123,0.4972902,0.4389872,0.70649505,1.8005334,3.2786856,3.6936657,0.5761707,0.4355576,0.26064864,0.31209245,0.6927767,1.3581166,2.2052248,3.1140654,3.0317552,1.8073926,0.2194936,0.17833854,0.15433143,0.15090185,0.14061308,0.061732575,0.01371835,0.36010668,1.4953002,3.426158,5.7822843,4.9008803,3.882293,3.5359046,4.8288593,8.8929205,11.465111,8.285883,4.197815,1.9068506,1.9754424,2.8499873,4.187526,6.691125,9.9801,12.600305,10.621432,8.299602,7.606825,8.882631,10.837497,13.454271,15.62863,15.018164,11.900668,9.170717,7.6274023,7.1266828,9.280463,13.598314,17.487467,20.138538,23.921373,29.827122,36.034676,37.896942,33.856888,28.76395,25.008553,23.883648,25.564144,27.066305,28.146624,28.558174,28.088322,26.555296,28.472435,28.304386,26.822803,25.478405,26.407824,28.232365,26.69248,23.791048,21.386908,21.160555,22.415783,20.265432,16.029892,11.640019,9.640571,8.934075,9.349055,13.004995,18.972477,23.297188,22.487804,19.833303,15.937293,11.89038,9.239308,10.131001,8.580828,7.4181976,7.5450926,7.9463544,6.8626046,8.848335,10.738038,10.988399,9.685155,10.175586,10.659158,10.539123,10.738038,13.694343,14.781522,15.556609,15.388559,13.786942,10.398509,9.39707,10.377932,11.002116,10.350495,8.934075,9.89093,10.844356,11.417097,10.902658,8.255017,7.222711,6.927767,6.7494283,6.677407,7.3221693,7.764586,8.128122,7.795452,6.773435,5.693115,5.411889,4.245829,3.1312134,2.277246,1.1763484,0.71678376,0.3566771,0.18862732,0.22635277,0.4081209,0.21263443,0.20234565,0.18519773,0.1097468,0.06859175,0.07545093,0.10288762,0.18519773,0.28122616,0.29151493,0.29151493,0.3018037,0.33266997,0.37039545,0.39440256,0.50757897,0.5453044,0.58302987,0.64133286,0.6824879,0.4938606,0.28122616,0.13375391,0.06859175,0.041155048,0.037725464,0.030866288,0.030866288,0.041155048,0.044584636,0.07888051,0.11317638,0.1371835,0.14747226,0.14747226,0.16119061,0.116605975,0.08573969,0.06859175,0.01371835,0.29837412,0.5658819,0.47671264,0.20577525,0.44927597,0.36010668,0.31895164,0.2709374,0.18862732,0.082310095,0.017147938,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.01371835,0.030866288,0.0274367,0.024007112,0.06859175,0.19548649,0.25378948,0.18176813,0.041155048,0.030866288,0.15090185,0.22978236,0.2194936,0.16119061,0.18519773,0.216064,0.17147937,0.09259886,0.020577524,0.010288762,0.08573969,0.15433143,0.2469303,0.32581082,0.26750782,0.28808534,0.47671264,0.5796003,0.6824879,1.2380811,0.6379033,0.490431,0.58302987,0.66191036,0.42869842,0.67219913,0.9602845,1.7113642,3.9337368,9.239308,16.064188,19.397747,20.502073,19.764713,16.695232,17.778982,24.19917,34.018078,46.673256,62.994663,92.420525,115.5428,126.79185,126.12651,119.0204,99.40659,76.48666,56.677364,43.257385,36.40164,34.072952,35.362476,37.420227,37.07041,30.783978,20.406046,12.1921835,7.407909,6.1732574,7.466212,10.700313,11.958971,11.026124,8.327039,4.9420357,2.7470996,1.8245405,1.3649758,0.99801,0.805953,0.6756287,0.5521636,0.4629943,0.4424168,0.52472687,0.823101,1.2380811,1.371835,1.1763484,0.78194594,0.48700142,0.48700142,0.6241849,0.9842916,1.5673214,2.287535,1.8142518,1.7490896,2.1194851,2.7539587,3.2649672,3.9611735,4.4756117,4.846007,5.7754254,8.621983,16.506605,28.393555,37.64658,46.831017,67.70348,87.18697,75.872765,57.1335,43.373993,36.027817,35.537384,40.781223,46.127953,47.846176,44.087345,36.710304,31.974045,30.300406,30.900583,31.75455,33.476204,32.32043,27.169191,20.20027,16.890718,14.915276,12.524854,11.2421875,11.146159,10.878652,6.776865,4.681387,4.1635194,4.4550343,4.4550343,3.1243541,2.5893385,2.335549,1.961724,1.2072148,3.3781435,4.3521466,3.642222,3.3609958,8.193284,12.696333,13.989287,9.949233,3.6113555,3.1586502,2.4384367,2.3218307,2.8705647,3.8479972,4.715683,8.155559,6.334448,4.57164,4.7431192,5.2781353,4.0091877,3.7005248,3.57363,3.0557625,1.786815,0.9911508,0.84024894,0.8711152,0.91227025,1.0837497,1.3512574,1.786815,2.2909644,3.0317552,4.4104495,6.166398,5.535354,4.149801,3.1826572,3.340418,2.4007113,2.3218307,2.6887965,3.2889743,4.1189346,5.305572,5.0243454,4.180667,3.292404,2.486451,2.9151495,2.4898806,2.0508933,2.054323,2.5790498,2.0303159,2.6716487,3.2203827,3.4192986,4.029765,4.540774,4.5682106,4.506478,4.4584637,4.2252517,3.7519686,3.309552,2.836269,2.335549,1.9068506,1.821111,1.9480057,2.2841053,2.7230926,3.0523329,2.9288676,3.0454736,3.5461934,4.122364,4.012617,3.9508848,4.557922,4.5270553,3.5804894,2.4555845,1.7113642,1.4267083,1.5844694,2.1091962,2.8534167,1.961724,2.1057668,2.4967396,2.7882545,3.083199,2.5207467,2.5550427,2.585909,2.3424082,1.8931323,1.7216529,2.4212887,2.644212,2.2052248,2.061182,2.7573884,3.542764,3.8925817,3.806842,3.8308492,4.232111,5.120374,6.385892,7.5759587,7.905199,8.025234,7.8194594,7.6857057,7.864044,8.436785,9.4862385,10.398509,10.55284,10.511685,12.024134,12.243628,12.188754,10.5597,8.025234,7.233,7.0375133,6.7700057,7.380472,8.611694,9.002667,6.6225333,6.420188,8.1041155,10.593996,12.006986,10.017825,7.3427467,5.9640527,6.48535,8.131552,7.8023114,8.076678,7.1266828,4.8082814,2.6853669,2.1846473,3.1209247,4.1120753,4.0537724,2.136633,0.805953,0.5658819,0.51100856,0.30866286,0.19891608,0.45613512,0.47328308,0.29494452,0.06859175,0.030866288,0.10288762,0.09602845,0.09602845,0.116605975,0.09259886,0.07888051,0.15090185,0.18519773,0.17490897,0.19891608,0.19891608,0.14404267,0.06516216,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0274367,0.020577524,0.020577524,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.01371835,0.006859175,0.01371835,0.034295876,0.044584636,0.020577524,0.006859175,0.0548734,0.12689474,0.09259886,0.12689474,0.29151493,0.37725464,0.30866286,0.1371835,0.06516216,0.0274367,0.020577524,0.034295876,0.044584636,0.020577524,0.006859175,0.006859175,0.01371835,0.01371835,0.07545093,0.16462019,0.23664154,0.26407823,0.21263443,0.09259886,0.05144381,0.044584636,0.041155048,0.030866288,0.030866288,0.048014224,0.09259886,0.14404267,0.16804978,0.20577525,0.21263443,0.18176813,0.12346515,0.07545093,0.08916927,0.17490897,0.216064,0.21263443,0.274367,0.33609957,0.37725464,0.432128,0.48357183,0.47328308,0.20577525,0.2469303,0.37382504,0.4115505,0.22978236,0.13032432,0.07888051,0.048014224,0.048014224,0.12346515,0.14747226,0.22635277,0.5693115,0.9328478,0.64133286,0.922559,1.1283343,1.0734608,0.7442205,0.30523327,0.2194936,0.22635277,0.37725464,0.5624523,0.48700142,0.20920484,0.3566771,0.7339317,1.3992717,2.6545007,4.839148,5.7891436,5.1238036,3.2512488,1.3581166,0.65162164,0.5007198,0.42869842,0.28808534,0.274367,0.5418748,1.0048691,1.371835,1.6187652,1.9823016,3.5461934,2.8122618,1.4129901,0.39440256,0.19891608,0.19891608,0.14404267,0.13032432,0.29151493,0.7922347,0.85396725,0.84367853,1.313532,1.786815,0.7476501,0.28465575,0.24007112,0.5144381,1.0768905,1.9685832,2.884283,3.2683969,2.5790498,1.1111864,0.0,0.08573969,0.15090185,0.14061308,0.061732575,0.0,0.0,0.010288762,0.08916927,0.25378948,0.47328308,0.51100856,0.44584638,0.5144381,1.4953002,4.729401,5.2438393,3.9714622,2.4247184,1.3889829,0.90198153,1.3272504,3.841138,7.8331776,11.989838,14.29795,12.747777,10.666017,8.786603,7.8091707,8.4093485,11.629731,14.88098,16.026463,14.7369375,12.466551,11.050131,10.412228,9.997248,9.846346,10.590566,14.177915,19.54522,27.251501,34.978363,37.50597,33.42819,28.242653,24.044838,22.511812,24.915953,24.758192,25.313786,26.054577,26.164322,24.566135,25.982555,25.385807,23.571554,22.758743,26.565584,28.568464,26.476416,22.648996,19.099373,17.487467,19.36688,19.644676,16.702091,11.629731,8.224151,8.505377,12.812939,18.410025,23.554407,27.495003,26.43526,18.79757,13.145609,11.362224,8.652849,7.2604365,6.4990683,6.0052075,5.8234396,6.4098988,6.2144127,8.48137,11.231899,13.190193,13.762935,15.484588,15.107333,14.46257,14.376831,14.695783,16.475739,17.490896,17.03819,15.549749,14.572317,11.910957,12.315649,12.871242,12.061859,9.764035,8.289313,8.488229,8.700864,8.169277,7.034084,6.461343,6.7185616,6.2144127,5.576509,7.675417,8.529384,6.307011,5.15467,5.6793966,4.9591837,4.9351764,4.57164,3.4295874,1.762808,0.5178677,0.36010668,0.3018037,0.51100856,0.89855194,1.1283343,0.59331864,0.3566771,0.22292319,0.12689474,0.15090185,0.14061308,0.15433143,0.2469303,0.34981793,0.29151493,0.25378948,0.32581082,0.47328308,0.61389613,0.6241849,0.7099246,0.84367853,0.86082643,0.7682276,0.7339317,0.61046654,0.38754338,0.22978236,0.17833854,0.15090185,0.12689474,0.09602845,0.07545093,0.082310095,0.106317215,0.13032432,0.15433143,0.17833854,0.20920484,0.24350071,0.26750782,0.2194936,0.15090185,0.09602845,0.061732575,0.31895164,0.7099246,0.8265306,0.97400284,2.1812177,1.6942163,1.471293,1.2758065,0.91227025,0.22978236,0.044584636,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.017147938,0.0,0.0,0.01371835,0.01371835,0.010288762,0.006859175,0.030866288,0.030866288,0.10288762,0.12689474,0.07888051,0.030866288,0.09259886,0.13375391,0.23321195,0.3806842,0.5041494,0.5041494,0.4664239,0.30866286,0.09602845,0.044584636,0.082310095,0.082310095,0.08916927,0.08573969,0.0,0.0,0.12003556,0.40126175,0.6790583,0.5796003,0.31209245,0.40126175,0.4972902,0.45613512,0.31895164,0.65162164,0.66876954,1.0220171,2.5961976,6.5162163,12.373952,17.429163,20.097382,19.222837,14.085316,14.267084,11.595435,9.952662,10.786053,13.080446,24.898806,45.30485,67.91612,89.12469,108.093735,108.62875,98.5149,85.04691,71.969894,59.50677,45.335716,40.15361,39.930687,40.524006,37.704884,25.910534,14.970149,7.795452,5.086078,5.3570156,8.968371,12.96727,14.400838,12.144169,6.883182,2.9391565,1.4129901,0.96714365,0.82996017,0.7922347,0.78194594,0.5658819,0.36696586,0.28122616,0.30523327,2.1297739,2.3972816,2.7573884,3.2581081,3.5461934,2.843128,2.5413244,2.1640697,1.5433143,0.9911508,1.2998136,1.1934965,1.5227368,2.153781,2.860276,3.3129816,4.712253,6.118384,6.2898636,6.6053853,11.050131,22.930222,33.911762,37.0807,35.537384,42.386272,51.851933,51.917095,49.54039,46.46405,39.210472,35.75345,36.291893,39.16589,41.882122,41.14133,34.957787,30.83542,29.919722,31.120077,31.106358,29.01088,25.9414,22.796469,19.994495,17.477179,14.904987,13.13532,12.603734,12.061859,8.56025,6.138962,6.3893213,6.694555,5.8543057,4.0777793,3.8514268,3.1963756,2.3972816,1.6530612,1.0700313,1.3581166,1.3272504,1.3306799,2.3081124,5.7651367,4.65395,4.0880685,3.2306714,2.2978237,2.5619018,2.534465,7.140401,9.901219,9.650859,10.539123,6.23499,4.3007026,4.139512,4.6093655,4.0229063,3.525616,3.8102717,3.6936657,2.750529,1.3341095,1.2243627,0.9259886,0.7476501,0.9431366,1.7182233,1.99602,2.0817597,2.2600982,2.952875,4.7019644,5.6485305,4.2869844,3.0043187,2.6407824,2.486451,2.6304936,2.170929,2.270387,3.1449318,4.0846386,3.7725463,3.508468,3.2855449,3.0626216,2.7573884,2.7539587,2.6476414,2.294394,2.085189,2.9322972,2.4418662,2.6785078,2.9665933,3.2066643,3.9063,3.9714622,3.5564823,3.1586502,3.1072063,3.5804894,3.3266997,3.0386145,2.7333813,2.4212887,2.1023371,1.920569,1.9308578,2.1812177,2.5824795,2.942586,3.1517909,3.3438478,3.8137012,4.448175,4.7088237,4.32471,4.5682106,4.945465,5.0174866,4.372724,2.8945718,1.9342873,1.7216529,2.1297739,2.6579304,1.845118,1.5536032,1.5055889,1.5090185,1.4575747,1.5330256,1.9068506,2.1297739,2.0749004,1.9651536,2.1469216,2.301253,2.085189,1.6084765,1.4610043,1.8073926,2.1846473,2.4247184,2.568761,2.867135,3.0454736,3.6182148,4.1463714,4.482471,4.791134,6.475061,7.5519514,7.8091707,7.394191,6.8145905,7.6788464,9.798331,11.640019,12.38424,11.924676,9.030104,9.455373,9.866923,9.506817,10.199594,9.016385,8.457363,9.040393,9.990388,9.259886,7.0923867,6.931196,8.937505,12.055,13.999576,14.273943,12.099585,9.685155,8.251588,8.035523,8.008087,6.893471,5.6793966,4.530485,2.7951138,1.8554068,2.4041407,3.642222,4.629943,4.2835546,1.8519772,0.83681935,0.4046913,0.15776102,0.12346515,0.16804978,0.16119061,0.1097468,0.044584636,0.017147938,0.072021335,0.05144381,0.06859175,0.2194936,0.5693115,0.6241849,0.39440256,0.19891608,0.18176813,0.33266997,0.15776102,0.08573969,0.072021335,0.058302987,0.0,0.0034295875,0.017147938,0.0548734,0.08916927,0.061732575,0.030866288,0.017147938,0.006859175,0.0034295875,0.0034295875,0.006859175,0.0034295875,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0034295875,0.0,0.01371835,0.034295876,0.044584636,0.020577524,0.0274367,0.058302987,0.106317215,0.17833854,0.14404267,0.1920569,0.17490897,0.082310095,0.0274367,0.024007112,0.017147938,0.017147938,0.020577524,0.034295876,0.0274367,0.017147938,0.01371835,0.034295876,0.11317638,0.26064864,0.25378948,0.24007112,0.25721905,0.23664154,0.1371835,0.06516216,0.044584636,0.0548734,0.041155048,0.024007112,0.07888051,0.18519773,0.26407823,0.17833854,0.06859175,0.05144381,0.048014224,0.037725464,0.0274367,0.07888051,0.09945804,0.09602845,0.08916927,0.14061308,0.28808534,0.29494452,0.29151493,0.33952916,0.42526886,0.25378948,0.19548649,0.22978236,0.28465575,0.22978236,0.17147937,0.12689474,0.09602845,0.09259886,0.14747226,0.18176813,0.2194936,0.28122616,0.32238123,0.22635277,0.3018037,0.44927597,0.5453044,0.5796003,0.64819205,1.196926,0.9877212,0.59674823,0.3841138,0.48700142,0.2469303,0.15776102,0.2194936,0.432128,0.8128122,1.5227368,1.8828435,1.7593783,1.3272504,1.0768905,1.1797781,1.3272504,1.2003556,0.8471081,0.6893471,0.96714365,1.138623,1.2655178,1.3889829,1.5330256,1.9239986,2.1915064,1.9857311,1.3375391,0.6756287,2.7162333,2.527606,1.5193073,0.66191036,0.48700142,0.548734,0.939707,1.3546871,1.371835,0.42869842,0.42526886,1.2449403,2.3972816,3.175798,2.6407824,1.7182233,1.2346514,0.823101,0.39440256,0.12346515,0.19891608,0.1097468,0.16462019,0.37382504,0.4389872,0.08916927,0.0034295875,0.017147938,0.12003556,0.4355576,0.25721905,0.16804978,0.21263443,0.53844523,1.4095604,1.6393428,1.5776103,1.2586586,0.82996017,0.5453044,0.8745448,2.8980014,5.305572,8.052671,12.332796,12.274493,10.340206,8.656279,8.285883,9.225591,10.864933,12.322508,13.05301,13.039291,12.758065,11.530273,9.304471,7.829748,8.028665,10.0041065,12.6757555,17.062197,22.889067,28.93886,33.08866,33.404182,29.391565,23.94538,20.910194,25.053137,25.468117,26.01342,26.740494,27.251501,26.726774,26.726774,24.302057,21.585823,20.7833,24.171732,22.77589,22.597551,21.208569,18.45461,16.462019,17.422304,19.03764,17.833855,14.143619,12.106443,11.828648,14.915276,20.563807,26.733635,30.156363,22.690151,16.70552,12.854094,10.415657,7.298162,5.0929375,4.945465,6.451054,8.244728,7.970361,6.6705475,9.338767,12.867812,14.887839,13.762935,11.842365,11.14273,11.273054,11.674315,11.629731,13.677195,16.53404,16.328266,12.97413,10.203023,10.645439,11.204462,11.050131,9.997248,8.532814,7.3873315,6.3378778,5.9297566,6.1972647,6.6431108,6.927767,8.076678,7.8983397,6.5333643,6.468202,7.058091,5.0414934,3.525616,3.4467354,3.566771,3.6010668,3.2821152,3.0283258,2.6407824,1.2860953,0.85396725,0.5761707,0.52472687,0.65162164,0.77508676,0.85396725,1.3203912,1.2072148,0.5693115,0.50757897,0.29837412,0.20577525,0.24007112,0.3566771,0.45956472,0.5212973,0.70649505,0.91227025,1.0837497,1.2243627,1.0837497,1.1660597,1.1214751,0.90884066,0.7922347,0.7990939,0.65162164,0.4424168,0.28808534,0.31209245,0.28808534,0.22292319,0.1920569,0.20920484,0.25378948,0.22978236,0.2709374,0.30523327,0.30523327,0.29151493,0.29837412,0.22978236,0.14747226,0.10288762,0.13375391,0.116605975,0.216064,0.58988905,1.0631721,1.1214751,1.0425946,1.1694894,1.2209331,0.9774324,0.31552204,0.15090185,0.058302987,0.01371835,0.01371835,0.06516216,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.037725464,0.024007112,0.010288762,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.006859175,0.11317638,0.10288762,0.06516216,0.05144381,0.09259886,0.11317638,0.09602845,0.20234565,0.432128,0.61389613,0.5144381,0.5796003,0.6893471,0.70306545,0.44927597,0.3566771,0.2469303,0.16804978,0.13375391,0.09602845,0.07888051,0.08916927,0.16462019,0.26750782,0.28808534,0.20234565,0.3018037,0.36010668,0.31209245,0.23664154,0.6927767,1.1214751,1.9102802,3.9646032,8.724871,11.996697,16.101913,19.726988,20.718138,16.098484,9.513676,7.222711,8.47451,10.72432,9.609704,12.922686,19.658396,28.599329,39.453976,52.84651,61.43077,64.93238,72.01448,82.56389,87.71856,69.92243,53.19976,43.758106,41.347107,39.279064,26.93941,15.978448,8.827758,5.830299,5.2575574,6.7802944,11.612583,15.947581,16.341984,9.712592,3.4844608,1.2037852,0.66876954,0.5727411,0.53844523,0.48700142,0.34981793,0.23664154,0.18862732,0.18176813,11.893809,18.139088,23.050257,23.376068,18.193962,8.906639,8.471081,7.4936485,5.9640527,4.1017866,2.3629858,2.4658735,2.7162333,3.199805,3.7039545,3.7108135,4.787704,6.48535,6.7322803,6.427047,9.441654,17.185663,23.671013,26.075153,25.869379,28.798246,34.635403,39.467693,43.994747,46.45719,42.64349,39.3991,36.7446,36.154713,36.864635,35.91121,32.817722,30.50961,29.648783,29.5116,27.995722,25.289778,23.228596,22.237446,21.225718,17.597214,13.900118,12.123591,11.249047,10.151579,7.613684,7.1884155,7.2535777,6.550512,5.079219,4.1120753,4.729401,3.5359046,2.294394,2.1846473,3.7931237,8.340756,6.574519,4.605936,4.976331,6.667118,4.256118,2.9974594,2.5481834,2.6750782,3.2546785,6.636252,8.573969,8.471081,7.8331776,10.254466,6.8728933,5.4496145,4.671098,3.8720043,3.0214665,2.7093742,2.8396983,2.901431,2.5413244,1.587899,1.2517995,1.1214751,1.2998136,1.7422304,2.2600982,2.1915064,2.0131679,2.551613,3.8342788,5.06893,5.3878818,4.249259,3.275256,3.2135234,3.940596,3.4535947,3.1620796,3.642222,4.619654,4.9523244,4.787704,4.5784993,4.214963,3.8205605,3.7382503,3.7451096,3.9508848,3.6456516,3.1449318,3.7794054,3.882293,4.1600895,4.338428,4.3452873,4.297273,3.9474552,3.1449318,2.4487255,2.2086544,2.5481834,2.7059445,2.5413244,2.4452958,2.4452958,2.2326615,1.961724,1.8348293,1.9239986,2.2258022,2.6476414,2.8019729,2.9220085,3.1860867,3.5359046,3.683377,3.525616,3.6593697,4.0023284,4.3109913,4.173808,3.1380725,2.1983654,2.0063086,2.417859,2.5001693,1.5947582,1.2449403,1.0700313,0.90541106,0.8162418,1.097468,1.4061309,1.5364552,1.4747226,1.4061309,1.5158776,1.4747226,1.3443983,1.1797781,1.0185875,0.9842916,1.0700313,1.2655178,1.5227368,1.762808,1.8999915,2.452155,3.1209247,3.683377,3.957744,4.386442,5.394741,6.0875177,6.1904054,6.042933,6.9552035,8.783174,10.693454,11.921246,11.784062,9.506817,9.9698105,11.019264,11.784062,12.672326,10.525404,9.427936,8.868914,8.618553,8.711152,8.128122,7.5450926,7.7542973,9.554831,13.7526455,14.867262,12.703192,10.076128,8.700864,9.174147,10.47396,9.349055,7.589677,6.042933,4.588788,2.726522,2.668219,3.1380725,3.3369887,2.952875,1.4438564,0.6859175,0.39440256,0.32238123,0.24350071,0.18862732,0.13032432,0.09259886,0.09259886,0.16119061,0.106317215,0.22292319,0.6001778,0.9431366,0.5761707,0.7682276,0.47328308,0.19548649,0.12689474,0.16462019,0.09259886,0.044584636,0.030866288,0.044584636,0.072021335,0.030866288,0.048014224,0.072021335,0.06859175,0.030866288,0.024007112,0.017147938,0.010288762,0.0,0.0,0.006859175,0.024007112,0.044584636,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.037725464,0.09945804,0.116605975,0.12689474,0.15433143,0.216064,0.25721905,0.24350071,0.15776102,0.037725464,0.0,0.0034295875,0.006859175,0.006859175,0.010288762,0.020577524,0.0274367,0.020577524,0.024007112,0.0548734,0.14747226,0.3018037,0.25378948,0.20577525,0.20920484,0.16119061,0.1097468,0.044584636,0.030866288,0.058302987,0.0548734,0.05144381,0.13032432,0.20577525,0.20920484,0.09259886,0.048014224,0.044584636,0.044584636,0.041155048,0.07888051,0.12689474,0.09945804,0.061732575,0.0548734,0.13375391,0.14404267,0.18862732,0.30523327,0.4698535,0.58645946,0.4389872,0.31895164,0.28808534,0.30523327,0.23664154,0.19548649,0.16462019,0.14747226,0.14747226,0.14404267,0.13032432,0.12003556,0.116605975,0.14747226,0.30523327,0.41840968,0.41498008,0.41840968,0.48700142,0.6310441,1.4267083,1.2655178,0.77508676,0.39097297,0.33266997,0.18862732,0.106317215,0.09602845,0.15433143,0.24007112,0.39097297,0.4698535,0.5555932,0.7956643,1.4095604,1.4438564,1.3958421,1.2998136,1.2072148,1.1866373,1.1763484,1.0220171,0.980862,1.1214751,1.3443983,1.9720128,1.9720128,1.6427724,1.1592005,0.58302987,2.1229146,2.1880767,1.6324836,1.1420527,1.2175035,1.0734608,1.2620882,1.2860953,1.0048691,0.6241849,0.8025235,1.5604624,2.3389788,2.620205,1.9548649,1.2860953,0.85739684,0.5658819,0.35324752,0.19891608,0.19891608,0.16119061,0.26750782,0.48700142,0.58645946,0.48357183,0.23321195,0.07888051,0.09259886,0.17147937,0.07888051,0.12689474,0.35324752,0.6927767,1.0117283,1.3238207,1.5570327,1.6324836,1.6221949,1.7593783,1.7559488,2.1263442,3.1517909,5.192395,8.683716,8.611694,7.874333,8.049242,9.6645775,12.212761,12.528283,12.024134,11.739478,12.103014,12.922686,13.9309845,13.855534,13.471419,13.210771,13.179905,13.049581,15.453721,20.237995,25.667032,28.410702,28.818823,27.114319,24.418663,22.94394,25.982555,26.815945,26.826233,26.34266,26.071724,27.11089,25.073713,22.374628,20.258574,19.61724,21.013083,20.457489,20.875898,20.821026,19.69955,17.778982,17.165085,19.672113,20.29287,18.001905,15.776102,14.658057,16.976458,21.109112,25.056566,26.455837,21.678423,17.36057,13.821238,10.751757,7.2158523,5.717122,6.4544835,8.388771,10.024684,9.39707,8.779744,10.796341,13.409687,15.021593,14.459141,13.056439,12.075578,12.048141,12.641459,12.6757555,12.38767,13.22106,12.397959,9.822338,8.1041155,8.618553,8.076678,6.9071894,5.5559316,4.4516044,3.9165888,3.4776018,3.457024,3.940596,4.7602673,6.046363,7.7097125,7.781734,6.341307,5.5319247,6.6225333,4.9248877,3.1826572,2.5378947,2.5138876,3.1072063,2.9700227,2.7745364,2.568761,1.7833855,1.4781522,1.1008976,0.89169276,0.90198153,0.97057325,1.2312219,1.4438564,1.3032433,0.939707,0.90541106,0.77508676,0.70306545,0.6859175,0.7339317,0.8779744,0.8025235,0.84367853,0.89855194,0.96371406,1.1249046,1.2895249,1.1694894,1.0254467,0.94656616,0.864256,0.89169276,0.7956643,0.61046654,0.44927597,0.5144381,0.4629943,0.3841138,0.31895164,0.28465575,0.28122616,0.26750782,0.3566771,0.40126175,0.3566771,0.28808534,0.36010668,0.29494452,0.19891608,0.13032432,0.09602845,0.048014224,0.08916927,0.29837412,0.61389613,0.8265306,1.0185875,1.1866373,1.155771,0.90541106,0.5453044,0.29837412,0.14747226,0.061732575,0.0274367,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.024007112,0.020577524,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0548734,0.11317638,0.116605975,0.08573969,0.116605975,0.061732575,0.041155048,0.09259886,0.24007112,0.4938606,0.548734,0.70306545,0.8265306,0.78537554,0.42183927,0.30523327,0.25721905,0.22635277,0.20920484,0.21263443,0.2777966,0.36010668,0.37382504,0.3841138,0.6173257,0.65162164,0.5521636,0.4389872,0.4115505,0.53501564,1.1317638,1.5501735,2.435007,4.2869844,7.48336,8.344186,12.061859,15.597764,16.46888,12.764925,6.9860697,5.926327,7.805741,10.079557,9.403929,11.773774,14.38026,16.911295,20.255144,26.527859,32.296425,37.272755,50.277752,69.0033,79.99856,69.877846,63.87607,58.326996,51.87251,45.421455,33.640823,19.78872,9.757176,5.4187484,4.629943,5.7925735,11.084427,17.95389,20.965069,11.80464,4.6745276,1.5261664,0.53844523,0.432128,0.44584638,0.4081209,0.28122616,0.16119061,0.09945804,0.07888051,11.434244,19.973917,30.814844,33.77458,25.667032,10.30591,9.918367,8.549961,6.9689217,5.3261495,3.1552205,3.1517909,3.1277838,3.4604537,4.0674906,4.400161,3.923448,5.3501563,6.1629686,6.15268,7.4353456,11.46854,13.577737,15.584045,18.941612,24.723896,29.981453,35.211575,40.493137,44.1285,42.64692,40.331947,37.447666,35.25616,33.784866,31.816282,30.060333,28.746801,27.9237,27.200058,25.749342,23.173723,21.548098,21.009653,20.11453,15.837835,12.847235,11.766914,10.799771,9.22902,7.431916,7.6342616,7.0272245,5.785714,4.6402316,4.897451,5.689686,4.307562,2.9734523,4.0434837,9.9869585,20.423193,15.426285,9.174147,8.025234,10.508256,9.853205,9.325048,8.882631,7.9463544,5.394741,8.193284,7.5279446,5.73427,5.178677,8.23444,7.3187394,6.0737996,4.4927597,3.100347,2.9734523,2.5996273,2.4452958,2.3767042,2.2086544,1.6770682,1.2758065,1.2312219,1.5090185,1.9994495,2.5413244,2.2566686,2.136633,3.0420442,4.537344,4.897451,5.305572,4.4447455,3.4878905,3.2992632,4.4413157,4.232111,4.2389703,4.6882463,5.3227196,5.3673043,5.4736214,5.3673043,5.099797,4.852866,4.945465,4.90431,5.020916,4.6745276,4.0880685,4.3109913,4.588788,5.2266912,5.7308407,5.796003,5.2987127,4.557922,3.2992632,2.2429502,1.7456601,1.7902447,1.9411465,1.99602,2.2292318,2.527606,2.3732746,1.9239986,1.6839274,1.6221949,1.7422304,2.0646117,2.1983654,2.3218307,2.4761622,2.6236343,2.644212,2.6785078,2.7539587,2.8911421,3.0489032,3.1140654,2.6853669,2.1160555,1.9514352,2.1126258,1.8897027,1.2312219,1.0151579,0.86082643,0.65848076,0.5590228,0.7339317,0.83338976,0.8471081,0.85396725,1.0288762,1.1420527,1.0837497,1.0357354,1.0117283,0.85396725,0.59331864,0.548734,0.65162164,0.805953,0.90884066,1.1832076,1.6976458,2.3218307,2.8877127,3.1895163,3.1140654,3.8925817,4.6608095,5.0757895,5.3227196,6.1492505,7.284444,8.745448,10.127572,10.604284,9.325048,9.695444,11.015835,12.641459,14.006435,11.921246,10.521975,8.906639,7.48336,7.970361,8.615124,8.573969,8.64942,9.647429,12.394529,13.735497,11.753197,9.863494,9.438225,9.791472,11.444533,10.6488695,9.002667,7.449064,6.3001523,4.698535,4.184097,3.5564823,2.8088322,3.093488,1.762808,1.0425946,0.7407909,0.6036074,0.32924038,0.26407823,0.18176813,0.12346515,0.1371835,0.3018037,0.17147937,0.29151493,0.66876954,0.9602845,0.4972902,0.7407909,0.44584638,0.16804978,0.09945804,0.06859175,0.041155048,0.01371835,0.006859175,0.05144381,0.18862732,0.10288762,0.14404267,0.1371835,0.048014224,0.0,0.006859175,0.017147938,0.01371835,0.0,0.0,0.0274367,0.06516216,0.106317215,0.11317638,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.0274367,0.006859175,0.0,0.0,0.0,0.017147938,0.072021335,0.16119061,0.2503599,0.2469303,0.15776102,0.116605975,0.14404267,0.16119061,0.20234565,0.17833854,0.1097468,0.034295876,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.010288762,0.020577524,0.034295876,0.058302987,0.106317215,0.17147937,0.28808534,0.20920484,0.15433143,0.17147937,0.14404267,0.13375391,0.072021335,0.041155048,0.058302987,0.0548734,0.05144381,0.11317638,0.14404267,0.11317638,0.061732575,0.12003556,0.1371835,0.10288762,0.06516216,0.1097468,0.1371835,0.09602845,0.058302987,0.072021335,0.15776102,0.0548734,0.12346515,0.32238123,0.53844523,0.58645946,0.48357183,0.40126175,0.39097297,0.4081209,0.32924038,0.23321195,0.18862732,0.17833854,0.17490897,0.12003556,0.1097468,0.14404267,0.21263443,0.3566771,0.65848076,0.5761707,0.4424168,0.44584638,0.65162164,1.0151579,1.5158776,1.2586586,0.7373613,0.3018037,0.15433143,0.10288762,0.08916927,0.1097468,0.16462019,0.22978236,0.21263443,0.19891608,0.4115505,0.94999576,1.786815,1.4404267,1.1111864,1.0528834,1.2380811,1.3443983,1.1626302,0.9328478,0.89512235,1.1420527,1.6153357,2.6064866,2.170929,1.3924125,0.8162418,0.48357183,1.5124481,1.9823016,1.8931323,1.5433143,1.5158776,1.3375391,1.3958421,1.2723769,0.94999576,0.8093826,1.0906088,1.4267083,1.5981878,1.5261664,1.2723769,1.0082988,0.8128122,0.6241849,0.42869842,0.2469303,0.2709374,0.28808534,0.32924038,0.4081209,0.52472687,0.58988905,0.34295875,0.15433143,0.116605975,0.041155048,0.034295876,0.14747226,0.4389872,0.85396725,1.2312219,1.2449403,1.3546871,1.5158776,1.8073926,2.435007,2.4247184,1.8245405,2.5893385,4.98662,7.6205435,6.385892,6.327589,7.970361,10.88894,13.666906,13.351384,12.22648,11.543991,11.952112,13.485138,16.12249,17.336565,17.333136,16.407146,14.946142,13.05301,14.335675,18.276272,22.731306,23.931662,23.85964,24.161444,24.442669,24.720467,25.444109,25.334362,24.576424,23.674442,23.177153,23.671013,20.841602,19.661825,18.567787,17.075916,15.80011,16.235666,18.591793,20.11453,19.819586,18.506054,18.334574,20.217419,21.462358,21.016512,19.469769,16.54433,18.214539,21.877338,24.86108,24.422092,21.006224,16.03675,11.89038,9.403929,7.8983397,7.9772205,9.1981535,10.549411,11.293632,10.981539,11.286773,11.674315,12.751206,14.009865,13.848674,13.437123,12.590015,12.048141,11.873232,11.458252,10.072699,9.102125,8.114404,7.0203657,6.077229,5.720552,4.4996185,3.1723683,2.170929,1.6084765,1.6290541,1.8142518,2.1812177,2.7951138,3.7794054,4.9248877,6.464772,6.509357,5.2609873,5.007198,6.0497923,5.038064,3.542764,2.4795918,2.0989075,2.784825,2.784825,2.5756202,2.4075704,2.318401,2.411,1.9102802,1.5055889,1.4507155,1.5673214,1.5604624,1.471293,1.3546871,1.2380811,1.1249046,1.1694894,1.2106444,1.1729189,1.0837497,1.08032,1.097468,0.97057325,0.82996017,0.805953,1.0460242,1.2586586,1.0666018,0.9294182,0.94999576,0.8745448,0.85739684,0.823101,0.70306545,0.5555932,0.58988905,0.52472687,0.45956472,0.38754338,0.32238123,0.30523327,0.31895164,0.38754338,0.40126175,0.34295875,0.274367,0.38754338,0.32581082,0.22978236,0.14747226,0.06859175,0.0274367,0.1097468,0.2194936,0.37039545,0.66191036,0.88826317,0.99801,0.90541106,0.70649505,0.6756287,0.34638834,0.20234565,0.12346515,0.058302987,0.041155048,0.006859175,0.0034295875,0.024007112,0.044584636,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.041155048,0.17490897,0.09259886,0.05144381,0.020577524,0.0,0.0,0.0,0.072021335,0.09602845,0.06516216,0.072021335,0.01371835,0.010288762,0.024007112,0.08573969,0.28808534,0.51100856,0.6310441,0.69963586,0.6790583,0.42869842,0.33266997,0.30866286,0.28465575,0.25378948,0.26750782,0.35324752,0.5007198,0.5418748,0.5453044,0.83681935,0.9328478,0.77851635,0.6241849,0.7339317,1.3821237,1.7250825,1.961724,2.6990852,4.2355404,6.550512,6.725421,9.122703,11.533703,12.109874,9.39021,6.39961,6.341307,9.126132,12.788932,13.516005,13.13189,12.97413,13.320518,14.606613,17.439453,19.936192,22.494663,33.469345,51.097424,63.52282,60.36417,62.44936,65.77949,66.86667,62.723724,45.366585,26.061436,12.854094,7.606825,6.0086374,6.8728933,12.339656,18.663815,21.078245,13.817808,6.924337,2.510458,0.59331864,0.41840968,0.4629943,0.4355576,0.29494452,0.14747226,0.0548734,0.030866288,1.2723769,6.060081,18.351723,24.322634,18.917604,5.871454,5.579939,4.7191124,4.0434837,3.6868064,3.1792276,3.3678548,3.6285036,3.6182148,3.6627994,4.7602673,2.860276,3.6353626,5.130663,6.2830043,6.931196,9.568549,9.39707,10.182446,14.740367,24.92624,29.899143,34.103817,37.708313,39.944405,39.107586,37.2316,36.110126,34.525658,32.17982,29.703657,27.326952,25.684181,24.871368,24.6896,24.658733,21.94936,19.497204,17.878439,16.37285,12.977559,12.109874,12.298501,11.760056,9.952662,7.56567,7.1232533,6.258997,5.3878818,4.99005,5.597087,6.1286726,5.2575574,4.506478,6.560801,15.254805,27.073164,20.310017,12.250486,10.964391,15.316538,15.635489,15.88242,15.834405,14.092175,8.090397,6.835168,6.1629686,5.4941993,5.3501563,7.3358874,6.9792104,5.305572,3.508468,2.5790498,3.292404,2.935727,2.7985435,2.4898806,1.99602,1.6599203,1.6942163,1.6599203,1.6256244,1.8005334,2.527606,2.486451,2.603057,3.316411,4.2218223,4.0503426,5.099797,4.3041325,3.2786856,2.9803114,3.7348208,4.5442033,4.7534084,4.7602673,4.7842746,4.863155,4.73969,4.7979927,5.0277753,5.3570156,5.6485305,5.5147767,5.3432975,4.955754,4.4756117,4.2938433,4.190956,5.096367,6.090947,6.6225333,6.495639,5.6245236,4.0023284,2.551613,1.7216529,1.5261664,1.2929544,1.488441,1.9548649,2.3732746,2.2566686,1.7490896,1.5021594,1.3478279,1.2483698,1.3238207,1.5398848,1.7388009,1.9239986,2.0714707,2.1332035,2.1640697,2.177788,2.16064,2.1057668,2.0406046,1.9068506,1.7353712,1.5398848,1.3169615,1.0425946,0.83338976,0.7442205,0.64133286,0.490431,0.3566771,0.32581082,0.2709374,0.25378948,0.38754338,0.85739684,1.1077567,1.1626302,1.0837497,0.939707,0.8128122,0.5418748,0.48357183,0.4629943,0.432128,0.48357183,0.90541106,1.4472859,1.7799559,1.8759843,2.0303159,2.8122618,3.6319332,4.170378,4.400161,4.57507,5.178677,5.90575,6.914048,7.949784,8.357904,7.332458,7.8434668,9.534253,11.828648,13.9309845,12.775213,11.406808,9.465661,7.654839,7.7680154,8.549961,9.640571,11.190743,12.229909,10.662587,12.096155,10.734609,10.024684,10.580277,10.179015,10.88551,10.1652975,9.098696,8.176137,7.2878733,7.082098,6.3893213,5.1992545,4.3281393,5.4153185,3.1655092,2.1434922,1.5981878,1.1111864,0.58645946,0.5555932,0.39783216,0.2469303,0.20234565,0.33609957,0.25378948,0.274367,0.28122616,0.28808534,0.45613512,0.58302987,0.32238123,0.11317638,0.09602845,0.116605975,0.034295876,0.061732575,0.09259886,0.12689474,0.28808534,0.20234565,0.25721905,0.2194936,0.072021335,0.020577524,0.05144381,0.05144381,0.030866288,0.0034295875,0.0,0.06516216,0.11317638,0.16119061,0.15776102,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.09259886,0.044584636,0.0,0.0034295875,0.01371835,0.01371835,0.048014224,0.14747226,0.30523327,0.4629943,0.30866286,0.106317215,0.024007112,0.058302987,0.05144381,0.010288762,0.0,0.0034295875,0.010288762,0.0,0.0034295875,0.006859175,0.010288762,0.006859175,0.0034295875,0.017147938,0.0548734,0.106317215,0.15433143,0.18519773,0.24007112,0.14747226,0.09945804,0.16119061,0.26750782,0.2777966,0.20920484,0.1371835,0.09602845,0.072021335,0.030866288,0.037725464,0.048014224,0.06516216,0.12346515,0.22635277,0.23664154,0.16804978,0.09259886,0.12346515,0.12689474,0.08573969,0.061732575,0.08916927,0.15776102,0.058302987,0.09945804,0.26064864,0.42869842,0.3841138,0.3806842,0.4046913,0.45270553,0.4938606,0.48357183,0.35324752,0.26750782,0.22292319,0.18519773,0.09602845,0.14061308,0.25378948,0.4355576,0.69963586,1.0768905,0.5041494,0.30523327,0.45613512,0.89169276,1.5124481,1.4610043,1.0425946,0.52472687,0.13032432,0.041155048,0.041155048,0.058302987,0.11317638,0.20577525,0.33609957,0.25721905,0.23664154,0.5658819,1.2415106,1.9582944,1.3101025,0.8128122,0.7339317,0.9774324,1.097468,1.0117283,0.96714365,1.0700313,1.430138,2.177788,3.3266997,2.5584722,1.4575747,0.85739684,0.8265306,1.9308578,2.5653315,2.4761622,1.8382589,1.2415106,1.1729189,1.3203912,1.3375391,1.1317638,0.8711152,1.1077567,1.0563129,0.9362774,0.89169276,0.9842916,0.764798,0.69963586,0.59331864,0.4115505,0.2709374,0.41840968,0.4389872,0.3566771,0.29494452,0.4629943,0.42183927,0.3018037,0.20234565,0.17147937,0.17833854,0.14747226,0.18176813,0.32238123,0.5727411,0.90198153,0.44927597,0.40126175,0.5693115,0.9568549,1.7593783,1.99602,1.6496316,3.083199,6.478491,9.877212,7.6274023,6.725421,8.131552,11.026124,12.812939,12.55915,12.099585,11.856084,12.418536,14.544881,17.233677,17.700102,16.846134,15.4914465,14.359683,12.816368,14.05102,17.04505,20.03908,20.53294,20.687271,21.897917,23.389786,24.106571,22.731306,20.841602,19.476627,19.305147,19.600092,18.231688,15.827546,16.170506,15.573756,12.932974,9.750318,9.73317,13.937843,16.86671,17.315987,18.3723,20.917053,21.139977,21.37662,22.179142,22.350622,17.559488,18.708399,23.005672,26.747353,25.306927,19.44576,12.758065,8.340756,7.4353456,9.431366,11.080997,12.092726,12.212761,11.914387,12.425395,13.227919,12.195613,11.818358,12.367092,11.876661,11.489118,11.105004,10.158438,8.772884,7.7783046,7.1541195,6.334448,5.9228973,5.6828265,4.5442033,3.3678548,2.1297739,1.3443983,1.1317638,1.2209331,1.5741806,1.8485477,2.2806756,3.0283258,4.15323,4.420738,5.1066556,4.7362604,3.7519686,4.530485,5.103226,5.0106273,4.1429415,2.867135,2.0028791,2.3252604,2.3904223,2.3732746,2.4315774,2.7402403,3.1140654,2.6064866,2.1400626,2.0817597,2.2429502,1.7388009,1.6290541,1.5604624,1.3889829,1.2037852,1.313532,1.4610043,1.4438564,1.2380811,1.0254467,1.2620882,1.1180456,0.8848336,0.8093826,1.0837497,1.0460242,0.9431366,0.922559,0.9602845,0.88826317,0.7922347,0.83681935,0.78194594,0.61389613,0.5521636,0.50757897,0.47328308,0.42869842,0.3841138,0.38754338,0.4081209,0.37725464,0.35324752,0.35324752,0.34295875,0.3841138,0.31209245,0.2194936,0.15090185,0.09259886,0.0274367,0.16119061,0.3566771,0.490431,0.44584638,0.5590228,0.58988905,0.5178677,0.4389872,0.5418748,0.2469303,0.18519773,0.14747226,0.08573969,0.1097468,0.030866288,0.01371835,0.048014224,0.08916927,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06859175,0.34638834,0.23321195,0.17833854,0.12003556,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.058302987,0.08916927,0.1371835,0.432128,0.432128,0.44927597,0.548734,0.5418748,0.5041494,0.44584638,0.36696586,0.29837412,0.28122616,0.25721905,0.37725464,0.4698535,0.52815646,0.6962063,0.90198153,0.9431366,0.91569984,1.1180456,2.061182,1.9514352,2.0440342,2.4898806,3.625074,5.9812007,7.2604365,8.213862,9.338767,9.767465,7.2638664,6.3207297,7.164408,11.406808,17.226818,19.377169,13.207341,9.355915,9.499957,12.850664,16.160215,18.578075,19.332584,25.420103,37.56084,50.19887,50.421795,50.346344,60.007492,76.706154,85.01261,61.293587,34.779446,17.79613,12.034423,8.556821,8.371623,12.517994,15.518884,15.402277,13.701202,8.289313,3.3198407,0.77508676,0.58988905,0.66191036,0.58302987,0.39097297,0.1920569,0.058302987,0.0274367,1.1763484,1.2346514,1.7182233,2.5138876,2.9185789,1.6496316,1.2072148,2.8465576,3.4467354,2.8259802,3.7519686,5.8165803,8.134981,6.8111606,3.1380725,3.6010668,3.333559,3.4021509,4.746549,6.917478,8.100685,6.893471,6.756287,8.069819,12.123591,21.1194,23.952238,29.364128,32.98234,34.066093,35.50652,33.58938,32.85545,31.884874,30.118637,27.84825,26.126596,23.85621,22.299177,21.839613,21.973368,19.312008,16.925014,14.88098,13.224489,11.979549,11.489118,11.924676,11.509696,9.81205,7.7371492,7.2364297,6.2692857,5.267846,4.523626,4.180667,4.938606,5.1992545,6.0840883,7.9086285,10.179015,11.105004,10.762046,12.555719,16.170506,17.562918,11.629731,9.671436,9.599416,9.849775,9.383351,8.381912,7.9120584,8.210432,8.886061,8.9100685,7.421627,5.0895076,3.210094,2.3046827,2.1194851,2.1469216,2.5996273,2.7951138,2.6133456,2.503599,3.1140654,3.4124396,3.199805,2.6476414,2.318401,3.1483612,3.1380725,2.6785078,2.3424082,2.8534167,4.245829,3.6696587,3.3884325,4.029765,4.5784993,4.187526,4.482471,4.6848164,4.448175,3.875434,3.3026927,3.6079261,4.0709205,4.4275975,4.866585,5.1238036,5.2609873,5.07236,4.5853586,4.07435,3.707384,4.091498,4.9420357,5.98463,6.9723516,6.7048435,5.2747054,3.5461934,2.16064,1.5261664,1.1832076,1.0151579,1.0906088,1.2792361,1.2655178,1.3169615,1.3272504,1.155771,0.8848336,0.823101,0.922559,1.0563129,1.2037852,1.3512574,1.5090185,1.6084765,1.6770682,1.704505,1.6393428,1.4198492,1.2860953,1.2243627,1.2003556,1.1283343,0.8848336,0.5693115,0.37039545,0.2469303,0.17490897,0.1371835,0.12346515,0.11317638,0.11317638,0.12346515,0.1371835,0.26064864,0.6207553,0.7339317,0.5555932,0.45613512,0.32238123,0.23664154,0.22978236,0.31209245,0.45613512,0.7133542,1.7936742,2.5447538,2.4795918,1.786815,2.4212887,3.210094,3.758828,4.0503426,4.4413157,5.0620713,5.950334,6.40304,6.2727156,5.967482,5.562791,6.8557453,8.940934,11.050131,12.528283,11.869802,10.569988,9.126132,8.268735,8.940934,9.026674,9.688584,10.439664,10.528833,8.940934,10.443094,10.021255,9.791472,10.731179,12.696333,12.511135,11.423956,10.124143,8.985519,8.056101,8.594546,7.8949103,7.6857057,7.8434668,6.3790326,4.2183924,3.5393343,3.0386145,2.270387,1.646202,1.6359133,1.1489118,0.65848076,0.37382504,0.21263443,0.39783216,0.53501564,0.45956472,0.2709374,0.31895164,0.1371835,0.0548734,0.030866288,0.041155048,0.09259886,0.07888051,0.31552204,0.3806842,0.2503599,0.274367,0.28808534,0.24350071,0.17833854,0.12003556,0.106317215,0.25378948,0.18862732,0.07888051,0.01371835,0.0,0.12346515,0.17833854,0.16804978,0.09602845,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.01371835,0.061732575,0.072021335,0.058302987,0.044584636,0.037725464,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.017147938,0.041155048,0.01371835,0.041155048,0.072021335,0.10288762,0.12346515,0.1371835,0.11317638,0.05144381,0.034295876,0.15776102,0.548734,0.548734,0.51100856,0.39783216,0.24350071,0.18176813,0.061732575,0.01371835,0.024007112,0.08916927,0.19891608,0.2709374,0.24350071,0.20234565,0.19548649,0.24350071,0.2194936,0.14061308,0.07888051,0.072021335,0.12346515,0.061732575,0.044584636,0.12346515,0.2503599,0.274367,0.39783216,0.44584638,0.4389872,0.44584638,0.5796003,0.66533995,0.53844523,0.36353627,0.216064,0.106317215,0.14404267,0.18176813,0.34981793,0.7339317,1.3581166,0.34638834,0.1097468,0.32238123,0.65848076,0.7922347,0.67219913,0.5693115,0.39783216,0.17833854,0.030866288,0.030866288,0.041155048,0.082310095,0.18862732,0.39783216,0.29837412,0.26407823,0.59674823,1.2758065,1.9823016,1.3238207,0.764798,0.5418748,0.6241849,0.7339317,0.8779744,1.0700313,1.2586586,1.6187652,2.534465,4.2183924,2.6613598,1.313532,1.3992717,1.937717,2.3767042,2.3767042,2.3046827,2.1572106,1.5707511,1.3169615,1.3992717,1.3615463,1.1489118,1.1146159,0.78537554,0.6276145,0.59674823,0.607037,0.53501564,0.88826317,1.039165,0.85739684,0.4664239,0.26064864,0.45613512,0.53158605,0.4938606,0.47671264,0.7339317,0.6241849,0.40126175,0.26407823,0.29151493,0.47328308,0.40126175,0.30866286,0.18176813,0.048014224,0.0,0.072021335,0.12003556,0.15433143,0.18519773,0.19891608,0.2469303,0.6241849,2.335549,6.1561093,12.648318,11.746337,8.05953,6.914048,9.287323,11.825217,11.862943,11.732618,11.982979,13.152468,15.776102,17.658945,17.569777,16.45173,15.21365,14.723219,14.88441,15.656067,17.658945,19.847023,19.5315,19.421753,20.28258,21.019941,20.728426,18.677534,16.417435,15.121051,15.556609,16.852993,16.510035,13.810948,11.866373,10.412228,8.920357,6.5779486,5.562791,6.025785,8.021805,12.195613,19.775002,25.121729,24.699888,22.70044,21.668133,22.5221,18.296848,19.411465,22.957659,25.60187,23.574984,16.921585,12.284782,9.897789,9.932085,12.4974165,14.582606,14.778092,13.197053,11.482259,12.80265,13.9481325,13.999576,12.600305,10.679735,10.436234,9.911508,9.781183,8.89635,7.582818,7.6445503,7.010077,7.675417,7.840037,7.1198235,6.5470824,4.5201964,2.6956558,1.7250825,1.5981878,1.646202,2.0989075,2.6613598,3.216953,3.7622573,4.4104495,5.1066556,4.3178506,3.1209247,2.4795918,3.234101,4.4927597,5.0174866,4.6436615,3.357566,1.2826657,1.7696671,1.9754424,2.1469216,2.3389788,2.411,2.3252604,2.3321195,2.4418662,2.5619018,2.486451,1.7182233,1.6187652,1.4815818,1.2380811,1.4335675,1.2517995,1.3443983,1.3684053,1.2312219,1.097468,1.0117283,1.1111864,1.0494537,0.8162418,0.71678376,0.8162418,0.7476501,0.8093826,1.0117283,1.0837497,0.94999576,1.0357354,0.97400284,0.7339317,0.6241849,0.58988905,0.58988905,0.58302987,0.5590228,0.53501564,0.4972902,0.37725464,0.40126175,0.5624523,0.61046654,0.4389872,0.29494452,0.19891608,0.15090185,0.15090185,0.07888051,0.216064,0.4115505,0.53158605,0.45613512,0.59331864,0.4424168,0.28465575,0.20234565,0.09259886,0.07888051,0.058302987,0.041155048,0.048014224,0.12346515,0.061732575,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09259886,0.2503599,0.3806842,0.38754338,0.24350071,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1097468,0.18862732,0.19891608,0.19891608,0.45613512,0.44584638,0.3841138,0.3806842,0.4424168,0.5521636,0.5521636,0.51100856,0.45270553,0.36696586,0.15776102,0.13375391,0.23664154,0.37725464,0.42869842,1.0254467,1.3409687,1.4129901,1.2792361,0.9602845,0.99801,1.1729189,1.2517995,1.3924125,2.136633,4.870014,7.366754,8.790032,8.021805,3.6627994,4.173808,7.133542,11.423956,16.177364,20.766151,12.723769,7.881192,8.333898,12.583157,15.549749,17.977898,18.272842,20.165974,25.979126,36.638283,42.972733,40.170757,46.70412,67.374245,93.33622,80.41011,46.254845,21.688711,14.208781,8.056101,6.1046658,4.928317,5.161529,6.293293,6.684266,4.4756117,2.136633,0.9534253,1.0151579,1.2346514,0.980862,0.6036074,0.274367,0.07545093,0.01371835,0.8196714,1.2723769,0.8779744,0.66533995,1.2620882,2.8945718,1.6153357,1.6496316,2.1023371,3.018037,5.3878818,4.856296,8.134981,9.798331,8.069819,4.822,3.5873485,2.7573884,3.350707,5.051782,6.1972647,4.3452873,3.8205605,4.461893,6.6568294,11.317638,14.393978,18.12537,21.462358,24.250612,27.244642,28.667921,28.729654,27.618467,26.068295,25.368658,24.459818,22.662714,21.290878,20.773012,20.642687,18.440891,15.861842,13.834956,12.6757555,12.075578,12.878101,15.436573,15.748666,13.526293,12.202472,10.151579,7.7920227,6.228131,5.610805,5.1340923,5.295283,5.164959,5.0655007,4.8837323,4.0880685,5.1409516,6.2692857,9.661148,13.999576,14.476289,8.951223,8.443645,9.427936,9.674867,8.224151,8.042382,7.8023114,7.3084507,6.697984,6.4098988,5.895461,4.262977,2.8568463,2.2395205,2.1812177,2.510458,3.0454736,3.5530527,3.9440255,4.2835546,5.2472687,5.192395,4.5956473,3.9165888,3.625074,4.07435,3.426158,2.9734523,3.1723683,3.6456516,3.858286,3.5702004,3.5187566,3.9440255,4.602506,5.120374,6.543653,6.725421,5.638242,5.377593,5.7994323,5.8337283,5.5662203,5.504488,6.5882373,7.500508,7.2158523,6.8145905,6.7219915,6.6876955,6.495639,6.420188,6.3001523,6.262427,6.7048435,6.416758,5.411889,4.201245,3.1483612,2.452155,1.9754424,1.4507155,1.1043272,1.0528834,1.3169615,1.762808,1.611906,1.2620882,0.91569984,0.5796003,0.53158605,0.5693115,0.6379033,0.71678376,0.8265306,0.89512235,0.9294182,0.922559,0.8779744,0.78537554,0.78537554,0.8196714,0.8471081,0.8265306,0.6893471,0.490431,0.29837412,0.16119061,0.09259886,0.07545093,0.12346515,0.13375391,0.12689474,0.12346515,0.1371835,0.20234565,0.29151493,0.3566771,0.4081209,0.50757897,0.42183927,0.37382504,0.35324752,0.36696586,0.44584638,0.90541106,1.9857311,2.6647894,2.6922262,2.603057,2.369845,2.6922262,3.3609958,4.3041325,5.610805,5.8817425,5.3501563,4.880303,4.7808447,4.8082814,4.2081037,4.650521,6.1732574,8.354475,10.329918,10.978109,9.904649,8.416207,7.449064,7.5759587,8.529384,9.825768,9.911508,8.868914,8.405919,9.253027,8.7317295,8.632272,9.764035,11.962401,12.55229,12.679185,11.653738,9.709162,8.018375,7.922347,7.915488,7.7268605,7.2638664,6.608815,5.778855,4.2595477,3.1140654,2.5653315,2.0028791,1.3855534,1.7422304,2.0234566,1.8348293,1.4232788,2.0920484,2.301253,1.6770682,0.6344737,0.37039545,0.36353627,0.4698535,0.61046654,0.66191036,0.44584638,0.4424168,0.84024894,0.85396725,0.4081209,0.14061308,0.28122616,0.15090185,0.041155048,0.034295876,0.020577524,0.061732575,0.072021335,0.058302987,0.034295876,0.01371835,0.106317215,0.14061308,0.10288762,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.017147938,0.017147938,0.030866288,0.061732575,0.024007112,0.020577524,0.041155048,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.041155048,0.082310095,0.07545093,0.082310095,0.10288762,0.12346515,0.12689474,0.09945804,0.07545093,0.037725464,0.01371835,0.037725464,0.13375391,0.22292319,0.23664154,0.17833854,0.12003556,0.19548649,0.10288762,0.037725464,0.020577524,0.0548734,0.12346515,0.13032432,0.1371835,0.15090185,0.16119061,0.12346515,0.19548649,0.16804978,0.12003556,0.13032432,0.31895164,0.30523327,0.22292319,0.15433143,0.15776102,0.2503599,0.31209245,0.33266997,0.29837412,0.26750782,0.37382504,0.7407909,0.65848076,0.4664239,0.30866286,0.13032432,0.14747226,0.22978236,0.45956472,0.9259886,1.7250825,0.8471081,0.29494452,0.17833854,0.33266997,0.32924038,0.33609957,0.29837412,0.2503599,0.19548649,0.12689474,0.12689474,0.106317215,0.14747226,0.28122616,0.5178677,0.45956472,0.45956472,0.7099246,1.3478279,2.4487255,2.0028791,1.4027013,1.0254467,0.9431366,0.9294182,0.7133542,0.84367853,1.097468,1.3375391,1.5330256,2.170929,1.5776103,1.1934965,1.4335675,1.670209,1.8073926,1.7971039,1.8691251,1.9857311,1.8279701,1.5536032,1.7833855,1.6633499,1.0597426,0.5658819,0.6173257,0.5555932,0.48700142,0.47328308,0.5453044,0.90198153,1.4267083,1.5501735,1.1420527,0.5041494,0.72707254,0.70306545,0.6859175,0.72707254,0.67219913,0.5624523,0.39440256,0.29494452,0.30866286,0.36353627,0.28122616,0.20234565,0.13032432,0.07888051,0.061732575,0.12346515,0.2709374,0.29837412,0.20920484,0.20920484,0.082310095,0.3018037,1.5021594,4.705394,11.30735,15.100473,12.442543,8.759167,6.927767,7.2604365,8.477941,9.489669,11.105004,13.375391,15.570327,16.249386,15.54632,14.658057,14.1299,13.858963,14.30138,15.765814,17.62465,19.010202,18.79757,18.084215,18.396307,18.115082,16.911295,15.758954,15.923574,16.702091,18.073925,19.027351,17.573206,14.757515,10.569988,7.8331776,7.2707253,7.517656,4.0503426,4.170378,7.0889573,11.780633,16.969599,22.851341,25.005123,24.302057,22.508383,22.2786,19.253704,19.013634,21.565247,23.842491,19.716698,13.046151,14.472859,16.369421,15.3302555,12.178465,14.4317045,15.121051,15.748666,15.566897,11.592006,16.345413,15.484588,12.476839,10.113853,10.521975,9.880642,9.208443,8.375052,7.455923,6.7048435,7.3873315,6.910619,6.691125,7.0272245,7.1061053,5.147811,4.2115335,3.3781435,2.5241764,2.318401,2.7813954,3.0523329,3.2718265,3.5359046,3.9097297,4.9077396,4.8768735,4.057202,3.093488,3.0386145,4.033195,4.3590055,4.3109913,3.9097297,2.9185789,2.3424082,1.5981878,1.3546871,1.6530612,1.9239986,2.2978237,2.6716487,2.976882,3.1620796,3.2066643,2.1743584,1.6770682,1.3375391,1.0425946,0.94656616,0.9294182,1.0700313,1.1626302,1.097468,0.8676856,1.1214751,0.9774324,0.78537554,0.6824879,0.59674823,0.7510797,0.7956643,0.85396725,0.97400284,1.0940384,1.0117283,0.94656616,0.86082643,0.75450927,0.6756287,0.6859175,0.66191036,0.59674823,0.4938606,0.34981793,0.39097297,0.3806842,0.40126175,0.45613512,0.47671264,0.37382504,0.26064864,0.17833854,0.13032432,0.09259886,0.116605975,0.31552204,0.5693115,0.72021335,0.5796003,0.53844523,0.47671264,0.3806842,0.26064864,0.14061308,0.08916927,0.058302987,0.1097468,0.17490897,0.061732575,0.116605975,0.20920484,0.2194936,0.12689474,0.0,0.048014224,0.07545093,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.06516216,0.07888051,0.13032432,0.31552204,0.4664239,0.48700142,0.32924038,0.23321195,0.14747226,0.08573969,0.048014224,0.048014224,0.010288762,0.030866288,0.044584636,0.041155048,0.041155048,0.16804978,0.28808534,0.2777966,0.22635277,0.4424168,0.47328308,0.3806842,0.40126175,0.51100856,0.42869842,0.25721905,0.216064,0.4938606,1.0597426,1.6359133,0.7682276,0.53501564,0.548734,0.607037,0.6790583,1.0494537,1.3512574,1.4575747,1.4267083,1.4781522,2.1400626,4.383013,7.4113383,8.529384,3.1380725,3.6696587,7.3564653,10.882081,12.651748,12.809509,9.774324,7.7680154,7.5553813,8.899779,10.556271,13.893259,13.543441,13.437123,16.431154,24.343212,33.140102,30.324413,32.26213,45.918747,68.8764,70.86214,48.30917,25.286348,12.648318,8.056101,3.9337368,2.3424082,3.093488,4.945465,5.610805,4.972902,2.8568463,1.5776103,1.6873571,2.0063086,1.9651536,1.7971039,1.529596,1.0734608,0.22292319,0.29151493,1.0323058,0.53158605,0.09602845,0.3841138,1.4369972,1.3752645,1.4267083,1.3581166,1.5570327,3.0146074,3.2512488,11.06042,18.475187,18.61923,5.7308407,3.7485392,3.4021509,3.6079261,4.07435,5.2815647,5.627953,6.3721733,7.2295704,7.857185,7.8674736,8.213862,10.343636,13.906977,17.720678,19.78529,21.69214,22.36091,21.541239,20.231136,20.666695,21.064526,20.515793,20.53294,21.27716,21.53781,17.521763,14.579176,13.395968,13.193623,11.71547,15.254805,20.251715,20.676983,16.19794,12.175035,10.751757,8.573969,6.81802,6.0635104,6.3138704,5.5559316,5.435896,6.601956,7.1781263,2.784825,4.016047,5.9743414,8.076678,9.290752,8.134981,6.64997,7.3427467,7.864044,7.250148,5.919468,5.885172,5.3844523,4.695105,4.0537724,3.6593697,3.1552205,2.386993,1.9720128,2.0920484,2.4727325,2.7299516,3.1072063,3.3198407,3.391862,3.6593697,4.5682106,4.4996185,4.2389703,4.108646,3.9611735,3.8617156,3.3061223,3.1483612,3.4398763,3.4433057,2.9974594,2.486451,2.3629858,2.7093742,3.216953,4.1429415,5.518206,5.8234396,5.15467,5.212973,5.2164025,4.979761,4.664239,4.588788,5.2335505,7.0786686,7.747438,7.459353,6.807731,6.7528577,7.3084507,7.442205,7.3427467,7.291303,7.6616983,7.3050213,6.2075534,5.020916,4.033195,3.1723683,2.3664153,1.6393428,1.0666018,0.7339317,0.7407909,1.1660597,1.6359133,1.6359133,1.1900668,0.84024894,0.72364295,0.6344737,0.5041494,0.37039545,0.37382504,0.42526886,0.4698535,0.5007198,0.5178677,0.5144381,0.5521636,0.5796003,0.58988905,0.5693115,0.4938606,0.39783216,0.29151493,0.19548649,0.12003556,0.06859175,0.10288762,0.1097468,0.11317638,0.12003556,0.12003556,0.116605975,0.11317638,0.15090185,0.24350071,0.39097297,0.3841138,0.3841138,0.37039545,0.3566771,0.39783216,0.65162164,1.2963841,2.136633,2.719663,2.3046827,2.5790498,2.7230926,3.0043187,3.5633414,4.448175,4.866585,4.65395,4.0263357,3.4398763,3.5564823,3.4947495,4.091498,5.302142,6.999788,8.964942,9.547972,8.529384,7.2021337,6.3790326,6.3893213,7.051232,8.436785,8.940934,8.64599,9.342196,9.784613,10.196163,10.432805,10.63858,11.2593355,12.682614,13.858963,13.4474125,11.4376745,9.153569,8.985519,8.573969,7.764586,7.5588107,10.110424,8.31332,6.217842,4.7191124,3.7794054,2.4487255,1.371835,1.6427724,2.0268862,1.9102802,1.3032433,1.5604624,1.488441,1.1934965,0.90884066,0.9774324,0.91912943,0.64476246,0.5041494,0.50757897,0.31552204,0.32924038,0.50757897,0.4938606,0.2469303,0.041155048,0.12689474,0.07545093,0.034295876,0.037725464,0.017147938,0.1097468,0.17833854,0.20920484,0.17833854,0.05144381,0.07888051,0.13375391,0.13375391,0.072021335,0.0,0.0,0.020577524,0.020577524,0.0034295875,0.017147938,0.034295876,0.048014224,0.041155048,0.041155048,0.12346515,0.024007112,0.0034295875,0.020577524,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05144381,0.11317638,0.044584636,0.034295876,0.05144381,0.09945804,0.1371835,0.0548734,0.041155048,0.044584636,0.058302987,0.072021335,0.06516216,0.030866288,0.020577524,0.017147938,0.020577524,0.020577524,0.058302987,0.072021335,0.061732575,0.06859175,0.17147937,0.09259886,0.034295876,0.006859175,0.017147938,0.041155048,0.037725464,0.044584636,0.058302987,0.072021335,0.0548734,0.116605975,0.116605975,0.116605975,0.16804978,0.32924038,0.39440256,0.28465575,0.15433143,0.11317638,0.216064,0.39097297,0.44927597,0.3806842,0.29151493,0.4115505,0.6756287,0.45956472,0.2709374,0.35324752,0.6790583,1.4815818,1.728512,1.4850113,1.0906088,1.155771,0.5624523,0.18176813,0.07888051,0.15433143,0.13032432,0.19548649,0.24007112,0.24007112,0.22635277,0.2709374,0.34638834,0.34638834,0.4046913,0.6241849,1.08032,1.2072148,1.1763484,1.1489118,1.2929544,1.7593783,1.7113642,1.4061309,1.2517995,1.3032433,1.2586586,0.7956643,0.7922347,1.039165,1.3786942,1.7113642,2.3835633,2.085189,1.6393428,1.4472859,1.5090185,1.7559488,1.6564908,1.6667795,1.8313997,1.7902447,1.5604624,1.6770682,1.5330256,1.0734608,0.78537554,0.864256,0.8162418,0.61389613,0.40126175,0.51100856,0.86082643,1.1523414,1.3443983,1.3409687,1.0117283,0.96714365,0.9568549,1.0117283,1.0734608,0.9774324,0.65505123,0.40126175,0.26750782,0.24007112,0.23664154,0.37039545,0.33266997,0.24007112,0.17490897,0.18519773,0.20234565,0.25721905,0.4389872,0.6790583,0.7442205,0.5521636,0.432128,0.91912943,2.9391565,7.795452,14.29452,13.169616,9.619993,6.9380555,6.5230756,7.267296,9.5033865,12.240198,14.29452,14.30138,13.032433,13.118172,13.265644,12.88839,12.103014,12.212761,13.395968,15.035312,16.513464,17.178804,16.88386,16.37971,15.337115,14.006435,13.227919,13.7697935,15.083325,16.424294,17.086205,16.400288,13.958421,9.784613,6.7802944,5.844017,5.857735,4.6265135,4.8425775,7.2707253,10.933525,13.097594,14.575747,20.11453,22.882208,21.02337,17.658945,16.6335,17.319416,19.613811,21.472647,18.907316,16.582056,19.823015,23.022821,22.570116,16.842705,15.71094,14.445422,13.96185,14.071597,13.488567,17.772121,15.896138,12.950122,11.238758,10.288762,9.616563,8.440215,7.5039372,7.1781263,7.449064,8.748878,8.1487,7.3358874,6.9826403,6.7802944,5.6519604,4.602506,3.7005248,3.0489032,2.7882545,3.340418,3.4295874,3.223812,3.0626216,3.4535947,4.602506,4.7019644,4.232111,3.673088,3.5050385,3.6627994,3.4124396,3.2546785,3.3609958,3.5633414,3.0146074,1.9171394,1.6530612,2.1674993,1.9651536,2.4007113,2.9734523,3.3815732,3.415869,2.976882,2.534465,2.0165975,1.4232788,0.9328478,0.91569984,1.08032,1.2072148,1.1454822,0.99801,1.1283343,1.0597426,0.8162418,0.6207553,0.5555932,0.5727411,0.66533995,0.66876954,0.7305021,0.8676856,0.980862,0.8471081,0.77508676,0.78537554,0.8196714,0.7613684,0.64476246,0.5624523,0.51100856,0.4629943,0.37725464,0.38754338,0.3841138,0.4046913,0.45613512,0.53501564,0.41840968,0.31895164,0.24007112,0.17833854,0.13032432,0.22978236,0.5007198,0.6859175,0.6893471,0.58302987,0.65848076,0.7476501,0.66533995,0.4081209,0.16119061,0.072021335,0.048014224,0.07545093,0.1097468,0.082310095,0.29837412,0.66191036,0.7442205,0.44584638,0.0,0.024007112,0.07545093,0.06516216,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.037725464,0.06859175,0.061732575,0.14747226,0.26750782,0.37725464,0.4389872,0.4629943,0.35324752,0.20234565,0.082310095,0.024007112,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.13375391,0.22978236,0.18176813,0.07545093,0.17833854,0.33609957,0.28808534,0.2709374,0.37039545,0.53501564,0.6036074,0.3018037,0.28808534,0.70306545,1.1694894,0.6310441,0.29151493,0.19548649,0.26750782,0.29837412,0.48700142,0.65505123,0.823101,0.91912943,0.7888051,0.85739684,2.4452958,5.0757895,6.842027,4.40702,4.3281393,6.852316,9.208443,9.935514,8.886061,6.210983,6.3653145,7.4456344,8.275595,8.4093485,12.055,12.977559,12.394529,13.310229,20.52951,28.59247,26.610168,24.840502,31.908882,54.839104,73.86988,64.10585,39.06986,14.928994,10.501397,12.891819,14.092175,11.032983,5.809721,5.717122,5.442755,3.5804894,2.3252604,2.3424082,2.7642474,2.8054025,2.136633,2.4555845,2.9288676,0.20920484,0.0,0.5590228,0.34295875,0.082310095,0.06859175,0.16804978,0.6927767,1.3546871,1.1660597,0.4355576,0.7682276,1.6016173,9.283894,17.412016,18.61923,4.557922,3.1449318,3.2855449,3.3678548,3.1483612,3.7553983,4.866585,6.358455,7.5382333,8.008087,7.6651278,5.552502,6.0052075,9.3079,13.749216,15.621771,15.278812,16.616352,17.240536,17.137648,18.670673,21.328604,18.986197,18.392878,20.855322,22.227156,19.19197,18.173384,16.863281,14.483148,11.784062,15.13134,18.9519,18.71526,14.342535,10.192734,9.990388,8.591117,8.303031,9.5205345,10.72089,8.488229,6.7940125,7.0923867,7.8537555,4.5647807,6.077229,7.5416627,7.5416627,6.0532217,4.431027,5.8405876,6.636252,6.416758,5.4839106,4.822,4.5819287,3.765687,3.000889,2.4658735,1.8965619,1.2758065,1.0323058,1.1626302,1.5364552,1.8862731,1.9857311,2.3561265,2.5961976,2.5481834,2.287535,2.784825,2.9322972,3.2786856,3.8891523,4.314421,3.9063,3.4913201,3.3952916,3.3815732,2.6545007,2.177788,1.7490896,1.6667795,1.9308578,2.2292318,3.0969174,4.029765,4.314421,4.040054,4.0880685,3.6216443,3.316411,3.2203827,3.2958336,3.4021509,5.113515,6.475061,6.883182,6.543653,6.468202,7.2467184,7.5210853,7.534804,7.5931067,8.042382,7.9257765,7.0203657,5.919468,4.9008803,3.9165888,2.9082901,2.0508933,1.3615463,0.84024894,0.4664239,0.5693115,1.0837497,1.2346514,0.91912943,0.6790583,0.58988905,0.48700142,0.3566771,0.24007112,0.23664154,0.2194936,0.23321195,0.2777966,0.33266997,0.36353627,0.4046913,0.4355576,0.4355576,0.40126175,0.34295875,0.3018037,0.26407823,0.216064,0.15433143,0.07545093,0.06859175,0.072021335,0.07888051,0.08916927,0.07545093,0.0548734,0.044584636,0.061732575,0.12689474,0.24350071,0.30523327,0.35324752,0.36696586,0.36010668,0.3841138,0.4938606,0.71678376,1.3752645,2.1194851,1.9239986,2.3321195,2.3767042,2.3561265,2.4795918,2.867135,3.4467354,3.9508848,3.9474552,3.5942078,3.6525106,4.081209,4.8117113,5.6210938,6.5367937,7.8606143,7.953213,7.140401,6.258997,5.7925735,5.8645945,6.183546,7.222711,8.217292,9.105555,10.511685,10.878652,12.092726,13.001566,12.9981365,12.044711,13.090735,14.589465,14.788382,13.162757,10.405369,10.360784,9.012956,7.6205435,7.73029,11.180455,9.469091,8.001227,6.1904054,4.184097,2.8568463,2.3218307,2.5721905,2.8019729,2.5653315,1.7593783,1.7525192,1.2723769,0.9877212,1.0940384,1.3238207,1.0425946,0.70649505,0.52472687,0.4972902,0.4355576,0.4424168,0.34638834,0.2194936,0.106317215,0.024007112,0.044584636,0.07545093,0.08916927,0.082310095,0.09602845,0.17147937,0.21263443,0.21263443,0.16462019,0.044584636,0.037725464,0.09602845,0.1371835,0.116605975,0.030866288,0.010288762,0.0274367,0.024007112,0.0034295875,0.017147938,0.08573969,0.08573969,0.0548734,0.041155048,0.12003556,0.058302987,0.037725464,0.041155048,0.05144381,0.041155048,0.072021335,0.037725464,0.01371835,0.01371835,0.0,0.0,0.037725464,0.12689474,0.20577525,0.12003556,0.09602845,0.07888051,0.09259886,0.10288762,0.017147938,0.0034295875,0.0,0.006859175,0.020577524,0.0274367,0.010288762,0.020577524,0.034295876,0.05144381,0.058302987,0.07888051,0.12003556,0.116605975,0.07545093,0.09259886,0.048014224,0.01371835,0.017147938,0.048014224,0.06859175,0.05144381,0.05144381,0.048014224,0.041155048,0.048014224,0.072021335,0.07545093,0.11317638,0.1920569,0.29837412,0.42526886,0.25721905,0.1097468,0.1371835,0.33952916,0.6001778,0.6276145,0.47671264,0.29494452,0.29494452,0.3841138,0.18862732,0.07888051,0.26407823,0.7922347,1.5433143,1.6839274,1.3032433,0.7133542,0.44927597,0.1920569,0.061732575,0.048014224,0.08916927,0.07545093,0.13375391,0.20577525,0.2469303,0.2777966,0.4115505,0.45270553,0.432128,0.47328308,0.6859175,1.1660597,1.4198492,1.4198492,1.3272504,1.2620882,1.2758065,1.3306799,1.2380811,1.2483698,1.3512574,1.2860953,0.91227025,0.84024894,0.9568549,1.2517995,1.8348293,2.5756202,2.3972816,1.8348293,1.3786942,1.4918705,1.786815,1.6221949,1.5124481,1.6016173,1.6633499,1.3752645,1.4953002,1.3821237,0.99801,0.89512235,1.0837497,1.039165,0.7476501,0.41840968,0.48700142,0.7990939,0.9431366,1.1077567,1.2620882,1.1351935,0.89855194,0.90884066,1.0014396,1.0288762,0.8676856,0.53844523,0.32924038,0.2709374,0.39097297,0.72364295,1.471293,1.5913286,1.2689474,0.7510797,0.34981793,0.2503599,0.24350071,0.48357183,0.89855194,1.1900668,0.99801,0.7613684,0.8196714,1.6907866,4.064061,8.913498,9.043822,7.599966,6.5950966,6.9071894,7.040943,8.834618,11.135871,12.651748,11.945253,9.914937,10.1481495,10.741467,10.64201,9.644,10.100135,11.406808,12.915827,14.345964,15.80011,16.221949,15.536031,14.328816,13.049581,12.0309925,12.020704,13.4645605,14.908417,15.577187,15.374841,14.421415,12.0138445,9.030104,6.9071894,7.654839,9.445084,8.64942,8.549961,10.189304,12.360233,11.495977,16.6335,19.771572,18.355152,15.289101,14.5243025,15.422854,17.065628,18.482046,18.62266,18.506054,23.249174,28.023159,28.93886,23.057117,17.346853,13.745787,11.900668,12.178465,15.656067,18.44775,15.937293,13.227919,11.818358,9.609704,8.889491,7.9189177,7.0718093,6.708273,7.181556,8.268735,7.7028537,6.756287,6.138962,5.9983487,4.99005,3.841138,3.0866287,2.8637056,2.8980014,3.1037767,3.4398763,3.415869,3.1895163,3.5530527,4.3521466,4.32471,4.1292233,4.0503426,4.0091877,3.5530527,2.9117198,2.5619018,2.6956558,3.2409601,3.1449318,2.3149714,2.1229146,2.5447538,2.1469216,2.3767042,2.819121,3.2203827,3.2581081,2.5550427,2.719663,2.3081124,1.611906,1.0563129,1.214074,1.4164196,1.3752645,1.1694894,1.0117283,1.2517995,0.9842916,0.7510797,0.5624523,0.47328308,0.5727411,0.5453044,0.52815646,0.6036074,0.7613684,0.88826317,0.71678376,0.6756287,0.7373613,0.8196714,0.78537554,0.61046654,0.490431,0.44584638,0.45270553,0.4389872,0.41498008,0.37382504,0.37039545,0.42183927,0.51100856,0.51100856,0.4698535,0.38754338,0.28465575,0.18519773,0.25721905,0.5007198,0.61389613,0.5590228,0.5590228,0.85396725,0.9774324,0.84367853,0.5144381,0.20920484,0.116605975,0.106317215,0.15433143,0.20577525,0.19891608,0.52472687,0.84024894,0.82996017,0.4629943,0.0,0.020577524,0.0548734,0.044584636,0.0,0.0,0.037725464,0.020577524,0.0,0.010288762,0.05144381,0.041155048,0.07545093,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.020577524,0.030866288,0.072021335,0.16462019,0.30523327,0.4115505,0.34638834,0.22978236,0.12346515,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.23321195,0.24007112,0.12346515,0.0,0.0,0.23664154,0.19548649,0.12003556,0.17490897,0.4355576,0.5041494,0.20920484,0.06516216,0.22978236,0.48357183,0.4081209,0.1920569,0.07545093,0.09602845,0.072021335,0.08916927,0.12346515,0.2503599,0.40126175,0.37382504,0.37382504,1.1043272,2.6545007,4.5956473,5.994919,5.096367,5.7719955,7.675417,9.403929,8.508806,5.6656785,7.010077,9.283894,10.666017,10.779194,16.45859,17.130789,15.892709,16.21509,21.976797,30.331272,27.618467,21.644127,22.223726,41.182487,59.222115,57.10263,38.401093,16.496315,14.579176,25.93111,24.86451,17.079346,8.683716,6.210983,5.6210938,3.9543142,2.8225505,2.750529,3.1689389,2.9803114,1.9514352,2.0886188,2.644212,0.15090185,0.0,0.07888051,0.15776102,0.1371835,0.044584636,0.024007112,0.0034295875,0.9431366,1.0528834,0.25721905,0.17833854,0.5418748,3.5118976,7.191845,8.443645,2.8739944,2.74367,2.3424082,2.2120838,2.4761622,2.8294096,2.1126258,2.8294096,3.8274195,4.962613,7.0958166,5.0483527,4.664239,6.835168,10.703742,13.677195,11.7086115,13.430264,15.172495,16.077906,18.1288,22.477516,17.014183,14.373401,17.597214,20.152256,20.519222,22.470657,20.721567,15.409137,12.085866,12.298501,12.332796,11.640019,10.175586,8.381912,9.023245,8.906639,10.717461,13.910407,14.71636,12.127021,8.875772,6.756287,6.3961806,7.2467184,8.467651,8.601405,7.3050213,5.3330083,4.537344,6.1801167,6.279575,5.703404,5.1238036,4.979761,4.461893,3.542764,2.6990852,2.0303159,1.2586586,0.7442205,0.6207553,0.6962063,0.8025235,0.7888051,0.85739684,1.4267083,2.085189,2.335549,1.5707511,1.5844694,1.8691251,2.4898806,3.3541365,4.2526884,4.016047,3.7382503,3.5359046,3.1346428,1.8759843,1.8279701,1.8588364,1.9445761,2.0440342,2.1057668,2.633923,3.2683969,3.4295874,3.0866287,2.7539587,2.369845,2.2566686,2.4041407,2.6064866,2.4624438,3.1106358,4.314421,5.504488,6.2830043,6.4064693,6.9346256,7.143831,7.082098,7.034084,7.5279446,7.7440085,7.366754,6.6122446,5.6828265,4.787704,3.7862647,2.8328393,2.0577524,1.4335675,0.77508676,0.4664239,0.33609957,0.28122616,0.22978236,0.12346515,0.09602845,0.07888051,0.12346515,0.22978236,0.34981793,0.22292319,0.15433143,0.15433143,0.1920569,0.2194936,0.2469303,0.29837412,0.31552204,0.28465575,0.23321195,0.22292319,0.20577525,0.1920569,0.16804978,0.08916927,0.05144381,0.048014224,0.048014224,0.041155048,0.030866288,0.030866288,0.030866288,0.037725464,0.06859175,0.1371835,0.22292319,0.30866286,0.37039545,0.4081209,0.44584638,0.5590228,0.5727411,0.7476501,1.1626302,1.7182233,1.6907866,1.7250825,1.728512,1.762808,2.020027,2.5996273,3.6147852,4.6127954,5.2644167,5.329579,5.7651367,6.193835,6.5333643,6.8214493,7.208993,6.7494283,6.2144127,5.7719955,5.5147767,5.4633327,5.9743414,6.8454566,8.032094,9.373062,10.590566,11.211322,12.737488,14.359683,15.059319,13.605173,13.317088,14.490007,15.254805,14.407697,11.38966,10.868362,8.711152,7.3255987,7.706283,9.431366,9.3079,8.549961,6.252138,3.4398763,3.069481,3.6696587,3.940596,3.923448,3.5633414,2.7059445,2.7128036,2.0474637,1.4472859,1.1934965,1.0940384,0.7133542,0.6859175,0.6962063,0.65505123,0.6859175,0.65848076,0.4629943,0.24007112,0.08573969,0.06859175,0.12003556,0.17833854,0.17833854,0.14747226,0.2194936,0.18176813,0.15090185,0.106317215,0.058302987,0.041155048,0.0274367,0.058302987,0.10288762,0.12689474,0.08573969,0.037725464,0.020577524,0.017147938,0.01371835,0.010288762,0.1371835,0.106317215,0.048014224,0.0274367,0.041155048,0.07545093,0.106317215,0.13375391,0.14747226,0.12003556,0.15090185,0.07888051,0.034295876,0.034295876,0.0,0.0548734,0.12003556,0.17147937,0.1920569,0.15433143,0.16462019,0.13032432,0.09259886,0.061732575,0.024007112,0.0274367,0.024007112,0.017147938,0.010288762,0.006859175,0.0274367,0.082310095,0.09945804,0.09259886,0.16462019,0.33952916,0.4389872,0.33952916,0.106317215,0.0,0.0,0.01371835,0.10288762,0.2194936,0.22292319,0.15776102,0.1371835,0.11317638,0.072021335,0.072021335,0.07888051,0.07888051,0.12689474,0.216064,0.30523327,0.4389872,0.2503599,0.106317215,0.17490897,0.4424168,0.7133542,0.67219913,0.4698535,0.22635277,0.044584636,0.13032432,0.13375391,0.08573969,0.09259886,0.34638834,0.24350071,0.106317215,0.034295876,0.041155048,0.041155048,0.041155048,0.041155048,0.0548734,0.072021335,0.061732575,0.07545093,0.13032432,0.19891608,0.29151493,0.44584638,0.39097297,0.31209245,0.28808534,0.3841138,0.6344737,0.86082643,0.980862,1.1180456,1.2826657,1.371835,1.214074,1.1043272,1.0700313,1.0563129,0.91912943,0.8711152,0.83681935,0.8162418,0.9294182,1.4129901,1.903421,1.8245405,1.5090185,1.3101025,1.5810398,1.7902447,1.6736387,1.5055889,1.4541451,1.5913286,1.2037852,1.3855534,1.3101025,0.881404,0.7133542,1.1180456,1.097468,0.83338976,0.5658819,0.59674823,0.9774324,1.2003556,1.2483698,1.1249046,0.83338976,0.6001778,0.5693115,0.607037,0.5727411,0.32924038,0.23664154,0.21263443,0.37382504,0.9294182,2.153781,3.8034124,4.1292233,3.4295874,2.1743584,1.0082988,0.5041494,0.36353627,0.4424168,0.69963586,1.1660597,1.0254467,0.94999576,1.0014396,1.1763484,1.4198492,2.0886188,2.7333813,3.5942078,4.8014226,6.4064693,6.90033,7.332458,8.114404,8.97866,8.968371,7.8983397,7.473071,7.438775,7.3873315,6.7528577,8.014946,9.774324,11.197603,12.277924,13.824667,14.774663,14.606613,13.958421,13.13189,12.068718,11.63659,13.416546,15.700651,17.04162,16.245956,16.818697,16.492886,13.612033,10.302481,12.459691,15.738377,13.649758,11.06042,11.207891,15.704081,15.309678,16.935303,17.45317,16.510035,16.523752,15.309678,15.107333,15.436573,16.492886,19.133669,17.902447,22.919933,28.630196,30.880005,26.93941,18.427174,14.243076,12.744347,13.601744,17.78927,18.053349,15.289101,12.9707,11.818358,9.788043,8.793462,8.165848,7.3255987,6.355026,6.0086374,6.427047,5.658819,5.0106273,4.955754,5.144381,3.40901,2.651071,2.4418662,2.5447538,2.8945718,2.3424082,2.9151495,3.4124396,3.5118976,3.7725463,3.9303071,3.799983,3.8617156,4.15323,4.245829,3.6010668,2.9665933,2.5756202,2.469303,2.486451,2.7539587,2.5447538,2.4315774,2.49331,2.2978237,2.2669573,2.4007113,2.7128036,2.8808534,2.2463799,2.5001693,2.253239,1.7833855,1.4541451,1.7216529,1.8313997,1.5844694,1.3375391,1.2312219,1.1832076,0.9911508,0.7990939,0.6036074,0.4698535,0.5555932,0.4424168,0.45956472,0.548734,0.67219913,0.8025235,0.67219913,0.66533995,0.70306545,0.72707254,0.7099246,0.58645946,0.4698535,0.42869842,0.44584638,0.4355576,0.41498008,0.34981793,0.31552204,0.32924038,0.36010668,0.53844523,0.58302987,0.5144381,0.37039545,0.19891608,0.16462019,0.28465575,0.36696586,0.39097297,0.50757897,0.939707,1.0460242,0.94999576,0.72707254,0.41840968,0.26407823,0.20920484,0.28122616,0.3841138,0.28465575,0.5624523,0.5796003,0.42183927,0.1920569,0.0274367,0.082310095,0.09259886,0.06859175,0.030866288,0.0,0.08916927,0.0548734,0.017147938,0.030866288,0.08573969,0.11317638,0.18862732,0.15090185,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.07888051,0.15090185,0.15433143,0.15433143,0.15090185,0.09259886,0.024007112,0.0034295875,0.0,0.0,0.0,0.274367,0.216064,0.07888051,0.0,0.0,0.16462019,0.082310095,0.0,0.030866288,0.15776102,0.044584636,0.006859175,0.0,0.037725464,0.18176813,0.13032432,0.07545093,0.030866288,0.010288762,0.05144381,0.07545093,0.07545093,0.07888051,0.12003556,0.23321195,0.20920484,0.24350071,0.8471081,2.7299516,6.783724,5.178677,4.7774153,7.3701835,11.351934,11.746337,8.615124,10.2236,12.782072,14.661487,16.383139,24.27805,25.20061,24.706749,24.919382,24.504402,32.58451,29.467016,21.181131,16.667795,27.807095,31.363577,30.530188,24.284908,16.973028,18.331144,32.17982,25.114868,15.7966795,11.427385,7.7748747,6.2384195,4.1943855,2.9254382,2.7573884,3.0626216,2.5173173,1.5364552,0.83338976,0.5212973,0.106317215,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.12003556,0.21263443,0.15090185,0.7613684,2.8122618,4.417309,5.0586414,5.5833683,5.1821065,2.4898806,1.4541451,3.292404,6.5162163,3.3301294,1.9548649,1.8142518,2.1503513,2.0303159,3.8479972,5.4667625,5.8371577,6.0497923,9.3079,12.932974,13.821238,12.686044,11.122152,11.598865,13.564018,10.8958,9.112414,10.203023,12.620882,12.9981365,13.999576,14.627191,14.003006,11.351934,9.839486,9.424506,10.600855,11.619442,8.467651,9.225591,11.694893,12.860953,11.46854,8.025234,9.770895,10.161868,9.630281,8.738589,8.162418,7.1369715,6.7528577,6.101236,5.1855364,4.928317,5.8680243,5.9297566,5.453044,4.7602673,4.149801,3.5050385,2.8019729,2.0989075,1.4267083,0.7922347,0.47671264,0.41498008,0.5007198,0.6927767,1.0220171,1.3169615,2.0097382,2.6750782,2.976882,2.6716487,2.633923,2.469303,2.2600982,2.0646117,1.9068506,2.3835633,2.8499873,3.0351849,2.74367,1.8759843,2.3149714,2.4898806,2.4795918,2.311542,1.9823016,2.2292318,2.976882,3.275256,2.8259802,1.9823016,2.1194851,2.352697,2.6750782,2.877424,2.5481834,2.8156912,3.4604537,4.266407,5.0277753,5.5387836,6.526505,6.931196,6.910619,6.8454566,7.3084507,7.1129646,6.927767,6.615674,6.1801167,5.751418,4.8014226,3.8308492,2.9322972,2.1194851,1.313532,0.7990939,0.4698535,0.274367,0.17147937,0.12346515,0.08573969,0.058302987,0.08916927,0.216064,0.47328308,0.32581082,0.18176813,0.09602845,0.08573969,0.12346515,0.061732575,0.0548734,0.06859175,0.08573969,0.12346515,0.17147937,0.18176813,0.18862732,0.18519773,0.1371835,0.09945804,0.072021335,0.0548734,0.041155048,0.030866288,0.030866288,0.030866288,0.024007112,0.0274367,0.07545093,0.11317638,0.23321195,0.36696586,0.48357183,0.5796003,0.5555932,0.5212973,0.58988905,0.8025235,1.1454822,1.4987297,1.862266,2.0817597,2.1674993,2.287535,2.8396983,4.2835546,5.895461,7.1266828,7.613684,7.4936485,7.3701835,7.5759587,7.9772205,7.963502,6.6465406,6.0154963,5.3673043,4.4859004,3.6319332,4.914599,6.9380555,8.261876,8.464222,8.1487,9.3079,11.063849,12.730629,13.615462,13.032433,12.274493,13.183334,14.723219,15.22051,12.3911,9.582268,7.507367,7.1541195,8.354475,9.794902,10.30934,7.160979,3.998899,2.6064866,2.8980014,3.5461934,2.8568463,2.411,2.486451,2.061182,1.5947582,1.4438564,1.4061309,1.2037852,0.47328308,0.65505123,0.490431,0.26064864,0.11317638,0.07545093,0.041155048,0.041155048,0.041155048,0.041155048,0.09259886,0.31209245,0.36696586,0.31209245,0.24350071,0.30523327,0.25721905,0.25378948,0.28465575,0.29837412,0.21263443,0.14061308,0.14061308,0.14747226,0.13375391,0.12346515,0.072021335,0.041155048,0.048014224,0.06859175,0.044584636,0.106317215,0.058302987,0.010288762,0.006859175,0.030866288,0.006859175,0.1371835,0.2709374,0.3018037,0.16804978,0.034295876,0.010288762,0.020577524,0.024007112,0.0,0.26750782,0.22635277,0.10288762,0.034295876,0.044584636,0.17833854,0.29494452,0.32581082,0.25721905,0.12346515,0.13375391,0.12003556,0.08916927,0.0548734,0.030866288,0.09259886,0.28122616,0.26750782,0.12689474,0.33609957,0.90884066,1.0425946,0.66533995,0.08573969,0.0,0.0,0.072021335,0.34295875,0.6241849,0.4424168,0.26064864,0.16804978,0.106317215,0.061732575,0.061732575,0.09602845,0.09602845,0.15090185,0.26750782,0.36696586,0.45270553,0.4629943,0.31895164,0.08916927,0.01371835,0.29494452,0.37382504,0.33266997,0.22978236,0.106317215,0.5212973,0.6173257,0.37382504,0.01371835,0.01371835,0.0034295875,0.017147938,0.0548734,0.07888051,0.030866288,0.030866288,0.020577524,0.01371835,0.01371835,0.0,0.024007112,0.06859175,0.09602845,0.12689474,0.21263443,0.274367,0.18862732,0.10288762,0.08573969,0.12346515,0.18176813,0.4355576,0.8505377,1.2723769,1.4198492,1.1763484,0.94999576,0.8025235,0.6859175,0.4424168,0.5041494,0.5453044,0.6859175,0.84024894,0.71678376,0.97400284,0.7888051,0.9294182,1.4472859,1.6770682,1.99602,2.1023371,2.0165975,1.821111,1.6633499,1.4438564,1.2415106,1.1146159,1.0082988,0.7613684,1.1283343,1.1214751,0.9911508,0.9294182,1.039165,1.8691251,2.0028791,1.6839274,1.1626302,0.6859175,0.490431,0.32238123,0.2194936,0.17147937,0.12346515,0.14747226,0.216064,0.64476246,1.8862731,4.547633,6.975781,7.346176,6.385892,4.7671266,3.083199,1.4953002,0.72364295,0.44927597,0.432128,0.5178677,0.50757897,0.58645946,0.83681935,1.0048691,0.5041494,0.48014224,0.78537554,1.2655178,2.085189,3.707384,6.2212715,7.6651278,8.093826,7.6033955,6.3310184,7.0889573,6.9209075,5.597087,3.9337368,3.799983,4.5819287,5.5559316,6.7219915,7.8434668,8.453933,9.493098,9.73317,10.31277,11.399949,12.1921835,12.47341,14.867262,18.849012,22.021381,20.141968,19.483486,19.171394,16.832415,13.437123,13.289652,15.817257,15.340545,15.066177,16.777542,20.841602,18.183672,19.147387,19.569225,18.344864,17.439453,19.661825,18.852442,17.79613,18.766703,23.5304,21.966507,20.258574,21.211998,24.000254,24.171732,18.176813,17.38115,18.78042,20.560377,22.11055,15.71437,12.593445,12.288212,13.38911,13.533153,11.739478,9.764035,7.949784,6.776865,6.852316,6.9860697,5.874883,5.223262,5.219832,4.547633,2.4590142,2.5070283,3.1826572,3.5873485,3.4192986,2.270387,1.8828435,1.9994495,2.369845,2.7470996,2.7093742,2.6819375,3.175798,3.9886103,4.197815,3.415869,3.0557625,2.9322972,2.8054025,2.3664153,2.5241764,2.719663,2.8225505,2.750529,2.4555845,2.4555845,2.5378947,2.7299516,2.7230926,1.8931323,1.5021594,1.5673214,1.8073926,2.0646117,2.318401,2.3801336,2.2292318,1.9994495,1.7456601,1.4644338,1.1351935,0.88826317,0.70649505,0.5796003,0.5178677,0.44584638,0.5007198,0.5555932,0.5590228,0.53501564,0.5693115,0.6344737,0.64819205,0.6001778,0.5658819,0.42869842,0.37725464,0.3841138,0.40126175,0.34981793,0.33952916,0.33609957,0.31209245,0.274367,0.274367,0.33609957,0.38754338,0.38754338,0.30866286,0.1371835,0.06516216,0.06516216,0.11317638,0.20234565,0.33609957,0.64133286,0.97400284,1.3203912,1.4678634,0.9911508,0.5144381,0.20577525,0.106317215,0.1371835,0.07545093,0.05144381,0.12003556,0.15090185,0.12346515,0.1371835,0.22292319,0.29837412,0.274367,0.14747226,0.0,0.061732575,0.07545093,0.082310095,0.1097468,0.18176813,0.23321195,0.18176813,0.13032432,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.0548734,0.09259886,0.10288762,0.07888051,0.072021335,0.09259886,0.09259886,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.030866288,0.0,0.0,0.0,0.072021335,0.037725464,0.0,0.01371835,0.07545093,0.08916927,0.1097468,0.08573969,0.037725464,0.061732575,0.048014224,0.0548734,0.17833854,1.4850113,6.025785,4.0503426,5.0312047,9.174147,14.980438,19.239986,12.367092,13.708061,16.081335,17.470318,21.009653,25.859089,34.99894,41.552883,39.361374,22.978235,22.796469,25.817934,23.249174,17.981327,24.597002,29.43272,27.42641,23.393215,20.176264,18.660385,16.894148,11.074138,8.224151,9.97324,12.572867,9.033533,5.0895076,2.7230926,2.2806756,2.486451,2.0234566,1.1489118,0.4629943,0.16804978,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.041155048,0.030866288,1.5981878,1.5330256,1.255229,1.4953002,2.3149714,3.6696587,2.9322972,1.6324836,1.0528834,2.2429502,2.1915064,2.510458,2.627064,2.5653315,2.9220085,3.5770597,4.931747,4.650521,3.07634,3.2306714,5.3913116,7.3187394,7.085528,5.3673043,5.446185,6.8728933,6.708273,7.2192817,8.745448,9.688584,10.302481,12.833516,15.175924,16.822126,18.87302,13.1593275,12.0309925,15.107333,18.293419,13.766364,9.757176,9.952662,10.220171,9.050681,7.56224,8.683716,9.942374,9.6988735,8.097256,7.06495,5.9126086,5.744559,5.6793966,5.363875,4.99005,5.518206,5.669108,5.206114,4.3178506,3.6010668,3.0111778,2.318401,1.6324836,1.0323058,0.5727411,0.35324752,0.39097297,0.7339317,1.2758065,1.7422304,1.7730967,2.2463799,3.6216443,5.171818,5.0003386,3.5290456,3.4227283,3.4810312,3.2889743,3.2375305,3.3129816,2.7299516,2.369845,2.3424082,1.9754424,2.5207467,3.1620796,3.391862,3.1346428,2.726522,3.0797696,3.6216443,4.2081037,4.523626,4.0846386,3.4947495,4.479041,5.0895076,4.914599,5.0620713,5.9743414,6.759717,6.852316,6.509357,6.7974424,7.874333,8.1212635,7.517656,6.543653,6.1972647,6.5024977,6.4544835,6.3481665,6.2727156,6.118384,5.5559316,4.773986,3.8514268,2.8739944,1.9239986,1.1934965,0.70306545,0.39440256,0.22292319,0.13375391,0.106317215,0.09602845,0.16804978,0.34981793,0.64476246,0.53501564,0.40126175,0.29151493,0.2503599,0.31895164,0.22635277,0.12689474,0.0548734,0.030866288,0.037725464,0.048014224,0.072021335,0.1097468,0.15776102,0.19891608,0.16119061,0.12003556,0.07545093,0.041155048,0.030866288,0.020577524,0.017147938,0.017147938,0.020577524,0.041155048,0.048014224,0.08573969,0.19891608,0.34638834,0.3841138,0.48700142,0.47671264,0.5453044,0.71678376,0.864256,1.0220171,1.3306799,1.5433143,1.546744,1.3375391,1.9925903,3.3781435,5.1992545,6.9963584,8.1384115,8.759167,9.355915,9.589127,9.355915,8.80718,7.380472,6.3207297,5.7651367,5.4324665,4.5956473,5.1855364,6.2727156,6.975781,7.143831,7.3427467,8.237869,9.266746,10.840926,12.3533745,12.175035,10.796341,10.398509,11.375941,12.607163,11.4754,10.172156,10.096705,10.744898,11.269625,10.504827,8.889491,6.5162163,4.835718,4.280125,4.290414,2.7711067,1.8245405,1.3786942,1.2963841,1.3752645,1.762808,1.3238207,0.78537554,0.45613512,0.24007112,0.41498008,0.24007112,0.082310095,0.07545093,0.1371835,0.13032432,0.09259886,0.07888051,0.14404267,0.34638834,0.26407823,0.28122616,0.31895164,0.31552204,0.2194936,0.26750782,0.22292319,0.1371835,0.1097468,0.29837412,0.25378948,0.28465575,0.32924038,0.31209245,0.13375391,0.15433143,0.09602845,0.037725464,0.01371835,0.010288762,0.14747226,0.14061308,0.06859175,0.020577524,0.10288762,0.07888051,0.16804978,0.21263443,0.15776102,0.034295876,0.017147938,0.020577524,0.0274367,0.034295876,0.048014224,0.12346515,0.082310095,0.041155048,0.034295876,0.010288762,0.06516216,0.16804978,0.20920484,0.15776102,0.072021335,0.16462019,0.14747226,0.07545093,0.01371835,0.017147938,0.030866288,0.16462019,0.216064,0.23321195,0.5178677,0.7133542,0.50757897,0.2194936,0.030866288,0.01371835,0.01371835,0.13032432,0.26064864,0.29837412,0.12346515,0.058302987,0.048014224,0.041155048,0.030866288,0.061732575,0.16462019,0.15433143,0.23321195,0.4424168,0.64819205,0.5761707,0.41840968,0.21263443,0.037725464,0.0034295875,0.40126175,0.6276145,0.61389613,0.45956472,0.42526886,0.9774324,0.9568549,0.5178677,0.01371835,0.01371835,0.01371835,0.024007112,0.034295876,0.041155048,0.030866288,0.030866288,0.0274367,0.0274367,0.034295876,0.061732575,0.14404267,0.12003556,0.09259886,0.12003556,0.22635277,0.26750782,0.16119061,0.06859175,0.041155048,0.048014224,0.07888051,0.22978236,0.5007198,0.8093826,1.0048691,1.1008976,0.85739684,0.5521636,0.32238123,0.18519773,0.26750782,0.4389872,0.65162164,0.805953,0.75450927,0.9431366,0.90198153,1.0048691,1.2723769,1.3992717,1.4815818,1.5227368,1.488441,1.4335675,1.4815818,1.2792361,1.155771,1.0631721,0.9877212,0.9568549,1.6359133,1.704505,1.4953002,1.2758065,1.2586586,1.1111864,1.097468,1.1934965,1.2346514,0.89512235,0.48357183,0.2777966,0.16804978,0.1097468,0.1097468,0.11317638,0.17833854,0.5727411,1.762808,4.4241676,7.459353,8.2310095,7.8091707,6.924337,5.9640527,2.5207467,1.0734608,0.72364295,0.8093826,0.8848336,0.7373613,0.5453044,0.5693115,0.6756287,0.37039545,0.33609957,0.50757897,0.8471081,1.5810398,3.1963756,5.672538,7.706283,8.292743,7.373613,5.8200097,7.2707253,6.8866115,5.5319247,4.1120753,3.566771,3.234101,3.7108135,4.139512,4.6093655,6.159539,6.6705475,7.421627,8.676856,10.134431,10.947243,10.943813,12.435684,16.101913,20.409475,21.606401,17.401728,15.649208,14.706071,13.759505,12.80265,12.908967,12.30193,12.857523,15.031882,17.864721,19.023922,19.03078,18.097933,17.182234,17.977898,22.04539,23.808197,20.567236,15.429714,17.29198,18.101362,18.135658,19.11652,20.361462,18.773561,17.027903,16.79126,16.890718,16.53747,15.337115,12.308789,13.920695,16.94902,18.482046,15.913286,11.962401,9.510246,8.81747,9.3936405,10.010965,8.182996,6.4579134,5.6210938,5.5387836,5.1683884,3.5804894,3.450165,3.7794054,3.782835,2.867135,2.3664153,2.0886188,2.0028791,2.0886188,2.318401,2.486451,2.4590142,2.5447538,2.7813954,2.9391565,2.568761,2.4041407,2.6167753,2.9048605,2.5241764,2.5550427,2.7128036,2.5893385,2.301253,2.4555845,3.3438478,3.3061223,2.7333813,1.9925903,1.4164196,1.5124481,1.5330256,1.728512,2.0920484,2.369845,2.0680413,2.061182,1.937717,1.587899,1.2209331,1.0768905,0.90541106,0.66876954,0.42526886,0.32238123,0.31895164,0.3841138,0.44927597,0.47328308,0.44927597,0.52472687,0.53844523,0.5796003,0.6036074,0.42869842,0.37382504,0.37039545,0.37382504,0.33266997,0.216064,0.19548649,0.18176813,0.16804978,0.17147937,0.2503599,0.34981793,0.4115505,0.3566771,0.216064,0.11317638,0.058302987,0.06516216,0.1097468,0.216064,0.45613512,0.7339317,0.8676856,0.96714365,1.0837497,1.2106444,0.91227025,0.47671264,0.17147937,0.072021335,0.041155048,0.044584636,0.06859175,0.058302987,0.024007112,0.0274367,0.17147937,0.2194936,0.17490897,0.10288762,0.12346515,0.11317638,0.09259886,0.106317215,0.14061308,0.08573969,0.14404267,0.10288762,0.072021335,0.06859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.030866288,0.116605975,0.12003556,0.09259886,0.072021335,0.06859175,0.07888051,0.058302987,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.0274367,0.034295876,0.024007112,0.006859175,0.01371835,0.020577524,0.024007112,0.09259886,0.490431,1.6804979,1.8039631,4.664239,8.64256,12.411677,14.932424,13.978998,14.671775,17.466888,22.669573,30.458166,34.75887,42.773815,45.23969,38.33936,23.674442,16.081335,20.385468,20.073376,14.04759,16.602633,33.359596,30.567913,25.094292,22.885637,18.979338,15.206791,10.443094,7.610255,7.4044795,8.275595,5.919468,3.7348208,2.4795918,2.1434922,1.9514352,1.2517995,0.77165717,0.45270553,0.2469303,0.106317215,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.90541106,0.9568549,0.59331864,0.44927597,1.3409687,2.0577524,1.5810398,0.7407909,0.216064,0.53501564,1.1351935,1.2723769,1.1797781,1.2243627,1.8897027,2.7813954,3.673088,3.3781435,2.16064,1.7353712,3.391862,4.863155,4.73969,3.7965534,4.996909,7.6514096,9.386781,9.39021,8.447074,8.947794,7.970361,8.210432,10.127572,14.044161,20.128248,17.28512,13.738928,13.71492,15.806969,12.994707,9.602845,9.829198,9.383351,7.8091707,8.460793,7.442205,7.654839,7.8263187,7.5039372,7.0375133,6.036074,6.258997,6.509357,6.118384,4.9694724,4.787704,4.756838,4.273266,3.4021509,2.877424,2.6545007,2.061182,1.4027013,0.8745448,0.5453044,0.42526886,0.65162164,1.2449403,2.1263442,3.1415021,2.9220085,2.750529,3.2718265,4.064061,3.6456516,2.860276,3.7451096,4.48933,4.6573796,5.192395,4.6608095,4.262977,3.9543142,3.6868064,3.3987212,4.1429415,4.7431192,4.856296,4.623084,4.671098,4.57507,4.1463714,3.8171308,3.7759757,3.974892,3.6182148,3.7211025,3.882293,4.0949273,4.756838,5.305572,5.7377,5.909179,6.025785,6.6636887,7.284444,7.332458,6.708273,5.717122,5.051782,4.8905916,5.0312047,5.0449233,4.938606,5.1409516,4.938606,4.523626,3.9303071,3.1826572,2.294394,1.4781522,0.8676856,0.4664239,0.24350071,0.1371835,0.09945804,0.082310095,0.12003556,0.24007112,0.48357183,0.64476246,0.67219913,0.59674823,0.4972902,0.5041494,0.37039545,0.20920484,0.08573969,0.0274367,0.006859175,0.006859175,0.017147938,0.044584636,0.07888051,0.10288762,0.1097468,0.08573969,0.058302987,0.034295876,0.020577524,0.017147938,0.010288762,0.006859175,0.010288762,0.020577524,0.01371835,0.024007112,0.09602845,0.20920484,0.30866286,0.4629943,0.5007198,0.5418748,0.61389613,0.64819205,0.6893471,0.7579388,0.7956643,0.77165717,0.6790583,1.097468,1.9137098,3.0900583,4.6127954,6.468202,7.915488,9.448513,10.213311,10.062409,9.547972,8.762596,7.6274023,6.526505,5.627953,4.8905916,4.6127954,4.9248877,5.2266912,5.4907694,6.252138,7.3530354,8.172707,9.15014,10.209882,10.734609,10.566559,9.846346,10.076128,11.194174,11.585147,11.688034,12.133881,12.133881,11.427385,10.278474,8.31332,7.39762,6.2727156,4.839148,4.1635194,2.6579304,1.7182233,1.2380811,1.0631721,1.0220171,1.196926,0.83681935,0.50757897,0.39783216,0.3566771,0.432128,0.47328308,0.36353627,0.16804978,0.15090185,0.18862732,0.20234565,0.18519773,0.16462019,0.2194936,0.216064,0.20920484,0.2194936,0.20577525,0.07888051,0.1097468,0.08573969,0.041155048,0.09259886,0.4664239,0.26064864,0.2469303,0.22978236,0.15776102,0.09259886,0.106317215,0.058302987,0.01371835,0.0,0.0,0.20234565,0.18519773,0.08573969,0.017147938,0.048014224,0.216064,0.22292319,0.14747226,0.058302987,0.010288762,0.006859175,0.041155048,0.07545093,0.1371835,0.33609957,0.28122616,0.22635277,0.24350071,0.2503599,0.0,0.01371835,0.0548734,0.072021335,0.0548734,0.024007112,0.07545093,0.20920484,0.2777966,0.216064,0.024007112,0.037725464,0.30866286,0.44927597,0.39440256,0.39097297,0.37039545,0.24007112,0.14404267,0.12346515,0.116605975,0.058302987,0.072021335,0.09602845,0.08916927,0.0274367,0.034295876,0.0548734,0.061732575,0.058302987,0.07888051,0.22978236,0.3806842,0.34295875,0.19548649,0.28808534,0.24350071,0.16119061,0.07888051,0.017147938,0.0,0.26750782,0.42183927,0.39097297,0.24350071,0.20234565,0.4355576,0.41840968,0.22292319,0.010288762,0.024007112,0.017147938,0.01371835,0.020577524,0.030866288,0.041155048,0.061732575,0.06859175,0.24007112,0.47328308,0.37039545,0.17490897,0.09259886,0.13032432,0.22292319,0.23664154,0.23664154,0.1371835,0.048014224,0.020577524,0.020577524,0.037725464,0.106317215,0.26064864,0.4938606,0.7442205,0.91912943,0.82996017,0.548734,0.22292319,0.08573969,0.20920484,0.4115505,0.61046654,0.7099246,0.607037,0.8162418,0.864256,0.9842916,1.2209331,1.4267083,1.546744,1.529596,1.3924125,1.2723769,1.4438564,1.8348293,1.488441,1.0460242,0.84024894,0.88826317,1.4610043,1.488441,1.371835,1.2929544,1.1934965,0.94999576,0.9328478,1.1111864,1.2895249,1.1283343,0.5624523,0.2777966,0.14404267,0.08916927,0.07888051,0.07888051,0.14747226,0.41498008,1.1626302,2.8294096,5.24041,7.140401,7.8846216,7.281014,5.576509,2.4830213,1.255229,1.3066728,1.8999915,2.1469216,1.6804979,1.1008976,0.72364295,0.6001778,0.5178677,0.805953,0.8779744,0.8196714,0.9774324,1.99602,4.1463714,6.200694,7.3839016,7.15069,5.206114,5.7239814,5.641671,5.192395,4.7671266,4.9180284,3.8102717,3.0043187,2.726522,3.234101,4.8254294,6.0978065,6.8214493,7.4936485,8.2310095,8.786603,10.875222,12.109874,14.788382,18.770132,21.496655,17.189093,14.599753,13.5503,13.351384,12.79922,13.516005,13.845244,13.718349,13.783512,15.415996,19.908754,20.683842,20.001354,19.425184,19.823015,24.134007,26.822803,24.662163,19.229696,16.921585,18.941612,20.882757,22.902784,23.739605,20.69413,19.387459,16.564907,15.049029,15.254805,15.169065,14.757515,16.87014,19.078794,19.332584,15.9613,12.946692,13.323947,13.756075,13.066729,12.250486,10.662587,8.169277,6.2727156,5.9331865,7.5588107,5.888602,4.40702,3.998899,4.07435,2.5653315,2.9631636,3.0900583,2.49331,1.529596,1.3889829,1.7902447,1.9925903,2.287535,2.6304936,2.6167753,2.4212887,2.2052248,2.2635276,2.5241764,2.5447538,2.8739944,2.9734523,2.6613598,2.2395205,2.4555845,3.1792276,3.210094,2.7333813,2.0817597,1.7353712,1.546744,1.8656956,2.335549,2.5790498,2.170929,2.095478,2.0920484,1.9582944,1.6599203,1.3341095,1.2449403,1.0117283,0.6859175,0.39783216,0.33952916,0.34295875,0.32581082,0.36353627,0.4389872,0.44584638,0.44927597,0.4046913,0.41498008,0.4629943,0.41498008,0.34295875,0.31895164,0.29837412,0.24007112,0.12003556,0.116605975,0.12346515,0.11317638,0.1097468,0.17147937,0.22292319,0.26064864,0.21263443,0.106317215,0.07888051,0.037725464,0.034295876,0.0548734,0.1097468,0.23321195,0.5590228,0.91227025,0.94999576,0.7305021,0.71678376,0.5555932,0.33952916,0.17147937,0.08916927,0.058302987,0.061732575,0.061732575,0.037725464,0.017147938,0.082310095,0.19548649,0.23664154,0.18519773,0.08916927,0.061732575,0.08916927,0.0548734,0.044584636,0.08573969,0.15090185,0.24350071,0.19548649,0.12346515,0.06859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.11317638,0.12003556,0.09945804,0.061732575,0.024007112,0.030866288,0.024007112,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0034295875,0.006859175,0.030866288,0.106317215,0.2469303,0.6756287,2.9117198,5.6073756,7.747438,8.656279,13.9481325,18.139088,19.764713,20.893047,27.138325,30.859428,37.269325,40.89783,37.012108,21.606401,12.377381,11.05356,10.021255,8.052671,10.299051,25.622448,27.42641,25.817934,27.385256,35.215004,35.702007,27.292658,18.4649,13.63604,13.197053,7.9257765,4.431027,2.7745364,2.270387,1.4953002,0.84024894,0.5521636,0.48014224,0.4355576,0.18519773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.0548734,0.0,0.0,0.18176813,0.50757897,0.4698535,0.2709374,0.8196714,0.8779744,0.42869842,0.072021335,0.030866288,0.12003556,0.6036074,0.4355576,0.17147937,0.18176813,0.66191036,1.5810398,2.0989075,1.9445761,1.430138,1.4541451,3.6319332,4.4756117,3.882293,3.3712845,6.0703697,9.760606,11.197603,10.268185,8.779744,10.460241,8.556821,7.888051,9.249598,12.63803,17.230247,16.770683,13.577737,11.4754,11.163307,10.230459,8.97866,10.628291,10.299051,7.9429245,8.327039,6.684266,6.2247014,6.5710897,7.160979,7.274155,6.6293926,7.023795,7.298162,6.7322803,5.0655007,4.15323,4.9831905,4.8082814,3.3747141,2.901431,2.942586,2.4590142,1.879414,1.5021594,1.4918705,1.3032433,1.4541451,1.9823016,2.9631636,4.5201964,3.210094,2.4007113,2.4075704,2.8294096,2.534465,2.6716487,3.7622573,4.355576,4.3007026,4.746549,4.32471,4.5647807,4.681387,4.465323,4.290414,5.23698,5.9297566,6.355026,6.5539417,6.6122446,5.0312047,3.9337368,3.1860867,2.8465576,3.1517909,3.0043187,2.609916,2.6133456,3.175798,4.0023284,4.3624353,4.537344,4.763697,5.1683884,5.751418,6.341307,6.307011,5.7925735,5.06893,4.537344,3.9063,3.8308492,3.7691166,3.6593697,3.9200184,3.8514268,3.6387923,3.316411,2.8808534,2.277246,1.5604624,0.9534253,0.52472687,0.28122616,0.15433143,0.09602845,0.072021335,0.072021335,0.16462019,0.4972902,1.0082988,1.1351935,1.0185875,0.8093826,0.6790583,0.4972902,0.274367,0.1097468,0.0274367,0.006859175,0.0,0.0,0.006859175,0.017147938,0.017147938,0.041155048,0.034295876,0.0274367,0.020577524,0.010288762,0.01371835,0.010288762,0.0034295875,0.0034295875,0.010288762,0.0034295875,0.006859175,0.034295876,0.09602845,0.1920569,0.32924038,0.3841138,0.4046913,0.4081209,0.39097297,0.40126175,0.3566771,0.31552204,0.3018037,0.32924038,0.4972902,0.8162418,1.3306799,2.2120838,3.7451096,5.2987127,7.040943,8.309891,8.858624,8.882631,8.64942,7.939495,6.9071894,5.8543057,5.219832,4.623084,4.6676683,4.698535,4.6436615,4.996909,6.1492505,6.9620624,7.5931067,8.203573,8.954653,9.362774,9.451943,9.784613,10.398509,10.81006,11.197603,11.502836,11.533703,11.286773,10.930096,8.97523,8.169277,7.2432885,5.8508763,4.5647807,2.8088322,1.8759843,1.4953002,1.3684053,1.1763484,0.980862,0.69963586,0.58302987,0.8505377,1.6804979,1.6530612,1.1351935,0.58302987,0.28465575,0.33609957,0.3566771,0.34981793,0.26064864,0.13032432,0.06859175,0.116605975,0.106317215,0.09259886,0.072021335,0.0,0.0,0.0,0.0,0.06859175,0.33952916,0.22635277,0.3018037,0.24007112,0.048014224,0.08573969,0.05144381,0.017147938,0.0,0.020577524,0.09602845,0.22292319,0.19548649,0.10288762,0.017147938,0.0,0.22292319,0.19548649,0.11317638,0.09259886,0.17833854,0.08573969,0.06859175,0.072021335,0.12003556,0.31209245,0.26064864,0.22292319,0.24007112,0.23321195,0.0,0.0,0.030866288,0.041155048,0.034295876,0.041155048,0.14404267,0.2469303,0.29494452,0.24350071,0.061732575,0.12003556,0.37382504,0.47671264,0.36353627,0.2503599,0.22635277,0.24007112,0.24007112,0.19891608,0.13375391,0.06516216,0.024007112,0.006859175,0.01371835,0.01371835,0.058302987,0.07545093,0.06859175,0.0548734,0.061732575,0.19891608,0.34638834,0.25378948,0.0,0.0,0.08916927,0.1371835,0.09602845,0.01371835,0.0,0.09602845,0.14747226,0.116605975,0.037725464,0.006859175,0.006859175,0.006859175,0.006859175,0.01371835,0.024007112,0.01371835,0.006859175,0.010288762,0.020577524,0.034295876,0.06516216,0.11317638,0.37039545,0.66533995,0.45956472,0.13375391,0.058302987,0.14747226,0.26407823,0.21263443,0.17833854,0.106317215,0.044584636,0.020577524,0.010288762,0.020577524,0.048014224,0.13032432,0.28808534,0.53158605,0.77508676,0.8505377,0.64476246,0.2777966,0.07888051,0.16119061,0.3018037,0.41840968,0.490431,0.53501564,0.83338976,0.9294182,1.0185875,1.1763484,1.3615463,1.5638919,1.5673214,1.4061309,1.2586586,1.4507155,2.020027,1.605047,1.0871792,0.86082643,0.84024894,1.1111864,1.1180456,1.1694894,1.2826657,1.2037852,0.97057325,1.0254467,1.1489118,1.1763484,0.9877212,0.51100856,0.29494452,0.18519773,0.11317638,0.08573969,0.18862732,0.216064,0.28808534,0.5624523,1.2415106,2.651071,4.715683,5.874883,5.4633327,3.7005248,1.7902447,1.1043272,1.4267083,2.335549,3.2032347,2.8637056,2.0714707,1.3443983,1.0700313,1.5124481,1.7250825,1.5330256,1.0151579,0.6344737,1.2277923,2.9734523,4.5819287,5.778855,6.2487082,5.627953,5.9400454,5.686256,5.2781353,5.0449233,5.254128,4.4687524,3.0386145,2.1915064,2.5824795,4.3109913,5.950334,6.831738,7.39762,7.8263187,7.997798,10.353925,11.506266,13.176475,15.896138,18.993055,17.597214,14.819247,12.902108,12.47341,12.562579,13.516005,14.826107,14.424845,13.107883,14.527733,19.925903,21.44521,21.60983,21.825895,22.388348,23.76361,24.730755,24.144297,22.343761,21.163984,22.830763,24.387796,25.708187,25.571005,21.678423,21.019941,17.175373,14.483148,14.610043,16.55119,19.60695,20.183123,18.879879,16.273392,12.898679,13.828096,18.187103,19.360022,16.314548,13.598314,13.183334,11.561139,9.671436,8.738589,10.261326,8.354475,6.0737996,4.722542,4.0777793,2.4007113,3.1860867,3.391862,2.7230926,1.5364552,0.83338976,1.0597426,1.6599203,2.1229146,2.2841053,2.3046827,2.2223728,2.0646117,2.1126258,2.428148,2.8259802,3.3541365,3.4947495,2.9974594,2.2600982,2.3458378,2.503599,2.5481834,2.4418662,2.2429502,2.1091962,1.646202,1.9308578,2.3149714,2.3424082,1.7662375,2.1846473,2.1160555,1.8348293,1.5433143,1.3889829,1.3821237,1.0460242,0.66876954,0.432128,0.4115505,0.37382504,0.34638834,0.36696586,0.41498008,0.39097297,0.37725464,0.31895164,0.28808534,0.31209245,0.3841138,0.28122616,0.23321195,0.216064,0.18862732,0.09602845,0.09259886,0.1097468,0.116605975,0.11317638,0.14747226,0.14747226,0.16462019,0.13375391,0.072021335,0.0548734,0.0274367,0.017147938,0.024007112,0.041155048,0.06859175,0.29837412,0.6756287,0.7682276,0.5624523,0.45956472,0.31552204,0.25721905,0.20920484,0.15090185,0.12003556,0.1097468,0.07888051,0.0548734,0.0548734,0.082310095,0.15776102,0.19891608,0.17490897,0.08916927,0.0,0.07545093,0.037725464,0.0,0.024007112,0.12689474,0.2194936,0.21263443,0.15433143,0.07545093,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06516216,0.12003556,0.11317638,0.06859175,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.05144381,0.4115505,1.5673214,2.8911421,4.3007026,6.262427,12.13731,15.079896,15.391989,15.988737,22.419212,22.727877,28.002583,32.567364,30.34156,14.826107,7.48336,3.7622573,2.6545007,3.350707,5.254128,13.341095,18.420315,21.904776,27.786518,42.64006,43.205944,33.534508,23.19087,17.079346,15.446862,9.211872,5.0414934,2.8534167,1.9685832,1.097468,0.77508676,0.65505123,0.6927767,0.70649505,0.36353627,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1097468,0.1097468,0.0,0.0,0.0,0.072021335,0.12346515,0.13375391,0.17833854,0.3841138,0.2194936,0.048014224,0.0274367,0.11317638,0.4629943,0.45956472,0.274367,0.09259886,0.09602845,0.41840968,0.7682276,0.8196714,0.69963586,0.9877212,3.5804894,4.15323,3.275256,2.860276,6.15268,9.740028,9.606275,8.625413,9.050681,12.517994,10.635151,11.303921,12.281353,12.490558,12.010415,11.7257595,11.197603,9.685155,7.781734,7.442205,7.623973,10.340206,10.645439,8.093826,6.7185616,6.3481665,6.258997,6.557371,7.040943,7.1884155,6.7974424,6.9517736,6.9860697,6.420188,4.976331,3.8925817,5.98463,6.3893213,4.537344,4.15666,4.396731,4.1943855,3.875434,3.7039545,3.882293,3.316411,3.1449318,3.340418,4.040054,5.5147767,3.069481,2.1503513,2.4487255,3.2032347,3.2032347,3.5153272,3.9474552,3.9646032,3.5633414,3.2855449,3.0077481,3.3644254,3.9028704,4.280125,4.2526884,5.528495,6.4236174,7.377043,8.134981,7.740579,4.32471,3.0969174,2.6613598,2.369845,2.301253,2.170929,2.153781,2.4247184,2.959734,3.532475,4.1360826,4.4275975,4.623084,4.8288593,5.0414934,6.252138,6.3001523,5.768566,5.147811,4.822,4.166949,3.6525106,3.340418,3.2135234,3.1723683,2.9906003,2.74367,2.49331,2.2463799,1.9582944,1.4781522,0.97400284,0.58645946,0.35324752,0.21263443,0.13375391,0.09945804,0.082310095,0.18176813,0.6241849,1.3203912,1.4747226,1.3786942,1.1797781,0.89169276,0.64133286,0.32924038,0.106317215,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.0,0.010288762,0.01371835,0.010288762,0.0034295875,0.0,0.0034295875,0.006859175,0.010288762,0.017147938,0.041155048,0.11317638,0.15433143,0.16119061,0.14747226,0.13032432,0.15090185,0.16462019,0.17490897,0.1920569,0.20920484,0.2503599,0.37039545,0.5624523,0.8471081,1.2620882,2.194936,3.340418,4.6745276,5.926327,6.5985265,6.667118,6.7219915,6.56766,6.1561093,5.5902276,5.164959,5.23698,5.137522,4.664239,4.0880685,4.773986,5.4941993,6.1492505,6.691125,7.14726,7.0546613,8.165848,9.2153015,9.530824,9.043822,8.889491,8.886061,9.616563,10.837497,11.47197,9.798331,8.4093485,7.6651278,7.1198235,5.5319247,3.1963756,2.2806756,2.0817597,2.0474637,1.7593783,1.4987297,1.1523414,0.9534253,1.3512574,3.018037,2.9151495,1.611906,0.5727411,0.3806842,0.72021335,0.5418748,0.44927597,0.29151493,0.09259886,0.041155048,0.030866288,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.18176813,0.40126175,0.36353627,0.12689474,0.1097468,0.030866288,0.006859175,0.0034295875,0.044584636,0.216064,0.17147937,0.16804978,0.12003556,0.0274367,0.0,0.09602845,0.09602845,0.09602845,0.16804978,0.34295875,0.16462019,0.072021335,0.020577524,0.0,0.0,0.030866288,0.030866288,0.01371835,0.0,0.0,0.0,0.061732575,0.09945804,0.09602845,0.1097468,0.28122616,0.20577525,0.10288762,0.08573969,0.15433143,0.216064,0.26064864,0.24007112,0.19891608,0.26407823,0.3566771,0.37382504,0.3018037,0.16804978,0.048014224,0.030866288,0.020577524,0.020577524,0.020577524,0.01371835,0.05144381,0.0548734,0.034295876,0.01371835,0.01371835,0.07888051,0.06516216,0.0274367,0.0034295875,0.0,0.31209245,0.39783216,0.2469303,0.01371835,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.01371835,0.017147938,0.024007112,0.01371835,0.006859175,0.006859175,0.006859175,0.0034295875,0.01371835,0.034295876,0.12003556,0.29494452,0.42869842,0.24350071,0.061732575,0.048014224,0.13375391,0.22635277,0.18519773,0.12346515,0.07888051,0.048014224,0.024007112,0.0034295875,0.01371835,0.030866288,0.082310095,0.19548649,0.4115505,0.8093826,0.9911508,0.805953,0.3806842,0.11317638,0.12346515,0.14404267,0.16119061,0.25378948,0.58988905,0.939707,1.0460242,1.0734608,1.1077567,1.1420527,1.4267083,1.5227368,1.4404267,1.3203912,1.4335675,1.6427724,1.371835,1.097468,0.9774324,0.84024894,0.82996017,0.9431366,1.1592005,1.3478279,1.2689474,0.9534253,1.0700313,1.138623,0.96714365,0.65162164,0.5007198,0.5178677,0.4115505,0.1920569,0.15090185,0.41498008,0.4081209,0.30523327,0.25378948,0.39783216,0.9568549,2.0680413,2.7333813,2.5756202,1.8382589,1.1043272,0.8676856,1.1077567,1.8897027,3.3541365,3.6868064,3.1072063,2.3664153,2.1846473,3.2615378,2.8808534,2.1332035,1.2380811,0.65848076,1.0940384,2.435007,3.4021509,4.0194764,4.7602673,6.5230756,7.455923,6.7357097,5.7479887,5.1238036,4.7362604,4.6916757,3.4673128,2.2806756,2.1880767,4.098357,5.302142,6.715132,8.196714,9.249598,9.043822,9.174147,10.566559,12.120162,13.591455,15.611482,17.88873,16.13278,13.7697935,12.655178,13.05301,13.145609,14.153908,13.7697935,12.648318,14.407697,17.947031,19.13024,20.155685,21.891056,23.897366,21.225718,19.054789,18.927893,21.129688,24.682741,26.915403,28.09518,27.553307,24.795918,19.486916,19.37031,16.763824,14.006435,13.200482,16.21509,22.10712,20.989075,16.46888,11.537132,8.591117,13.502286,20.087093,21.585823,17.53548,13.749216,14.099034,14.637479,14.150477,12.747777,11.866373,9.788043,7.7783046,5.8645945,4.1360826,2.7402403,2.9665933,2.9288676,2.726522,2.2395205,1.1214751,0.72364295,1.4987297,1.8656956,1.5776103,1.7525192,1.8005334,1.845118,2.1023371,2.585909,3.1072063,3.525616,3.724532,3.2032347,2.2841053,2.1023371,1.8588364,1.7936742,1.9274281,2.1400626,2.170929,1.862266,1.8897027,1.7765263,1.4781522,1.3889829,2.136633,2.0508933,1.6084765,1.2243627,1.2449403,1.3272504,0.9877212,0.65162164,0.4938606,0.44927597,0.38754338,0.44927597,0.48014224,0.41840968,0.31895164,0.37382504,0.33952916,0.274367,0.24007112,0.31209245,0.21263443,0.15090185,0.15090185,0.17490897,0.12003556,0.09602845,0.10288762,0.12003556,0.1371835,0.15433143,0.15433143,0.18176813,0.17833854,0.12346515,0.05144381,0.037725464,0.024007112,0.030866288,0.058302987,0.08916927,0.1097468,0.25378948,0.41840968,0.5453044,0.61046654,0.490431,0.42869842,0.3566771,0.28122616,0.2777966,0.22292319,0.16462019,0.16119061,0.16804978,0.05144381,0.058302987,0.08916927,0.106317215,0.07888051,0.010288762,0.07888051,0.041155048,0.0034295875,0.0034295875,0.010288762,0.058302987,0.11317638,0.12003556,0.072021335,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13375391,0.13375391,0.08573969,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0,0.0034295875,0.0,0.0,0.006859175,0.01371835,0.041155048,0.15090185,0.61046654,1.2106444,1.7010754,2.942586,6.9071894,9.259886,8.045813,7.8126,10.981539,17.837284,14.496866,18.62609,21.843042,18.831865,7.3118806,2.3424082,0.78537554,0.72364295,1.1077567,1.7319417,3.1792276,7.781734,13.834956,21.407484,32.32386,29.748241,24.60729,20.244854,17.518333,14.805529,8.580828,4.650521,2.4247184,1.3581166,0.9568549,0.9945804,0.9534253,0.94999576,0.91227025,0.5796003,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09259886,0.5418748,0.44584638,0.19548649,0.0274367,0.01371835,0.01371835,0.061732575,0.14061308,0.20577525,0.16804978,0.06859175,0.37382504,1.0048691,1.4781522,0.91569984,1.4644338,1.8862731,2.2155135,2.819121,4.3933015,6.800872,7.274155,7.3530354,8.405919,11.626302,8.796892,9.578837,8.934075,6.3824625,6.029215,7.8331776,6.8866115,5.878313,5.5147767,4.5030484,4.8185706,5.6485305,5.844017,5.3398676,5.1580997,5.693115,6.029215,6.4990683,6.883182,6.4098988,5.6142344,5.1409516,4.746549,4.3178506,3.8925817,4.07435,5.2472687,6.001778,6.1458206,6.684266,7.548522,8.207003,8.56025,8.495089,7.874333,6.5196457,6.1629686,6.1492505,6.135532,6.0875177,4.90431,5.038064,5.453044,5.4736214,4.791134,4.437886,4.9248877,6.029215,7.010077,6.6053853,4.2389703,3.0248961,3.450165,4.6402316,4.3487167,6.385892,6.914048,7.390761,7.9943686,7.630832,3.8925817,2.503599,1.8691251,1.3615463,1.313532,1.6427724,1.8348293,2.0406046,2.287535,2.4555845,3.0420442,3.8205605,4.5784993,5.23698,5.857735,7.8606143,8.069819,7.3427467,6.3481665,5.552502,5.3090014,4.9180284,4.338428,3.683377,3.2203827,2.8534167,2.5619018,2.2806756,1.9823016,1.6770682,1.371835,0.9945804,0.66533995,0.44584638,0.33609957,0.22635277,0.16119061,0.12346515,0.13375391,0.24350071,0.61046654,0.9294182,1.3203912,1.587899,1.2209331,0.84367853,0.39097297,0.1097468,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.01371835,0.024007112,0.0,0.01371835,0.034295876,0.0274367,0.0034295875,0.01371835,0.041155048,0.044584636,0.041155048,0.034295876,0.044584636,0.044584636,0.044584636,0.06516216,0.09602845,0.12346515,0.14747226,0.216064,0.29494452,0.37382504,0.45613512,0.86082643,1.3649758,2.0714707,2.8980014,3.5702004,4.2046742,4.9214582,5.56965,5.8474464,5.3090014,4.6882463,4.338428,4.3590055,4.554492,4.4550343,4.016047,4.280125,4.835718,5.377593,5.7068334,5.6348124,5.9812007,6.831738,7.7851634,7.98065,8.1041155,7.747438,7.4936485,7.613684,8.1041155,8.237869,8.9100685,8.429926,6.667118,5.0826488,4.139512,3.566771,3.3609958,3.199805,2.4555845,2.4075704,1.9548649,1.4747226,1.1763484,1.1146159,0.9431366,0.72707254,0.4938606,0.48700142,1.1592005,0.41498008,0.34638834,0.31895164,0.1371835,0.07545093,0.12346515,0.09945804,0.058302987,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.12346515,0.14404267,0.22292319,0.29151493,0.061732575,0.01371835,0.017147938,0.024007112,0.034295876,0.106317215,0.020577524,0.09259886,0.1097468,0.037725464,0.0,0.0,0.044584636,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.08573969,0.15776102,0.12346515,0.048014224,0.020577524,0.044584636,0.14404267,0.34981793,0.216064,0.1371835,0.1371835,0.23664154,0.45613512,0.5796003,0.37382504,0.13375391,0.01371835,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.017147938,0.024007112,0.01371835,0.0,0.6824879,0.6344737,0.29837412,0.01371835,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.01371835,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.0,0.01371835,0.01371835,0.034295876,0.048014224,0.0,0.01371835,0.061732575,0.15776102,0.26064864,0.26064864,0.1371835,0.06859175,0.041155048,0.0274367,0.01371835,0.01371835,0.024007112,0.08573969,0.25378948,0.59674823,1.1694894,1.4232788,1.1043272,0.4424168,0.1371835,0.2469303,0.16462019,0.12689474,0.2709374,0.6241849,0.77165717,0.864256,0.9568549,1.0425946,1.0666018,1.5673214,1.7388009,1.6187652,1.3855534,1.371835,1.3855534,1.1317638,0.88826317,0.75450927,0.65505123,0.607037,0.9877212,1.3615463,1.4164196,0.9774324,0.8676856,0.96714365,1.0151579,0.9431366,0.8711152,1.1008976,1.3512574,1.0220171,0.32238123,0.274367,0.5693115,0.6790583,0.5693115,0.34638834,0.274367,0.34638834,0.77851635,1.1008976,1.1797781,1.1900668,1.3375391,1.2072148,1.1660597,1.4747226,2.3046827,3.426158,3.6525106,3.5873485,3.8342788,5.020916,3.9954693,2.3732746,1.2449403,0.90884066,0.8848336,1.786815,2.3424082,2.7539587,3.5564823,5.6313825,5.861165,5.7274113,5.844017,6.2247014,6.2864337,5.284994,3.981751,2.7539587,2.2292318,3.2821152,4.122364,6.1286726,8.862054,11.043272,10.542552,8.81061,11.592006,15.055889,16.671225,15.182784,17.830425,19.390888,18.646667,16.688372,16.921585,16.993607,14.79867,12.562579,11.63659,12.466551,12.624311,12.041282,13.7697935,17.86815,21.407484,19.270851,16.026463,14.781522,16.112202,18.067066,27.124607,34.99208,35.369335,27.84825,17.899017,13.55373,11.122152,10.010965,10.2921915,12.710052,16.20137,14.812388,11.852654,9.249598,7.5519514,10.628291,14.006435,15.748666,15.004445,12.037852,11.355364,12.850664,13.88297,13.207341,10.984968,8.848335,7.455923,6.3618846,5.353586,4.4241676,3.059192,3.0900583,3.309552,3.0729103,2.3046827,1.1934965,1.2003556,1.4129901,1.4335675,1.371835,1.5673214,1.6633499,1.8519772,2.1674993,2.4727325,2.568761,2.5378947,2.551613,2.4555845,1.786815,1.786815,1.5844694,1.5947582,1.8416885,1.937717,2.2566686,2.6716487,2.270387,1.3512574,1.4507155,1.8142518,1.9342873,1.611906,1.0871792,1.039165,1.0014396,0.9568549,0.8162418,0.59674823,0.4115505,0.4972902,0.64819205,0.67219913,0.548734,0.42869842,0.5624523,0.5041494,0.37039545,0.26407823,0.274367,0.21263443,0.12346515,0.082310095,0.09602845,0.106317215,0.082310095,0.07545093,0.06516216,0.044584636,0.044584636,0.082310095,0.20234565,0.25721905,0.19891608,0.07545093,0.05144381,0.037725464,0.041155048,0.07545093,0.1371835,0.15090185,0.25378948,0.37039545,0.4629943,0.548734,0.82996017,0.77165717,0.6310441,0.5693115,0.65505123,0.48357183,0.432128,0.45613512,0.45613512,0.26064864,0.05144381,0.037725464,0.037725464,0.010288762,0.044584636,0.010288762,0.010288762,0.010288762,0.010288762,0.044584636,0.044584636,0.044584636,0.05144381,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18176813,0.16462019,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.006859175,0.07888051,0.33609957,0.72707254,1.1900668,1.6187652,2.1194851,3.0351849,6.893471,11.190743,11.567999,8.05953,5.0826488,5.8645945,6.910619,7.8674736,8.556821,8.971801,3.07634,0.7133542,0.14747226,0.29151493,0.71678376,1.3752645,3.57363,6.228131,8.776315,11.170166,14.599753,19.5315,24.127148,26.10945,22.765602,9.506817,3.5839188,1.6564908,1.3958421,1.4815818,1.3821237,1.039165,0.823101,0.7888051,0.64133286,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.1097468,0.08916927,0.072021335,0.07888051,0.0274367,0.006859175,0.01371835,0.058302987,0.12003556,0.13032432,0.05144381,0.09945804,0.22635277,0.32238123,0.2194936,0.53501564,0.9774324,1.371835,1.9342873,3.2821152,4.928317,4.7191124,4.938606,5.675967,4.8151407,3.6936657,5.144381,6.2075534,6.6293926,8.882631,8.570539,6.307011,4.650521,4.3795834,4.48933,4.0949273,4.417309,5.813151,7.407909,7.099246,5.7891436,5.164959,5.0895076,5.178677,4.8082814,4.1326528,3.5942078,3.3747141,3.433017,3.525616,3.981751,4.629943,5.2918534,5.950334,6.7322803,7.394191,7.750868,8.128122,8.529384,8.628842,7.490219,6.416758,6.0154963,6.48535,7.6274023,7.798882,8.580828,9.431366,9.702303,8.635701,6.944915,6.0806584,5.8371577,5.8645945,5.6656785,5.2335505,5.0277753,5.2472687,6.0326443,7.4970784,7.8091707,6.0497923,4.8185706,4.756838,4.5647807,3.9954693,3.3712845,2.318401,1.1111864,0.6893471,0.764798,0.7339317,0.66191036,0.6001778,0.5658819,0.70306545,1.1249046,1.7353712,2.3458378,2.6853669,3.8377085,5.0277753,6.0395036,6.759717,7.1781263,7.8331776,7.5931067,6.7494283,5.6176643,4.537344,3.6627994,3.2306714,2.9151495,2.534465,2.0337453,1.6290541,1.2346514,0.8848336,0.61389613,0.44584638,0.31552204,0.22635277,0.17490897,0.15776102,0.17147937,0.4972902,0.64133286,1.0117283,1.4781522,1.3684053,1.4678634,0.922559,0.35324752,0.058302987,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.0034295875,0.006859175,0.024007112,0.041155048,0.037725464,0.030866288,0.037725464,0.0274367,0.0034295875,0.01371835,0.07888051,0.1097468,0.082310095,0.030866288,0.034295876,0.044584636,0.05144381,0.061732575,0.07888051,0.12346515,0.106317215,0.1371835,0.19891608,0.2709374,0.34638834,0.52472687,0.78194594,1.1351935,1.5158776,1.786815,2.1194851,3.2306714,4.3109913,4.8151407,4.4447455,3.7622573,3.3987212,3.4433057,3.7485392,3.9543142,3.683377,3.5770597,3.7725463,4.2218223,4.7191124,4.8494368,4.671098,4.880303,5.7377,7.06495,6.8145905,6.677407,7.0958166,8.06639,9.139851,9.908078,9.6817255,8.182996,6.4716315,6.924337,7.0478024,5.8474464,4.6402316,3.899441,3.2615378,2.9974594,2.6407824,2.4795918,2.486451,2.2978237,1.5604624,1.6564908,1.8725548,1.7456601,1.0494537,0.71678376,0.53844523,0.40126175,0.26750782,0.19891608,0.1097468,0.058302987,0.030866288,0.020577524,0.037725464,0.017147938,0.0034295875,0.0,0.017147938,0.08573969,0.072021335,0.072021335,0.07545093,0.058302987,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.017147938,0.06859175,0.4629943,0.24350071,0.020577524,0.006859175,0.0,0.0,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.030866288,0.024007112,0.020577524,0.044584636,0.13032432,0.26064864,0.40126175,0.45270553,0.36010668,0.31895164,0.42526886,0.65162164,0.48357183,0.20920484,0.037725464,0.01371835,0.01371835,0.0034295875,0.0034295875,0.006859175,0.010288762,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.14747226,0.13032432,0.058302987,0.0034295875,0.01371835,0.12003556,0.1097468,0.12346515,0.4424168,1.4815818,0.7682276,0.23664154,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0034295875,0.034295876,0.106317215,0.20234565,0.26064864,0.22635277,0.12003556,0.041155048,0.017147938,0.01371835,0.01371835,0.024007112,0.061732575,0.17147937,0.4355576,0.77508676,0.90541106,0.66876954,0.28122616,0.30866286,0.29151493,0.1920569,0.15433143,0.26407823,0.5418748,0.6001778,0.61046654,0.72021335,0.94999576,1.1763484,1.4438564,1.8416885,1.8999915,1.5844694,1.2895249,1.3203912,1.0117283,0.7990939,0.77508676,0.71678376,0.66876954,1.1454822,1.6290541,1.7730967,1.3924125,1.1832076,1.0700313,1.0563129,1.1592005,1.4061309,1.3272504,1.08032,0.64819205,0.23664154,0.28808534,0.490431,0.70306545,0.7305021,0.61389613,0.6276145,0.45613512,0.44584638,0.51100856,0.64476246,0.922559,1.097468,1.1317638,1.1111864,1.3958421,2.5961976,4.081209,5.1580997,5.720552,5.878313,5.960623,4.7774153,2.8259802,1.6187652,1.3889829,1.08032,1.3786942,2.0234566,2.819121,4.0537724,6.509357,5.950334,5.8371577,6.0703697,6.2727156,5.785714,4.8254294,3.3609958,2.4041407,2.411,3.3061223,4.8905916,7.6651278,9.815479,10.340206,9.067829,8.213862,10.364213,13.570878,15.927004,15.560039,18.063637,19.21255,18.396307,16.894148,17.899017,16.849564,14.562028,13.176475,13.13532,13.173045,12.181894,10.988399,10.436234,11.22161,13.900118,16.060759,17.816708,18.79414,18.732407,17.494326,23.808197,32.629097,33.97349,25.9414,14.723219,13.183334,12.627741,15.933864,22.041958,25.989414,20.646116,15.9921665,12.984418,11.533703,10.532263,10.501397,11.14273,11.592006,11.396519,10.501397,10.676306,10.47396,11.331357,12.614022,11.619442,8.790032,6.3310184,4.588788,3.799983,4.0846386,3.9371665,3.2203827,2.767677,2.9048605,3.4638834,1.6976458,0.939707,1.1111864,1.7113642,1.8382589,1.3581166,1.2037852,1.4369972,1.9308578,2.3732746,2.2566686,1.879414,1.6667795,1.670209,1.5638919,1.4095604,1.4164196,1.5947582,2.085189,3.1723683,2.5001693,2.2498093,1.9582944,1.5673214,1.3992717,1.3478279,1.5604624,1.5673214,1.2689474,0.9294182,0.9294182,0.8505377,0.7442205,0.65848076,0.6310441,0.75450927,0.8779744,0.8848336,0.764798,0.6241849,0.58988905,0.50757897,0.39440256,0.30523327,0.28808534,0.26407823,0.17833854,0.09602845,0.058302987,0.06859175,0.12346515,0.13032432,0.106317215,0.10288762,0.1920569,0.30866286,0.34981793,0.32581082,0.2503599,0.1371835,0.09259886,0.06516216,0.058302987,0.072021335,0.11317638,0.1920569,0.21263443,0.1920569,0.19548649,0.32924038,0.5041494,0.42526886,0.29151493,0.21263443,0.24007112,0.18862732,0.17833854,0.22978236,0.29837412,0.30866286,0.061732575,0.030866288,0.034295876,0.01371835,0.020577524,0.034295876,0.044584636,0.0548734,0.07888051,0.15433143,0.09602845,0.24350071,0.28465575,0.14747226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15433143,0.09259886,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.006859175,0.006859175,0.030866288,0.14061308,0.4424168,0.7956643,1.2106444,1.8073926,2.8294096,3.357566,3.3129816,2.6853669,1.7799559,1.2243627,1.7696671,2.7813954,4.108646,6.2075534,10.120712,3.0214665,0.5590228,0.116605975,0.21263443,0.47328308,0.94656616,1.9102802,3.8685746,6.584808,9.095266,11.372512,17.607502,24.994833,30.029469,28.489584,13.642899,5.6793966,2.369845,1.6256244,1.5158776,1.0563129,0.72364295,0.6173257,0.6893471,0.7373613,0.0,0.0,0.0,0.0,0.024007112,0.11317638,0.09602845,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06859175,0.20577525,0.34295875,0.082310095,0.006859175,0.01371835,0.037725464,0.048014224,0.020577524,0.01371835,0.01371835,0.06859175,0.3018037,0.77165717,1.2998136,1.7490896,2.1812177,2.867135,3.3678548,3.0660512,2.8054025,2.9220085,3.2306714,3.7725463,4.9523244,6.2864337,7.6925645,9.469091,10.6488695,10.484249,8.597976,5.8234396,4.2286816,3.7211025,3.7348208,5.2438393,7.3873315,7.4936485,5.3981705,4.262977,3.82399,3.7108135,3.457024,3.0969174,3.0283258,3.3952916,4.0434837,4.540774,5.3741636,5.669108,6.0875177,6.694555,6.9654922,7.2295704,7.706283,8.436785,9.153569,9.249598,7.8983397,6.9380555,6.944915,7.939495,9.3936405,9.510246,9.688584,9.794902,9.523964,8.416207,6.420188,5.164959,4.5819287,4.5030484,4.671098,5.1683884,5.895461,6.4133286,6.5710897,6.4819202,5.24041,3.5976372,2.5996273,2.417859,2.3424082,2.9151495,2.8568463,2.1229146,1.0700313,0.4698535,0.44584638,0.37039545,0.26407823,0.15433143,0.082310095,0.08573969,0.2709374,0.6276145,0.9534253,0.8848336,1.3341095,2.294394,3.6319332,5.305572,7.3839016,9.294182,9.554831,8.920357,7.9875093,7.191845,6.125243,5.2987127,4.547633,3.82399,3.199805,2.393852,1.7216529,1.2072148,0.84367853,0.61046654,0.44584638,0.32581082,0.24350071,0.19891608,0.17147937,0.28465575,0.3018037,0.6344737,1.1866373,1.3581166,1.1832076,0.64133286,0.22978236,0.09259886,0.05144381,0.030866288,0.017147938,0.010288762,0.006859175,0.0,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.0,0.010288762,0.020577524,0.041155048,0.09945804,0.08916927,0.061732575,0.037725464,0.030866288,0.041155048,0.1097468,0.16119061,0.14061308,0.06859175,0.041155048,0.044584636,0.048014224,0.0548734,0.06516216,0.08573969,0.0548734,0.061732575,0.13032432,0.2469303,0.3566771,0.44927597,0.5178677,0.65848076,0.89169276,1.1489118,1.3409687,1.879414,2.4315774,2.7642474,2.7333813,2.6819375,2.4898806,2.4624438,2.6304936,2.7573884,2.6064866,2.702515,2.8122618,3.000889,3.6113555,4.0194764,4.1017866,4.256118,4.671098,5.305572,5.9983487,6.375603,6.4373355,6.5230756,7.3118806,9.170717,9.277034,8.416207,7.98065,9.983529,8.735159,6.0703697,4.2938433,4.1292233,4.7259717,4.6436615,4.098357,3.9268777,4.0777793,3.6113555,2.510458,2.6853669,2.8259802,2.4041407,1.6804979,1.039165,0.66191036,0.52815646,0.4938606,0.274367,0.07888051,0.020577524,0.010288762,0.13375391,0.65162164,0.13375391,0.0034295875,0.0,0.006859175,0.041155048,0.024007112,0.020577524,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.22978236,0.11317638,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.07545093,0.18519773,0.29837412,0.39097297,0.48357183,0.7510797,0.4698535,0.22978236,0.23321195,0.28122616,0.18176813,0.06859175,0.006859175,0.006859175,0.006859175,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.1371835,0.19891608,0.16462019,0.06516216,0.0,0.0034295875,0.0034295875,0.006859175,0.08573969,0.35324752,0.52472687,0.4355576,0.5144381,0.9911508,1.8725548,0.7339317,0.17833854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.010288762,0.044584636,0.09945804,0.15090185,0.23321195,0.12689474,0.034295876,0.024007112,0.01371835,0.024007112,0.05144381,0.06516216,0.09602845,0.22292319,0.3806842,0.40126175,0.28808534,0.15090185,0.22292319,0.16804978,0.13375391,0.18176813,0.3566771,0.70306545,0.65848076,0.58302987,0.6962063,0.9911508,1.2415106,1.471293,1.7010754,1.6839274,1.4369972,1.2380811,1.0700313,0.77165717,0.6001778,0.6207553,0.6962063,0.78537554,1.2929544,1.4815818,1.3101025,1.4507155,1.7456601,1.6324836,1.3512574,1.1489118,1.2586586,1.0185875,0.71678376,0.41840968,0.23664154,0.30866286,0.5727411,0.70306545,0.66533995,0.5418748,0.53501564,0.5007198,0.36010668,0.28808534,0.3841138,0.6790583,1.1351935,0.9842916,0.8676856,1.155771,1.9651536,3.6044965,5.521636,6.8626046,7.226141,6.6705475,4.870014,2.9460156,1.8725548,1.7902447,1.9994495,2.1229146,2.7745364,3.6970954,4.7602673,5.9880595,5.2301207,5.360445,5.453044,5.06893,4.232111,3.6970954,3.2581081,2.9940298,2.9288676,3.000889,5.0277753,7.6685576,9.06097,8.748878,7.7097125,7.5416627,8.934075,11.413667,14.280802,16.588915,19.500635,20.570665,19.922474,18.46147,17.878439,15.902997,14.452282,13.704632,13.097594,11.317638,11.502836,11.413667,10.408798,9.410788,10.88894,13.63261,15.6869335,16.918156,17.655516,18.684393,20.855322,23.93852,23.36235,19.267422,16.513464,17.099922,15.028452,16.088194,20.975357,25.303495,19.651537,15.700651,14.212211,14.013294,12.017275,10.539123,9.736599,10.14129,11.245617,11.489118,11.602294,11.441104,12.754636,14.393978,12.312219,8.793462,5.960623,3.875434,2.8396983,3.3747141,3.474172,3.3815732,2.9391565,2.6236343,3.5530527,2.3424082,1.3478279,2.136633,4.1943855,4.928317,3.1895163,1.5536032,0.9911508,1.5536032,2.3595562,1.9171394,1.5707511,1.3821237,1.3546871,1.4541451,1.4061309,1.5364552,1.7833855,2.1332035,2.6373527,1.8519772,1.5021594,1.430138,1.4369972,1.2689474,1.5810398,1.9857311,1.8039631,1.1283343,0.83681935,1.0254467,0.97400284,0.84024894,0.7442205,0.77851635,0.78194594,0.8128122,0.8676856,0.8676856,0.66191036,0.52472687,0.4698535,0.4115505,0.31209245,0.20920484,0.216064,0.24007112,0.19548649,0.09259886,0.05144381,0.082310095,0.08916927,0.09945804,0.1371835,0.23664154,0.32238123,0.33266997,0.2777966,0.18519773,0.09602845,0.072021335,0.05144381,0.041155048,0.05144381,0.08916927,0.28122616,0.32924038,0.28465575,0.22292319,0.22978236,0.37382504,0.36010668,0.2469303,0.13032432,0.12003556,0.1371835,0.15090185,0.17147937,0.18519773,0.17490897,0.041155048,0.01371835,0.01371835,0.020577524,0.06859175,0.06516216,0.06859175,0.106317215,0.14061308,0.072021335,0.044584636,0.18176813,0.20920484,0.082310095,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.05144381,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14061308,0.06859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.01371835,0.0,0.0,0.0034295875,0.0034295875,0.006859175,0.037725464,0.14747226,0.33952916,0.6790583,1.1420527,1.605047,1.371835,0.7579388,0.29494452,0.16119061,0.15776102,0.48700142,0.94656616,1.821111,5.960623,18.811287,5.6348124,1.0185875,0.1371835,0.20234565,0.45613512,0.6001778,1.0700313,3.1106358,6.667118,10.371073,9.753747,12.836946,17.566347,21.150267,20.073376,11.393089,5.7068334,2.8054025,1.8656956,1.4438564,0.84367853,0.548734,0.5041494,0.6173257,0.77165717,0.0,0.0,0.0,0.0,0.020577524,0.106317215,0.09602845,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.19548649,0.36696586,0.08916927,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.1097468,0.5041494,1.2106444,1.587899,1.7010754,1.7147937,1.8999915,2.1503513,2.4555845,2.3218307,2.2429502,3.6970954,4.763697,5.271276,5.9914894,7.010077,7.7131424,8.570539,9.6988735,8.824328,6.15268,4.383013,3.0626216,2.7299516,3.6285036,5.06893,5.40503,4.166949,3.789694,3.5599117,3.1860867,2.784825,2.8122618,3.5393343,4.897451,6.625963,8.292743,9.455373,8.862054,8.06639,7.723431,7.6033955,7.7131424,7.9292064,8.285883,8.64599,8.687145,7.874333,7.6857057,8.14527,8.913498,9.294182,8.831187,8.529384,8.165848,7.613684,6.848886,5.970912,5.518206,5.192395,4.7499785,4.0057583,4.07435,4.6882463,5.1855364,5.0895076,4.108646,2.7333813,1.8348293,1.3478279,1.1866373,1.2449403,1.8416885,2.1263442,1.8348293,1.097468,0.432128,0.29151493,0.20234565,0.1371835,0.082310095,0.044584636,0.037725464,0.09259886,0.216064,0.31209245,0.16462019,0.20920484,0.71678376,1.704505,3.2375305,5.429037,7.7885933,8.779744,8.776315,8.423067,8.639131,8.213862,7.442205,6.4133286,5.3673043,4.695105,3.7279615,2.7368107,1.9274281,1.3649758,0.9945804,0.69963586,0.4972902,0.36010668,0.26750782,0.20234565,0.17833854,0.16119061,0.6344737,1.3924125,1.546744,0.90884066,0.39783216,0.14061308,0.09602845,0.06859175,0.041155048,0.024007112,0.01371835,0.01371835,0.0,0.006859175,0.0034295875,0.0,0.0,0.006859175,0.0,0.006859175,0.010288762,0.024007112,0.082310095,0.07888051,0.0548734,0.034295876,0.034295876,0.0548734,0.106317215,0.16804978,0.18176813,0.13375391,0.06859175,0.05144381,0.041155048,0.044584636,0.0548734,0.061732575,0.034295876,0.024007112,0.07545093,0.17490897,0.26064864,0.31895164,0.34981793,0.4424168,0.6207553,0.84367853,0.9568549,0.99801,1.0357354,1.1180456,1.2517995,1.5433143,1.587899,1.6187652,1.6976458,1.7079345,1.6393428,1.8073926,1.903421,2.0680413,2.884283,3.1346428,3.5702004,4.012617,4.372724,4.629943,5.3844523,5.809721,5.6210938,5.1066556,5.127233,6.931196,7.3393173,7.3050213,7.8434668,10.045261,8.899779,6.3721733,4.705394,4.664239,5.521636,5.579939,4.5647807,4.012617,4.0949273,3.6113555,2.7745364,2.8122618,2.7162333,2.2463799,1.9514352,1.2037852,0.66876954,0.42869842,0.3841138,0.24350071,0.048014224,0.0,0.0,0.12689474,0.6310441,0.12689474,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.07545093,0.18519773,0.2777966,0.33609957,0.4046913,0.5796003,0.30866286,0.082310095,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.010288762,0.041155048,0.13375391,0.32581082,0.51100856,0.64819205,0.59331864,0.09602845,0.17147937,0.26407823,0.32924038,0.42183927,0.66533995,0.7373613,0.51100856,0.48357183,0.77851635,1.1351935,0.35324752,0.061732575,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.030866288,0.05144381,0.14061308,0.082310095,0.030866288,0.0274367,0.020577524,0.08573969,0.18176813,0.15776102,0.0548734,0.08916927,0.13375391,0.1097468,0.072021335,0.061732575,0.09602845,0.05144381,0.06859175,0.17490897,0.39783216,0.7579388,0.7133542,0.65162164,0.6859175,0.85739684,1.1214751,1.5261664,1.5398848,1.3375391,1.1180456,1.1180456,0.89512235,0.6893471,0.52815646,0.4698535,0.6276145,0.864256,1.2209331,1.2346514,1.097468,1.6324836,2.0165975,1.7559488,1.2758065,0.88826317,0.823101,0.6276145,0.4629943,0.35324752,0.3018037,0.2709374,0.5144381,0.58302987,0.548734,0.45956472,0.34981793,0.39097297,0.30866286,0.24350071,0.30866286,0.6001778,1.0117283,0.7613684,0.6173257,0.8265306,1.1351935,2.2292318,4.290414,6.2041235,7.2192817,6.9517736,4.2355404,2.6785078,2.1400626,2.4144297,3.2306714,3.5804894,3.998899,4.681387,5.422178,5.6210938,4.7945633,4.513337,4.2046742,3.683377,3.1415021,2.4007113,2.3492675,2.4212887,2.3732746,2.2669573,3.9508848,6.0806584,7.5450926,7.8777623,7.2638664,7.058091,7.881192,9.743458,12.432255,15.532601,19.329155,20.817596,20.803877,19.95334,18.79757,16.568336,14.654627,13.306799,12.205902,10.4533825,11.55428,11.96926,11.180455,10.179015,11.461681,12.830087,14.335675,15.415996,16.088194,16.945591,16.88729,16.904436,16.403717,16.770683,21.393766,24.075705,22.161995,19.888178,18.879879,18.142517,17.309128,16.88043,16.564907,15.453721,12.024134,10.031544,9.431366,10.710602,12.843805,13.3033695,12.939834,13.073587,14.671775,15.940722,12.312219,8.584257,6.0635104,4.2115335,3.0351849,3.1072063,2.8054025,3.0454736,3.0969174,2.959734,3.350707,2.8122618,2.2223728,3.3438478,5.675967,6.4544835,4.787704,2.1434922,0.8711152,1.4129901,2.2909644,1.6599203,1.4953002,1.5433143,1.7010754,1.9925903,2.0165975,1.8759843,1.9274281,2.1263442,2.037175,1.4747226,1.3889829,1.3443983,1.2689474,1.4335675,1.8554068,2.2978237,1.9171394,0.980862,0.8848336,1.1592005,1.0563129,0.85396725,0.7407909,0.8025235,0.75450927,0.7579388,0.82996017,0.881404,0.7305021,0.4972902,0.48014224,0.48014224,0.39097297,0.18176813,0.18862732,0.2503599,0.25721905,0.18862732,0.12003556,0.07888051,0.072021335,0.09602845,0.15776102,0.2503599,0.2503599,0.22978236,0.17490897,0.10288762,0.048014224,0.048014224,0.037725464,0.034295876,0.05144381,0.08916927,0.29151493,0.5144381,0.7373613,0.8505377,0.6310441,0.64476246,0.607037,0.4629943,0.274367,0.20920484,0.22635277,0.1920569,0.14404267,0.1097468,0.08916927,0.09945804,0.06859175,0.030866288,0.020577524,0.06859175,0.05144381,0.048014224,0.082310095,0.106317215,0.017147938,0.037725464,0.14061308,0.15090185,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.082310095,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1097468,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.048014224,0.058302987,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.061732575,0.24007112,0.48357183,0.6173257,0.65848076,0.50757897,0.34295875,0.23664154,0.17833854,0.30866286,0.33609957,0.89512235,4.8494368,17.28512,5.6073756,1.2175035,0.18176813,0.16462019,0.42183927,0.37725464,0.8128122,2.983741,6.7940125,10.765475,10.882081,11.739478,13.241637,14.7026415,14.853543,11.585147,7.606825,4.4996185,2.7916842,1.9685832,1.313532,0.78537554,0.53844523,0.61389613,0.9362774,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.0548734,0.072021335,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.1097468,0.44584638,1.2003556,1.3889829,1.0631721,0.6036074,0.72707254,1.9685832,2.6716487,2.784825,2.7642474,3.5976372,4.232111,4.3041325,4.249259,4.297273,4.461893,3.3266997,4.5682106,5.5319247,5.2815647,4.623084,2.5447538,1.8382589,1.7902447,1.9274281,2.0337453,2.3801336,3.2992632,3.7005248,3.4981792,3.5976372,3.5942078,4.7328305,6.7185616,9.170717,11.657167,12.768354,11.417097,9.561689,8.40249,8.40249,8.471081,7.98065,7.380472,7.040943,7.2535777,7.6342616,8.405919,9.019815,8.903209,7.449064,6.776865,6.6568294,6.3207297,5.65539,5.223262,5.8508763,6.509357,6.5710897,5.6519604,3.6079261,2.7368107,2.644212,2.8465576,2.935727,2.5790498,2.0989075,1.605047,1.2175035,1.039165,1.1351935,1.587899,2.4658735,2.760818,2.1194851,0.85396725,0.29151493,0.06859175,0.010288762,0.0,0.0,0.020577524,0.048014224,0.082310095,0.12346515,0.18519773,0.13375391,0.41840968,0.94656616,1.6736387,2.5961976,4.40702,5.936616,6.660259,6.9723516,8.186425,8.683716,8.440215,7.6033955,6.560801,5.960623,5.1821065,4.029765,2.9494452,2.1503513,1.5913286,1.0768905,0.7579388,0.5624523,0.4389872,0.33266997,0.28808534,0.2777966,0.86082643,1.7456601,1.7765263,0.9774324,0.47328308,0.1920569,0.07545093,0.061732575,0.024007112,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.0,0.010288762,0.020577524,0.017147938,0.010288762,0.041155048,0.072021335,0.13032432,0.17490897,0.18176813,0.106317215,0.058302987,0.034295876,0.030866288,0.041155048,0.0548734,0.041155048,0.024007112,0.0274367,0.0548734,0.06859175,0.10288762,0.19548649,0.31552204,0.42526886,0.4938606,0.5453044,0.5144381,0.4355576,0.37382504,0.432128,0.5761707,0.78537554,0.97057325,1.08032,1.0940384,1.0768905,1.0666018,1.1180456,1.4164196,2.2909644,2.2498093,2.8499873,3.5770597,4.214963,4.8425775,4.73969,4.8082814,4.846007,4.6848164,4.1943855,4.972902,5.254128,5.3570156,5.717122,6.8797526,7.298162,6.39961,5.3878818,4.8905916,4.945465,5.0277753,3.7931237,2.9288676,2.8259802,2.5893385,2.3835633,2.153781,1.8176813,1.488441,1.4541451,1.1146159,0.64819205,0.23321195,0.05144381,0.26407823,0.09259886,0.08573969,0.11317638,0.09602845,0.037725464,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.106317215,0.17147937,0.22978236,0.07545093,0.01371835,0.0,0.0,0.0,0.0,0.020577524,0.034295876,0.037725464,0.037725464,0.08573969,0.09259886,0.082310095,0.07545093,0.106317215,0.08573969,0.0548734,0.0548734,0.12689474,0.28808534,0.5418748,0.9294182,1.2449403,1.155771,0.21263443,0.37382504,0.5521636,0.65848076,0.6756287,0.6379033,0.548734,0.26064864,0.061732575,0.020577524,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.0,0.0034295875,0.010288762,0.017147938,0.017147938,0.017147938,0.01371835,0.020577524,0.024007112,0.0274367,0.0274367,0.16804978,0.32581082,0.26407823,0.0548734,0.05144381,0.05144381,0.034295876,0.020577524,0.01371835,0.0274367,0.017147938,0.037725464,0.1371835,0.32581082,0.6001778,0.6962063,0.7407909,0.6824879,0.6310441,0.8779744,1.4610043,1.4061309,1.0940384,0.84367853,0.9294182,0.88826317,0.77508676,0.5727411,0.4046913,0.5418748,0.8711152,0.96371406,1.0254467,1.2415106,1.7593783,1.7730967,1.3101025,0.84367853,0.59331864,0.5007198,0.4355576,0.4046913,0.4081209,0.37725464,0.20577525,0.30866286,0.37725464,0.45270553,0.4664239,0.24007112,0.19548649,0.2194936,0.24350071,0.31895164,0.6173257,0.72021335,0.6173257,0.5418748,0.5624523,0.5727411,0.7407909,2.411,4.5167665,6.138962,6.5299344,3.3438478,2.3252604,2.3835633,3.1380725,4.90431,5.90575,5.73427,5.562791,5.720552,5.7102633,4.8117113,3.6353626,2.8396983,2.609916,2.6853669,1.4232788,0.9259886,0.85396725,1.0254467,1.4095604,2.3046827,3.981751,6.1286726,7.7714453,7.281014,6.701414,7.281014,8.687145,10.542552,12.421966,16.979887,19.483486,20.467777,20.457489,19.980776,18.019053,14.88441,12.641459,11.900668,11.808069,13.063298,12.785502,12.05157,12.000127,13.831526,13.9481325,15.182784,16.012743,15.419425,12.88496,12.823228,14.188204,16.03675,19.006773,25.303495,30.643364,31.415022,28.204927,21.918493,13.80066,17.315987,20.19341,19.52807,15.409137,10.902658,8.738589,9.040393,11.163307,13.653188,14.263655,14.123041,14.949572,16.479168,16.71238,11.938394,8.279024,6.3138704,4.9214582,3.806842,3.4776018,3.1415021,3.0454736,3.4055803,3.8274195,3.3026927,3.0351849,3.2821152,4.2526884,5.4187484,5.521636,4.887162,2.469303,1.1832076,1.646202,2.1469216,1.4747226,1.5330256,1.9754424,2.5001693,2.8534167,2.867135,2.2978237,1.9582944,2.0165975,2.0131679,1.5981878,1.7388009,1.6153357,1.2792361,1.6667795,1.8348293,2.0817597,1.6736387,0.88826317,0.9842916,1.2072148,1.0323058,0.8025235,0.70306545,0.7510797,0.7373613,0.7956643,0.83681935,0.83338976,0.82996017,0.5590228,0.53158605,0.5555932,0.5007198,0.28808534,0.28122616,0.25721905,0.25721905,0.26750782,0.21263443,0.14404267,0.12689474,0.14404267,0.1920569,0.2709374,0.18519773,0.12003556,0.07545093,0.05144381,0.034295876,0.044584636,0.041155048,0.058302987,0.09259886,0.12346515,0.22635277,0.6310441,1.2449403,1.7079345,1.3821237,1.1900668,1.0117283,0.77851635,0.5418748,0.4698535,0.4115505,0.28122616,0.17833854,0.15776102,0.22292319,0.26064864,0.20234565,0.116605975,0.05144381,0.044584636,0.034295876,0.034295876,0.0274367,0.017147938,0.041155048,0.09259886,0.20234565,0.2194936,0.11317638,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.072021335,0.061732575,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072021335,0.058302987,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.09259886,0.10288762,0.08573969,0.0274367,0.017147938,0.006859175,0.0,0.0,0.006859175,0.020577524,0.037725464,0.037725464,0.07888051,0.29151493,0.6824879,0.7442205,0.59674823,0.39097297,0.29837412,0.29494452,0.24007112,0.8093826,2.4967396,5.6519604,2.6133456,0.980862,0.28122616,0.13375391,0.29151493,0.23321195,0.7579388,2.7402403,6.2727156,10.652299,13.584596,14.812388,15.038741,15.169065,16.307688,15.090185,11.763485,8.038953,5.103226,3.625074,2.5961976,1.5021594,0.8162418,0.7442205,1.2243627,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.3841138,1.0597426,1.1626302,0.8471081,1.313532,4.2046742,3.1620796,1.4232788,0.64476246,0.90198153,1.5844694,2.1572106,2.085189,1.5570327,1.4953002,2.411,6.0635104,8.018375,6.7459984,3.6456516,3.6593697,2.8396983,1.8554068,1.1043272,0.70306545,0.9842916,1.4267083,2.1674993,3.7313912,7.06495,5.7719955,5.7411294,6.447624,7.1781263,7.0203657,7.2021337,7.267296,7.5519514,8.097256,8.621983,8.097256,7.1061053,6.3173003,6.118384,6.608815,7.486789,8.628842,9.167287,8.47451,6.1801167,6.5710897,7.034084,6.2041235,4.3590055,3.4192986,3.4776018,3.5393343,3.5770597,3.4604537,2.959734,2.7162333,3.1689389,3.7348208,3.957744,3.4947495,2.8945718,2.3081124,1.9171394,1.7079345,1.4644338,2.5996273,5.2918534,6.958633,6.138962,2.503599,0.8162418,0.20577525,0.044584636,0.0,0.0,0.09602845,0.24007112,0.4115505,0.5521636,0.5658819,0.6001778,0.8025235,1.1489118,1.6221949,2.1812177,3.2306714,4.372724,5.3261495,6.101236,7.0032177,7.0889573,7.1849856,7.0443726,6.680836,6.3618846,5.802862,4.8185706,3.7862647,2.9117198,2.2292318,1.5090185,1.097468,0.90884066,0.83338976,0.7476501,0.6241849,0.5212973,0.58988905,0.8848336,1.371835,1.1420527,0.5796003,0.18176813,0.08573969,0.061732575,0.024007112,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.041155048,0.017147938,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0274367,0.058302987,0.09945804,0.13032432,0.106317215,0.058302987,0.0274367,0.01371835,0.017147938,0.030866288,0.017147938,0.006859175,0.006859175,0.020577524,0.044584636,0.06859175,0.09602845,0.12346515,0.15090185,0.15090185,0.16462019,0.16804978,0.1371835,0.09259886,0.09259886,0.17833854,0.28122616,0.40126175,0.53158605,0.64133286,0.65162164,0.66533995,0.65162164,0.66876954,0.84024894,1.5090185,2.2086544,2.7402403,3.1346428,3.6456516,3.865145,4.057202,4.413879,4.8905916,5.219832,5.9400454,6.1458206,5.4187484,4.290414,4.2423997,3.7553983,3.340418,2.9974594,2.8088322,2.9288676,3.199805,3.0729103,2.8705647,2.7230926,2.5619018,2.428148,1.9274281,1.3066728,0.7682276,0.48700142,0.7579388,0.805953,0.47671264,0.14061308,0.70306545,0.33609957,0.4355576,0.5590228,0.47671264,0.18176813,0.13375391,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.12346515,0.25378948,0.29151493,0.058302987,0.0,0.0,0.0,0.0,0.0,0.09945804,0.17833854,0.19548649,0.18176813,0.42869842,0.4698535,0.4081209,0.36353627,0.47328308,0.37382504,0.21263443,0.17147937,0.2503599,0.274367,0.8128122,1.5124481,1.3786942,0.50757897,0.09259886,0.16462019,0.12689474,0.061732575,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.01371835,0.01371835,0.020577524,0.030866288,0.030866288,0.006859175,0.0,0.006859175,0.01371835,0.01371835,0.1371835,0.22292319,0.1920569,0.07545093,0.01371835,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.06859175,0.17490897,0.3806842,0.7099246,0.8676856,0.85396725,0.7682276,0.7922347,1.1111864,1.1797781,1.0597426,0.8711152,0.8093826,0.9911508,0.7442205,0.48357183,0.39440256,0.4424168,0.83338976,0.82996017,0.7990939,0.881404,0.9911508,1.1008976,0.91912943,0.7476501,0.6962063,0.67219913,0.53844523,0.51100856,0.4698535,0.36353627,0.22978236,0.216064,0.24007112,0.34638834,0.4115505,0.16804978,0.14404267,0.16462019,0.20920484,0.28808534,0.45613512,0.6790583,0.86082643,0.805953,0.5727411,0.48700142,0.48700142,2.2360911,4.1429415,5.212973,5.0655007,3.199805,2.5310357,2.3835633,3.426158,7.675417,9.860064,8.656279,6.619104,5.305572,5.295283,4.513337,3.192946,2.177788,1.7696671,1.7079345,1.2586586,0.89855194,0.7579388,0.86082643,1.1283343,1.9342873,3.590778,5.5833683,6.9037595,6.0737996,6.108095,6.694555,7.3564653,8.220721,10.041832,14.1299,18.28313,20.20027,19.576086,18.11165,16.170506,14.393978,13.88297,14.38369,14.29795,16.520323,15.470869,14.147048,14.0750265,15.319967,16.736387,16.383139,15.920145,15.227368,12.421966,11.921246,13.121602,15.265094,18.11165,21.956219,31.08921,33.699127,33.33902,30.643364,23.345201,22.95423,24.02083,21.04052,14.198492,9.352485,6.8763227,6.557371,7.939495,10.30934,12.7272,15.193072,18.87302,20.412905,18.238546,12.572867,8.385342,6.3310184,4.7019644,3.4295874,4.0880685,5.7754254,5.579939,4.914599,4.3281393,3.508468,3.1552205,4.15666,5.0483527,5.1409516,4.530485,3.2135234,2.061182,1.7730967,2.1332035,1.9994495,1.2415106,1.5913286,2.4590142,3.1449318,2.8534167,2.9631636,2.5961976,1.9685832,1.5638919,2.136633,1.5124481,1.2655178,1.4061309,1.5913286,1.1283343,1.4815818,1.4164196,1.0254467,0.64133286,0.823101,1.0185875,1.0494537,0.9774324,0.86082643,0.7613684,0.64133286,0.77508676,0.83681935,0.7682276,0.7922347,0.65848076,0.53501564,0.45956472,0.45613512,0.5178677,0.5796003,0.42183927,0.25721905,0.17833854,0.15090185,0.20234565,0.24007112,0.26064864,0.2709374,0.31895164,0.17490897,0.072021335,0.030866288,0.034295876,0.044584636,0.044584636,0.06516216,0.12003556,0.18519773,0.19891608,0.22292319,0.5041494,1.1077567,1.7490896,1.786815,1.5536032,1.2106444,0.89855194,0.7510797,0.8848336,0.7373613,0.5658819,0.47328308,0.5144381,0.6859175,0.490431,0.36010668,0.26407823,0.1920569,0.16804978,0.15433143,0.14404267,0.106317215,0.0548734,0.030866288,0.09259886,0.26407823,0.31209245,0.18176813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.1097468,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072021335,0.14747226,0.14747226,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.044584636,0.082310095,0.1371835,0.1371835,0.08916927,0.030866288,0.0,0.006859175,0.030866288,0.0548734,0.16119061,0.1371835,0.048014224,0.24350071,0.67219913,0.823101,0.65162164,0.33609957,0.274367,0.2503599,0.31895164,0.58645946,1.1111864,1.8931323,1.2929544,0.86082643,0.5178677,0.26407823,0.16804978,0.034295876,0.3841138,1.8485477,5.9297566,14.997586,14.363112,16.503176,17.566347,16.2974,14.037301,14.832966,15.001016,13.080446,9.534253,6.773435,4.3692946,2.585909,1.471293,1.0666018,1.4198492,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.07545093,0.32238123,0.42526886,0.34981793,0.33609957,1.5398848,1.1077567,0.548734,0.47671264,0.607037,0.52815646,0.58988905,0.5624523,0.42869842,0.39783216,3.8137012,7.06495,7.31531,4.763697,2.6716487,2.2429502,1.8313997,1.3375391,0.85396725,0.66533995,0.6241849,0.6962063,1.6633499,3.8445675,7.0889573,5.5422134,4.90431,4.822,4.928317,4.846007,6.327589,8.584257,10.281903,10.7586155,10.014396,9.750318,9.403929,8.735159,8.038953,8.155559,8.597976,9.301042,9.897789,9.595985,7.191845,6.351596,6.385892,6.310441,5.7411294,4.870014,3.9851806,3.391862,3.1826572,3.1792276,2.9220085,2.668219,2.74367,2.9906003,3.223812,3.2375305,3.2649672,3.059192,2.6647894,2.1915064,1.8313997,2.4590142,3.6970954,4.386442,3.8925817,2.0989075,0.90198153,0.37382504,0.13375391,0.0,0.0,0.020577524,0.048014224,0.16119061,0.31209245,0.34638834,0.37039545,0.52815646,0.7579388,1.1146159,1.7559488,2.7368107,3.6696587,4.506478,5.206114,5.7582774,5.717122,5.627953,5.7308407,6.0497923,6.385892,5.9331865,5.0277753,4.1429415,3.4398763,2.7642474,1.9582944,1.5193073,1.2895249,1.1454822,0.9911508,0.8025235,0.7099246,0.6927767,0.72707254,0.7888051,0.61389613,0.35324752,0.17490897,0.116605975,0.072021335,0.0548734,0.044584636,0.034295876,0.0274367,0.037725464,0.0274367,0.017147938,0.01371835,0.01371835,0.01371835,0.041155048,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.017147938,0.017147938,0.024007112,0.044584636,0.058302987,0.0274367,0.010288762,0.0034295875,0.0034295875,0.006859175,0.01371835,0.01371835,0.01371835,0.020577524,0.034295876,0.0274367,0.044584636,0.06516216,0.07545093,0.06859175,0.058302987,0.06516216,0.06859175,0.072021335,0.09259886,0.08916927,0.106317215,0.14404267,0.20577525,0.28808534,0.32924038,0.3566771,0.37382504,0.39097297,0.4355576,0.6276145,0.89512235,1.3546871,2.020027,2.767677,3.6216443,4.557922,5.1100855,5.219832,5.267846,5.4976287,5.2781353,4.266407,3.0454736,3.093488,3.3987212,3.457024,3.4055803,3.2135234,2.7093742,2.959734,3.4227283,3.6799474,3.40901,2.3801336,2.1400626,2.037175,1.8725548,1.5055889,0.85396725,0.6824879,0.5796003,0.5453044,0.5761707,0.6276145,0.34981793,0.4081209,0.4698535,0.4629943,0.548734,0.13032432,0.2503599,0.34981793,0.23664154,0.1097468,0.07888051,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.048014224,0.0,0.0,0.01371835,0.030866288,0.05144381,0.058302987,0.010288762,0.0,0.010288762,0.0274367,0.037725464,0.15433143,0.5178677,0.66191036,0.5178677,0.42869842,0.66191036,0.45270553,0.30523327,0.29837412,0.09602845,0.07545093,0.058302987,0.22978236,0.50757897,0.5418748,0.6893471,0.58302987,0.35324752,0.12003556,0.017147938,0.034295876,0.024007112,0.01371835,0.0034295875,0.0034295875,0.0,0.0,0.034295876,0.20577525,0.6824879,0.72364295,0.32238123,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.010288762,0.010288762,0.0034295875,0.01371835,0.01371835,0.01371835,0.017147938,0.017147938,0.017147938,0.01371835,0.0034295875,0.0,0.0034295875,0.0034295875,0.048014224,0.082310095,0.07888051,0.034295876,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.006859175,0.01371835,0.034295876,0.09602845,0.23664154,0.5144381,0.77508676,0.8505377,0.84367853,1.1111864,1.0768905,0.94999576,0.8676856,0.91912943,1.1489118,1.0906088,0.8676856,0.6344737,0.50757897,0.5761707,0.64476246,0.5453044,0.47328308,0.5007198,0.6001778,0.6344737,0.6207553,0.7373613,0.91227025,0.8162418,0.53844523,0.4629943,0.42526886,0.33952916,0.216064,0.17490897,0.14747226,0.15433143,0.16462019,0.106317215,0.11317638,0.14747226,0.17490897,0.20577525,0.29837412,0.64476246,0.9911508,1.0014396,0.7682276,0.8162418,0.6036074,1.529596,2.9906003,4.2766957,4.588788,3.4535947,2.2806756,2.0303159,3.542764,7.5279446,10.621432,10.2236,8.244728,6.3653145,6.0395036,5.970912,5.4736214,4.57507,3.2615378,1.4541451,0.90198153,1.1420527,1.4507155,1.8382589,3.0454736,3.7142432,4.2252517,5.099797,6.2727156,7.0752387,7.130112,7.64798,8.05953,8.340756,9.026674,11.866373,16.263103,19.507494,20.45063,19.504065,17.679523,17.662374,18.910746,19.579515,16.506605,16.191082,17.53891,18.46147,18.118511,16.942162,17.031332,18.639809,20.471207,20.793589,17.436022,13.704632,15.110763,17.61779,21.174273,29.696798,34.470783,36.25074,33.48992,26.85367,19.233126,16.479168,14.688923,12.027563,9.253027,9.709162,9.047252,8.06296,8.385342,10.943813,15.947581,19.692692,18.108221,16.554619,16.407146,15.038741,14.582606,13.227919,9.849775,5.7994323,4.8940215,5.826869,5.381023,4.6436615,4.2698364,4.4859004,3.673088,3.7965534,4.629943,5.5147767,5.3741636,3.4878905,3.4604537,3.1689389,2.1057668,1.3752645,1.5570327,2.1640697,2.4898806,2.2635276,1.670209,1.6633499,1.6907866,1.6324836,1.5604624,1.7319417,1.4438564,1.3649758,1.4918705,1.6187652,1.3478279,1.2449403,1.155771,0.91912943,0.6036074,0.5418748,0.7888051,1.0048691,0.9911508,0.77851635,0.64133286,0.5761707,0.66191036,0.7442205,0.7510797,0.64819205,0.5521636,0.4355576,0.36353627,0.3566771,0.4081209,0.45956472,0.44584638,0.37382504,0.2709374,0.18862732,0.16119061,0.19548649,0.21263443,0.18519773,0.1371835,0.07888051,0.044584636,0.041155048,0.061732575,0.082310095,0.072021335,0.07545093,0.11317638,0.23664154,0.5041494,0.50757897,0.70306545,1.1283343,1.7182233,2.311542,2.1846473,1.6359133,1.1694894,0.9877212,0.9945804,1.4747226,1.6153357,1.529596,1.3101025,1.039165,0.85396725,0.5521636,0.30523327,0.21263443,0.2777966,0.2469303,0.11317638,0.08573969,0.14747226,0.0548734,0.09602845,0.2194936,0.2469303,0.14404267,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.058302987,0.07888051,0.1097468,0.072021335,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.12346515,0.16804978,0.11317638,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.0274367,0.07888051,0.15090185,0.16119061,0.17147937,0.106317215,0.07888051,0.12346515,0.17833854,0.20234565,0.26407823,0.31209245,0.29151493,0.14747226,0.31895164,0.5178677,0.5007198,0.29494452,0.22635277,0.30866286,0.28465575,0.39440256,0.66533995,0.9294182,0.53501564,0.25378948,0.19548649,0.39440256,0.8162418,0.29837412,0.16804978,1.0700313,3.5359046,7.956643,17.271402,21.013083,21.263443,18.883308,13.488567,14.692352,15.405707,16.859852,17.12393,11.084427,6.090947,3.3747141,2.0989075,1.6976458,1.8965619,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.09945804,0.11317638,0.1097468,0.45956472,0.29494452,0.14747226,0.18519773,0.23321195,0.14061308,0.12689474,0.11317638,0.07545093,0.058302987,2.7951138,4.170378,3.7108135,2.4041407,2.6990852,4.0537724,2.651071,1.2175035,0.7682276,0.61046654,0.48014224,0.6241849,1.8005334,3.875434,5.796003,3.590778,3.3541365,3.806842,4.1360826,3.974892,5.9640527,7.4456344,7.874333,7.363324,6.691125,7.2192817,7.390761,7.006647,6.4098988,6.495639,7.438775,8.182996,8.841476,8.875772,7.099246,6.118384,5.9571934,6.3961806,6.8900414,6.5710897,5.3090014,4.1429415,3.5702004,3.532475,3.4192986,3.0523329,2.901431,2.8980014,2.9734523,3.0626216,3.4535947,3.2409601,2.6819375,2.0474637,1.6221949,1.7250825,1.903421,1.8725548,1.4987297,0.7990939,0.37039545,0.16804978,0.061732575,0.0,0.0,0.0,0.017147938,0.0548734,0.10288762,0.116605975,0.15433143,0.23664154,0.36696586,0.59331864,0.9877212,1.5501735,2.1846473,2.7813954,3.2889743,3.707384,3.9200184,4.1772375,4.5853586,5.1066556,5.56965,5.4496145,5.003768,4.4241676,3.799983,3.1380725,2.417859,1.8999915,1.5433143,1.2895249,1.0528834,1.0151579,0.939707,0.8745448,0.83681935,0.823101,0.83338976,0.77851635,0.64476246,0.45613512,0.26064864,0.18862732,0.14404267,0.12346515,0.1097468,0.09945804,0.08916927,0.082310095,0.06859175,0.048014224,0.024007112,0.034295876,0.020577524,0.010288762,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0034295875,0.01371835,0.037725464,0.0274367,0.010288762,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.01371835,0.006859175,0.024007112,0.037725464,0.037725464,0.017147938,0.01371835,0.020577524,0.030866288,0.037725464,0.044584636,0.05144381,0.058302987,0.061732575,0.06859175,0.09602845,0.12346515,0.14404267,0.15776102,0.16804978,0.18176813,0.22292319,0.29494452,0.490431,0.8265306,1.2312219,2.2806756,3.9954693,5.40503,5.861165,5.0243454,4.729401,4.2218223,3.6319332,3.1655092,3.100347,2.884283,4.016047,4.3795834,3.4878905,2.4898806,2.7059445,3.340418,3.426158,2.8568463,2.3904223,2.9048605,2.942586,2.5207467,1.7765263,0.97400284,0.85396725,0.8505377,0.8676856,0.89169276,0.9842916,0.9568549,0.8505377,0.61389613,0.36696586,0.40126175,0.25721905,0.42183927,0.48700142,0.3566771,0.25721905,0.2194936,0.15433143,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.030866288,0.037725464,0.037725464,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.18176813,0.59331864,0.8848336,0.70649505,0.24007112,0.19548649,0.28808534,0.17833854,0.1097468,0.12346515,0.06516216,0.048014224,0.030866288,0.20234565,0.5212973,0.7099246,0.38754338,0.16119061,0.044584636,0.010288762,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.041155048,0.33609957,0.71678376,1.0220171,1.138623,0.89512235,0.36353627,0.030866288,0.0034295875,0.010288762,0.0034295875,0.006859175,0.010288762,0.010288762,0.01371835,0.010288762,0.006859175,0.006859175,0.006859175,0.006859175,0.01371835,0.010288762,0.010288762,0.01371835,0.01371835,0.024007112,0.020577524,0.01371835,0.006859175,0.0,0.010288762,0.024007112,0.0274367,0.017147938,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.0034295875,0.0034295875,0.01371835,0.048014224,0.12346515,0.29151493,0.47671264,0.5418748,0.5555932,0.805953,0.64133286,0.61046654,0.6927767,0.84024894,0.99801,0.9259886,0.84024894,0.72707254,0.6379033,0.7099246,0.69963586,0.5453044,0.42526886,0.42183927,0.5041494,0.5658819,0.58988905,0.6824879,0.77851635,0.6241849,0.4389872,0.5727411,0.66191036,0.5658819,0.34295875,0.2194936,0.19891608,0.18519773,0.14404267,0.1097468,0.13032432,0.15433143,0.16462019,0.17833854,0.26064864,0.50757897,0.8128122,0.8779744,0.7682276,0.881404,1.2449403,2.311542,3.4776018,4.32128,4.6093655,3.6936657,2.3149714,1.8828435,3.3026927,6.9792104,11.118723,11.55771,10.192734,8.344186,6.756287,5.627953,5.717122,5.40503,4.125794,2.386993,1.4232788,1.6393428,2.1057668,2.5310357,3.2306714,3.0317552,3.216953,3.8274195,4.866585,6.2727156,6.3310184,6.584808,6.8043017,7.0615206,7.720001,9.3764925,12.188754,15.357693,18.139088,19.833303,22.04539,24.4461,25.841942,24.819925,19.723558,18.886738,19.312008,20.255144,20.508932,18.410025,15.728088,15.6869335,17.46003,19.322296,18.636377,16.21852,17.103354,21.006224,27.810524,37.543694,38.624016,36.56626,31.888304,25.752771,19.970488,16.80155,15.391989,13.090735,10.497967,11.451392,10.967821,9.160428,8.591117,10.1481495,13.035862,14.904987,15.100473,14.695783,14.616901,15.666355,17.885298,16.760393,12.898679,8.165848,5.693115,5.1821065,4.4275975,3.9337368,3.782835,3.6147852,2.8911421,2.6064866,3.4433057,4.856296,5.07236,3.4844608,3.2649672,3.1655092,3.0386145,3.8205605,5.003768,4.5442033,3.0660512,1.5844694,1.4918705,1.587899,1.3958421,1.2517995,1.2689474,1.3478279,1.2449403,1.2517995,1.5261664,1.8313997,1.5604624,1.3409687,1.214074,0.9568549,0.6173257,0.5453044,0.65505123,0.7373613,0.7339317,0.65505123,0.5727411,0.48014224,0.5178677,0.5727411,0.5796003,0.51100856,0.53501564,0.5144381,0.47328308,0.44584638,0.4629943,0.45270553,0.432128,0.37725464,0.29151493,0.216064,0.20577525,0.2469303,0.25721905,0.20577525,0.12003556,0.05144381,0.044584636,0.06859175,0.09945804,0.09945804,0.082310095,0.15433143,0.2709374,0.41840968,0.6173257,0.8711152,1.313532,1.821111,2.2738166,2.551613,2.7093742,2.294394,1.728512,1.2998136,1.1489118,1.5364552,1.7250825,1.8142518,1.8073926,1.5947582,1.5021594,1.2037852,0.9259886,0.7099246,0.4046913,0.28122616,0.16119061,0.1371835,0.17490897,0.116605975,0.2194936,0.4664239,0.53844523,0.33952916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.048014224,0.0548734,0.09259886,0.0548734,0.037725464,0.072021335,0.12346515,0.048014224,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10288762,0.15433143,0.116605975,0.07545093,0.06516216,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.07888051,0.106317215,0.14061308,0.15776102,0.15433143,0.11317638,0.12689474,0.21263443,0.29494452,0.2469303,0.22978236,0.29151493,0.34981793,0.20577525,0.25721905,0.53844523,0.5555932,0.26750782,0.12346515,0.15776102,0.12346515,0.18176813,0.3566771,0.51100856,0.4046913,0.15090185,0.048014224,0.19891608,0.53844523,0.3806842,0.33609957,0.72707254,1.8142518,3.7691166,8.916927,14.140189,22.885637,30.766829,25.571005,31.384155,30.578201,22.755312,12.88839,11.345076,7.1849856,5.1580997,3.7211025,2.4795918,2.170929,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.072021335,0.12003556,0.07545093,0.030866288,0.024007112,0.030866288,0.06516216,0.09602845,0.08916927,0.044584636,0.010288762,1.1626302,1.3752645,1.039165,0.91227025,2.1194851,3.7553983,2.3492675,0.96714365,0.6927767,0.6036074,0.48357183,1.0906088,2.2052248,3.3644254,3.841138,2.6236343,2.9803114,4.201245,4.962613,3.3129816,4.3178506,4.5270553,4.016047,3.2135234,2.8980014,3.5839188,4.0057583,3.9440255,3.6010668,3.5702004,4.715683,5.5250654,6.0737996,6.1904054,5.4324665,4.9214582,4.8597255,5.429037,6.279575,6.5230756,5.717122,4.633373,4.0194764,3.8788633,3.4913201,2.9700227,2.7368107,2.6133456,2.5001693,2.3561265,2.6476414,2.393852,1.8725548,1.3203912,0.96714365,0.8025235,0.59674823,0.37382504,0.16804978,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.017147938,0.0,0.0,0.030866288,0.05144381,0.10288762,0.19891608,0.32924038,0.5041494,0.8025235,1.1008976,1.3821237,1.7559488,2.1983654,2.6887965,3.2306714,3.7965534,4.3178506,4.6882463,4.8151407,4.7259717,4.461893,4.0709205,3.4055803,2.7642474,2.2600982,1.9068506,1.6256244,1.5741806,1.4404267,1.2826657,1.1489118,1.0666018,1.2277923,1.4335675,1.4404267,1.1763484,0.7407909,0.5178677,0.39097297,0.3018037,0.22978236,0.1920569,0.20920484,0.216064,0.20234565,0.16119061,0.10288762,0.07545093,0.05144381,0.030866288,0.020577524,0.020577524,0.010288762,0.0034295875,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0034295875,0.006859175,0.017147938,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.006859175,0.01371835,0.017147938,0.01371835,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.0274367,0.05144381,0.05144381,0.034295876,0.017147938,0.030866288,0.037725464,0.041155048,0.041155048,0.058302987,0.10288762,0.09945804,0.10288762,0.14747226,0.2469303,0.9259886,2.287535,3.6525106,4.482471,4.383013,4.623084,4.297273,4.091498,4.1600895,4.15666,3.549623,4.389872,4.5647807,3.5873485,2.5824795,2.568761,2.6853669,2.4795918,1.9891608,1.7490896,2.4727325,2.7642474,2.5001693,1.8519772,1.2860953,1.2106444,1.1489118,1.138623,1.1832076,1.2792361,1.1523414,0.9328478,0.6241849,0.34295875,0.31895164,0.45270553,0.6001778,0.58988905,0.4629943,0.4698535,0.8128122,0.59331864,0.34638834,0.2503599,0.12689474,0.030866288,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.0034295875,0.017147938,0.020577524,0.01371835,0.037725464,0.01371835,0.0034295875,0.024007112,0.048014224,0.0,0.0,0.006859175,0.0548734,0.18862732,0.45270553,0.67219913,0.6859175,0.4115505,0.037725464,0.01371835,0.0034295875,0.0,0.0,0.01371835,0.06516216,0.058302987,0.10288762,0.21263443,0.36353627,0.48014224,0.13375391,0.09259886,0.07545093,0.0034295875,0.0,0.0,0.006859175,0.024007112,0.048014224,0.048014224,0.15776102,0.5418748,0.8848336,0.9911508,0.7956643,0.53158605,0.23664154,0.106317215,0.1371835,0.106317215,0.030866288,0.01371835,0.01371835,0.010288762,0.010288762,0.01371835,0.010288762,0.010288762,0.01371835,0.006859175,0.01371835,0.017147938,0.030866288,0.08916927,0.24007112,0.42869842,0.33266997,0.14747226,0.006859175,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.006859175,0.0034295875,0.006859175,0.024007112,0.05144381,0.14061308,0.24007112,0.28465575,0.31209245,0.45613512,0.32924038,0.36696586,0.5007198,0.6756287,0.83338976,0.7476501,0.66876954,0.6379033,0.6824879,0.8162418,0.8025235,0.59674823,0.4355576,0.42526886,0.5521636,0.70306545,0.78537554,0.8093826,0.75450927,0.5521636,0.4972902,0.71678376,0.89512235,0.8471081,0.5178677,0.31209245,0.25378948,0.21263443,0.14747226,0.1097468,0.14747226,0.15090185,0.15090185,0.16804978,0.19891608,0.30866286,0.48357183,0.5555932,0.5555932,0.7339317,1.903421,3.6387923,4.681387,4.7362604,4.4859004,3.5702004,2.5481834,2.836269,4.3041325,5.2781353,8.838047,9.750318,9.342196,8.330468,6.848886,5.65539,6.060081,5.8817425,4.482471,2.7711067,1.9342873,2.3972816,3.210094,3.673088,3.3301294,2.5001693,2.6236343,3.2786856,4.2766957,5.6793966,6.375603,6.9620624,7.4010496,7.682276,7.8434668,8.076678,9.626852,12.055,15.093615,18.643238,22.724447,25.872808,27.241213,26.400965,23.334913,22.261452,21.04395,20.978786,21.407484,19.730417,15.244516,13.245067,13.992717,16.695232,19.53493,19.675543,21.256582,25.663603,32.046066,37.32763,37.862644,34.926918,30.948597,26.486704,20.237995,19.586374,17.960749,14.445422,10.984968,12.38767,11.694893,9.431366,8.378482,9.091836,9.89436,9.911508,13.55373,16.654078,16.986746,14.280802,15.6869335,15.892709,13.786942,10.017825,6.9723516,5.9126086,4.5270553,3.74168,3.5153272,2.843128,2.0817597,1.9754424,2.8534167,4.190956,4.5853586,3.9783216,4.064061,4.3041325,4.7019644,5.768566,6.0635104,5.4839106,4.07435,2.9185789,4.1360826,3.4055803,2.2841053,1.4095604,1.0837497,1.2895249,1.1694894,1.7182233,2.2635276,2.301253,1.529596,1.471293,1.2998136,1.0185875,0.77851635,0.85739684,0.8848336,0.72364295,0.58988905,0.6001778,0.7922347,0.6276145,0.64476246,0.6962063,0.7339317,0.83338976,0.64133286,0.5212973,0.4972902,0.52815646,0.52472687,0.48700142,0.41498008,0.33952916,0.2777966,0.216064,0.19891608,0.22635277,0.25378948,0.24350071,0.18519773,0.082310095,0.0548734,0.07888051,0.116605975,0.12346515,0.09259886,0.19891608,0.5796003,1.2380811,2.0577524,2.1126258,1.9651536,1.9857311,2.2258022,2.411,2.760818,2.7882545,2.4452958,1.8656956,1.371835,1.4644338,1.7696671,2.1057668,2.318401,2.2841053,2.218943,1.8005334,1.4232788,1.1454822,0.6927767,0.42526886,0.24007112,0.17147937,0.20234565,0.274367,0.4389872,0.78194594,0.8196714,0.4629943,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05144381,0.12003556,0.09259886,0.09945804,0.05144381,0.024007112,0.044584636,0.072021335,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08573969,0.11317638,0.06859175,0.044584636,0.07888051,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07888051,0.106317215,0.106317215,0.116605975,0.18862732,0.25378948,0.22978236,0.22292319,0.26750782,0.32581082,0.24350071,0.18862732,0.21263443,0.26750782,0.216064,0.23321195,0.42869842,0.41840968,0.17833854,0.037725464,0.030866288,0.010288762,0.048014224,0.14747226,0.28122616,0.274367,0.1097468,0.0,0.030866288,0.15776102,0.25721905,0.29837412,0.4389872,0.89855194,1.9857311,2.8259802,6.848886,17.237106,29.08633,29.412142,34.144974,29.467016,18.005335,6.948344,8.025234,6.4887795,6.125243,5.288424,3.7176728,2.5413244,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.058302987,0.037725464,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.034295876,0.048014224,0.05144381,0.0274367,0.08573969,0.16462019,0.17490897,0.10288762,0.0,0.06859175,0.26407823,0.37039545,0.44584638,0.8025235,0.94999576,0.7133542,0.77851635,1.0871792,0.85396725,0.7990939,3.0351849,4.040054,3.0043187,1.8279701,2.7299516,3.7211025,4.9591837,5.284994,2.2086544,1.6633499,1.3341095,1.0734608,0.84367853,0.72364295,0.89169276,1.2620882,1.4232788,1.2723769,1.0357354,1.7182233,2.3492675,2.6407824,2.6476414,2.7573884,2.7813954,2.9563043,3.3850029,4.0057583,4.588788,4.5647807,4.1155047,3.8274195,3.6216443,2.7539587,2.1057668,1.8965619,1.786815,1.5570327,1.1214751,1.0734608,0.90884066,0.66191036,0.40126175,0.23321195,0.09602845,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.07888051,0.17833854,0.45270553,0.8848336,1.2723769,1.7113642,2.2360911,2.8259802,3.6079261,4.1429415,4.5339146,4.8185706,4.962613,4.506478,3.9303071,3.457024,3.1415021,2.9048605,2.6716487,2.411,2.1057668,1.7593783,1.3992717,1.4747226,1.821111,1.9994495,1.8005334,1.2209331,0.864256,0.64476246,0.4698535,0.32581082,0.274367,0.32581082,0.34295875,0.33952916,0.31895164,0.2709374,0.21263443,0.14747226,0.09259886,0.0548734,0.041155048,0.024007112,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0034295875,0.01371835,0.0274367,0.020577524,0.006859175,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.010288762,0.034295876,0.044584636,0.030866288,0.0,0.017147938,0.020577524,0.01371835,0.006859175,0.024007112,0.08916927,0.072021335,0.048014224,0.061732575,0.11317638,0.18176813,0.3806842,0.7956643,1.6221949,3.1860867,4.5613513,5.0449233,5.0243454,4.8905916,5.0346346,4.7774153,4.249259,3.8377085,3.508468,2.8019729,2.4967396,2.07833,1.8691251,1.7353712,1.0666018,1.1694894,1.5501735,1.7902447,1.8073926,1.8588364,1.6770682,1.3581166,1.2895249,1.4232788,1.2895249,0.9911508,0.75450927,0.5761707,0.4629943,0.4664239,0.6344737,0.7442205,0.72707254,0.64819205,0.7339317,1.4781522,1.1008976,0.7407909,0.70306545,0.4664239,0.19548649,0.12346515,0.08573969,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.037725464,0.006859175,0.0,0.0,0.0,0.0034295875,0.020577524,0.010288762,0.05144381,0.09945804,0.0,0.0274367,0.06516216,0.31895164,0.77851635,1.2243627,0.65848076,0.23664154,0.106317215,0.16119061,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.020577524,0.17490897,0.23664154,0.14747226,0.037725464,0.07888051,0.25721905,0.24350071,0.041155048,0.0,0.0034295875,0.0274367,0.058302987,0.07888051,0.1097468,0.30866286,0.45613512,0.38754338,0.15433143,0.041155048,0.09602845,0.15433143,0.26407823,0.34981793,0.22635277,0.06859175,0.017147938,0.006859175,0.0,0.0,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.030866288,0.06516216,0.1920569,0.53501564,0.9259886,0.69963586,0.29151493,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0034295875,0.01371835,0.01371835,0.07888051,0.15776102,0.20577525,0.23321195,0.30523327,0.29837412,0.2709374,0.31895164,0.47671264,0.7407909,0.6036074,0.44584638,0.45270553,0.6344737,0.83681935,0.8025235,0.5761707,0.42183927,0.4629943,0.6824879,0.9602845,1.2072148,1.2312219,1.0151579,0.70649505,0.6927767,0.78537554,0.9431366,1.0014396,0.66876954,0.45270553,0.32238123,0.22978236,0.14747226,0.10288762,0.16462019,0.15090185,0.14404267,0.15090185,0.10288762,0.13032432,0.17833854,0.20234565,0.25721905,0.4938606,2.1332035,4.712253,5.8234396,5.079219,4.1120753,3.1963756,2.7333813,4.197815,5.9914894,3.4467354,4.448175,5.2815647,5.751418,5.909179,6.0806584,6.375603,6.852316,6.358455,4.6676683,2.4761622,2.1674993,3.0557625,4.180667,4.6402316,3.6044965,2.7059445,2.8019729,3.5599117,4.7259717,6.121814,7.720001,9.033533,9.89093,10.045261,9.184435,8.347616,9.554831,11.173596,13.046151,16.489456,19.552078,22.096832,23.849352,25.042849,26.394106,24.44953,22.216867,21.04052,20.814167,19.9602,16.407146,14.510585,14.21564,15.933864,20.53637,23.242313,27.080023,31.044626,33.544796,32.41989,33.89461,33.14696,31.631084,28.359259,19.925903,20.982216,17.53548,12.47341,9.331907,12.284782,12.236768,10.1652975,8.841476,8.97523,9.1981535,8.951223,14.517444,20.2037,21.139977,13.293081,11.108434,12.411677,12.775213,10.984968,9.040393,7.9943686,6.060081,4.5270553,3.666229,2.7230926,1.903421,2.270387,2.9974594,3.6559403,4.232111,4.5784993,5.2747054,5.7651367,5.909179,5.9914894,4.5956473,4.9694724,5.23698,5.3741636,7.1952744,5.6005163,3.7759757,2.2498093,1.4232788,1.5913286,1.4129901,2.7162333,3.5770597,3.069481,1.2723769,1.3958421,1.2106444,0.9774324,0.89512235,1.1077567,1.2209331,1.0288762,0.75450927,0.66191036,1.0563129,0.85739684,0.89169276,0.9774324,1.1077567,1.4815818,0.9568549,0.5658819,0.45270553,0.5521636,0.5796003,0.5521636,0.4355576,0.33609957,0.2777966,0.22635277,0.16119061,0.14061308,0.18176813,0.24350071,0.2469303,0.12689474,0.06859175,0.072021335,0.11317638,0.15433143,0.12003556,0.19548649,0.78537554,2.0131679,3.7005248,3.2512488,2.177788,1.4781522,1.5124481,2.0028791,2.352697,2.7985435,2.8637056,2.4075704,1.6187652,1.6804979,2.16064,2.6407824,2.942586,3.117495,2.976882,2.1743584,1.5570327,1.3615463,1.2106444,0.82996017,0.47671264,0.29151493,0.33266997,0.5590228,0.77165717,1.0631721,0.97057325,0.48014224,0.024007112,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.006859175,0.072021335,0.14061308,0.072021335,0.01371835,0.020577524,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058302987,0.058302987,0.0,0.0,0.037725464,0.058302987,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07545093,0.082310095,0.06516216,0.07888051,0.19548649,0.37039545,0.36353627,0.31552204,0.31209245,0.3806842,0.31895164,0.216064,0.14747226,0.12689474,0.12346515,0.14061308,0.13032432,0.09945804,0.05144381,0.0,0.0,0.0,0.0034295875,0.0274367,0.08573969,0.017147938,0.0,0.0,0.006859175,0.024007112,0.044584636,0.020577524,0.14404267,0.6036074,1.5810398,2.452155,3.5564823,7.349606,13.831526,20.560377,19.102802,11.640019,5.7136927,3.8548563,3.6319332,4.540774,5.926327,6.1801167,4.979761,3.2889743,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.06859175,0.106317215,0.106317215,0.06859175,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.07545093,0.1371835,0.01371835,0.11317638,0.33952916,0.39440256,0.2194936,0.0,0.0,0.010288762,0.041155048,0.082310095,0.106317215,0.16804978,0.274367,1.5433143,3.0283258,1.7079345,1.8313997,8.453933,10.007536,4.6608095,0.29151493,1.3889829,3.5393343,3.1860867,0.7099246,0.42869842,0.32924038,0.18519773,0.082310095,0.05144381,0.07545093,0.1371835,0.26407823,0.37725464,0.40126175,0.22978236,0.32581082,0.45270553,0.5418748,0.59674823,0.65505123,0.6790583,0.8711152,1.2346514,1.7833855,2.503599,2.2841053,2.2360911,2.311542,2.201795,1.371835,0.72707254,0.59331864,0.548734,0.36696586,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15776102,0.31895164,0.48357183,0.70306545,1.0666018,1.8005334,2.294394,2.7162333,3.2032347,3.875434,4.3761535,4.5099077,4.57164,4.6402316,4.5784993,4.383013,4.029765,3.5564823,2.9151495,1.9994495,1.4850113,1.3478279,1.3478279,1.2826657,0.9774324,0.7579388,0.5555932,0.39097297,0.28808534,0.274367,0.28808534,0.28122616,0.31209245,0.39440256,0.5041494,0.5041494,0.36696586,0.23321195,0.15090185,0.09259886,0.041155048,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.0274367,0.01371835,0.01371835,0.030866288,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.044584636,0.034295876,0.01371835,0.0,0.024007112,0.048014224,0.08573969,0.1371835,0.19891608,0.19891608,0.23664154,0.37382504,0.6824879,1.2209331,2.3321195,4.2286816,4.6402316,3.5839188,3.3884325,3.998899,3.5564823,3.2855449,3.2786856,2.4727325,2.2635276,2.9185789,3.3198407,3.0557625,2.393852,1.8965619,1.3032433,1.1077567,1.5055889,2.3972816,2.1640697,1.704505,1.4781522,1.4472859,1.0666018,1.5810398,1.3512574,0.9602845,0.7099246,0.6241849,0.6756287,0.7407909,0.8711152,1.0014396,0.9774324,1.0494537,0.9945804,0.97057325,1.0151579,1.0528834,0.6756287,0.58988905,0.42526886,0.13375391,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.05144381,0.034295876,0.01371835,0.01371835,0.0,0.13375391,0.26064864,1.1146159,2.49331,3.2512488,1.7490896,0.6859175,0.3566771,0.4389872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09945804,0.106317215,0.024007112,0.061732575,0.26750782,0.58645946,0.53844523,0.15776102,0.0,0.01371835,0.06859175,0.06516216,0.048014224,0.24350071,0.36696586,0.22292319,0.08916927,0.09259886,0.21263443,0.48357183,0.4389872,0.39783216,0.3841138,0.15090185,0.041155048,0.006859175,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.01371835,0.01371835,0.05144381,0.15433143,0.34981793,0.4972902,0.34295875,0.13375391,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.14404267,0.18176813,0.17147937,0.24350071,0.30523327,0.23664154,0.22635277,0.31552204,0.4115505,0.34981793,0.35324752,0.4389872,0.5796003,0.70306545,0.5796003,0.44927597,0.45956472,0.64819205,0.91569984,1.3684053,1.8931323,1.9480057,1.4610043,0.84024894,0.7305021,0.66533995,0.7442205,0.864256,0.71678376,0.65505123,0.5693115,0.432128,0.274367,0.15090185,0.21263443,0.22978236,0.19891608,0.14061308,0.09259886,0.07888051,0.06859175,0.06859175,0.12689474,0.33609957,1.5433143,4.8940215,6.3035817,5.0757895,3.8925817,3.1346428,2.469303,3.683377,5.641671,4.2869844,1.821111,2.0097382,2.6647894,3.1860867,4.5784993,6.2487082,6.667118,6.327589,5.2472687,2.976882,2.4624438,2.884283,3.3781435,3.4467354,2.9460156,2.2120838,2.386993,3.3678548,5.0346346,7.233,8.625413,9.849775,10.569988,10.539123,9.613133,9.527394,10.367643,11.574858,13.008426,14.939283,18.722118,22.306036,24.61072,25.869379,27.60475,24.085993,21.53438,19.805868,18.557497,17.226818,18.44775,20.11796,19.329155,17.21653,18.934752,25.053137,31.442457,35.82547,37.58142,37.766617,35.82547,34.58739,33.465916,30.84914,24.123718,17.641798,12.55229,9.73317,9.760606,12.908967,15.54632,14.363112,12.343085,11.005547,10.405369,11.4205265,16.37971,19.044498,18.214539,17.700102,12.97413,10.933525,10.432805,10.834066,11.993267,9.3079,7.9600725,6.2487082,3.9680326,2.3801336,2.393852,2.836269,2.750529,2.486451,3.707384,3.7313912,3.1517909,3.3541365,4.513337,5.6005163,5.857735,6.23156,6.135532,5.353586,4.0606318,4.4859004,4.1635194,3.4776018,2.7128036,2.0303159,2.1160555,3.3541365,4.4584637,4.1292233,1.0528834,0.9294182,0.84367853,0.6790583,0.4972902,0.53501564,0.91227025,1.2895249,1.2312219,0.8128122,0.64133286,0.5796003,0.65505123,0.75450927,0.9911508,1.7250825,1.6016173,1.1146159,0.6927767,0.5693115,0.7613684,0.7133542,0.5727411,0.432128,0.34638834,0.33609957,0.2503599,0.18176813,0.15776102,0.17490897,0.19891608,0.1371835,0.08573969,0.072021335,0.106317215,0.16804978,0.1920569,0.20920484,0.37725464,0.85396725,1.7696671,1.5398848,1.3512574,1.2003556,1.2072148,1.6496316,1.879414,2.085189,2.2258022,2.194936,1.8142518,2.510458,2.8396983,3.1209247,3.5461934,4.180667,3.9131594,2.5001693,1.5398848,1.5536032,1.9685832,1.6256244,1.155771,0.7956643,0.70649505,0.9602845,1.2415106,1.3409687,1.1214751,0.6344737,0.12346515,0.17147937,0.072021335,0.0,0.0,0.0,0.0,0.037725464,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08573969,0.041155048,0.0,0.0,0.0,0.09602845,0.15776102,0.23664154,0.4046913,0.7476501,0.6859175,0.34295875,0.08573969,0.024007112,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.1097468,0.4081209,0.94656616,1.1523414,2.1229146,4.4756117,7.8777623,11.002116,9.280463,7.3221693,4.8185706,2.620205,2.7162333,3.5942078,5.65539,6.217842,5.1100855,4.6676683,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.020577524,0.037725464,0.041155048,0.030866288,0.01371835,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.0034295875,0.030866288,0.08573969,0.10288762,0.06516216,0.0,0.106317215,0.13032432,0.17490897,0.2469303,0.24007112,0.20577525,0.37382504,2.3664153,4.32128,0.90198153,1.2689474,4.4756117,6.680836,6.094377,2.976882,2.568761,2.7642474,1.9171394,0.32581082,0.23321195,0.13375391,0.058302987,0.017147938,0.010288762,0.01371835,0.0274367,0.05144381,0.07545093,0.07888051,0.044584636,0.06516216,0.08916927,0.1097468,0.15433143,0.31552204,0.22292319,0.19891608,0.2469303,0.53844523,1.4027013,1.2243627,0.94656616,0.82996017,0.7613684,0.274367,0.14404267,0.12003556,0.1097468,0.072021335,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.06516216,0.09602845,0.14061308,0.21263443,0.6036074,0.94656616,1.2517995,1.5810398,2.0577524,2.4487255,2.8499873,3.2135234,3.4981792,3.6627994,3.8479972,3.9508848,3.8171308,3.3884325,2.7059445,2.020027,1.6599203,1.4507155,1.214074,0.78194594,0.44584638,0.28808534,0.25721905,0.28122616,0.2503599,0.32924038,0.34981793,0.36010668,0.38754338,0.42869842,0.42869842,0.35324752,0.26064864,0.18519773,0.10288762,0.0548734,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.07545093,0.058302987,0.0,0.0034295875,0.01371835,0.020577524,0.0274367,0.0274367,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.12346515,0.19891608,0.106317215,0.020577524,0.0034295875,0.0,0.01371835,0.05144381,0.06516216,0.0548734,0.07545093,0.09602845,0.2777966,0.4938606,0.6310441,0.5727411,1.0220171,1.903421,2.287535,2.1846473,2.5584722,2.620205,2.510458,2.095478,1.5158776,1.1763484,1.3203912,1.4918705,1.5673214,1.6153357,1.8828435,1.6359133,1.1077567,0.7990939,0.94656616,1.5055889,1.821111,1.728512,1.4953002,1.2415106,0.97057325,1.1317638,1.1077567,1.0425946,0.9877212,0.89512235,1.3924125,1.4918705,1.5844694,1.7662375,1.8176813,2.1846473,1.6256244,1.2963841,1.2998136,0.66191036,0.35324752,0.7613684,1.3512574,1.4781522,0.36696586,0.10288762,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.0274367,0.030866288,0.06516216,0.17147937,0.58988905,1.1660597,1.7113642,1.8691251,1.1146159,0.5007198,0.16804978,0.072021335,0.08916927,0.0,0.0,0.0,0.0034295875,0.017147938,0.037725464,0.06516216,0.058302987,0.034295876,0.0548734,0.20920484,0.28808534,0.22978236,0.12689474,0.07888051,0.18176813,0.36010668,0.38754338,0.31895164,0.24007112,0.26750782,0.116605975,0.044584636,0.072021335,0.18176813,0.32238123,0.5624523,0.7099246,0.5212973,0.15433143,0.17833854,0.59331864,0.72021335,0.59674823,0.31895164,0.037725464,0.010288762,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.010288762,0.061732575,0.216064,0.29494452,0.18176813,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.01371835,0.030866288,0.05144381,0.09602845,0.16462019,0.25721905,0.25721905,0.22978236,0.20234565,0.20920484,0.2777966,0.32581082,0.37725464,0.42869842,0.47328308,0.50757897,0.4629943,0.432128,0.4355576,0.5212973,0.7682276,1.3169615,1.8245405,1.879414,1.4507155,0.8745448,0.65848076,0.64819205,0.8093826,0.9877212,0.89855194,0.65505123,0.52472687,0.41498008,0.29494452,0.20234565,0.24350071,0.28122616,0.25721905,0.1920569,0.20234565,0.14061308,0.08573969,0.05144381,0.07545093,0.21263443,1.0597426,3.5461934,5.6828265,6.420188,5.6348124,4.5682106,3.1655092,3.0454736,3.981751,3.8857226,1.8382589,1.3066728,1.3101025,1.6256244,2.784825,4.3109913,5.31929,5.7102633,5.4804807,4.7328305,3.7794054,2.760818,2.2086544,2.1126258,1.8965619,2.3629858,3.1689389,4.4275975,6.4304767,9.623423,11.05699,10.909517,10.045261,9.318189,9.551401,9.644,10.275044,11.787492,13.924125,15.854982,17.058767,18.488907,20.7833,23.300617,24.137436,22.419212,20.687271,19.456049,18.70497,17.87501,18.879879,21.270302,21.767591,20.172834,19.377169,24.885086,31.226395,35.033237,35.451645,34.141544,31.360147,29.919722,32.224403,34.878906,28.6885,19.246845,16.684942,15.9750185,14.932424,14.21564,12.857523,12.55915,12.545431,12.140739,10.762046,10.47396,13.197053,15.22051,15.069608,13.502286,11.382801,10.206452,9.47595,8.985519,8.80718,6.883182,5.871454,5.970912,5.9331865,3.07634,2.8739944,2.9700227,3.1860867,3.8137012,5.610805,4.3178506,3.0489032,3.0557625,4.280125,5.3673043,6.036074,6.210983,5.909179,5.219832,4.3281393,4.773986,4.396731,4.3487167,4.7842746,4.8734436,4.3041325,4.1360826,4.2081037,3.666229,0.9431366,0.52815646,0.4115505,0.33266997,0.21263443,0.18176813,0.30523327,0.52472687,0.6379033,0.61389613,0.5796003,0.64476246,0.65162164,0.6310441,0.7442205,1.2723769,1.4232788,1.4953002,1.3478279,1.0528834,0.89855194,0.66191036,0.5555932,0.45956472,0.36010668,0.34638834,0.41840968,0.4115505,0.3841138,0.34638834,0.2709374,0.17147937,0.116605975,0.09945804,0.11317638,0.14404267,0.18862732,0.20920484,0.24007112,0.33266997,0.52472687,0.4972902,0.47328308,0.5796003,0.8779744,1.3684053,1.6290541,1.7662375,1.8005334,1.7525192,1.6564908,2.0989075,2.393852,2.3081124,2.0440342,2.2395205,2.4315774,2.1057668,1.8897027,2.0646117,2.5653315,2.3218307,2.0817597,1.8725548,1.7593783,1.8416885,2.1812177,2.7882545,2.3801336,1.0323058,0.20920484,0.18862732,0.13032432,0.082310095,0.058302987,0.048014224,0.06859175,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.037725464,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.07545093,0.034295876,0.0,0.0034295875,0.01371835,0.020577524,0.030866288,0.1097468,0.24350071,0.33266997,0.18519773,0.072021335,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.01371835,0.061732575,0.20577525,0.5693115,1.255229,1.99602,3.350707,5.6039457,8.769455,8.628842,6.8385973,4.7808447,3.210094,2.2635276,2.7333813,3.2683969,3.5873485,3.666229,3.7553983,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.017147938,0.006859175,0.024007112,0.020577524,0.01371835,0.006859175,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.017147938,0.0274367,0.024007112,0.017147938,0.024007112,0.017147938,0.020577524,0.024007112,0.0,0.09602845,0.16804978,0.36010668,0.6344737,0.7613684,0.83681935,2.1126258,4.012617,4.5784993,0.48357183,1.5398848,3.4878905,5.209543,5.518206,3.1346428,2.177788,1.9685832,1.6153357,1.0048691,0.823101,0.4046913,0.12003556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09259886,0.041155048,0.01371835,0.0,0.08916927,0.45270553,0.3841138,0.2503599,0.18176813,0.16119061,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12346515,0.30523327,0.44584638,0.5693115,0.8162418,1.1008976,1.4472859,1.8039631,2.1297739,2.4075704,2.6819375,3.1552205,3.457024,3.4467354,3.2032347,2.49331,1.961724,1.5981878,1.3101025,0.89855194,0.44927597,0.20577525,0.116605975,0.12346515,0.16119061,0.25378948,0.3566771,0.45270553,0.5041494,0.47671264,0.36696586,0.26407823,0.19548649,0.15776102,0.12346515,0.09259886,0.06516216,0.044584636,0.034295876,0.0274367,0.020577524,0.034295876,0.030866288,0.010288762,0.010288762,0.010288762,0.0034295875,0.0,0.0034295875,0.010288762,0.082310095,0.16462019,0.14404267,0.0548734,0.0548734,0.030866288,0.017147938,0.01371835,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.017147938,0.07888051,0.15090185,0.07888051,0.024007112,0.037725464,0.082310095,0.10288762,0.106317215,0.07545093,0.030866288,0.037725464,0.082310095,0.216064,0.35324752,0.45270553,0.5212973,0.7373613,1.2380811,1.4438564,1.3478279,1.5090185,1.8588364,2.428148,2.9151495,2.8396983,1.5124481,1.2620882,1.08032,1.0563129,1.2209331,1.5433143,1.5090185,1.2175035,0.9328478,0.8128122,0.90541106,1.1180456,1.255229,1.2895249,1.1866373,0.9362774,0.9294182,1.0185875,1.0871792,1.1592005,1.3924125,1.862266,1.8691251,1.7765263,1.7799559,1.9102802,1.8965619,1.6324836,1.4678634,1.4027013,1.0940384,1.2346514,1.4850113,1.8862731,2.1434922,1.6016173,0.9431366,0.48700142,0.22635277,0.11317638,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.044584636,0.020577524,0.0,0.0,0.0,0.0274367,0.09259886,0.18519773,0.3018037,0.45270553,1.1729189,1.587899,1.6084765,1.2517995,0.64476246,0.28122616,0.082310095,0.006859175,0.0,0.0,0.05144381,0.041155048,0.0274367,0.030866288,0.0548734,0.048014224,0.07545093,0.14061308,0.20920484,0.20920484,0.14747226,0.058302987,0.034295876,0.10288762,0.22978236,0.4355576,0.4972902,0.39783216,0.216064,0.14747226,0.044584636,0.017147938,0.082310095,0.216064,0.37039545,0.5144381,0.47671264,0.29151493,0.10288762,0.17490897,0.45270553,0.53158605,0.40126175,0.16119061,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.08573969,0.34638834,0.45270553,0.2709374,0.082310095,0.006859175,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.006859175,0.010288762,0.017147938,0.048014224,0.116605975,0.22292319,0.23321195,0.19891608,0.15090185,0.14404267,0.26407823,0.45956472,0.6379033,0.67219913,0.58302987,0.5212973,0.39440256,0.33609957,0.31895164,0.35324752,0.5041494,0.8779744,1.3032433,1.4095604,1.1420527,0.7476501,0.5624523,0.53158605,0.6173257,0.7442205,0.77165717,0.61046654,0.50757897,0.42183927,0.33609957,0.2503599,0.3018037,0.31209245,0.33952916,0.4046913,0.5041494,0.24007112,0.106317215,0.058302987,0.07545093,0.1371835,0.5658819,1.8691251,3.549623,4.938606,5.223262,4.602506,3.6353626,2.784825,2.3218307,2.3389788,1.4507155,1.2963841,1.3203912,1.4541451,2.1160555,2.9288676,3.974892,4.523626,4.496189,4.4584637,3.1483612,2.8054025,2.4247184,1.903421,2.0646117,2.5378947,3.6044965,4.629943,5.826869,8.22758,9.8429165,10.456812,10.31277,9.856634,9.729739,9.619993,9.901219,10.909517,12.456262,13.810948,14.13333,15.354263,17.161655,18.945042,19.78186,19.565796,19.353163,19.089085,18.965618,19.435472,20.35803,23.214878,24.94339,24.562706,23.1943,28.558174,35.66085,38.541702,36.09298,32.035778,29.806545,29.43615,30.444448,30.75654,26.709627,20.635828,19.562366,19.589804,18.358582,15.018164,11.1393,10.38479,10.38479,10.504827,11.828648,12.103014,12.0138445,11.712041,11.489118,11.736049,12.109874,11.14273,10.034973,9.253027,8.505377,6.574519,5.353586,5.6348124,6.5779486,5.7411294,5.212973,4.962613,4.976331,5.130663,5.192395,3.018037,2.170929,3.4535947,6.307011,8.80718,6.375603,5.164959,4.619654,4.307562,3.9097297,4.0674906,3.9680326,4.0023284,4.3349986,4.880303,5.223262,4.938606,4.506478,3.7485392,1.8313997,0.69963586,0.31552204,0.216064,0.15090185,0.09945804,0.12346515,0.21263443,0.31895164,0.38754338,0.3806842,0.3841138,0.36353627,0.36010668,0.45613512,0.78537554,1.0323058,1.2346514,1.2346514,1.0460242,0.84024894,0.70649505,0.6824879,0.6790583,0.61046654,0.42526886,0.61389613,0.66191036,0.5624523,0.3806842,0.22635277,0.13032432,0.07888051,0.06516216,0.072021335,0.082310095,0.116605975,0.13375391,0.14061308,0.14404267,0.14061308,0.14404267,0.1920569,0.39097297,0.72364295,1.039165,1.1934965,1.2449403,1.2826657,1.3341095,1.3992717,1.7250825,2.1263442,2.2326615,2.0886188,2.1297739,2.2223728,2.3424082,2.3561265,2.287535,2.3149714,2.4898806,2.4315774,2.3458378,2.3904223,2.6819375,3.1963756,3.3678548,2.633923,1.2792361,0.4115505,0.3018037,0.23321195,0.16462019,0.09602845,0.061732575,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.030866288,0.01371835,0.0,0.006859175,0.041155048,0.037725464,0.01371835,0.030866288,0.082310095,0.09259886,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.024007112,0.058302987,0.037725464,0.05144381,0.0548734,0.041155048,0.030866288,0.082310095,0.13375391,0.08916927,0.041155048,0.061732575,0.18862732,0.548734,1.0185875,1.8519772,3.5770597,6.999788,7.599966,6.1801167,4.0434837,2.2463799,1.6016173,1.821111,2.0131679,2.218943,2.5001693,2.9494452,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.017147938,0.0274367,0.0274367,0.024007112,0.024007112,0.020577524,0.030866288,0.041155048,0.006859175,0.05144381,0.14404267,0.33952916,0.58988905,0.7476501,1.0700313,3.4467354,4.7671266,3.6696587,0.53158605,2.3801336,3.8205605,4.2595477,3.566771,2.095478,1.4164196,1.1351935,1.1317638,1.1934965,1.0082988,0.53844523,0.16804978,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.09259886,0.106317215,0.19891608,0.31895164,0.47328308,0.6790583,0.9328478,1.2346514,1.4850113,1.9068506,2.2600982,2.4418662,2.503599,2.1915064,1.8073926,1.5364552,1.3889829,1.1900668,0.75450927,0.40126175,0.16119061,0.048014224,0.06516216,0.116605975,0.20920484,0.32924038,0.41498008,0.37382504,0.2777966,0.19548649,0.14061308,0.116605975,0.13032432,0.11317638,0.082310095,0.06859175,0.07888051,0.07545093,0.041155048,0.041155048,0.034295876,0.017147938,0.020577524,0.020577524,0.01371835,0.006859175,0.006859175,0.010288762,0.072021335,0.1371835,0.12689474,0.06859175,0.06859175,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0034295875,0.017147938,0.0548734,0.041155048,0.048014224,0.1097468,0.22292319,0.13375391,0.08916927,0.05144381,0.017147938,0.017147938,0.0548734,0.10288762,0.16804978,0.28122616,0.48357183,0.53501564,0.7407909,0.7956643,0.6824879,0.6790583,1.3272504,1.9651536,2.8705647,3.7965534,3.9783216,3.059192,2.0097382,1.3924125,1.2620882,1.1660597,1.4164196,1.4232788,1.3066728,1.1111864,0.7956643,1.0220171,1.2346514,1.313532,1.2243627,1.0151579,0.881404,0.9602845,1.0940384,1.2415106,1.5090185,1.8897027,1.9582944,1.8245405,1.728512,2.0577524,1.8862731,2.0268862,2.0817597,2.0920484,2.5653315,2.901431,2.4555845,2.253239,2.585909,3.0043187,2.7368107,2.177788,1.6187652,1.1146159,0.4972902,0.20234565,0.06859175,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.010288762,0.044584636,0.020577524,0.0,0.0034295875,0.01371835,0.09259886,0.2503599,0.4046913,0.59331864,1.0082988,1.7593783,2.0097382,1.7971039,1.2792361,0.7305021,0.2709374,0.072021335,0.01371835,0.034295876,0.116605975,0.12689474,0.07888051,0.0548734,0.06859175,0.072021335,0.07545093,0.19891608,0.29151493,0.28808534,0.18862732,0.07545093,0.024007112,0.037725464,0.09259886,0.16119061,0.33266997,0.3841138,0.29151493,0.13032432,0.07888051,0.058302987,0.05144381,0.116605975,0.24350071,0.34638834,0.35324752,0.216064,0.12003556,0.11317638,0.13032432,0.18862732,0.18862732,0.1097468,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.08916927,0.31895164,0.39783216,0.24350071,0.07545093,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.061732575,0.13032432,0.15433143,0.13375391,0.09602845,0.08916927,0.19548649,0.41840968,0.6344737,0.69963586,0.61389613,0.4972902,0.33266997,0.24350071,0.20920484,0.22292319,0.30866286,0.5041494,0.8025235,0.9602845,0.90541106,0.7339317,0.53844523,0.42869842,0.42183927,0.4972902,0.6001778,0.5418748,0.48014224,0.42183927,0.36010668,0.24350071,0.37725464,0.32238123,0.32581082,0.4629943,0.6379033,0.32924038,0.14747226,0.082310095,0.08916927,0.09602845,0.21263443,0.64476246,1.5021594,2.6990852,3.9646032,4.033195,3.9268777,3.2821152,2.270387,1.5913286,1.3409687,1.3684053,1.4232788,1.5055889,1.8691251,2.277246,2.9734523,3.4124396,3.5873485,4.0434837,3.3472774,3.5290456,3.216953,2.4967396,2.942586,2.8945718,3.5530527,4.331569,5.1821065,6.6053853,7.5107965,8.886061,10.556271,11.832077,11.478829,10.933525,10.635151,10.871792,11.516555,12.017275,12.274493,13.642899,14.946142,15.717799,16.194511,17.37772,18.248835,18.499195,18.855871,21.061096,23.101702,25.080574,27.076593,28.6885,29.034887,33.77115,40.541153,41.100178,34.892624,29.031458,28.51702,28.136335,27.285797,25.59844,22.94394,19.61724,18.975908,18.941612,17.861292,14.479718,11.499407,10.367643,9.692014,9.6817255,12.133881,12.850664,11.077567,9.146709,8.625413,10.316199,11.489118,10.830637,9.863494,9.259886,8.834618,7.5725293,6.3961806,6.1629686,6.8283086,7.438775,7.8023114,7.390761,6.5813785,5.669108,4.8734436,3.8274195,4.331569,6.759717,10.010965,11.537132,6.866034,4.6916757,4.0503426,3.9371665,3.309552,2.9220085,2.9288676,2.9700227,3.2512488,4.557922,5.439326,5.0312047,4.122364,3.093488,1.9102802,0.6893471,0.29494452,0.22292319,0.1920569,0.14404267,0.12346515,0.13032432,0.16462019,0.19891608,0.18519773,0.15090185,0.13375391,0.15090185,0.216064,0.37039545,0.548734,0.72021335,0.8196714,0.8162418,0.7099246,0.61046654,0.5727411,0.5624523,0.5178677,0.31552204,0.45613512,0.5007198,0.41498008,0.2503599,0.12346515,0.06516216,0.034295876,0.030866288,0.041155048,0.041155048,0.0548734,0.06859175,0.08573969,0.10288762,0.1097468,0.09602845,0.20234565,0.4081209,0.66191036,0.85739684,0.9568549,1.0254467,1.097468,1.1763484,1.2517995,1.4850113,1.8519772,2.1126258,2.177788,2.0920484,2.2395205,2.585909,2.7573884,2.6545007,2.4487255,2.6613598,2.4247184,2.3561265,2.7333813,3.4707425,4.07435,3.2855449,2.1812177,1.3546871,0.91227025,0.52472687,0.26407823,0.12346515,0.06516216,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.037725464,0.01371835,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.006859175,0.010288762,0.006859175,0.0548734,0.1371835,0.18176813,0.2503599,0.20577525,0.116605975,0.05144381,0.09602845,0.1371835,0.07888051,0.020577524,0.0,0.0,0.08573969,0.3806842,0.91569984,2.2086544,5.2781353,6.492209,5.0003386,2.8705647,1.4164196,1.1797781,1.4198492,1.5193073,1.5193073,1.605047,2.1126258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.010288762,0.010288762,0.006859175,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0274367,0.05144381,0.058302987,0.01371835,0.030866288,0.12346515,0.16804978,0.16119061,0.20920484,0.823101,4.149801,4.7191124,2.1091962,0.97057325,3.789694,4.3521466,3.4638834,2.277246,2.2669573,1.4953002,0.66876954,0.3806842,0.5693115,0.5178677,0.33952916,0.116605975,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.010288762,0.0,0.048014224,0.17833854,0.40126175,0.59331864,0.6859175,0.75450927,0.84024894,0.94656616,1.1694894,1.1420527,1.138623,1.2655178,1.4507155,1.2415106,0.88826317,0.51100856,0.20577525,0.037725464,0.006859175,0.0,0.0548734,0.13032432,0.12346515,0.15090185,0.14404267,0.106317215,0.06859175,0.09602845,0.08916927,0.0548734,0.058302987,0.09259886,0.106317215,0.044584636,0.010288762,0.0034295875,0.01371835,0.024007112,0.0274367,0.017147938,0.01371835,0.01371835,0.0034295875,0.010288762,0.020577524,0.024007112,0.0274367,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0034295875,0.0,0.0,0.024007112,0.06859175,0.14747226,0.28122616,0.07545093,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0548734,0.15776102,0.25721905,0.15090185,0.06516216,0.06516216,0.14061308,0.22292319,0.77851635,1.0082988,1.5604624,3.0146074,5.888602,4.636802,2.9391565,1.8039631,1.430138,1.2346514,1.6736387,1.6907866,1.7902447,1.9137098,1.4369972,1.5227368,1.6324836,1.5055889,1.196926,1.0837497,0.91569984,0.94999576,1.0940384,1.2346514,1.214074,1.546744,1.9754424,2.2155135,2.287535,2.49331,2.6887965,3.0866287,3.1620796,3.1895163,4.2183924,4.3692946,3.433017,2.8088322,3.0866287,4.057202,4.5647807,4.266407,3.673088,2.8637056,1.488441,0.864256,0.53158605,0.3018037,0.11317638,0.044584636,0.0274367,0.01371835,0.0034295875,0.0,0.0034295875,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.06516216,0.12689474,0.10288762,0.21263443,0.39097297,0.548734,0.7956643,1.4369972,1.9823016,2.2600982,2.1332035,1.5673214,0.65162164,0.17490897,0.11317638,0.1371835,0.14061308,0.26064864,0.16804978,0.09602845,0.09602845,0.14404267,0.14061308,0.16804978,0.32924038,0.36696586,0.26750782,0.23321195,0.14061308,0.06516216,0.030866288,0.030866288,0.05144381,0.1920569,0.22635277,0.21263443,0.22978236,0.36010668,0.23664154,0.13375391,0.14404267,0.22978236,0.24007112,0.16119061,0.106317215,0.09602845,0.09945804,0.061732575,0.061732575,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.041155048,0.08916927,0.08916927,0.058302987,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.006859175,0.017147938,0.0274367,0.048014224,0.05144381,0.044584636,0.041155048,0.06516216,0.17490897,0.31209245,0.4115505,0.432128,0.33609957,0.24007112,0.17490897,0.14061308,0.14747226,0.2194936,0.32581082,0.490431,0.65505123,0.764798,0.7888051,0.5761707,0.41498008,0.37039545,0.432128,0.4972902,0.44927597,0.40126175,0.36010668,0.30523327,0.1920569,0.3841138,0.28122616,0.216064,0.31552204,0.52472687,0.34295875,0.17490897,0.09259886,0.09259886,0.072021335,0.061732575,0.12346515,0.34638834,1.0220171,2.6476414,3.4467354,4.091498,4.232111,3.673088,2.386993,2.0303159,1.7593783,1.6221949,1.6736387,1.9514352,2.3492675,2.5001693,2.6990852,3.210094,4.2698364,4.7534084,4.3624353,3.5393343,2.976882,3.6353626,3.2649672,3.223812,3.8720043,5.051782,6.0978065,6.094377,7.8331776,11.026124,14.068168,14.05102,12.994707,12.113303,11.88352,12.103014,11.89038,12.123591,13.306799,14.308239,14.55174,14.023583,15.868701,17.21653,17.761833,18.468328,21.585823,25.114868,26.095732,28.218645,32.306713,36.33648,39.48141,42.95901,39.75235,30.790836,24.963966,25.800787,24.6896,23.482386,22.347193,19.761284,16.904436,15.964729,15.422854,14.393978,12.644889,12.531713,11.821788,11.067279,10.909517,12.061859,11.862943,9.8429165,7.81603,7.0615206,8.320179,8.855195,8.834618,8.615124,8.567109,9.06097,9.139851,8.361334,7.6445503,7.3873315,7.459353,8.831187,8.371623,7.0203657,5.785714,5.7274113,6.725421,8.357904,10.484249,11.866373,10.192734,6.1286726,4.2286816,3.724532,3.57363,2.4761622,1.7559488,1.6907866,1.8005334,2.287535,4.0709205,4.5442033,3.806842,2.6304936,1.5673214,0.9294182,0.37382504,0.25721905,0.26407823,0.24350071,0.1920569,0.15090185,0.13375391,0.12003556,0.106317215,0.09602845,0.09259886,0.09259886,0.09259886,0.09602845,0.12346515,0.15776102,0.26064864,0.40126175,0.5178677,0.52815646,0.36353627,0.2469303,0.17833854,0.14061308,0.07545093,0.06516216,0.06859175,0.06516216,0.048014224,0.0274367,0.017147938,0.01371835,0.020577524,0.0274367,0.0274367,0.034295876,0.058302987,0.09602845,0.13375391,0.15433143,0.15433143,0.32581082,0.52815646,0.7133542,0.9534253,1.1317638,1.2209331,1.2895249,1.3684053,1.4781522,1.5364552,1.762808,2.1434922,2.4795918,2.369845,2.4315774,2.836269,3.1449318,3.1655092,2.942586,2.8465576,2.352697,2.4007113,3.2272418,4.389872,5.0003386,3.0660512,1.5193073,1.2998136,1.3649758,0.6344737,0.18176813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.024007112,0.06516216,0.16462019,0.3018037,0.4115505,0.32238123,0.18176813,0.07545093,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.09945804,0.34981793,0.6824879,1.4438564,3.391862,5.562791,4.2218223,2.3904223,1.4404267,1.0666018,1.3992717,1.2723769,1.0117283,0.91227025,1.2483698,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.058302987,0.0274367,0.01371835,0.0274367,0.01371835,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.0274367,0.01371835,0.09945804,0.22292319,0.20577525,0.07545093,0.07545093,0.9431366,5.826869,5.7377,1.0563129,1.5570327,6.036074,4.4927597,3.4535947,5.0757895,7.1266828,3.6113555,1.3855534,0.31209245,0.041155048,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072021335,0.16462019,0.2194936,0.22635277,0.21263443,0.2503599,0.28808534,0.42183927,0.75450927,1.3889829,1.7182233,1.6084765,1.2106444,0.6824879,0.18176813,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.044584636,0.020577524,0.006859175,0.0,0.0,0.0,0.01371835,0.006859175,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.09945804,0.65162164,1.0666018,1.2037852,1.3752645,0.8745448,0.85739684,1.1249046,1.7250825,2.9460156,2.9940298,2.1743584,2.3252604,3.340418,3.1586502,1.6324836,1.4438564,1.2895249,0.864256,0.84024894,0.9842916,1.1317638,1.1763484,1.1180456,1.0666018,1.1660597,2.253239,3.5393343,4.105216,2.884283,3.666229,4.355576,4.184097,3.5702004,4.1189346,4.0949273,4.245829,4.0503426,3.765687,4.4241676,4.3624353,4.3487167,4.4584637,4.2835546,2.9288676,2.393852,1.9651536,1.3238207,0.5693115,0.22978236,0.13032432,0.061732575,0.017147938,0.0034295875,0.01371835,0.0274367,0.020577524,0.010288762,0.0,0.0,0.024007112,0.07545093,0.33266997,0.6173257,0.39783216,0.34638834,0.25378948,0.4115505,0.7407909,0.77851635,1.255229,1.5021594,1.2998136,0.7099246,0.07545093,0.2469303,0.53844523,0.59674823,0.3806842,0.1371835,0.07545093,0.09602845,0.17147937,0.26407823,0.33609957,0.23664154,0.24007112,0.26407823,0.29151493,0.36696586,0.25721905,0.1097468,0.024007112,0.01371835,0.01371835,0.18519773,0.40126175,0.6036074,0.86082643,1.371835,0.8128122,0.34295875,0.09259886,0.044584636,0.044584636,0.082310095,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.082310095,0.072021335,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0034295875,0.01371835,0.041155048,0.06516216,0.07545093,0.07888051,0.09259886,0.10288762,0.08916927,0.082310095,0.09602845,0.12346515,0.15776102,0.24007112,0.32581082,0.4081209,0.5178677,0.53158605,0.50757897,0.51100856,0.5212973,0.4115505,0.31552204,0.22635277,0.14061308,0.09602845,0.16804978,0.14404267,0.12689474,0.13375391,0.19548649,0.36696586,0.19548649,0.07888051,0.041155048,0.061732575,0.061732575,0.048014224,0.044584636,0.11317638,0.47328308,1.5090185,3.2203827,4.187526,4.6127954,4.619654,4.2423997,3.875434,3.5633414,3.234101,2.9391565,2.8534167,2.9871707,2.5824795,2.3801336,2.976882,4.804852,5.31929,3.6627994,2.0989075,1.8039631,2.8534167,3.1586502,3.1620796,3.5599117,4.547633,5.830299,7.133542,10.189304,13.015285,14.538021,14.586036,13.1593275,12.205902,12.425395,13.293081,13.059869,12.620882,13.481709,14.387119,14.400838,12.922686,13.21763,15.241087,17.19938,18.46147,19.54522,22.196291,25.6053,30.231813,36.60399,45.332287,45.918747,41.288803,33.81573,26.294647,21.911634,20.923914,21.428062,21.321745,19.761284,17.134218,16.13621,14.839825,13.46799,12.044711,10.422516,10.299051,10.844356,11.897239,13.087306,13.855534,10.912948,8.961512,7.689135,6.8043017,6.012067,6.5367937,7.181556,7.8537555,8.669997,9.962952,10.597425,9.9869585,9.318189,8.7283,7.3255987,6.276145,5.545643,5.874883,6.9620624,7.4627824,7.6685576,8.076678,7.442205,5.394741,2.4418662,1.4027013,1.0528834,0.91912943,0.8025235,0.77851635,0.84024894,1.0014396,1.0734608,1.08032,1.2517995,1.1797781,0.7922347,0.41498008,0.20920484,0.18176813,0.24350071,0.26064864,0.25378948,0.22978236,0.16804978,0.15433143,0.15090185,0.16462019,0.17833854,0.16804978,0.15433143,0.15090185,0.15090185,0.14747226,0.12346515,0.09602845,0.09945804,0.14404267,0.19891608,0.19891608,0.15090185,0.12689474,0.16462019,0.19891608,0.07545093,0.07545093,0.058302987,0.041155048,0.0274367,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.05144381,0.13375391,0.2194936,0.26407823,0.22978236,0.26407823,0.5212973,0.764798,0.9877212,1.4027013,1.7593783,1.5638919,1.5090185,1.8416885,2.3801336,2.0989075,2.4247184,3.4981792,4.8117113,5.2026844,3.7519686,3.7176728,3.7965534,3.3678548,2.503599,2.5138876,2.5893385,3.3061223,4.6093655,5.844017,6.5882373,3.532475,1.3375391,1.2037852,0.90198153,0.17833854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.034295876,0.044584636,0.044584636,0.044584636,0.058302987,0.09602845,0.14747226,0.16462019,0.09259886,0.017147938,0.0,0.0,0.0,0.0,0.01371835,0.26407823,0.50757897,0.764798,1.3272504,5.0620713,6.0497923,4.5990767,2.07833,0.9294182,0.9431366,0.58988905,0.3018037,0.28465575,0.5041494,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.017147938,0.048014224,0.082310095,0.08916927,0.1097468,0.12003556,0.08916927,0.1371835,0.53844523,0.1097468,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.010288762,0.006859175,0.0034295875,0.006859175,0.01371835,0.1097468,0.41840968,0.39440256,0.116605975,0.2709374,2.5550427,8.519095,7.641121,1.0425946,1.4815818,3.590778,3.4604537,3.5839188,4.5956473,5.2575574,2.5824795,0.9328478,0.2469303,0.15433143,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.034295876,0.044584636,0.044584636,0.041155048,0.05144381,0.058302987,0.08573969,0.19548649,0.51100856,0.82996017,1.1111864,1.2586586,1.1489118,0.65848076,0.2777966,0.072021335,0.0,0.0,0.0,0.0,0.0,0.024007112,0.048014224,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.048014224,0.09945804,0.01371835,0.0034295875,0.0,0.0,0.006859175,0.0274367,0.024007112,0.024007112,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.072021335,0.13032432,0.024007112,0.01371835,0.0034295875,0.017147938,0.037725464,0.024007112,0.024007112,0.048014224,0.041155048,0.0034295875,0.0,0.010288762,0.034295876,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0034295875,0.31209245,0.5624523,0.607037,0.48014224,0.39783216,0.2469303,0.23321195,0.4389872,0.864256,1.430138,2.1434922,2.668219,3.3438478,3.7691166,2.8054025,2.194936,1.5981878,1.2175035,1.1626302,1.4507155,1.7147937,1.8588364,2.054323,2.5001693,3.4467354,3.74168,3.6525106,3.642222,3.683377,3.2615378,3.4467354,3.6147852,3.8445675,4.016047,3.8137012,4.4721823,4.6265135,4.3624353,4.040054,4.290414,4.3178506,4.2286816,4.554492,5.2472687,5.689686,5.0243454,4.9591837,4.880303,4.461893,3.6696587,3.1243541,1.7696671,0.83338976,0.6344737,0.58988905,0.26750782,0.15776102,0.1371835,0.14404267,0.18176813,0.20920484,0.22978236,0.4046913,0.6173257,0.50757897,0.36010668,0.2469303,0.805953,1.5981878,1.1077567,1.2826657,1.2998136,1.0151579,0.5727411,0.4046913,0.4389872,0.36010668,0.23321195,0.13375391,0.11317638,0.14061308,0.14747226,0.14061308,0.1371835,0.15090185,0.12346515,0.11317638,0.12346515,0.1371835,0.12346515,0.072021335,0.0274367,0.06516216,0.19548649,0.3806842,0.65162164,0.71678376,0.65162164,0.64476246,0.9842916,0.99801,0.6276145,0.2709374,0.10288762,0.082310095,0.061732575,0.037725464,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.0548734,0.072021335,0.037725464,0.017147938,0.0034295875,0.0,0.0,0.0034295875,0.0,0.006859175,0.006859175,0.006859175,0.01371835,0.034295876,0.048014224,0.0548734,0.058302987,0.05144381,0.058302987,0.061732575,0.07545093,0.09259886,0.10288762,0.08573969,0.08573969,0.09945804,0.11317638,0.09602845,0.09602845,0.14747226,0.20234565,0.23664154,0.2503599,0.2709374,0.36010668,0.5418748,0.7373613,0.75450927,0.42183927,0.25378948,0.17833854,0.14747226,0.14404267,0.07888051,0.08573969,0.1097468,0.14747226,0.23321195,0.12003556,0.041155048,0.05144381,0.1097468,0.061732575,0.037725464,0.0548734,0.14061308,0.548734,1.7422304,2.8054025,3.0420442,3.3609958,4.1189346,5.096367,4.417309,4.180667,4.214963,4.266407,4.0263357,3.2718265,2.644212,2.428148,2.627064,2.9631636,2.3732746,1.6187652,1.2346514,1.4918705,2.4144297,3.391862,4.5613513,6.0566516,7.829748,9.637141,12.037852,13.498857,15.114192,17.086205,18.739265,16.410576,13.900118,13.21763,14.147048,14.256795,13.63261,15.494876,17.487467,18.169954,17.024471,16.108772,16.80155,17.754974,18.396307,18.934752,20.052797,21.839613,24.957108,29.569902,35.34876,35.708866,33.06465,29.539038,26.52443,24.669024,24.120289,24.096281,22.95423,20.508932,18.04992,16.46545,14.562028,13.039291,11.835506,10.151579,9.054111,8.97523,10.371073,11.941824,10.621432,9.746887,9.527394,9.201583,8.621983,8.258447,8.862054,10.028113,10.871792,11.598865,13.516005,15.107333,14.538021,13.2862215,11.900668,9.997248,8.556821,7.613684,6.927767,6.3618846,5.874883,5.994919,4.938606,3.5016088,2.2258022,1.3924125,1.1729189,1.0871792,1.1077567,1.2449403,1.5227368,1.7593783,1.6427724,1.4472859,1.3443983,1.3992717,0.805953,0.44584638,0.28465575,0.2469303,0.23321195,0.26407823,0.2709374,0.26407823,0.2469303,0.216064,0.19548649,0.17490897,0.18519773,0.22292319,0.22978236,0.23664154,0.23664154,0.22978236,0.19891608,0.14747226,0.10288762,0.12346515,0.1371835,0.13032432,0.15090185,0.16804978,0.2469303,0.3018037,0.29494452,0.22292319,0.13375391,0.07888051,0.048014224,0.030866288,0.0274367,0.017147938,0.14747226,0.42869842,0.6893471,0.5521636,0.37382504,0.30866286,0.41840968,0.70649505,1.1214751,1.3238207,1.2620882,1.6221949,2.3252604,2.5138876,2.469303,2.1126258,2.0303159,2.3149714,2.5893385,2.551613,2.4727325,2.9563043,3.8445675,4.214963,4.029765,3.765687,3.3781435,2.9254382,2.5756202,2.352697,2.7093742,4.173808,5.8062916,5.1855364,3.6147852,2.9494452,3.093488,3.0626216,0.94999576,0.18862732,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.024007112,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.010288762,0.020577524,0.01371835,0.020577524,0.030866288,0.034295876,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.1097468,0.274367,0.5007198,0.77851635,2.170929,2.7916842,2.3424082,1.2860953,0.8711152,0.75450927,0.5658819,0.53501564,0.8265306,1.5638919,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.041155048,0.09945804,0.09259886,0.26064864,0.4081209,0.4389872,0.37382504,0.16462019,0.05144381,0.024007112,0.037725464,0.041155048,0.05144381,0.058302987,0.044584636,0.06859175,0.26750782,0.0548734,0.0034295875,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.01371835,0.010288762,0.010288762,0.024007112,0.07888051,0.2194936,0.29494452,0.2709374,0.35324752,0.980862,4.8254294,8.378482,6.6293926,1.5158776,1.9137098,2.452155,2.7402403,2.8980014,2.9151495,2.6407824,1.2723769,0.61389613,0.32581082,0.16804978,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.116605975,0.24350071,0.4389872,0.7407909,1.0254467,1.0082988,0.6927767,0.39783216,0.1920569,0.072021335,0.0,0.0,0.0,0.034295876,0.08573969,0.082310095,0.05144381,0.017147938,0.0,0.0,0.0,0.0,0.020577524,0.061732575,0.08573969,0.041155048,0.024007112,0.01371835,0.006859175,0.0034295875,0.01371835,0.020577524,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058302987,0.2709374,0.45613512,0.17833854,0.048014224,0.006859175,0.006859175,0.017147938,0.01371835,0.01371835,0.024007112,0.020577524,0.01371835,0.0274367,0.06859175,0.048014224,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14747226,0.216064,0.19548649,0.12689474,0.09602845,0.13032432,0.18519773,0.28465575,0.42869842,0.5761707,0.89855194,1.2072148,1.7388009,2.3252604,2.3972816,2.352697,1.6942163,1.3615463,1.5330256,1.6221949,1.5981878,1.670209,1.862266,2.3046827,3.2272418,3.7382503,3.7725463,3.8479972,4.1189346,4.389872,4.8837323,5.038064,5.130663,5.2781353,5.4496145,5.6073756,5.754848,5.5319247,5.055212,4.9077396,4.8254294,4.822,5.1238036,5.672538,6.138962,6.046363,6.310441,6.39961,6.159539,5.813151,5.658819,5.0449233,4.2115335,3.1655092,1.6736387,0.922559,0.6344737,0.53158605,0.4664239,0.44927597,0.52472687,0.6241849,0.6173257,0.5144381,0.4424168,0.28465575,0.45956472,1.2106444,1.9925903,1.4747226,1.0940384,0.83338976,0.6344737,0.5144381,0.5521636,0.4046913,0.38754338,0.30523327,0.16119061,0.15090185,0.1371835,0.13375391,0.106317215,0.058302987,0.05144381,0.041155048,0.044584636,0.0548734,0.0548734,0.024007112,0.017147938,0.09945804,0.33266997,0.6241849,0.7373613,0.5624523,0.42526886,0.31209245,0.2777966,0.41840968,0.4972902,0.34981793,0.16804978,0.061732575,0.082310095,0.061732575,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.034295876,0.041155048,0.0548734,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.017147938,0.034295876,0.06516216,0.09259886,0.08916927,0.082310095,0.07545093,0.07545093,0.08916927,0.116605975,0.09259886,0.08916927,0.1097468,0.14061308,0.14747226,0.14747226,0.17490897,0.18176813,0.16804978,0.15433143,0.16462019,0.24007112,0.38754338,0.6241849,0.9568549,0.64133286,0.38754338,0.2194936,0.13032432,0.082310095,0.05144381,0.06859175,0.09945804,0.12003556,0.106317215,0.061732575,0.037725464,0.05144381,0.082310095,0.041155048,0.034295876,0.058302987,0.2194936,0.7990939,2.2566686,3.3369887,3.690236,3.9371665,4.32471,4.7431192,4.712253,5.442755,6.478491,6.989499,5.7925735,4.016047,2.7951138,2.2155135,2.0817597,1.8965619,1.3101025,1.0117283,1.2929544,2.4624438,4.8494368,7.870903,10.556271,12.624311,13.759505,13.629181,13.598314,13.526293,14.616901,16.667795,18.04649,15.9921665,14.229359,13.900118,14.767803,15.189643,15.755525,17.720678,19.102802,19.089085,18.03277,18.554068,18.821575,18.818146,19.222837,21.421204,22.035099,22.889067,24.85422,28.0163,31.689388,33.702557,31.483612,28.338682,26.229485,25.807646,24.394655,23.238884,21.626978,19.36688,16.798119,13.927555,11.893809,10.882081,10.497967,9.736599,8.203573,7.675417,8.176137,8.97523,8.567109,10.151579,11.0981455,10.696883,9.582268,9.736599,10.422516,11.784062,12.775213,13.509145,15.247946,17.274832,16.61292,16.005884,15.412566,12.003556,9.80519,9.318189,8.669997,7.3290286,6.090947,5.662249,4.5784993,3.6936657,3.1209247,2.2463799,1.529596,1.0700313,0.9328478,1.0700313,1.3066728,1.587899,1.7353712,1.6907866,1.4541451,1.1043272,0.5453044,0.30866286,0.24350071,0.24007112,0.24350071,0.26064864,0.2709374,0.26407823,0.24350071,0.2194936,0.20234565,0.19548649,0.216064,0.2469303,0.25378948,0.26407823,0.26750782,0.26064864,0.23321195,0.17147937,0.13032432,0.15090185,0.15776102,0.1371835,0.14747226,0.2503599,0.38754338,0.4389872,0.36353627,0.22292319,0.12689474,0.072021335,0.058302987,0.072021335,0.08573969,0.2777966,0.5178677,0.72364295,0.83681935,0.83338976,1.2380811,1.3101025,1.1694894,1.0768905,1.4335675,1.5981878,1.7765263,2.085189,2.4898806,2.8294096,3.275256,3.0146074,2.8396983,3.1277838,3.8377085,3.8342788,3.5118976,3.2718265,3.3609958,3.858286,3.5976372,3.6799474,3.3644254,2.7059445,2.5756202,2.7779658,3.8137012,4.9660425,5.223262,3.2718265,2.6750782,3.3781435,4.0057583,3.5702004,1.4815818,0.3841138,0.044584636,0.020577524,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0274367,0.09602845,0.2503599,0.53158605,1.3375391,1.5330256,1.471293,1.4438564,1.6976458,2.1503513,1.6770682,1.0323058,0.7442205,1.0906088,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.041155048,0.09945804,0.09259886,0.26064864,0.4046913,0.4355576,0.3806842,0.16804978,0.058302987,0.01371835,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.08573969,0.09259886,0.061732575,0.034295876,0.09259886,0.19548649,0.14404267,0.25721905,0.7990939,1.9925903,8.213862,7.956643,5.0483527,2.8911421,4.4275975,4.0263357,3.6044965,2.9460156,2.0886188,1.3341095,0.70306545,0.4389872,0.26750782,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.23321195,0.5453044,0.8162418,0.78537554,0.61389613,0.39783216,0.19548649,0.041155048,0.006859175,0.0,0.05144381,0.15433143,0.26064864,0.20920484,0.18862732,0.22978236,0.31552204,0.3841138,0.15090185,0.14061308,0.2194936,0.29837412,0.31895164,0.10288762,0.0274367,0.010288762,0.0034295875,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.23321195,0.39097297,0.16462019,0.041155048,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.06516216,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.116605975,0.216064,0.31209245,0.38754338,0.4115505,0.36696586,0.31895164,0.5212973,0.96371406,1.371835,1.4507155,1.1626302,1.2517995,1.646202,1.4541451,1.5227368,1.6564908,1.7765263,1.9651536,2.4898806,2.7333813,3.0283258,3.4707425,4.057202,4.6779575,5.5319247,5.778855,5.751418,5.9983487,7.2947326,7.0546613,7.040943,6.9792104,6.7322803,6.3173003,6.3653145,6.468202,6.5059276,6.478491,6.495639,6.6636887,6.8591747,6.989499,7.085528,7.3084507,7.15069,7.301592,6.8214493,5.394741,3.3472774,2.393852,1.6770682,1.2072148,0.9568549,0.84367853,0.8265306,0.90884066,0.86082643,0.7099246,0.71678376,0.53158605,0.7922347,1.3581166,1.762808,1.2243627,0.7442205,0.4938606,0.42869842,0.4698535,0.4972902,0.42526886,0.44927597,0.44584638,0.34981793,0.17147937,0.09602845,0.10288762,0.08916927,0.048014224,0.07545093,0.08916927,0.1371835,0.15090185,0.11317638,0.048014224,0.048014224,0.17833854,0.45613512,0.71678376,0.61046654,0.274367,0.11317638,0.061732575,0.06859175,0.09945804,0.12003556,0.13032432,0.10288762,0.061732575,0.058302987,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.0034295875,0.017147938,0.048014224,0.07888051,0.09602845,0.082310095,0.06516216,0.06859175,0.09945804,0.14747226,0.1371835,0.12003556,0.14404267,0.19891608,0.2194936,0.2469303,0.24007112,0.19891608,0.14747226,0.14404267,0.13375391,0.15776102,0.22292319,0.3806842,0.7133542,0.5418748,0.36010668,0.20577525,0.10288762,0.05144381,0.05144381,0.08573969,0.106317215,0.08916927,0.034295876,0.0274367,0.037725464,0.05144381,0.0548734,0.030866288,0.041155048,0.07888051,0.25378948,0.7922347,2.0337453,3.2272418,4.091498,4.5647807,4.6265135,4.297273,4.3692946,5.435896,6.848886,7.6171136,6.40304,4.3452873,2.8637056,2.0097382,1.670209,1.5433143,1.3992717,1.7559488,3.8479972,8.213862,14.7095,19.397747,20.721567,19.70298,17.230247,14.027013,12.188754,12.082437,13.704632,15.841265,16.060759,14.1299,13.807519,13.982429,14.270514,15.004445,17.106783,19.03764,19.78529,19.305147,18.516342,19.243416,19.198832,19.229696,20.255144,23.262892,24.723896,26.154034,27.584171,29.161781,31.157803,33.22584,31.397873,28.523878,26.44212,25.985985,23.917942,21.428062,19.308577,17.573206,15.470869,11.739478,9.644,8.752307,8.639131,8.889491,8.385342,8.056101,7.8023114,7.716572,8.090397,11.087856,12.768354,12.291641,10.662587,10.731179,11.2421875,12.401388,13.368532,13.958421,14.637479,15.357693,14.7369375,14.688923,14.7197895,11.934964,9.829198,9.750318,9.47938,8.371623,7.3427467,6.9209075,6.018926,5.305572,4.5922174,2.8396983,1.605047,0.96371406,0.7407909,0.7442205,0.77508676,0.9328478,1.1763484,1.255229,1.0700313,0.67219913,0.3566771,0.24350071,0.22292319,0.22978236,0.23321195,0.24350071,0.25378948,0.2469303,0.22635277,0.20920484,0.19891608,0.20234565,0.2194936,0.24350071,0.25378948,0.2709374,0.2709374,0.26407823,0.24007112,0.18862732,0.15776102,0.17490897,0.17490897,0.15090185,0.15090185,0.2709374,0.39097297,0.4115505,0.32238123,0.20577525,0.13375391,0.116605975,0.1920569,0.33266997,0.4629943,0.6310441,0.9945804,1.0700313,0.86082643,0.85739684,1.4198492,1.6530612,1.762808,1.9308578,2.3321195,1.920569,2.1846473,2.4555845,2.6373527,3.2306714,3.6353626,3.216953,3.0043187,3.3266997,3.8137012,3.6696587,3.2272418,3.1449318,3.5976372,4.297273,3.4021509,3.642222,3.4433057,2.6167753,2.386993,3.117495,4.7671266,5.055212,3.7005248,2.393852,3.2066643,4.0229063,4.180667,3.357566,1.5433143,0.39783216,0.044584636,0.020577524,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.09602845,0.37725464,0.97057325,1.0117283,1.1832076,1.7593783,2.6133456,2.6956558,2.0406046,1.1420527,0.45270553,0.38754338,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.017147938,0.0,0.0,0.0,0.010288762,0.01371835,0.017147938,0.020577524,0.044584636,0.06516216,0.08916927,0.116605975,0.12346515,0.09259886,0.07888051,0.06516216,0.061732575,0.106317215,0.24007112,0.28122616,0.20577525,0.14061308,0.32924038,0.15776102,0.1371835,0.69963586,2.270387,5.2781353,13.234778,8.694004,4.9077396,6.1732574,7.8331776,8.868914,7.5039372,5.1683884,3.1037767,2.3664153,1.6016173,0.8162418,0.2777966,0.0548734,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.24350071,0.45956472,0.5178677,0.4424168,0.28465575,0.12346515,0.048014224,0.01371835,0.06516216,0.20577525,0.37382504,0.34638834,0.39440256,0.5418748,0.7305021,0.8505377,0.35324752,0.29837412,0.4664239,0.65505123,0.6790583,0.21263443,0.0548734,0.0274367,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.041155048,0.12689474,0.28808534,0.48014224,0.59674823,0.6379033,0.66533995,0.64476246,0.5178677,0.22635277,0.1371835,0.29494452,0.7682276,1.2312219,0.9842916,1.5810398,1.8108221,1.8142518,1.8108221,2.0920484,1.9651536,2.2566686,2.7299516,3.2512488,3.7862647,4.6779575,5.2506986,5.5559316,6.1492505,8.083538,7.840037,7.6205435,7.8091707,8.14527,7.73029,8.014946,8.217292,8.045813,7.6205435,7.449064,7.3598948,7.0923867,7.1129646,7.490219,7.888051,7.4113383,7.7371492,7.7440085,6.866034,5.096367,4.2389703,3.2581081,2.386993,1.7730967,1.4781522,1.2106444,1.2860953,1.5913286,1.8588364,1.6770682,1.313532,1.2380811,1.2860953,1.1934965,0.6001778,0.52472687,0.5178677,0.50757897,0.4629943,0.39097297,0.5212973,0.432128,0.4355576,0.48014224,0.16462019,0.09945804,0.12003556,0.1371835,0.1371835,0.16804978,0.1920569,0.26407823,0.28122616,0.22978236,0.18176813,0.14061308,0.18176813,0.30866286,0.3841138,0.14404267,0.06516216,0.044584636,0.0548734,0.07888051,0.09602845,0.08916927,0.116605975,0.12346515,0.09259886,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.006859175,0.0034295875,0.020577524,0.034295876,0.044584636,0.07888051,0.061732575,0.0548734,0.07888051,0.13375391,0.18176813,0.18176813,0.15776102,0.18862732,0.25721905,0.274367,0.30523327,0.25378948,0.17833854,0.13032432,0.1371835,0.13032432,0.13375391,0.16119061,0.20920484,0.2503599,0.216064,0.18862732,0.14747226,0.09259886,0.06516216,0.072021335,0.12003556,0.116605975,0.058302987,0.01371835,0.017147938,0.034295876,0.05144381,0.058302987,0.041155048,0.072021335,0.116605975,0.2194936,0.48357183,1.0837497,2.2155135,3.426158,4.2355404,4.431027,4.0674906,3.7485392,4.3521466,5.2164025,5.809721,5.7274113,4.1017866,2.7916842,1.8725548,1.4267083,1.5638919,2.0886188,4.1635194,10.371073,20.982216,33.956345,37.794052,33.08523,24.915953,17.04848,11.931535,10.782623,11.763485,13.876111,15.518884,14.510585,12.651748,13.231348,13.55373,13.310229,14.603184,17.586924,19.071936,19.332584,18.855871,18.313997,17.494326,17.267973,18.427174,20.70442,22.745024,25.162884,28.235794,30.269539,30.897154,31.099499,31.000042,29.59391,27.738503,25.972265,24.52498,22.46037,19.308577,16.96617,15.782962,14.562028,11.105004,8.851766,7.4353456,6.9380555,7.922347,9.167287,9.373062,8.968371,8.453933,8.4093485,11.231899,13.241637,13.255356,11.794352,11.111863,11.149589,12.003556,12.723769,12.847235,12.370522,11.4033785,10.63858,10.199594,10.034973,9.908078,8.738589,8.796892,8.81747,8.364764,7.822889,8.1041155,7.0546613,5.8371577,4.5956473,2.4452958,1.2792361,0.83681935,0.65162164,0.490431,0.36010668,0.36353627,0.4046913,0.432128,0.4115505,0.31895164,0.2194936,0.18519773,0.19548649,0.2194936,0.20920484,0.2194936,0.2194936,0.216064,0.20577525,0.1920569,0.18862732,0.19548649,0.20577525,0.22635277,0.25378948,0.26750782,0.25721905,0.24350071,0.23321195,0.20234565,0.17833854,0.18176813,0.17490897,0.15090185,0.15090185,0.21263443,0.2503599,0.23664154,0.1920569,0.19891608,0.18519773,0.2777966,0.53501564,0.88826317,1.1420527,1.0425946,1.4644338,1.4953002,1.0906088,1.0631721,1.2792361,1.5673214,2.1091962,2.8054025,3.2649672,2.3732746,2.5138876,2.7093742,2.8259802,3.5633414,3.940596,3.4810312,3.1792276,3.2272418,3.0043187,2.4658735,2.0406046,2.8019729,4.417309,5.137522,3.875434,3.865145,3.5016088,2.5961976,2.386993,3.2203827,4.5784993,4.1326528,2.4590142,3.0489032,4.0194764,3.9886103,3.5599117,2.7299516,0.89169276,0.17833854,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.048014224,0.037725464,0.037725464,0.048014224,0.034295876,0.0034295875,0.017147938,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.020577524,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.041155048,0.20920484,0.42526886,0.5453044,0.86082643,1.5433143,2.6476414,1.8142518,1.255229,0.70649505,0.20920484,0.07888051,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.017147938,0.0,0.0,0.0,0.010288762,0.01371835,0.034295876,0.106317215,0.17833854,0.22635277,0.34638834,0.52815646,0.6241849,0.4664239,0.40126175,0.32581082,0.26407823,0.34981793,0.4355576,0.5590228,0.51100856,0.5624523,1.4644338,0.59674823,0.31895164,1.862266,6.3893213,14.983868,20.426622,10.930096,7.874333,12.946692,8.162418,16.70895,16.071047,10.906088,5.895461,5.7377,4.3933015,2.5481834,1.0597426,0.28122616,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.15433143,0.22292319,0.19891608,0.16119061,0.061732575,0.037725464,0.09259886,0.09259886,0.15090185,0.26750782,0.4081209,0.4972902,0.4115505,0.26407823,0.31895164,0.4972902,0.65505123,0.59674823,0.26407823,0.1097468,0.072021335,0.08916927,0.07545093,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09259886,0.22978236,0.4115505,0.77851635,1.0631721,1.0185875,0.7133542,0.5178677,0.36010668,0.23664154,0.13375391,0.07888051,0.15433143,1.0940384,1.0357354,0.864256,1.0528834,1.6633499,2.3458378,2.7093742,2.7333813,2.5893385,2.6407824,3.3369887,5.103226,6.5127864,7.034084,7.034084,6.447624,6.3481665,6.824879,7.4970784,7.5210853,7.438775,7.8091707,8.083538,8.1212635,8.193284,7.888051,7.133542,6.608815,6.4716315,6.3618846,6.667118,7.3221693,8.47451,8.868914,5.830299,5.1580997,5.1100855,4.4927597,3.2581081,2.503599,2.0028791,2.5173173,3.841138,4.852866,3.508468,2.668219,1.8691251,1.3203912,1.0151579,0.7476501,1.0048691,0.9842916,0.8093826,0.61046654,0.548734,0.47671264,0.28465575,0.1920569,0.22635277,0.21263443,0.274367,0.25378948,0.3018037,0.36353627,0.16804978,0.09602845,0.06859175,0.07888051,0.17147937,0.42869842,0.30523327,0.1097468,0.006859175,0.034295876,0.106317215,0.15433143,0.15776102,0.14747226,0.13375391,0.12346515,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.030866288,0.017147938,0.034295876,0.05144381,0.06859175,0.09259886,0.0548734,0.09945804,0.15433143,0.18176813,0.18176813,0.13375391,0.15090185,0.1920569,0.23664154,0.274367,0.22635277,0.10288762,0.0548734,0.08916927,0.07545093,0.1371835,0.17833854,0.2469303,0.32238123,0.33609957,0.26407823,0.18862732,0.12346515,0.07545093,0.07545093,0.11317638,0.13032432,0.09945804,0.037725464,0.0,0.024007112,0.030866288,0.048014224,0.07888051,0.09259886,0.14061308,0.16119061,0.16119061,0.216064,0.47328308,1.3512574,2.1023371,2.702515,3.1655092,3.5564823,3.957744,4.506478,4.530485,4.3487167,5.2644167,3.8720043,2.6373527,1.6427724,1.097468,1.3443983,3.0043187,8.920357,22.230585,41.744938,61.93492,59.884026,44.14565,27.045727,15.9613,13.337666,14.959861,15.9613,15.96816,14.96329,13.289652,12.97413,13.077017,13.289652,14.064738,16.616352,18.900457,18.20768,16.7844,15.638919,14.5414505,13.2862215,13.80409,16.434584,19.668684,20.155685,20.875898,24.93996,29.480734,31.809423,29.405283,27.145185,24.806206,22.94394,21.424633,19.408035,17.394867,15.573756,14.555169,14.061309,12.939834,11.218181,8.766026,6.7494283,6.15268,7.750868,9.043822,9.030104,8.639131,8.22758,7.5690994,8.971801,10.844356,12.003556,11.842365,10.329918,9.791472,10.868362,11.183885,10.429376,10.329918,11.269625,9.242738,7.0478024,6.3207297,7.5519514,6.931196,7.133542,7.2364297,6.5642304,4.6848164,5.6005163,4.262977,3.018037,2.5310357,1.786815,1.1866373,0.864256,0.5693115,0.29837412,0.274367,0.3841138,0.39440256,0.33952916,0.25721905,0.18176813,0.13375391,0.14061308,0.16462019,0.18519773,0.19891608,0.19891608,0.18862732,0.18862732,0.1920569,0.16804978,0.15433143,0.18176813,0.216064,0.25378948,0.29151493,0.26407823,0.22292319,0.20920484,0.22635277,0.21263443,0.18862732,0.16462019,0.14747226,0.1371835,0.1371835,0.16119061,0.13032432,0.09945804,0.09945804,0.1371835,0.2709374,0.59674823,1.1489118,1.704505,1.8005334,1.605047,1.8416885,1.8759843,1.7833855,2.318401,2.7711067,2.983741,2.7470996,2.2292318,1.9823016,2.301253,2.6990852,2.486451,2.0028791,2.6236343,5.528495,6.3824625,5.6073756,4.396731,4.715683,3.3369887,3.1106358,4.012617,5.2815647,5.4153185,4.914599,4.5613513,3.6216443,2.644212,3.4467354,3.4604537,2.411,2.177788,3.0969174,3.9508848,3.2821152,2.3081124,1.8999915,1.6736387,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.044584636,0.037725464,0.18176813,0.19548649,0.24350071,0.16462019,0.017147938,0.09259886,0.16462019,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.106317215,0.08573969,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.061732575,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.058302987,0.22978236,0.65505123,0.8025235,0.39097297,0.09602845,0.10288762,0.09259886,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6344737,1.08032,0.7888051,0.048014224,0.0,0.0,0.06516216,0.07888051,0.044584636,0.072021335,0.06516216,0.041155048,0.017147938,0.0,0.0,0.010288762,0.0274367,0.024007112,0.06859175,0.33952916,0.12003556,0.0548734,0.07545093,0.13032432,0.19891608,0.19548649,0.16119061,0.11317638,0.07545093,0.082310095,0.29494452,0.9602845,1.0151579,0.4629943,0.39097297,0.4115505,0.7922347,1.9720128,4.081209,6.9517736,5.6793966,3.3129816,3.5359046,6.3618846,8.1384115,13.070158,12.627741,9.321619,5.885172,5.284994,4.7842746,3.4604537,2.3046827,1.6016173,0.9534253,0.4046913,0.106317215,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.072021335,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.044584636,0.041155048,0.030866288,0.01371835,0.006859175,0.017147938,0.017147938,0.030866288,0.06859175,0.106317215,0.12689474,0.12003556,0.06859175,0.11317638,0.21263443,0.30866286,0.31552204,0.17147937,0.11317638,0.1097468,0.12346515,0.09945804,0.048014224,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.072021335,0.16804978,0.4081209,0.7476501,0.94999576,0.939707,0.8128122,0.61389613,0.44584638,0.33266997,0.26750782,0.21263443,0.33266997,0.31895164,0.42183927,0.6207553,0.6241849,1.0666018,1.2860953,1.4541451,2.0989075,4.139512,4.046913,4.386442,4.8425775,5.271276,5.693115,6.4544835,6.8145905,6.948344,6.8454566,6.3035817,6.5779486,6.924337,7.1781263,7.284444,7.291303,7.5725293,6.941485,6.3790326,6.2864337,6.509357,6.7185616,7.3221693,7.8331776,7.905199,7.366754,7.829748,7.507367,6.807731,5.658819,3.5153272,2.760818,2.760818,2.901431,3.100347,3.789694,3.9543142,2.9906003,2.0474637,1.5570327,1.2586586,1.0768905,0.83338976,0.5555932,0.34981793,0.36696586,0.40126175,0.2503599,0.4081209,1.0220171,1.8965619,1.9480057,1.2517995,0.52472687,0.1371835,0.106317215,0.09259886,0.16119061,0.2194936,0.2503599,0.29151493,0.16119061,0.05144381,0.010288762,0.037725464,0.06859175,0.08916927,0.07888051,0.061732575,0.05144381,0.048014224,0.01371835,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.07545093,0.1371835,0.13032432,0.072021335,0.06859175,0.058302987,0.09945804,0.14747226,0.18862732,0.20920484,0.23664154,0.2777966,0.28808534,0.28808534,0.37382504,0.37382504,0.36353627,0.32581082,0.28122616,0.30866286,0.33952916,0.34638834,0.35324752,0.36353627,0.34638834,0.31209245,0.22978236,0.14061308,0.09602845,0.12346515,0.17147937,0.16462019,0.09945804,0.020577524,0.01371835,0.006859175,0.041155048,0.07888051,0.10288762,0.10288762,0.20234565,0.2777966,0.40126175,0.59331864,0.84024894,1.3958421,1.6770682,1.6942163,1.6736387,2.054323,2.9940298,4.184097,5.2575574,5.8543057,5.6176643,3.758828,2.4041407,1.5433143,1.3169615,2.0508933,6.883182,18.95533,36.21987,54.053726,65.27877,60.01778,46.199974,31.66881,21.832754,19.648108,21.0268,19.658396,16.160215,12.000127,9.517105,8.958082,9.630281,12.679185,17.487467,21.671564,20.495214,17.065628,13.927555,12.274493,11.928105,11.423956,12.812939,14.88098,16.825556,18.241976,20.141968,22.916504,25.564144,27.066305,26.400965,24.182022,21.740154,19.682402,18.094503,16.527182,14.55174,12.696333,12.065289,12.332796,11.766914,10.868362,9.870353,8.968371,8.556821,9.22902,8.364764,6.8214493,6.392751,7.2467184,7.936065,8.879202,10.364213,11.694893,12.123591,10.854645,10.299051,10.028113,10.089847,10.264755,10.048691,10.9198065,9.4862385,7.641121,6.3824625,5.8062916,5.439326,5.1855364,4.887162,4.4516044,3.8308492,3.1826572,2.335549,1.8554068,1.786815,1.6393428,1.3443983,0.96371406,0.6310441,0.44927597,0.48357183,0.59331864,0.52815646,0.37382504,0.216064,0.13375391,0.11317638,0.11317638,0.12003556,0.13032432,0.16119061,0.13375391,0.1371835,0.15776102,0.16804978,0.14404267,0.13032432,0.15433143,0.18862732,0.20920484,0.216064,0.22978236,0.22635277,0.22635277,0.23321195,0.2503599,0.23664154,0.19891608,0.18176813,0.1920569,0.20920484,0.17490897,0.15433143,0.15090185,0.18176813,0.2469303,0.33266997,0.61046654,1.0323058,1.6770682,2.7402403,3.7348208,4.554492,4.6779575,4.331569,4.4687524,3.3952916,3.1106358,2.884283,2.5721905,2.6304936,2.411,2.6853669,3.3815732,4.033195,3.7485392,4.4550343,4.8768735,4.756838,4.461893,4.996909,5.020916,4.482471,4.290414,4.506478,4.3178506,4.619654,4.331569,4.0709205,4.389872,5.7925735,4.3281393,2.2292318,1.3066728,1.8588364,2.6956558,2.435007,1.8554068,1.4953002,1.4438564,1.3546871,0.2709374,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.020577524,0.1097468,0.0548734,0.048014224,0.061732575,0.061732575,0.017147938,0.034295876,0.09602845,0.09602845,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08573969,0.12003556,0.06516216,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.017147938,0.08573969,0.2777966,0.2777966,0.29837412,0.4355576,0.65848076,0.8128122,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44927597,0.67219913,0.45956472,0.024007112,0.0,0.0,0.061732575,0.082310095,0.08573969,0.20920484,0.31552204,0.24350071,0.22635277,0.24007112,0.0,0.0034295875,0.034295876,0.034295876,0.034295876,0.16804978,0.044584636,0.017147938,0.024007112,0.034295876,0.037725464,0.058302987,0.09259886,0.16804978,0.24007112,0.19891608,0.18519773,0.4972902,0.59331864,0.432128,0.45270553,0.7613684,1.2415106,1.9480057,2.8259802,3.7176728,2.8808534,4.1943855,6.5059276,8.886061,10.6488695,13.1421795,13.368532,11.204462,7.966932,6.4098988,5.8817425,4.9077396,3.7931237,2.668219,1.4850113,0.5796003,0.14061308,0.0,0.0,0.0,0.0,0.034295876,0.09259886,0.15776102,0.20234565,0.15090185,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.017147938,0.006859175,0.024007112,0.058302987,0.09945804,0.116605975,0.08573969,0.082310095,0.10288762,0.12689474,0.116605975,0.07545093,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.041155048,0.14061308,0.35324752,0.58988905,0.78194594,0.8848336,0.7888051,0.6276145,0.48700142,0.38754338,0.3018037,0.22978236,0.20577525,0.26407823,0.42183927,0.65162164,0.5453044,0.58302987,0.83338976,1.4061309,2.4658735,2.4075704,2.5241764,3.1723683,4.15323,4.715683,5.7102633,5.5833683,5.576509,5.8543057,5.528495,5.3844523,5.5662203,5.7239814,5.761707,5.830299,5.9914894,5.8062916,5.675967,5.7994323,6.169828,6.464772,6.728851,6.8969,7.023795,7.284444,7.795452,7.06495,6.0497923,5.130663,4.125794,3.2649672,4.3521466,4.8117113,4.2046742,4.245829,4.9077396,4.8288593,3.9097297,2.8156912,2.9631636,1.6667795,1.0597426,0.7510797,0.6036074,0.70649505,0.58302987,0.67219913,1.0837497,1.6633499,1.961724,1.2346514,0.70649505,0.4081209,0.37039545,0.6310441,0.48357183,0.29837412,0.16462019,0.1097468,0.10288762,0.05144381,0.020577524,0.01371835,0.024007112,0.034295876,0.05144381,0.061732575,0.06516216,0.058302987,0.030866288,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.006859175,0.020577524,0.0274367,0.041155048,0.034295876,0.017147938,0.0034295875,0.01371835,0.10288762,0.14747226,0.13375391,0.09602845,0.09602845,0.07545093,0.08916927,0.12003556,0.14747226,0.15776102,0.22292319,0.33952916,0.37725464,0.32238123,0.29494452,0.34638834,0.36353627,0.4046913,0.4424168,0.37382504,0.3841138,0.37725464,0.38754338,0.40126175,0.37039545,0.2777966,0.19548649,0.14747226,0.14061308,0.14747226,0.14404267,0.12003556,0.07545093,0.024007112,0.024007112,0.020577524,0.041155048,0.061732575,0.08573969,0.14404267,0.15776102,0.39097297,0.7476501,1.2037852,1.8005334,1.821111,1.6153357,1.3821237,1.2380811,1.2209331,2.054323,3.450165,5.113515,6.200694,5.3398676,3.7279615,2.6647894,2.1126258,2.2635276,3.5290456,11.454823,26.661613,41.504868,51.14887,53.566727,49.78389,40.177616,29.295536,21.239435,19.678972,19.994495,17.37772,13.365103,9.705732,8.347616,8.207003,9.434795,13.025573,17.648657,19.637817,16.654078,13.004995,10.449953,9.506817,9.427936,9.249598,10.398509,11.674315,12.696333,13.934414,16.760393,19.377169,20.937632,21.510372,22.096832,20.03565,17.857862,16.184223,15.145059,14.38026,13.272504,12.339656,11.5645685,10.940384,10.477389,10.484249,10.22703,9.431366,8.477941,8.399059,7.4181976,5.9914894,5.312431,5.645101,6.2967224,7.720001,9.22216,10.545981,11.338216,11.170166,10.593996,9.746887,9.349055,9.523964,9.777754,10.089847,9.39707,8.522525,7.764586,6.910619,5.7102633,4.715683,3.8514268,3.1860867,2.9494452,2.2909644,1.7079345,1.3958421,1.3238207,1.2346514,1.3238207,1.155771,0.980862,0.922559,0.9568549,0.77851635,0.5658819,0.33952916,0.15776102,0.08573969,0.07888051,0.08573969,0.08916927,0.09259886,0.116605975,0.13032432,0.14747226,0.15090185,0.13375391,0.1097468,0.11317638,0.13375391,0.16119061,0.18176813,0.18862732,0.2194936,0.22292319,0.2194936,0.22292319,0.24007112,0.2503599,0.23321195,0.2194936,0.21263443,0.20234565,0.18176813,0.16119061,0.23664154,0.42869842,0.6790583,1.0494537,1.6839274,2.3492675,2.7402403,2.4624438,3.3609958,4.413879,4.681387,4.245829,4.2183924,3.532475,3.2718265,3.117495,2.877424,2.5001693,2.585909,2.9563043,3.4433057,3.6799474,3.1312134,3.9646032,4.6882463,4.8597255,4.6779575,4.9934793,5.055212,4.5819287,3.9097297,3.6627994,4.756838,5.127233,4.214963,4.232111,4.938606,3.6319332,2.1674993,1.5227368,1.313532,1.214074,0.9534253,0.9534253,0.91569984,0.8093826,0.823101,1.3546871,0.65162164,0.1920569,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.006859175,0.061732575,0.10288762,0.08916927,0.0,0.0,0.09945804,0.13375391,0.07545093,0.0548734,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.07545093,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.041155048,0.17490897,0.5041494,0.94999576,1.2826657,1.3272504,0.9294182,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13032432,0.13032432,0.06516216,0.0,0.0,0.0,0.034295876,0.05144381,0.072021335,0.18519773,0.29494452,0.22978236,0.2194936,0.2503599,0.048014224,0.010288762,0.020577524,0.024007112,0.006859175,0.010288762,0.010288762,0.0274367,0.034295876,0.0274367,0.0,0.01371835,0.082310095,0.2194936,0.36010668,0.36353627,0.2194936,0.19891608,0.30523327,0.5212973,0.8162418,0.9774324,1.2209331,1.762808,2.510458,3.069481,3.2478194,5.381023,8.862054,12.233338,13.169616,14.754086,14.534592,12.850664,10.405369,8.268735,7.56224,6.0978065,4.616225,3.3301294,1.8965619,0.7510797,0.18519773,0.0,0.0,0.0,0.0,0.15433143,0.31895164,0.4389872,0.5555932,0.5521636,0.3841138,0.16462019,0.0,0.0,0.0,0.020577524,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.024007112,0.044584636,0.07545093,0.09602845,0.09602845,0.06516216,0.030866288,0.010288762,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.08916927,0.24007112,0.45613512,0.6893471,0.7682276,0.7133542,0.59674823,0.4698535,0.37382504,0.31895164,0.2777966,0.26064864,0.32924038,0.59674823,0.35324752,0.38754338,0.6859175,1.0563129,1.1283343,1.4369972,1.4987297,1.9925903,2.9460156,3.7313912,4.8117113,4.605936,4.729401,5.2026844,4.461893,4.256118,4.32471,4.232111,4.0194764,4.2355404,4.57164,4.698535,4.8082814,5.038064,5.4804807,5.895461,5.936616,5.977771,6.1629686,6.39961,6.591667,6.101236,5.295283,4.647091,4.7431192,3.8479972,5.206114,5.7994323,4.962613,4.3624353,5.446185,5.970912,5.2575574,3.9508848,4.029765,2.253239,1.7456601,1.4815818,1.2689474,1.7730967,0.94656616,0.91912943,1.2655178,1.5433143,1.2655178,0.48014224,0.7476501,1.3306799,1.7216529,1.6187652,0.6790583,0.23664154,0.061732575,0.0,0.0,0.0034295875,0.044584636,0.08573969,0.09602845,0.020577524,0.030866288,0.058302987,0.08573969,0.082310095,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.041155048,0.01371835,0.017147938,0.020577524,0.034295876,0.0548734,0.07545093,0.106317215,0.09259886,0.05144381,0.017147938,0.034295876,0.15433143,0.1920569,0.16804978,0.116605975,0.10288762,0.09602845,0.13375391,0.16462019,0.17490897,0.16462019,0.2194936,0.36010668,0.41498008,0.36353627,0.34638834,0.32924038,0.38754338,0.45956472,0.4938606,0.4355576,0.37725464,0.3841138,0.4115505,0.41840968,0.3566771,0.22292319,0.15090185,0.14747226,0.18176813,0.19548649,0.17490897,0.13032432,0.082310095,0.05144381,0.07888051,0.09259886,0.061732575,0.037725464,0.05144381,0.12003556,0.08916927,0.37039545,0.90541106,1.7216529,2.9185789,3.0900583,2.6785078,2.061182,1.430138,0.7922347,1.4198492,2.9151495,4.722542,5.8165803,4.712253,3.4433057,2.620205,2.194936,2.527606,4.383013,14.565458,30.739393,41.079597,42.16335,38.9704,36.33305,28.856548,20.714708,15.227368,14.887839,14.339106,12.243628,9.602845,7.455923,6.9071894,7.226141,8.89635,12.199042,15.573756,15.638919,11.351934,8.196714,6.7631464,6.7871537,7.157549,7.257007,8.22758,9.043822,9.510246,10.261326,13.066729,15.261664,16.266533,16.558048,17.679523,16.571766,15.326826,14.393978,13.749216,12.895248,12.243628,12.144169,11.574858,10.47396,9.736599,9.863494,9.626852,8.796892,7.73029,7.39762,6.6636887,5.627953,4.846007,4.4927597,4.372724,5.4976287,6.6636887,7.73372,8.776315,10.052121,10.110424,9.403929,9.030104,9.3079,9.777754,9.170717,8.683716,8.615124,8.635701,7.7577267,5.9331865,4.5647807,3.4844608,2.719663,2.4898806,2.2429502,1.8828435,1.5776103,1.3786942,1.2106444,1.4027013,1.3992717,1.3649758,1.3546871,1.3203912,0.83338976,0.48700142,0.24350071,0.09602845,0.061732575,0.0548734,0.058302987,0.058302987,0.061732575,0.072021335,0.12346515,0.1371835,0.12003556,0.09602845,0.08573969,0.08916927,0.106317215,0.13032432,0.14747226,0.15776102,0.19548649,0.20234565,0.20234565,0.20920484,0.22292319,0.23664154,0.22978236,0.20920484,0.18176813,0.14747226,0.15776102,0.16462019,0.26750782,0.5418748,1.0734608,1.5055889,2.2120838,2.8945718,3.0866287,2.1572106,2.5447538,3.0969174,3.1860867,2.8156912,2.6236343,2.6236343,2.5961976,2.6853669,2.7230926,2.2292318,2.4144297,2.8019729,3.0420442,2.9803114,2.6373527,3.5530527,4.7019644,5.1169443,4.770556,4.5853586,4.588788,4.214963,3.9440255,4.170378,5.192395,4.9008803,4.297273,3.9646032,3.4467354,1.2517995,0.7956643,1.4198492,1.4610043,0.6790583,0.23664154,0.18519773,0.28808534,0.28465575,0.30523327,0.8745448,0.6276145,0.22635277,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.11317638,0.12003556,0.07888051,0.07888051,0.14747226,0.16462019,0.12003556,0.10288762,0.08916927,0.06859175,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05144381,0.25378948,0.8676856,1.4267083,1.7182233,1.5776103,0.8848336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.020577524,0.01371835,0.0274367,0.0274367,0.01371835,0.0034295875,0.020577524,0.09602845,0.020577524,0.0,0.0034295875,0.01371835,0.017147938,0.024007112,0.037725464,0.034295876,0.017147938,0.006859175,0.017147938,0.082310095,0.1920569,0.31552204,0.40126175,0.32238123,0.3018037,0.41498008,0.64819205,0.8711152,0.77851635,0.88826317,1.6873571,2.8534167,3.234101,2.767677,4.012617,7.5382333,12.003556,14.150477,14.946142,13.296511,11.667457,10.607714,8.755736,8.134981,6.138962,4.431027,3.3850029,2.095478,0.96714365,0.33266997,0.082310095,0.058302987,0.06859175,0.058302987,0.30866286,0.51100856,0.6036074,0.7476501,0.91569984,0.864256,0.5727411,0.21263443,0.14061308,0.10288762,0.13375391,0.12346515,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.034295876,0.048014224,0.048014224,0.030866288,0.017147938,0.006859175,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.048014224,0.14404267,0.33266997,0.5521636,0.65848076,0.64819205,0.5555932,0.45613512,0.39783216,0.35324752,0.31552204,0.28122616,0.22635277,0.2503599,0.39440256,0.66876954,0.9568549,1.0323058,1.5330256,1.4198492,1.3752645,1.8039631,2.8156912,4.297273,4.40359,4.5339146,4.6093655,3.0729103,3.2443898,3.2203827,2.8945718,2.5619018,2.9185789,3.7313912,3.8857226,3.9200184,4.139512,4.5922174,5.038064,5.161529,5.267846,5.411889,5.360445,5.4016004,5.693115,5.56965,5.1169443,5.192395,4.297273,4.804852,5.055212,4.5784993,4.1120753,5.2644167,5.638242,5.2472687,4.4721823,4.057202,2.7230926,2.6922262,2.4624438,1.978872,2.6545007,1.2826657,0.96714365,1.1008976,1.138623,0.58988905,0.61046654,1.6942163,2.6476414,2.8122618,2.054323,0.45956472,0.024007112,0.0,0.0,0.0,0.020577524,0.082310095,0.15776102,0.17147937,0.024007112,0.017147938,0.061732575,0.106317215,0.106317215,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09602845,0.16462019,0.048014224,0.058302987,0.07888051,0.08916927,0.09945804,0.12346515,0.14404267,0.1371835,0.09259886,0.041155048,0.0548734,0.19548649,0.26750782,0.2503599,0.16462019,0.082310095,0.116605975,0.19548649,0.2469303,0.25721905,0.26407823,0.26407823,0.33609957,0.37382504,0.38754338,0.51100856,0.4115505,0.51100856,0.5453044,0.48014224,0.52472687,0.3806842,0.39097297,0.41840968,0.39097297,0.31209245,0.1920569,0.1371835,0.14747226,0.20234565,0.2503599,0.24007112,0.18176813,0.116605975,0.08573969,0.14747226,0.16462019,0.082310095,0.024007112,0.0274367,0.048014224,0.05144381,0.2194936,0.7305021,1.7319417,3.3678548,4.5270553,4.5510626,3.6593697,2.2052248,0.6790583,1.1111864,2.6236343,4.3041325,5.1238036,3.9508848,2.8019729,2.054323,1.6187652,2.0165975,4.389872,14.812388,28.856548,34.84461,31.202387,26.448978,23.1943,16.170506,10.179015,7.630832,8.539673,8.169277,7.8777623,7.034084,5.7582774,4.9180284,5.3501563,7.281014,10.329918,13.042721,12.905538,7.73372,4.7259717,3.8274195,4.4241676,5.360445,5.7308407,6.759717,7.4765005,7.675417,7.9086285,9.856634,11.14273,11.941824,12.603734,13.656617,13.780083,13.570878,13.289652,12.730629,11.207891,10.405369,10.714031,10.854645,10.336777,9.445084,9.078118,8.433355,7.64798,6.9552035,6.6739774,5.936616,5.06893,4.4687524,4.0503426,3.2478194,3.2409601,3.6593697,4.2698364,5.288424,7.3839016,8.412778,8.31332,8.433355,9.033533,9.277034,8.114404,7.4010496,7.500508,7.829748,6.8557453,5.2438393,4.1600895,3.3266997,2.6750782,2.3595562,2.294394,2.1126258,1.903421,1.7113642,1.5330256,1.5913286,1.670209,1.6976458,1.6290541,1.430138,0.7510797,0.34981793,0.14404267,0.06859175,0.072021335,0.05144381,0.041155048,0.034295876,0.034295876,0.041155048,0.08916927,0.09259886,0.07545093,0.06859175,0.07888051,0.061732575,0.072021335,0.08916927,0.09945804,0.11317638,0.14404267,0.16462019,0.17833854,0.1920569,0.20234565,0.20234565,0.18862732,0.15776102,0.12346515,0.09602845,0.116605975,0.16804978,0.22978236,0.4424168,1.0940384,1.3375391,1.786815,2.1846473,2.311542,1.99602,2.1160555,1.8554068,1.5776103,1.3958421,1.1763484,1.3889829,1.5055889,1.8039631,2.1572106,2.0646117,2.0337453,2.270387,2.7813954,3.2066643,2.8259802,3.083199,4.1600895,4.616225,4.1635194,3.6353626,4.0263357,3.7039545,4.2218223,5.2987127,4.8185706,3.998899,4.3624353,3.2992632,1.0460242,0.6756287,1.4987297,1.9445761,1.3341095,0.26064864,0.58988905,0.3018037,0.17833854,0.13032432,0.18862732,0.5212973,0.26407823,0.07888051,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058302987,0.15776102,0.20920484,0.20234565,0.20920484,0.18519773,0.1371835,0.12346515,0.12689474,0.12689474,0.082310095,0.020577524,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.32924038,0.9431366,1.3752645,1.5536032,1.4335675,0.99801,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09259886,0.030866288,0.024007112,0.037725464,0.041155048,0.030866288,0.041155048,0.1371835,0.216064,0.25721905,0.30523327,0.24350071,0.2194936,0.4081209,0.6001778,0.19891608,0.28465575,0.9911508,2.2841053,3.4055803,2.867135,2.1983654,2.568761,4.3041325,7.6925645,13.015285,9.952662,7.7577267,6.2075534,5.1409516,4.4721823,4.3487167,4.0537724,3.4433057,2.5721905,1.6942163,1.1214751,0.6824879,0.4081209,0.29837412,0.33609957,0.29837412,0.32581082,0.29494452,0.20920484,0.19891608,0.5521636,1.0151579,1.2243627,1.0666018,0.70306545,0.5178677,0.44584638,0.40126175,0.29151493,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.07545093,0.2469303,0.47328308,0.6379033,0.6859175,0.6241849,0.53844523,0.4629943,0.3841138,0.29837412,0.21263443,0.18862732,0.2194936,0.28808534,0.37382504,0.45613512,0.48357183,0.52472687,0.96371406,1.7662375,2.486451,4.6608095,4.0777793,3.216953,2.8534167,2.061182,2.037175,1.6907866,1.605047,1.903421,2.2566686,2.9048605,2.9288676,3.0146074,3.3609958,3.6765177,3.957744,4.4413157,4.863155,4.996909,4.65395,5.0449233,5.6828265,5.8337283,5.360445,4.715683,3.8617156,4.232111,4.722542,4.6882463,3.9680326,3.858286,3.683377,3.8548563,4.2183924,4.057202,3.3884325,3.4192986,3.0420442,2.0817597,1.313532,1.2380811,1.3855534,1.8382589,2.0063086,0.6241849,1.1249046,2.0577524,1.6770682,0.2469303,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.048014224,0.024007112,0.0,0.0,0.0,0.01371835,0.106317215,0.18519773,0.17147937,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.20920484,0.41498008,0.18176813,0.13375391,0.16804978,0.17833854,0.15090185,0.1371835,0.08916927,0.12346515,0.116605975,0.0548734,0.030866288,0.10288762,0.23321195,0.32924038,0.31552204,0.106317215,0.13032432,0.15433143,0.19891608,0.2777966,0.4115505,0.31552204,0.24350071,0.25721905,0.35324752,0.48700142,0.5727411,0.59674823,0.58302987,0.5624523,0.548734,0.41498008,0.35324752,0.31895164,0.28808534,0.274367,0.21263443,0.17833854,0.16119061,0.16462019,0.21263443,0.16462019,0.13375391,0.116605975,0.1097468,0.12346515,0.061732575,0.0274367,0.0274367,0.048014224,0.061732575,0.072021335,0.07545093,0.22978236,0.75450927,1.937717,4.3178506,5.8200097,5.7102633,3.9028704,0.9602845,0.864256,2.085189,3.6970954,4.537344,3.2203827,1.961724,1.3169615,1.1900668,1.9582944,4.4859004,11.543991,17.645227,19.637817,17.364002,13.704632,10.285333,7.1884155,5.381023,5.07236,5.7068334,7.233,8.364764,7.98065,6.258997,4.6848164,4.746549,6.701414,9.80862,12.576297,12.771784,8.097256,4.5922174,3.1723683,3.5770597,4.3933015,4.7499785,5.2575574,5.693115,5.7822843,5.2335505,6.3824625,7.226141,8.069819,8.992378,9.873782,9.750318,9.253027,8.882631,8.56025,7.6445503,6.948344,7.6274023,8.4093485,8.724871,8.711152,8.491658,7.5690994,6.4990683,5.610805,4.99005,4.4756117,3.899441,3.7039545,3.758828,3.357566,2.976882,2.901431,2.976882,3.2855449,4.149801,5.188966,5.7136927,6.0978065,6.420188,6.4716315,6.420188,5.970912,5.4153185,4.8768735,4.3041325,3.7279615,3.5393343,3.100347,2.369845,1.9068506,1.6393428,1.4335675,1.4575747,1.605047,1.4953002,1.6427724,1.961724,2.085189,1.8588364,1.3581166,0.65162164,0.29837412,0.14747226,0.09602845,0.12346515,0.061732575,0.0548734,0.048014224,0.030866288,0.030866288,0.06859175,0.06859175,0.06859175,0.07888051,0.09259886,0.0548734,0.044584636,0.05144381,0.06516216,0.07545093,0.08916927,0.1097468,0.13375391,0.15090185,0.15090185,0.16462019,0.15776102,0.13375391,0.106317215,0.106317215,0.12003556,0.16804978,0.216064,0.274367,0.39783216,0.7373613,1.2003556,1.4507155,1.3855534,1.1283343,1.6770682,1.4953002,1.2998136,1.4232788,1.8005334,1.8245405,1.7216529,1.6667795,1.7216529,1.8313997,2.1229146,2.2155135,3.474172,4.863155,2.959734,2.7882545,2.6647894,2.3458378,1.961724,1.9994495,3.0351849,2.9117198,3.3198407,4.170378,3.5873485,4.07435,3.8857226,2.4555845,0.83338976,1.6633499,3.0043187,2.0131679,0.84367853,0.4424168,0.5658819,0.29494452,0.20234565,0.31895164,0.5453044,0.65505123,0.20577525,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072021335,0.19891608,0.26064864,0.20920484,0.18176813,0.1371835,0.09945804,0.1371835,0.15090185,0.106317215,0.08916927,0.10288762,0.09259886,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.12346515,0.5007198,1.0082988,1.3684053,1.4850113,1.4507155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.08573969,0.24350071,0.4424168,0.16804978,0.09945804,0.07888051,0.041155048,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.017147938,0.006859175,0.0034295875,0.006859175,0.01371835,0.030866288,0.041155048,0.08573969,0.18176813,0.3018037,0.39097297,0.4081209,0.42526886,0.41840968,0.33609957,0.09945804,0.216064,2.7916842,5.020916,5.038064,1.8931323,2.1194851,3.3301294,7.682276,13.248496,14.040731,8.241299,5.7891436,5.0757895,4.664239,3.2992632,2.3664153,1.7662375,1.3889829,1.1592005,1.0220171,1.0631721,1.3306799,1.5193073,1.5158776,1.3992717,1.039165,0.66191036,0.34638834,0.15090185,0.15090185,0.20234565,0.31895164,0.38754338,0.36696586,0.274367,0.34638834,0.30523327,0.29151493,0.31552204,0.25721905,0.18862732,0.06859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.12003556,0.16462019,0.16462019,0.14747226,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.1097468,0.28465575,0.48357183,0.66191036,0.7956643,0.6824879,0.5761707,0.45270553,0.31552204,0.20234565,0.19548649,0.24007112,0.31209245,0.3806842,0.4081209,0.4424168,0.5041494,0.7373613,1.0563129,1.1317638,1.6359133,1.7765263,1.6770682,1.5398848,1.646202,2.3732746,2.1640697,1.8005334,1.6976458,1.9171394,2.4967396,2.2155135,2.1846473,2.6579304,3.0557625,3.3541365,3.6456516,3.9303071,4.091498,3.8960114,4.57164,4.7808447,4.914599,4.98662,4.6402316,3.3198407,3.2306714,3.5770597,3.758828,3.3678548,3.7176728,3.5873485,3.391862,3.2958336,3.216953,3.4055803,4.2183924,4.108646,2.9220085,1.9102802,2.959734,2.9254382,2.3286898,1.704505,1.6153357,1.546744,1.1214751,0.53501564,0.048014224,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.6962063,0.59674823,0.26750782,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.28465575,0.5590228,0.41498008,0.26750782,0.18176813,0.18176813,0.2194936,0.19891608,0.13032432,0.09945804,0.07888051,0.061732575,0.06859175,0.1097468,0.216064,0.4424168,0.6241849,0.38754338,0.432128,0.32924038,0.26407823,0.3018037,0.38754338,0.4081209,0.48357183,0.52472687,0.4972902,0.41498008,0.75450927,0.58988905,0.432128,0.51100856,0.78194594,0.5796003,0.50757897,0.5041494,0.490431,0.36010668,0.24007112,0.21263443,0.216064,0.21263443,0.20234565,0.15090185,0.14404267,0.15090185,0.14747226,0.1097468,0.07888051,0.044584636,0.034295876,0.041155048,0.024007112,0.0274367,0.072021335,0.14747226,0.3018037,0.65505123,1.5604624,2.959734,4.0537724,4.1120753,2.4384367,1.4815818,1.5707511,2.8054025,4.2389703,3.865145,2.5790498,1.6290541,1.2072148,1.6016173,3.1792276,7.082098,9.832627,10.288762,8.587687,6.1458206,4.3795834,3.350707,3.5530527,4.712253,5.754848,5.6999745,5.638242,5.5902276,5.4804807,5.137522,4.4241676,6.560801,10.600855,14.743796,16.335125,9.002667,4.3692946,2.3424082,2.2258022,2.7230926,3.1072063,3.9371665,4.7499785,5.209543,5.099797,5.5250654,5.888602,6.1801167,6.3618846,6.3824625,5.9571934,5.65539,5.5593615,5.5319247,5.192395,4.8768735,4.681387,4.681387,4.911169,5.3673043,5.5490727,5.3913116,5.0757895,4.633373,3.9508848,3.223812,2.8225505,2.8911421,3.1209247,2.7470996,2.4452958,2.7642474,3.1586502,3.350707,3.309552,3.6044965,4.0674906,4.2218223,4.197815,4.7362604,5.0106273,4.9523244,4.822,4.557922,3.789694,2.8739944,2.4315774,1.9823016,1.4987297,1.3958421,1.3615463,1.3238207,1.5261664,1.8313997,1.7525192,2.5824795,3.2855449,3.2718265,2.7162333,2.5653315,0.9877212,0.37725464,0.20577525,0.17490897,0.2194936,0.12003556,0.09602845,0.072021335,0.0274367,0.017147938,0.0548734,0.034295876,0.034295876,0.06859175,0.07888051,0.041155048,0.034295876,0.034295876,0.041155048,0.05144381,0.06516216,0.07888051,0.09259886,0.106317215,0.116605975,0.14747226,0.14061308,0.12003556,0.10288762,0.09602845,0.12689474,0.15776102,0.1920569,0.23321195,0.28808534,0.41498008,0.90198153,1.3992717,1.5673214,1.0666018,0.9431366,0.922559,1.0494537,1.255229,1.3478279,1.4507155,1.5193073,1.5536032,1.5261664,1.3924125,1.9685832,2.9151495,2.983741,2.2052248,1.8725548,1.9582944,1.8725548,1.7182233,1.6221949,1.7662375,2.510458,2.5173173,2.6819375,3.1895163,3.5016088,4.7979927,3.758828,1.845118,0.3566771,0.4046913,0.8711152,0.64133286,0.45270553,0.5418748,0.6241849,0.3566771,0.25378948,0.33266997,0.4972902,0.5590228,0.274367,0.07888051,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.106317215,0.19891608,0.15776102,0.13032432,0.11317638,0.13375391,0.26064864,0.12346515,0.09602845,0.11317638,0.12003556,0.07888051,0.0548734,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.12003556,0.29837412,0.4698535,0.5796003,0.6310441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.09602845,0.20577525,0.50757897,0.8779744,0.8779744,0.72021335,0.3018037,0.058302987,0.058302987,0.006859175,0.0,0.0,0.0,0.0034295875,0.017147938,0.0548734,0.06516216,0.048014224,0.037725464,0.08573969,0.106317215,0.09259886,0.14404267,0.25378948,0.31895164,0.38754338,0.53158605,0.66533995,0.72021335,0.6344737,1.371835,3.3815732,4.2766957,3.357566,1.6221949,4.7088237,6.948344,9.115844,10.271614,7.7611566,4.647091,3.2409601,2.609916,2.1023371,1.3409687,0.8128122,0.4972902,0.45613512,0.6173257,0.7613684,0.864256,1.0666018,1.3821237,1.7319417,1.9480057,1.5501735,0.85739684,0.31895164,0.116605975,0.1371835,0.15090185,0.216064,0.33266997,0.48700142,0.65162164,0.7956643,0.7922347,0.7990939,0.8711152,0.9877212,1.0425946,0.8779744,0.6276145,0.39783216,0.26407823,0.1920569,0.13032432,0.10288762,0.09945804,0.0548734,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11317638,0.1920569,0.20920484,0.16462019,0.072021335,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.13032432,0.29151493,0.490431,0.6756287,0.66191036,0.61389613,0.51100856,0.36696586,0.24350071,0.22292319,0.24007112,0.28808534,0.34295875,0.37039545,0.39097297,0.42526886,0.53158605,0.66533995,0.6756287,0.7888051,1.0151579,1.1866373,1.3203912,1.6153357,2.1332035,1.9994495,1.6290541,1.3478279,1.3924125,1.6530612,1.5536032,1.5981878,1.9411465,2.386993,2.8877127,3.4055803,3.5770597,3.3644254,3.0214665,3.2683969,3.2786856,3.6285036,4.0091877,3.2409601,2.4247184,2.8122618,4.040054,4.835718,3.0351849,3.9337368,3.9680326,3.8034124,3.7451096,3.765687,3.6868064,3.8685746,3.7279615,3.175798,2.627064,2.633923,2.287535,1.8897027,1.6839274,1.879414,1.4438564,0.7990939,0.26407823,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.048014224,0.17833854,0.66876954,1.7113642,1.2277923,0.45613512,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.06516216,0.4115505,0.9877212,1.4164196,0.67219913,0.38754338,0.29151493,0.25721905,0.30523327,0.26750782,0.20920484,0.14061308,0.07888051,0.041155048,0.0548734,0.09945804,0.21263443,0.3566771,0.42183927,0.50757897,0.3806842,0.28465575,0.31209245,0.40126175,0.52815646,0.65505123,0.7099246,0.6824879,0.64476246,0.77508676,0.70649505,0.6173257,0.64476246,0.8848336,0.805953,0.71678376,0.58302987,0.4355576,0.36353627,0.25721905,0.24007112,0.2503599,0.23664154,0.15090185,0.14061308,0.1371835,0.19548649,0.26064864,0.16119061,0.09945804,0.11317638,0.12003556,0.08573969,0.024007112,0.030866288,0.07888051,0.13032432,0.18176813,0.25378948,0.4389872,1.0940384,1.9720128,2.7333813,2.952875,2.3458378,1.8828435,2.3252604,3.415869,3.8925817,2.860276,1.6667795,0.97057325,1.0734608,1.920569,3.8891523,5.346727,5.5730796,4.530485,2.8465576,2.218943,2.9631636,4.7774153,6.711703,7.1781263,5.796003,5.0003386,4.7774153,4.7499785,4.1772375,3.7279615,5.3707337,8.429926,11.588576,12.878101,8.186425,4.2081037,2.0646117,1.7147937,1.937717,2.1091962,2.7745364,3.4673128,3.8925817,3.9303071,4.15323,4.341858,4.3933015,4.3624353,4.4756117,4.125794,3.9440255,4.1429415,4.48933,4.2938433,3.8685746,3.4398763,3.199805,3.2409601,3.542764,3.4810312,3.724532,3.8925817,3.7794054,3.3541365,2.6887965,2.2600982,2.0989075,2.037175,1.704505,1.7182233,2.095478,2.603057,2.9631636,2.877424,2.3732746,2.2600982,2.177788,2.1434922,2.5447538,3.1277838,3.350707,3.532475,3.6868064,3.542764,2.5927682,1.8416885,1.371835,1.1832076,1.1934965,1.0940384,1.0940384,1.3066728,1.646202,1.8416885,2.5207467,3.2615378,3.4947495,3.1826572,2.8225505,1.3855534,0.5693115,0.20920484,0.13032432,0.13375391,0.08916927,0.08573969,0.06859175,0.041155048,0.05144381,0.058302987,0.05144381,0.041155048,0.041155048,0.07545093,0.061732575,0.037725464,0.024007112,0.034295876,0.044584636,0.058302987,0.06516216,0.072021335,0.082310095,0.07888051,0.1097468,0.11317638,0.09602845,0.06859175,0.06516216,0.08573969,0.12003556,0.15433143,0.18519773,0.21263443,0.28808534,0.5007198,0.85739684,1.1180456,0.7956643,0.86082643,1.1626302,1.3958421,1.4232788,1.2723769,1.3512574,1.2758065,1.1420527,1.0494537,1.1180456,1.7559488,2.3149714,2.1194851,1.4164196,1.3821237,1.6393428,1.6907866,1.5193073,1.3306799,1.5433143,2.136633,2.1880767,2.3252604,2.633923,2.6647894,2.8637056,2.287535,1.1660597,0.10288762,0.072021335,0.25721905,0.17833854,0.16804978,0.30523327,0.39440256,0.26407823,0.216064,0.274367,0.37382504,0.38754338,0.22292319,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.12689474,0.14404267,0.15433143,0.15433143,0.15433143,0.19891608,0.13032432,0.13032432,0.14747226,0.14747226,0.12346515,0.116605975,0.08573969,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.10288762,0.14747226,0.17147937,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.106317215,0.20577525,0.4664239,0.764798,0.6824879,0.64133286,0.25721905,0.020577524,0.037725464,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.1371835,0.4355576,0.38754338,0.058302987,0.07888051,0.1097468,0.09602845,0.12346515,0.2503599,0.5041494,0.47328308,0.61389613,0.97057325,1.2277923,0.70306545,1.7216529,2.6476414,2.5173173,1.903421,2.884283,6.108095,7.9875093,7.2878733,4.5510626,2.1160555,1.728512,1.3238207,0.7990939,0.28465575,0.1371835,0.06516216,0.017147938,0.106317215,0.29837412,0.42183927,0.4664239,0.51100856,0.7442205,1.1626302,1.5673214,1.3306799,0.71678376,0.26750782,0.16119061,0.22292319,0.26750782,0.32924038,0.4081209,0.5144381,0.65848076,0.7373613,0.7305021,0.7133542,0.7442205,0.86082643,0.94999576,0.84367853,0.6276145,0.39783216,0.26407823,0.1920569,0.13032432,0.10288762,0.09945804,0.0548734,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08916927,0.16119061,0.18176813,0.14747226,0.09259886,0.037725464,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.12689474,0.2709374,0.42526886,0.5144381,0.5521636,0.5178677,0.42526886,0.32238123,0.2777966,0.26407823,0.28122616,0.31209245,0.33952916,0.33952916,0.3566771,0.42526886,0.53501564,0.6310441,0.77165717,0.9294182,1.1111864,1.2998136,1.4610043,1.5810398,1.5330256,1.3478279,1.1489118,1.1283343,1.1694894,1.2175035,1.3341095,1.5604624,1.9239986,2.4452958,2.9494452,3.1209247,3.0214665,3.093488,3.1655092,2.935727,3.0111778,3.1483612,2.2326615,1.8897027,2.6304936,3.6868064,4.0434837,2.4144297,3.666229,3.7691166,3.799983,4.1360826,4.448175,3.7485392,3.3541365,3.1723683,3.0420442,2.74367,1.9239986,1.4610043,1.3821237,1.546744,1.6530612,0.9945804,0.4972902,0.16462019,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.0274367,0.048014224,0.48700142,2.218943,2.603057,1.4027013,0.34981793,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.05144381,0.38754338,1.1180456,2.201795,1.2655178,0.8848336,0.548734,0.21263443,0.28808534,0.30523327,0.26750782,0.22635277,0.17490897,0.034295876,0.020577524,0.017147938,0.037725464,0.11317638,0.30523327,0.4115505,0.37725464,0.33952916,0.34638834,0.3806842,0.4664239,0.6310441,0.7682276,0.83681935,0.8745448,0.85739684,0.8025235,0.7373613,0.69963586,0.7682276,0.77508676,0.6893471,0.5418748,0.4046913,0.39440256,0.31209245,0.29151493,0.2777966,0.23664154,0.13375391,0.16462019,0.15776102,0.20920484,0.29151493,0.24007112,0.20577525,0.216064,0.18176813,0.09945804,0.041155048,0.06516216,0.15433143,0.2777966,0.3566771,0.28465575,0.2194936,0.45613512,0.8711152,1.4575747,2.3081124,2.294394,1.9171394,1.8485477,2.3835633,3.4638834,2.7813954,1.5981878,0.8162418,0.7510797,1.1146159,2.0406046,3.0420442,3.357566,2.7745364,1.6324836,1.5398848,3.199805,5.7239814,7.6857057,7.116394,4.8117113,3.5873485,3.1312134,2.983741,2.5310357,2.4795918,3.3884325,4.9214582,6.540223,7.507367,5.809721,3.3026927,1.7250825,1.471293,1.6084765,1.6359133,1.9857311,2.3629858,2.603057,2.668219,2.8259802,2.959734,2.983741,2.9700227,3.1483612,3.0043187,2.935727,3.1826572,3.5599117,3.4878905,3.0386145,2.6304936,2.386993,2.311542,2.2909644,2.0131679,2.270387,2.5961976,2.7333813,2.627064,2.335549,2.037175,1.7456601,1.4610043,1.1797781,1.255229,1.4781522,1.8073926,2.1091962,2.1640697,1.5158776,1.1626302,0.9774324,0.922559,1.0323058,1.4953002,1.7765263,1.9754424,2.177788,2.4384367,1.9857311,1.3992717,1.0254467,0.94999576,1.0048691,0.864256,0.823101,0.922559,1.1626302,1.5330256,1.9651536,2.620205,2.9974594,2.8877127,2.369845,1.6427724,1.6221949,1.6496316,1.3409687,0.58645946,0.22978236,0.12346515,0.14061308,0.17147937,0.11317638,0.072021335,0.058302987,0.041155048,0.020577524,0.044584636,0.044584636,0.0274367,0.020577524,0.0274367,0.034295876,0.044584636,0.05144381,0.058302987,0.06516216,0.061732575,0.07545093,0.082310095,0.06859175,0.044584636,0.044584636,0.058302987,0.09259886,0.12689474,0.14404267,0.15776102,0.216064,0.4115505,0.77165717,1.08032,0.88826317,1.0768905,1.3615463,1.605047,1.6667795,1.4198492,1.4198492,1.1729189,0.89169276,0.7956643,1.097468,1.3512574,1.3855534,1.2963841,1.1832076,1.1694894,1.3032433,1.2929544,1.08032,0.83338976,0.939707,1.3786942,1.5981878,1.7490896,1.7662375,1.3752645,0.9328478,0.83338976,0.5041494,0.006859175,0.037725464,0.12346515,0.058302987,0.024007112,0.08573969,0.17490897,0.17147937,0.18176813,0.22978236,0.28465575,0.28465575,0.19891608,0.10288762,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0548734,0.12003556,0.16804978,0.19891608,0.20234565,0.17490897,0.15776102,0.15776102,0.16119061,0.16119061,0.15776102,0.16804978,0.14404267,0.08573969,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.01371835,0.0034295875,0.020577524,0.058302987,0.020577524,0.030866288,0.06516216,0.082310095,0.024007112,0.0548734,0.13032432,0.13375391,0.058302987,0.030866288,0.29494452,1.3238207,1.4027013,0.45270553,0.01371835,0.044584636,0.08573969,0.17833854,0.4046913,0.90541106,0.66533995,0.77165717,1.2517995,1.4850113,0.20577525,0.91569984,1.3238207,1.6290541,2.5927682,5.504488,6.3035817,6.5127864,4.07435,0.35324752,0.15433143,0.4115505,0.40126175,0.21263443,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.082310095,0.16119061,0.31895164,0.5727411,0.53501564,0.31895164,0.1920569,0.23664154,0.34638834,0.4081209,0.42526886,0.37382504,0.28122616,0.21263443,0.18862732,0.14404267,0.07888051,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058302987,0.106317215,0.14404267,0.23321195,0.116605975,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.08573969,0.17490897,0.28465575,0.37039545,0.41498008,0.41840968,0.3841138,0.34638834,0.33266997,0.33266997,0.33952916,0.34981793,0.3566771,0.38754338,0.45956472,0.5761707,0.70649505,0.8779744,0.9911508,1.0425946,1.0563129,1.0837497,1.0323058,1.08032,1.1214751,1.1317638,1.1592005,1.1832076,1.2072148,1.3203912,1.5193073,1.7182233,1.9823016,2.136633,2.335549,2.726522,3.4776018,3.8102717,3.4227283,3.0797696,3.000889,2.8396983,2.2463799,2.486451,2.270387,1.6187652,1.8862731,3.4227283,3.292404,3.210094,3.7622573,4.40702,3.673088,3.357566,3.100347,2.726522,2.2292318,1.6084765,1.2998136,1.2243627,1.2346514,1.1351935,0.45270553,0.11317638,0.0,0.0,0.0,0.0,0.0,0.037725464,0.07888051,0.020577524,0.0034295875,0.18176813,0.4629943,1.3409687,3.899441,3.000889,1.2277923,0.14747226,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.19891608,0.75450927,2.0097382,1.5193073,1.2758065,0.8505377,0.31209245,0.24350071,0.22292319,0.21263443,0.26064864,0.29151493,0.09602845,0.044584636,0.020577524,0.044584636,0.106317215,0.19891608,0.2777966,0.4424168,0.50757897,0.45270553,0.4424168,0.37039545,0.58645946,0.8265306,0.9774324,1.0871792,1.0254467,0.9294182,0.864256,0.7888051,0.5624523,0.5555932,0.48014224,0.44927597,0.4698535,0.47328308,0.42183927,0.39440256,0.33266997,0.23664154,0.16119061,0.20577525,0.20234565,0.20577525,0.24007112,0.31209245,0.33952916,0.29837412,0.18862732,0.06859175,0.058302987,0.1097468,0.26750782,0.48357183,0.6207553,0.45613512,0.34295875,0.58302987,0.7888051,0.8848336,1.1111864,1.3684053,1.3546871,1.214074,1.4164196,2.767677,2.5173173,1.5673214,0.864256,0.7407909,0.90541106,1.371835,2.037175,2.2978237,1.978872,1.3409687,1.3958421,3.0489032,5.1512403,6.341307,5.0277753,2.8465576,1.5364552,0.89855194,0.7613684,0.9602845,1.0494537,1.3443983,1.7353712,2.2909644,3.2581081,2.9254382,1.9445761,1.3238207,1.3306799,1.4850113,1.4610043,1.5261664,1.646202,1.7765263,1.8759843,1.8828435,1.9548649,2.0337453,2.0680413,1.99602,1.9651536,2.0063086,2.0680413,2.1332035,2.2292318,2.037175,1.7388009,1.5536032,1.4815818,1.2758065,1.0494537,1.1180456,1.3409687,1.5673214,1.6359133,1.7902447,1.7902447,1.6633499,1.4541451,1.2586586,1.155771,1.1934965,1.2689474,1.3272504,1.3786942,1.0563129,0.8779744,0.7339317,0.6001778,0.53158605,0.5521636,0.6859175,0.71678376,0.6824879,0.881404,1.1111864,1.0323058,0.8265306,0.66876954,0.72364295,0.65162164,0.5624523,0.5212973,0.6173257,0.96714365,1.4027013,1.9651536,2.2429502,2.1023371,1.6976458,1.6564908,2.901431,3.782835,3.4364467,1.7765263,0.8711152,0.4664239,0.35324752,0.33266997,0.20920484,0.12689474,0.072021335,0.037725464,0.020577524,0.006859175,0.0034295875,0.01371835,0.017147938,0.017147938,0.017147938,0.030866288,0.041155048,0.044584636,0.044584636,0.058302987,0.058302987,0.048014224,0.041155048,0.044584636,0.048014224,0.06516216,0.09259886,0.11317638,0.12003556,0.12346515,0.15090185,0.52472687,1.0494537,1.4164196,1.2003556,1.1934965,1.2243627,1.4335675,1.6839274,1.5398848,1.5570327,1.2620882,0.97400284,0.9259886,1.2655178,0.96714365,0.823101,0.8745448,1.039165,1.1146159,0.8848336,0.6207553,0.41498008,0.28465575,0.18176813,0.41840968,0.7990939,0.91227025,0.64819205,0.20920484,0.13032432,0.072021335,0.030866288,0.0,0.0,0.0,0.0,0.0,0.020577524,0.10288762,0.16119061,0.20234565,0.23664154,0.26750782,0.274367,0.22978236,0.17490897,0.09259886,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06859175,0.13375391,0.19891608,0.2469303,0.216064,0.19891608,0.17833854,0.16462019,0.16462019,0.17147937,0.18176813,0.16462019,0.116605975,0.0548734,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0034295875,0.0034295875,0.01371835,0.06516216,0.01371835,0.0,0.0,0.0034295875,0.0,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.048014224,0.12003556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.030866288,0.01371835,0.0,0.010288762,0.044584636,0.044584636,0.1097468,0.28808534,0.41498008,0.12346515,0.28122616,0.65848076,0.66533995,0.29837412,0.15090185,0.64133286,2.9048605,3.625074,2.0508933,0.0,0.01371835,0.116605975,0.40126175,0.7956643,1.0528834,0.6756287,1.1214751,1.5227368,1.2792361,0.044584636,0.29151493,1.0117283,2.9151495,5.7479887,8.299602,9.119273,8.097256,4.5613513,0.40126175,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.16119061,0.31895164,0.39440256,0.42183927,0.4081209,0.37382504,0.33609957,0.31209245,0.2503599,0.17147937,0.08573969,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.24350071,0.20920484,0.07888051,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.041155048,0.072021335,0.12689474,0.21263443,0.33609957,0.39783216,0.44927597,0.47328308,0.47328308,0.47328308,0.5453044,0.6001778,0.6310441,0.67219913,0.7922347,1.0631721,1.0014396,0.7922347,0.64476246,0.77851635,0.864256,0.9294182,0.9911508,1.0494537,1.097468,1.1592005,1.2380811,1.3375391,1.4610043,1.6324836,1.5364552,1.4472859,1.4541451,1.587899,1.8313997,2.270387,2.3252604,2.8122618,4.0366244,5.7822843,3.8308492,2.3629858,1.7147937,1.9342873,2.7779658,5.0483527,4.2046742,2.959734,2.6373527,3.1723683,4.0880685,4.245829,3.5564823,2.4247184,1.7559488,1.5707511,1.5364552,1.3958421,1.039165,0.48700142,0.15776102,0.030866288,0.0,0.0,0.0,0.0,0.0,0.18862732,0.38754338,0.044584636,0.010288762,0.90541106,2.311542,3.6079261,3.998899,2.6167753,1.5055889,0.6379033,0.08573969,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.10288762,0.274367,0.4698535,0.6824879,0.939707,1.039165,0.548734,0.20920484,0.12346515,0.17147937,0.24007112,0.22978236,0.12003556,0.082310095,0.09602845,0.16119061,0.31895164,0.31895164,0.7613684,0.881404,0.6756287,0.8711152,0.7476501,1.0185875,1.1900668,1.2209331,1.5261664,1.1214751,1.3169615,1.546744,1.4027013,0.61046654,0.5727411,0.5007198,0.45613512,0.47328308,0.53501564,0.5693115,0.5796003,0.4698535,0.28465575,0.19891608,0.17490897,0.20577525,0.24007112,0.274367,0.33609957,0.32238123,0.26407823,0.15433143,0.044584636,0.044584636,0.15433143,0.29151493,0.44584638,0.5796003,0.64133286,0.4081209,0.33266997,0.38754338,0.548734,0.7922347,0.805953,0.64476246,0.5041494,0.764798,1.9994495,2.452155,1.7216529,1.0185875,0.881404,1.1763484,1.4918705,1.7182233,1.8519772,1.8897027,1.8142518,2.1469216,3.316411,3.8960114,3.4776018,2.6716487,2.8054025,1.978872,0.97057325,0.31552204,0.29151493,0.33952916,0.432128,0.58645946,0.805953,1.097468,1.4781522,1.5158776,1.4987297,1.5227368,1.5090185,1.2312219,1.0940384,1.2312219,1.546744,1.7559488,1.4507155,1.3821237,1.4438564,1.4575747,1.1900668,1.0425946,1.097468,1.0323058,0.8471081,0.8848336,1.0563129,0.97057325,0.8848336,0.86082643,0.7613684,0.66533995,0.7407909,0.77851635,0.72021335,0.67219913,0.85396725,0.97400284,1.0837497,1.1729189,1.1592005,1.1489118,1.2346514,1.4815818,1.7319417,1.6496316,1.0014396,0.7579388,0.6824879,0.64133286,0.5796003,0.432128,0.39783216,0.45270553,0.58988905,0.8093826,0.980862,0.96714365,0.7956643,0.5658819,0.4424168,0.3806842,0.33952916,0.3018037,0.3566771,0.6859175,1.2963841,1.7799559,1.920569,1.7456601,1.5261664,1.4164196,2.3972816,3.6353626,4.266407,3.3884325,2.435007,1.5193073,0.7339317,0.26064864,0.3806842,0.30866286,0.18862732,0.09602845,0.0548734,0.030866288,0.017147938,0.024007112,0.024007112,0.017147938,0.030866288,0.041155048,0.044584636,0.041155048,0.034295876,0.044584636,0.044584636,0.037725464,0.030866288,0.037725464,0.061732575,0.08573969,0.09945804,0.106317215,0.1097468,0.12346515,0.12346515,0.19548649,0.548734,0.980862,0.8711152,0.7956643,1.0082988,1.1283343,1.1249046,1.2963841,1.6633499,1.471293,1.2517995,1.2415106,1.3889829,1.1694894,1.0597426,1.1694894,1.371835,1.2963841,0.78537554,0.40126175,0.2469303,0.24350071,0.12346515,0.12346515,0.20577525,0.22978236,0.14747226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.15090185,0.2503599,0.29151493,0.29837412,0.28808534,0.274367,0.2503599,0.19891608,0.13032432,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.12346515,0.16804978,0.16804978,0.22978236,0.23664154,0.216064,0.19548649,0.18176813,0.14747226,0.1371835,0.12003556,0.072021335,0.0,0.0,0.0,0.024007112,0.048014224,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.0,0.01371835,0.006859175,0.006859175,0.024007112,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.24007112,0.59674823,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.16462019,0.36010668,0.39097297,0.37382504,0.31895164,0.13032432,0.044584636,0.39440256,0.75450927,0.805953,0.31895164,0.29151493,0.35324752,0.29494452,0.1371835,0.12689474,0.16804978,0.90541106,1.2517995,0.89169276,0.30523327,0.51100856,1.5570327,2.9254382,3.683377,2.5070283,1.0220171,0.70306545,0.7305021,0.6379033,0.3018037,1.1317638,2.2326615,6.012067,10.816919,10.9369545,6.392751,3.5702004,1.605047,0.274367,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.06516216,0.22292319,0.18862732,0.18176813,0.18862732,0.21263443,0.274367,0.2503599,0.18862732,0.09945804,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.06859175,0.09945804,0.1097468,0.07888051,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.041155048,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.14747226,0.32924038,0.33609957,0.18519773,0.1371835,0.034295876,0.01371835,0.030866288,0.06859175,0.15090185,0.32238123,0.48014224,0.61046654,0.70649505,0.764798,0.7990939,0.8025235,0.8162418,0.86082643,0.90198153,0.8093826,0.67219913,0.59674823,0.6344737,0.77851635,0.84367853,0.89169276,0.9568549,1.0494537,1.1489118,1.2003556,1.2037852,1.2415106,1.2963841,1.2415106,1.2037852,1.2243627,1.2586586,1.2792361,1.2689474,1.5124481,1.7833855,2.6922262,3.7142432,3.1963756,3.0969174,3.3472774,3.3472774,3.083199,3.1072063,4.4413157,3.8685746,3.858286,4.8151407,5.0895076,3.7691166,2.8156912,2.0646117,1.5090185,1.3169615,1.6016173,1.8862731,1.7250825,1.08032,0.30523327,0.072021335,0.006859175,0.0,0.0,0.0,0.09602845,0.048014224,0.2194936,0.4389872,0.010288762,0.7339317,1.937717,2.668219,2.7230926,2.6545007,2.6716487,1.5330256,0.5144381,0.106317215,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.020577524,0.024007112,0.07888051,0.17833854,0.58645946,1.5055889,2.4007113,2.0028791,0.5178677,0.14061308,0.216064,0.39783216,0.6207553,0.64476246,0.5693115,0.42526886,0.274367,0.19891608,0.30523327,0.58988905,0.9602845,1.2963841,1.4438564,1.2929544,1.1249046,1.0357354,1.0837497,1.2826657,1.5055889,1.8005334,1.9068506,1.6907866,1.1729189,0.91227025,0.8025235,0.8128122,0.8505377,0.75450927,0.65505123,0.72364295,0.7442205,0.6859175,0.69963586,0.490431,0.32581082,0.28122616,0.33266997,0.3841138,0.35324752,0.26064864,0.19891608,0.17833854,0.12003556,0.24007112,0.37725464,0.42869842,0.4389872,0.6276145,0.7682276,0.548734,0.39097297,0.45270553,0.64819205,0.66876954,0.40126175,0.19548649,0.2469303,0.58302987,0.88826317,0.8676856,0.7133542,0.5555932,0.48014224,0.9431366,0.8848336,0.7922347,0.96714365,1.4987297,1.6221949,2.0337453,2.627064,2.8980014,1.9239986,2.469303,1.3924125,0.4389872,0.22978236,0.25378948,0.274367,0.35324752,0.5144381,0.7510797,1.0117283,1.08032,1.0906088,1.0700313,1.0528834,1.1214751,1.0837497,0.83338976,0.72021335,0.8676856,1.1797781,1.1008976,0.94999576,0.86082643,0.823101,0.6893471,0.5041494,0.4698535,0.4081209,0.30523327,0.31209245,0.47328308,0.5590228,0.5590228,0.490431,0.42183927,0.34295875,0.3566771,0.40126175,0.42526886,0.41498008,0.432128,0.42183927,0.41840968,0.432128,0.4389872,0.5555932,0.7990939,1.4061309,2.201795,2.6236343,1.937717,1.4061309,1.1077567,0.9911508,0.8711152,0.66876954,0.61046654,0.7956643,1.0700313,1.0151579,0.96371406,0.85739684,0.6859175,0.5144381,0.490431,0.45956472,0.41840968,0.3806842,0.37725464,0.4424168,1.0906088,2.527606,3.0111778,2.287535,1.5981878,1.8005334,2.5070283,2.7951138,2.5001693,2.2292318,2.5447538,2.0714707,1.3615463,0.8025235,0.61389613,0.47328308,0.4972902,0.45270553,0.31209245,0.2503599,0.33609957,0.548734,0.53844523,0.28122616,0.06859175,0.07888051,0.061732575,0.048014224,0.0548734,0.058302987,0.048014224,0.05144381,0.0548734,0.0548734,0.061732575,0.08573969,0.116605975,0.12689474,0.12003556,0.12346515,0.12346515,0.12346515,0.22292319,0.4389872,0.69963586,0.9774324,1.3649758,1.7250825,1.9445761,1.920569,2.177788,2.0028791,1.9137098,1.9480057,1.646202,1.2380811,0.9945804,1.0323058,1.196926,1.0666018,0.6310441,0.32581082,0.16804978,0.11317638,0.048014224,0.058302987,0.061732575,0.05144381,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.35324752,0.53844523,0.59331864,0.5590228,0.50757897,0.34638834,0.20920484,0.09259886,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.044584636,0.09602845,0.14747226,0.15090185,0.1371835,0.13032432,0.14747226,0.13032432,0.116605975,0.10288762,0.072021335,0.0,0.0,0.0,0.024007112,0.058302987,0.048014224,0.010288762,0.0034295875,0.0034295875,0.006859175,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.01371835,0.0034295875,0.030866288,0.030866288,0.01371835,0.061732575,0.01371835,0.030866288,0.048014224,0.048014224,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.037725464,0.020577524,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.6310441,1.6084765,1.8142518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.07888051,0.17833854,0.23321195,0.26407823,0.26064864,0.16119061,0.05144381,0.22635277,0.4355576,0.50757897,0.31895164,0.91227025,0.72707254,0.36010668,0.13375391,0.08573969,0.0274367,0.83338976,1.0528834,0.48357183,0.15090185,0.37382504,3.192946,5.4633327,5.576509,3.474172,2.5790498,1.8656956,1.5261664,1.6907866,2.4075704,3.6765177,4.434457,5.5662203,6.7494283,6.444195,2.983741,1.1454822,0.34638834,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.07888051,0.0548734,0.048014224,0.0548734,0.06859175,0.10288762,0.09259886,0.06859175,0.034295876,0.010288762,0.044584636,0.06859175,0.072021335,0.06859175,0.058302987,0.037725464,0.006859175,0.01371835,0.034295876,0.05144381,0.0548734,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.01371835,0.06516216,0.3806842,0.7888051,1.0597426,0.9568549,0.2503599,0.05144381,0.0,0.006859175,0.030866288,0.08916927,0.26750782,0.45613512,0.6036074,0.70649505,0.7922347,0.89169276,0.91227025,0.8848336,0.83338976,0.78537554,0.6756287,0.59674823,0.5761707,0.6241849,0.7407909,0.8471081,0.9294182,1.0151579,1.1077567,1.1489118,1.2517995,1.3203912,1.3169615,1.2175035,0.99801,0.980862,1.097468,1.1797781,1.1626302,1.0837497,1.2346514,1.6530612,2.1743584,2.4041407,1.704505,2.4761622,3.2409601,4.108646,4.8734436,5.020916,4.8940215,4.4550343,4.3590055,4.4275975,3.6456516,2.3389788,1.4987297,1.0151579,0.805953,0.8128122,1.039165,1.2277923,1.1351935,0.70649505,0.10288762,0.05144381,0.01371835,0.01371835,0.041155048,0.0548734,0.32238123,0.15776102,0.106317215,0.37382504,0.8162418,1.4232788,2.194936,2.5413244,2.1434922,0.9294182,1.0734608,0.7305021,0.37039545,0.16804978,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.034295876,0.06516216,0.07545093,0.037725464,0.006859175,0.0034295875,0.020577524,0.06516216,0.29151493,0.8025235,1.3341095,1.2586586,0.4389872,0.14404267,0.13375391,0.2469303,0.39783216,0.4938606,0.6173257,0.59331864,0.45613512,0.42526886,0.48357183,0.6241849,0.78537554,0.939707,1.0734608,1.1043272,1.1489118,1.3066728,1.4918705,1.4507155,1.6153357,1.7593783,1.8005334,1.6359133,1.155771,0.9431366,0.82996017,0.7922347,0.77851635,0.71678376,0.70649505,0.8025235,0.8779744,0.88826317,0.8505377,0.6036074,0.41498008,0.31552204,0.29151493,0.30523327,0.274367,0.25378948,0.26407823,0.28465575,0.2469303,0.33266997,0.5178677,0.64133286,0.6824879,0.77165717,0.77851635,0.548734,0.39783216,0.4389872,0.59331864,0.58645946,0.33266997,0.12689474,0.08573969,0.1371835,0.25378948,0.31895164,0.32238123,0.30866286,0.38754338,0.64476246,0.4938606,0.34638834,0.432128,0.77851635,0.764798,0.8505377,1.1523414,1.4541451,1.2072148,1.2929544,0.67219913,0.20234565,0.14404267,0.15090185,0.17833854,0.26064864,0.4046913,0.58645946,0.72707254,0.6927767,0.64819205,0.5727411,0.5007198,0.52815646,0.5453044,0.41840968,0.33266997,0.3806842,0.5624523,0.64819205,0.6962063,0.6379033,0.48700142,0.34638834,0.23664154,0.21263443,0.24007112,0.2469303,0.13032432,0.17147937,0.2194936,0.23664154,0.22635277,0.216064,0.18176813,0.16804978,0.16119061,0.18519773,0.29494452,0.23664154,0.19891608,0.16804978,0.14404267,0.14061308,0.20577525,0.31552204,0.6379033,1.3101025,2.428148,2.3767042,2.0406046,1.6187652,1.2895249,1.1832076,0.94999576,0.9362774,1.0906088,1.2792361,1.2895249,1.2655178,0.97400284,0.6962063,0.548734,0.47671264,0.48014224,0.44584638,0.39783216,0.36010668,0.34638834,0.7476501,1.5776103,2.0028791,1.8725548,1.728512,1.5776103,2.0337453,2.3664153,2.277246,1.920569,2.0989075,1.821111,1.4369972,1.1351935,0.94656616,0.53158605,0.41840968,0.3841138,0.37725464,0.5144381,0.764798,0.88826317,0.84024894,0.6310441,0.33266997,0.2194936,0.15776102,0.116605975,0.08573969,0.06859175,0.05144381,0.048014224,0.0548734,0.058302987,0.05144381,0.07545093,0.09945804,0.106317215,0.106317215,0.11317638,0.11317638,0.08916927,0.13375391,0.32581082,0.7305021,1.2655178,1.6324836,1.8073926,1.8073926,1.6907866,1.9514352,2.0508933,2.16064,2.1469216,1.5638919,1.0288762,0.67219913,0.5555932,0.58645946,0.5212973,0.29837412,0.17490897,0.106317215,0.06859175,0.048014224,0.030866288,0.020577524,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.09945804,0.19548649,0.31895164,0.6756287,0.8848336,0.881404,0.7442205,0.6756287,0.4424168,0.25721905,0.12689474,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.058302987,0.08573969,0.10288762,0.10288762,0.09259886,0.1097468,0.11317638,0.09259886,0.061732575,0.030866288,0.0,0.0,0.0,0.010288762,0.024007112,0.024007112,0.034295876,0.020577524,0.010288762,0.006859175,0.006859175,0.0,0.0,0.010288762,0.030866288,0.05144381,0.041155048,0.05144381,0.037725464,0.0034295875,0.024007112,0.034295876,0.061732575,0.082310095,0.08573969,0.06859175,0.044584636,0.037725464,0.020577524,0.0,0.0,0.020577524,0.010288762,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.31552204,0.8676856,1.2072148,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.18519773,0.3841138,0.44927597,0.7888051,1.6770682,1.7833855,1.2860953,1.8999915,2.6304936,1.9342873,1.1317638,0.7407909,0.45613512,0.31552204,1.1934965,1.3341095,0.6310441,0.6207553,1.2655178,4.108646,5.56965,4.633373,2.843128,3.3609958,2.877424,2.2086544,2.1469216,3.450165,4.32128,4.273266,3.340418,2.1229146,1.8039631,0.6962063,0.16804978,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.06859175,0.072021335,0.08916927,0.106317215,0.08573969,0.041155048,0.0274367,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.061732575,0.041155048,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06859175,0.33952916,0.6790583,0.9294182,0.864256,0.18176813,0.037725464,0.0,0.0034295875,0.020577524,0.06516216,0.19548649,0.31209245,0.39097297,0.4424168,0.53158605,0.6824879,0.75450927,0.7305021,0.6379033,0.5693115,0.5624523,0.5658819,0.5658819,0.5796003,0.66191036,0.78194594,0.8779744,0.9945804,1.1249046,1.2243627,1.3581166,1.3992717,1.2860953,1.0288762,0.71678376,0.7682276,0.91227025,1.0288762,1.0597426,1.0117283,1.1523414,1.587899,1.786815,1.5570327,1.039165,1.862266,2.6785078,4.0023284,5.5902276,6.39961,5.5422134,4.8185706,4.108646,3.216953,1.8828435,1.1111864,0.65505123,0.4424168,0.39440256,0.42183927,0.47671264,0.51100856,0.44927597,0.2709374,0.0,0.030866288,0.048014224,0.048014224,0.048014224,0.09259886,0.36010668,0.274367,0.42183927,1.0117283,1.8519772,2.0406046,2.5413244,2.6819375,2.0234566,0.35324752,0.16462019,0.22978236,0.30523327,0.26407823,0.10288762,0.058302987,0.0548734,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.010288762,0.0274367,0.058302987,0.082310095,0.07888051,0.030866288,0.0,0.0034295875,0.01371835,0.030866288,0.07545093,0.16119061,0.2709374,0.34638834,0.22292319,0.09602845,0.058302987,0.11317638,0.18862732,0.28808534,0.5007198,0.6207553,0.6173257,0.6207553,0.64476246,0.72707254,0.65848076,0.5178677,0.6790583,0.939707,1.2860953,1.605047,1.7250825,1.4267083,1.5090185,1.7765263,1.8656956,1.6427724,1.2003556,0.9877212,0.881404,0.8505377,0.8196714,0.66191036,0.6824879,0.7133542,0.7442205,0.7579388,0.7339317,0.548734,0.4081209,0.31209245,0.25721905,0.2503599,0.32924038,0.34638834,0.3566771,0.37039545,0.36353627,0.4081209,0.6276145,0.823101,0.91569984,0.9294182,0.6927767,0.5212973,0.48357183,0.5418748,0.5555932,0.47328308,0.28465575,0.12346515,0.058302987,0.06516216,0.07545093,0.09259886,0.2503599,0.4938606,0.5693115,0.6276145,0.5590228,0.40126175,0.26064864,0.28465575,0.26064864,0.32581082,0.42869842,0.5212973,0.5796003,0.42526886,0.24007112,0.14404267,0.13375391,0.12346515,0.18176813,0.22635277,0.29494452,0.3841138,0.45270553,0.34981793,0.2709374,0.19548649,0.13375391,0.12346515,0.13375391,0.116605975,0.10288762,0.11317638,0.17147937,0.28465575,0.42183927,0.41840968,0.2709374,0.15090185,0.09945804,0.08916927,0.14061308,0.18519773,0.07545093,0.0548734,0.044584636,0.05144381,0.06859175,0.082310095,0.07888051,0.06516216,0.041155048,0.05144381,0.16119061,0.106317215,0.08916927,0.07545093,0.048014224,0.037725464,0.044584636,0.041155048,0.08573969,0.39097297,1.2998136,1.6393428,2.1160555,2.3767042,2.3321195,2.16064,1.7593783,1.5124481,1.3992717,1.4164196,1.5570327,1.5604624,1.1797781,0.823101,0.64133286,0.5418748,0.5590228,0.53501564,0.48014224,0.4046913,0.3566771,0.4972902,0.6824879,0.90198153,1.1214751,1.2826657,1.0906088,1.4438564,1.9651536,2.2566686,1.920569,1.7490896,1.5501735,1.3272504,1.1283343,1.0666018,0.6962063,0.4938606,0.40126175,0.40126175,0.5212973,0.6790583,0.69963586,0.66533995,0.58645946,0.4046913,0.26750782,0.20577525,0.15433143,0.09945804,0.07545093,0.05144381,0.044584636,0.048014224,0.044584636,0.034295876,0.048014224,0.058302987,0.06516216,0.07545093,0.08916927,0.07545093,0.058302987,0.106317215,0.274367,0.59674823,1.1283343,1.4438564,1.5707511,1.5570327,1.4644338,1.7250825,1.903421,1.9720128,1.8142518,1.2277923,0.7339317,0.4046913,0.24350071,0.19891608,0.16119061,0.07545093,0.0548734,0.048014224,0.037725464,0.037725464,0.020577524,0.01371835,0.024007112,0.037725464,0.030866288,0.030866288,0.030866288,0.037725464,0.0548734,0.07888051,0.10288762,0.20234565,0.30523327,0.42869842,0.6756287,0.89855194,1.0357354,0.9842916,0.7922347,0.65162164,0.42183927,0.25378948,0.13032432,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.034295876,0.05144381,0.06859175,0.072021335,0.0548734,0.061732575,0.061732575,0.048014224,0.030866288,0.024007112,0.0034295875,0.0,0.0,0.0034295875,0.024007112,0.037725464,0.0274367,0.01371835,0.01371835,0.0,0.0034295875,0.0034295875,0.006859175,0.024007112,0.05144381,0.041155048,0.037725464,0.020577524,0.0,0.006859175,0.030866288,0.05144381,0.06516216,0.06516216,0.05144381,0.041155048,0.041155048,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.08573969,0.36353627,0.024007112,0.020577524,0.010288762,0.0034295875,0.0034295875,0.0,0.0,0.0,0.006859175,0.0274367,0.044584636,0.061732575,0.05144381,0.034295876,0.020577524,0.024007112,0.01371835,0.0034295875,0.216064,0.5693115,0.69963586,1.5124481,3.2786856,3.3952916,2.301253,3.4844608,3.7313912,2.7951138,2.020027,1.8554068,1.8382589,1.5158776,1.6496316,1.611906,1.471293,1.99602,2.8568463,3.858286,3.5221863,2.0577524,1.371835,2.7711067,2.7368107,1.9514352,1.4575747,2.668219,2.6956558,2.061182,1.2998136,0.64819205,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.09602845,0.09602845,0.06859175,0.0548734,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08916927,0.14747226,0.10288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.072021335,0.106317215,0.072021335,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.09602845,0.10288762,0.08916927,0.08916927,0.14747226,0.2777966,0.40126175,0.42869842,0.37382504,0.3806842,0.490431,0.5144381,0.50757897,0.50757897,0.5418748,0.65162164,0.764798,0.9259886,1.1420527,1.3581166,1.4644338,1.3821237,1.1111864,0.7339317,0.40126175,0.5453044,0.67219913,0.84024894,0.9945804,0.96371406,1.08032,1.3786942,1.5227368,1.3409687,0.83338976,1.2758065,1.9582944,3.0454736,4.3761535,5.4633327,4.8734436,3.9200184,2.901431,1.9548649,1.0597426,0.6790583,0.4081209,0.28122616,0.26064864,0.22292319,0.20234565,0.20577525,0.16462019,0.09602845,0.09602845,0.1097468,0.16119061,0.14747226,0.082310095,0.12346515,0.2503599,0.432128,1.1454822,2.2258022,2.867135,2.5824795,3.0214665,2.9940298,2.1194851,0.83681935,0.45613512,0.33609957,0.32238123,0.31552204,0.26407823,0.17147937,0.13032432,0.072021335,0.0,0.0,0.010288762,0.0034295875,0.0,0.0034295875,0.017147938,0.08573969,0.08573969,0.05144381,0.017147938,0.020577524,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.0274367,0.041155048,0.05144381,0.037725464,0.017147938,0.0034295875,0.0,0.0034295875,0.01371835,0.01371835,0.020577524,0.041155048,0.06516216,0.07545093,0.048014224,0.024007112,0.034295876,0.09602845,0.1920569,0.25721905,0.4046913,0.59331864,0.7373613,0.70649505,0.75450927,0.86082643,0.7407909,0.5007198,0.64133286,0.97057325,1.3752645,1.6256244,1.5947582,1.255229,1.4815818,2.020027,2.1332035,1.7319417,1.3752645,1.1111864,1.0631721,1.1111864,1.0631721,0.6756287,0.61046654,0.53501564,0.4629943,0.4355576,0.5212973,0.45270553,0.35324752,0.29494452,0.31552204,0.4115505,0.7099246,0.6344737,0.4938606,0.42526886,0.4081209,0.42526886,0.64476246,0.84367853,0.9259886,0.9259886,0.6276145,0.548734,0.607037,0.66191036,0.51100856,0.34981793,0.21263443,0.1097468,0.061732575,0.06859175,0.09602845,0.12689474,0.4081209,0.77508676,0.65162164,0.64476246,0.7476501,0.64476246,0.34638834,0.18519773,0.20920484,0.39097297,0.52472687,0.4972902,0.26064864,0.23664154,0.16462019,0.13375391,0.15776102,0.18519773,0.28465575,0.26750782,0.2194936,0.2194936,0.31895164,0.14061308,0.048014224,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.020577524,0.048014224,0.08916927,0.12689474,0.13032432,0.09945804,0.061732575,0.020577524,0.0034295875,0.0,0.0034295875,0.024007112,0.024007112,0.017147938,0.006859175,0.0,0.0,0.010288762,0.0034295875,0.0034295875,0.01371835,0.01371835,0.0034295875,0.006859175,0.01371835,0.010288762,0.0,0.0,0.0,0.0034295875,0.017147938,0.041155048,0.26407823,1.4129901,2.6853669,3.450165,3.2546785,2.6922262,2.07833,1.6530612,1.5364552,1.704505,1.6599203,1.3341095,0.97057325,0.71678376,0.6241849,0.65505123,0.65162164,0.58988905,0.48700142,0.4081209,0.39097297,0.44927597,0.5041494,0.53501564,0.5658819,0.7099246,1.0597426,1.5810398,2.0337453,1.9720128,1.728512,1.5501735,1.2860953,1.0117283,1.0220171,0.90884066,0.72364295,0.5453044,0.4046913,0.28465575,0.17490897,0.17833854,0.19548649,0.19891608,0.2194936,0.18176813,0.15433143,0.12346515,0.09259886,0.072021335,0.0548734,0.048014224,0.041155048,0.030866288,0.01371835,0.017147938,0.017147938,0.0274367,0.041155048,0.05144381,0.024007112,0.024007112,0.082310095,0.21263443,0.39440256,0.72707254,1.0014396,1.2655178,1.4438564,1.3443983,1.4987297,1.5398848,1.4438564,1.2037852,0.84367853,0.5658819,0.37039545,0.25721905,0.1920569,0.10288762,0.034295876,0.01371835,0.010288762,0.010288762,0.01371835,0.024007112,0.0274367,0.05144381,0.09602845,0.12689474,0.13375391,0.14747226,0.16804978,0.19891608,0.2469303,0.29494452,0.42526886,0.490431,0.53501564,0.77851635,0.8265306,0.8745448,0.82996017,0.6756287,0.45956472,0.29151493,0.18176813,0.082310095,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.048014224,0.0,0.0,0.030866288,0.0548734,0.058302987,0.048014224,0.010288762,0.0,0.0,0.010288762,0.048014224,0.030866288,0.017147938,0.01371835,0.010288762,0.0,0.010288762,0.0034295875,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.010288762,0.01371835,0.017147938,0.017147938,0.006859175,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.12346515,0.09602845,0.0548734,0.024007112,0.01371835,0.0,0.0,0.0,0.041155048,0.13032432,0.22978236,0.3018037,0.26407823,0.17490897,0.09602845,0.12346515,0.072021335,0.024007112,0.0,0.0034295875,0.01371835,0.0274367,0.01371835,0.030866288,0.09259886,0.15433143,0.31209245,0.8093826,1.5844694,2.8259802,4.972902,4.4859004,3.0283258,2.644212,3.474172,3.7519686,2.7882545,2.4830213,2.3321195,2.0680413,1.6770682,1.5810398,1.1900668,0.823101,0.7990939,1.4335675,1.6667795,1.7799559,1.6393428,1.1454822,0.22978236,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1097468,0.1097468,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.19548649,0.24350071,0.18519773,0.31895164,0.5761707,0.51100856,0.44584638,0.45613512,0.39783216,0.5555932,0.7956643,1.0700313,1.3101025,1.4198492,1.4198492,1.3375391,1.0117283,0.53844523,0.24350071,0.36696586,0.52472687,0.86082643,1.196926,1.039165,0.939707,0.9328478,0.8162418,0.6241849,0.6241849,0.83338976,1.0666018,1.2586586,1.2380811,0.764798,0.7373613,0.805953,0.67219913,0.44927597,0.65505123,0.89855194,0.6310441,0.37382504,0.29494452,0.19891608,0.19891608,0.30866286,0.41840968,0.47671264,0.48700142,0.548734,0.48357183,0.40126175,0.34638834,0.26064864,0.39440256,0.7373613,1.6496316,2.952875,3.9680326,3.07634,2.836269,2.5241764,1.786815,0.64133286,0.65162164,0.5178677,0.32238123,0.1920569,0.29151493,0.25378948,0.09602845,0.0,0.0,0.0,0.048014224,0.024007112,0.0,0.017147938,0.09259886,0.22635277,0.22292319,0.15090185,0.082310095,0.106317215,0.082310095,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.041155048,0.041155048,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.017147938,0.06859175,0.16804978,0.25378948,0.4115505,0.64476246,0.864256,0.89855194,0.9602845,1.0768905,1.0528834,0.89855194,0.823101,0.8128122,0.9294182,1.1523414,1.4267083,1.6324836,2.085189,2.2326615,2.0131679,1.5604624,1.2037852,1.0940384,1.2792361,1.3409687,1.1146159,0.6859175,0.61389613,0.5212973,0.40126175,0.32581082,0.47328308,0.5212973,0.41498008,0.36696586,0.53501564,1.0220171,1.5844694,1.2037852,0.6893471,0.42183927,0.33609957,0.31209245,0.5418748,0.7133542,0.6927767,0.53501564,0.5693115,0.6241849,0.6207553,0.548734,0.48700142,0.35324752,0.20234565,0.116605975,0.12003556,0.16804978,0.25378948,0.23664154,0.17833854,0.14061308,0.21263443,0.16462019,0.39097297,0.5624523,0.5041494,0.19891608,0.12346515,0.35324752,0.64133286,0.78537554,0.6241849,0.30866286,0.12003556,0.041155048,0.07545093,0.26064864,0.37039545,0.32238123,0.20920484,0.16119061,0.3806842,0.22292319,0.082310095,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.9842916,2.4727325,2.7162333,2.4487255,1.9857311,1.6496316,1.546744,1.5707511,1.5364552,1.2792361,0.9568549,0.65848076,0.42869842,0.58645946,0.607037,0.5418748,0.44584638,0.39783216,0.31209245,0.33609957,0.39783216,0.5144381,0.8093826,0.7956643,1.0597426,1.5913286,2.1194851,2.1057668,1.8725548,1.6221949,1.4472859,1.3409687,1.2037852,0.8265306,0.5761707,0.39440256,0.2469303,0.1371835,0.08916927,0.06859175,0.061732575,0.061732575,0.061732575,0.061732575,0.05144381,0.05144381,0.061732575,0.061732575,0.061732575,0.061732575,0.0548734,0.041155048,0.01371835,0.0274367,0.030866288,0.024007112,0.01371835,0.01371835,0.0274367,0.020577524,0.12346515,0.37039545,0.6859175,0.881404,1.0940384,1.2175035,1.1249046,0.6859175,0.5144381,0.64819205,0.7990939,0.83338976,0.7476501,0.7613684,0.6173257,0.42183927,0.23664154,0.09259886,0.041155048,0.048014224,0.0548734,0.05144381,0.07545093,0.07545093,0.07545093,0.09945804,0.17833854,0.33609957,0.36010668,0.42869842,0.45956472,0.4424168,0.4424168,0.42869842,0.4355576,0.4046913,0.34981793,0.34981793,0.40126175,0.4389872,0.4389872,0.38754338,0.29151493,0.18176813,0.106317215,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.01371835,0.017147938,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2929544,1.1317638,1.0185875,0.7305021,0.36696586,0.35324752,0.4115505,1.4095604,2.287535,2.2806756,0.91227025,0.84024894,0.78194594,0.8196714,0.922559,0.9259886,0.9877212,0.65505123,0.39783216,0.35324752,0.3566771,0.4081209,0.48357183,0.58302987,0.61389613,0.37382504,0.58988905,1.3958421,2.627064,4.0949273,5.5593615,5.7377,5.90232,5.809721,5.295283,4.280125,2.5138876,3.9337368,5.171818,4.513337,1.8862731,1.1626302,1.3855534,1.8554068,1.9651536,1.2037852,1.0837497,0.82996017,0.64133286,0.47328308,0.044584636,0.010288762,0.0,0.048014224,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.05144381,0.07888051,0.09602845,0.116605975,0.1371835,0.116605975,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16119061,0.38754338,0.42869842,0.26750782,0.1371835,0.31552204,0.32581082,0.28465575,0.2194936,0.07888051,0.22978236,0.48014224,1.0288762,1.488441,0.89512235,0.864256,0.7373613,0.4938606,0.24007112,0.23321195,0.34295875,0.5007198,0.7373613,0.9842916,1.0494537,1.6153357,1.4747226,0.939707,0.3806842,0.23664154,0.18862732,0.21263443,0.29494452,0.36353627,0.28808534,0.31209245,0.3018037,0.28122616,0.29837412,0.44927597,0.5658819,0.58645946,0.53501564,0.4355576,0.30866286,0.30866286,0.5555932,0.85396725,1.1214751,1.4267083,1.8313997,1.4987297,1.0906088,0.90884066,0.881404,1.7010754,1.3649758,1.430138,2.1194851,2.3321195,1.3615463,1.8416885,1.862266,1.0254467,0.432128,0.37725464,0.39440256,0.31552204,0.14747226,0.058302987,0.1371835,0.16462019,0.22978236,0.30866286,0.26750782,0.18176813,0.06516216,0.0,0.06516216,0.32238123,0.18519773,0.14061308,0.2777966,0.4664239,0.37382504,0.1371835,0.030866288,0.01371835,0.037725464,0.048014224,0.020577524,0.0034295875,0.01371835,0.037725464,0.048014224,0.020577524,0.0034295875,0.0034295875,0.01371835,0.01371835,0.017147938,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.017147938,0.0274367,0.044584636,0.09259886,0.15433143,0.28122616,0.42869842,0.4355576,0.4698535,0.64133286,0.9945804,1.2689474,0.922559,0.77165717,0.6927767,0.8162418,1.1626302,1.6324836,1.6530612,1.6393428,1.4953002,1.2312219,0.9362774,0.8745448,0.9259886,0.9945804,0.9842916,0.77165717,0.58988905,0.5624523,0.59674823,0.6962063,0.94999576,1.1351935,0.8779744,0.7476501,0.99801,1.5844694,1.8519772,1.1934965,0.5693115,0.37039545,0.42183927,0.44584638,0.6310441,0.69963586,0.6036074,0.53501564,0.8162418,0.70306545,0.5796003,0.58302987,0.61046654,0.4972902,0.22292319,0.08573969,0.18862732,0.45956472,0.4389872,0.24350071,0.14747226,0.20577525,0.2503599,0.10288762,0.106317215,0.16119061,0.20234565,0.20920484,0.09945804,0.106317215,0.17833854,0.2709374,0.3566771,0.20577525,0.07888051,0.020577524,0.030866288,0.08916927,0.13032432,0.13375391,0.12003556,0.116605975,0.16119061,0.09259886,0.037725464,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.20234565,0.52815646,0.66533995,0.8745448,1.0014396,1.0425946,0.99801,0.8745448,0.7305021,0.5521636,0.3806842,0.2503599,0.19548649,0.216064,0.21263443,0.18862732,0.16462019,0.16462019,0.16804978,0.18519773,0.24007112,0.32581082,0.39440256,0.53844523,0.823101,1.0425946,1.1111864,1.08032,1.4232788,1.6256244,1.5947582,1.5055889,1.7902447,1.5776103,1.371835,0.9568549,0.4355576,0.19891608,0.14061308,0.10288762,0.07545093,0.0548734,0.037725464,0.037725464,0.0274367,0.0274367,0.037725464,0.048014224,0.058302987,0.061732575,0.058302987,0.0548734,0.041155048,0.041155048,0.041155048,0.037725464,0.030866288,0.05144381,0.082310095,0.26407823,0.4629943,0.6344737,0.84367853,0.8848336,0.823101,0.7990939,0.78537554,0.58988905,0.7682276,1.2655178,1.5021594,1.3032433,0.89512235,0.94656616,0.6962063,0.42183927,0.26407823,0.22635277,0.17833854,0.18176813,0.16462019,0.1097468,0.07545093,0.16462019,0.24350071,0.26750782,0.2469303,0.2503599,0.216064,0.21263443,0.22978236,0.24350071,0.22292319,0.24007112,0.25378948,0.23321195,0.18519773,0.15433143,0.20577525,0.25721905,0.25721905,0.19891608,0.13032432,0.05144381,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.05144381,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058302987,0.058302987,0.044584636,0.030866288,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.017147938,0.0548734,0.034295876,0.006859175,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0034295875,0.010288762,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9362774,1.5330256,1.5330256,1.0323058,0.4424168,0.4972902,1.2655178,2.2395205,2.8156912,2.411,0.48014224,0.9568549,1.3238207,1.937717,2.4624438,1.8691251,2.0440342,2.9563043,4.0503426,4.647091,3.957744,3.4535947,2.867135,2.1194851,1.3443983,0.90198153,1.5741806,1.8313997,2.2395205,2.8225505,3.069481,3.923448,4.7431192,4.7362604,3.8514268,2.7711067,1.8965619,2.527606,3.0489032,2.6407824,1.2792361,1.138623,2.020027,2.2841053,1.5158776,0.48700142,0.40126175,0.2469303,0.15776102,0.12346515,0.010288762,0.0034295875,0.048014224,0.07545093,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.058302987,0.14061308,0.20234565,0.24007112,0.23664154,0.1920569,0.12003556,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.116605975,0.116605975,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07888051,0.17490897,0.18862732,0.11317638,0.037725464,0.09945804,0.11317638,0.09602845,0.06516216,0.0,0.058302987,0.22292319,0.4698535,0.61389613,0.30523327,0.29151493,0.23664154,0.14404267,0.07545093,0.12689474,0.20234565,0.42869842,0.66533995,0.7682276,0.6036074,0.7510797,0.64476246,0.38754338,0.12689474,0.0548734,0.010288762,0.0,0.020577524,0.058302987,0.06859175,0.082310095,0.072021335,0.106317215,0.20920484,0.34295875,0.39097297,0.48014224,0.4664239,0.34981793,0.29151493,0.31209245,0.47328308,0.67219913,0.86082643,1.039165,1.2517995,1.0563129,0.7442205,0.5658819,0.7442205,1.9239986,1.6530612,1.4472859,1.6221949,1.3169615,1.039165,1.196926,1.0254467,0.4938606,0.29837412,0.24007112,0.2777966,0.26750782,0.17490897,0.06516216,0.058302987,0.072021335,0.1371835,0.216064,0.22635277,0.30866286,0.24007112,0.18176813,0.1920569,0.22635277,0.22292319,0.28465575,0.42869842,0.5178677,0.24007112,0.08573969,0.13375391,0.14061308,0.07545093,0.12346515,0.12346515,0.116605975,0.08573969,0.072021335,0.17147937,0.061732575,0.024007112,0.082310095,0.15090185,0.041155048,0.01371835,0.010288762,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.020577524,0.041155048,0.08916927,0.15090185,0.17490897,0.21263443,0.3841138,0.6344737,0.8128122,0.65162164,0.5212973,0.37725464,0.3841138,0.6036074,1.0014396,1.0117283,1.0871792,1.1797781,1.1866373,0.9431366,0.7990939,0.8162418,0.85739684,0.8745448,0.922559,0.8093826,0.7407909,0.8162418,1.0837497,1.5158776,1.2003556,0.9945804,1.0048691,1.3032433,1.9445761,2.0577524,1.2483698,0.5007198,0.25721905,0.41498008,0.6276145,0.61046654,0.5041494,0.41840968,0.41498008,0.59674823,0.7888051,0.89169276,0.8745448,0.7682276,0.4389872,0.15776102,0.08573969,0.26750782,0.6344737,0.4115505,0.18176813,0.10288762,0.17490897,0.24007112,0.12003556,0.09259886,0.12003556,0.16119061,0.15776102,0.09602845,0.07888051,0.06859175,0.072021335,0.116605975,0.072021335,0.0274367,0.01371835,0.024007112,0.0274367,0.030866288,0.041155048,0.058302987,0.08573969,0.106317215,0.058302987,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.061732575,0.1920569,0.30866286,0.37725464,0.38754338,0.34638834,0.25378948,0.17490897,0.106317215,0.058302987,0.0548734,0.05144381,0.044584636,0.041155048,0.037725464,0.041155048,0.058302987,0.072021335,0.09945804,0.12689474,0.12346515,0.20577525,0.32581082,0.39440256,0.41498008,0.45613512,0.8128122,1.0460242,1.138623,1.2620882,1.762808,1.9239986,1.8554068,1.5158776,1.0666018,0.90884066,0.8196714,0.52815646,0.28122616,0.16804978,0.11317638,0.09259886,0.06516216,0.05144381,0.05144381,0.0548734,0.058302987,0.061732575,0.058302987,0.0548734,0.06516216,0.13032432,0.48014224,0.7682276,0.8711152,0.89512235,1.039165,1.2586586,1.4575747,1.5261664,1.3443983,1.1077567,1.0357354,1.1283343,1.2826657,1.2792361,1.7593783,2.0406046,1.8348293,1.2723769,0.8848336,1.1077567,0.9294182,0.6893471,0.64133286,0.97400284,0.8162418,0.52472687,0.26407823,0.11317638,0.058302987,0.116605975,0.16462019,0.19891608,0.20577525,0.18176813,0.15776102,0.14061308,0.16804978,0.2194936,0.23321195,0.2194936,0.216064,0.18519773,0.1371835,0.106317215,0.12689474,0.1371835,0.11317638,0.061732575,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06859175,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.072021335,0.09602845,0.082310095,0.07545093,0.044584636,0.020577524,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.030866288,0.037725464,0.006859175,0.0,0.0,0.0034295875,0.01371835,0.034295876,0.020577524,0.0034295875,0.0,0.006859175,0.01371835,0.010288762,0.006859175,0.0034295875,0.0,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3018037,0.9774324,1.0563129,0.72021335,0.31209245,0.31895164,1.0597426,1.646202,1.8519772,1.4164196,0.058302987,0.5693115,0.9602845,1.6770682,2.4658735,2.369845,2.335549,3.5016088,5.31929,6.7357097,6.2212715,5.4599032,3.8137012,2.633923,2.3561265,2.4967396,3.391862,4.448175,4.9248877,4.4516044,3.0077481,3.3815732,4.3281393,4.588788,3.7176728,2.0920484,1.7525192,1.6153357,1.4369972,1.1626302,0.91227025,1.0357354,1.786815,1.7971039,0.90541106,0.17490897,0.22292319,0.25378948,0.28808534,0.34295875,0.44927597,0.77165717,0.9534253,0.78194594,0.39097297,0.26750782,0.1920569,0.06859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041155048,0.20234565,0.25378948,0.26064864,0.18519773,0.06859175,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09259886,0.19548649,0.28122616,0.31895164,0.30866286,0.25378948,0.15433143,0.07545093,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.116605975,0.116605975,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.037725464,0.0,0.0,0.024007112,0.072021335,0.061732575,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.07888051,0.24007112,0.3841138,0.39440256,0.18176813,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.10288762,0.18176813,0.19891608,0.2503599,0.25378948,0.20920484,0.216064,0.2469303,0.30523327,0.3841138,0.4972902,0.66191036,0.67219913,0.6790583,0.58302987,0.5453044,1.0014396,2.393852,2.153781,1.5776103,1.2106444,0.8471081,1.0597426,1.0220171,0.77851635,0.4698535,0.31895164,0.216064,0.21263443,0.29151493,0.38754338,0.36353627,0.19548649,0.13032432,0.09259886,0.072021335,0.14747226,0.40126175,0.4664239,0.45270553,0.4046913,0.31209245,0.4389872,0.5007198,0.53158605,0.47328308,0.16804978,0.16462019,0.274367,0.26750782,0.15433143,0.15090185,0.15090185,0.17833854,0.14747226,0.09602845,0.17833854,0.12689474,0.10288762,0.14747226,0.20577525,0.13375391,0.07545093,0.030866288,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.06516216,0.13375391,0.18519773,0.14747226,0.2194936,0.31209245,0.37382504,0.39097297,0.28465575,0.17833854,0.14404267,0.22978236,0.48357183,0.6241849,0.7579388,0.91912943,1.0323058,0.91912943,0.7099246,0.69963586,0.71678376,0.7373613,0.8848336,0.85739684,0.7579388,0.8128122,1.0906088,1.4815818,0.9842916,0.89855194,1.0151579,1.2689474,1.7182233,1.7250825,1.0837497,0.50757897,0.35324752,0.59674823,0.70649505,0.5590228,0.41498008,0.39783216,0.47671264,0.45270553,0.65162164,0.7922347,0.77851635,0.6790583,0.4081209,0.24007112,0.21263443,0.33609957,0.61046654,0.37039545,0.15090185,0.06516216,0.106317215,0.16804978,0.106317215,0.09602845,0.13032432,0.17147937,0.16462019,0.18862732,0.3018037,0.28465575,0.116605975,0.0,0.0,0.0034295875,0.017147938,0.0274367,0.01371835,0.0034295875,0.006859175,0.024007112,0.048014224,0.07545093,0.05144381,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.041155048,0.06516216,0.041155048,0.024007112,0.010288762,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.006859175,0.017147938,0.020577524,0.017147938,0.010288762,0.017147938,0.017147938,0.034295876,0.072021335,0.13375391,0.32581082,0.5761707,0.91227025,1.2723769,1.5090185,1.7147937,1.8759843,1.7936742,1.4918705,1.2277923,1.1694894,0.864256,0.7339317,0.7956643,0.66191036,0.5727411,0.5555932,0.5590228,0.52472687,0.3841138,0.4629943,0.66191036,0.7476501,0.7373613,0.89855194,0.83338976,1.1866373,1.6633499,1.9891608,1.8999915,1.8416885,1.9411465,2.085189,2.1297739,1.8965619,1.762808,1.728512,1.903421,2.1469216,2.085189,2.551613,2.5241764,2.07833,1.4850113,1.2037852,1.4575747,1.4232788,1.214074,1.0666018,1.3101025,1.1077567,0.9431366,0.67219913,0.31895164,0.082310095,0.09602845,0.12689474,0.15090185,0.17147937,0.20920484,0.25721905,0.25378948,0.25721905,0.28465575,0.31209245,0.29837412,0.28465575,0.23321195,0.16462019,0.13032432,0.12689474,0.106317215,0.06516216,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.08573969,0.13032432,0.12003556,0.07888051,0.041155048,0.0274367,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.030866288,0.037725464,0.0274367,0.010288762,0.0034295875,0.010288762,0.020577524,0.020577524,0.01371835,0.006859175,0.0034295875,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.0,0.0,0.061732575,0.1097468,0.09602845,0.0,0.0,0.2194936,0.35324752,0.26750782,0.024007112,0.0034295875,0.0,0.26407823,0.90884066,1.9137098,1.5604624,1.7456601,2.9391565,4.540774,4.8905916,4.434457,2.3904223,1.7662375,3.192946,4.914599,4.955754,7.4524937,8.680285,7.363324,4.705394,4.0846386,5.4804807,6.4064693,5.56965,2.867135,2.1983654,1.9823016,1.8313997,1.5501735,1.1283343,0.82996017,0.90884066,0.91912943,0.7099246,0.432128,0.5521636,0.6824879,0.764798,0.84367853,1.0837497,1.9582944,2.4007113,2.1126258,1.3101025,0.7476501,0.48357183,0.18176813,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.017147938,0.08573969,0.432128,0.61046654,0.6824879,0.53844523,0.25721905,0.12346515,0.06516216,0.07888051,0.09602845,0.08916927,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.106317215,0.20234565,0.2777966,0.32238123,0.31895164,0.2469303,0.16119061,0.072021335,0.006859175,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072021335,0.072021335,0.0,0.0,0.048014224,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.10288762,0.12346515,0.15090185,0.15776102,0.19891608,0.33952916,0.65162164,0.65505123,0.7682276,0.83338976,0.9945804,1.6770682,3.1860867,2.8225505,1.7696671,0.91569984,0.8676856,1.1180456,1.2723769,1.1763484,0.85739684,0.5453044,0.34981793,0.26750782,0.39097297,0.6173257,0.65162164,0.37382504,0.29837412,0.20577525,0.106317215,0.23321195,0.490431,0.61389613,0.6207553,0.5693115,0.5555932,0.65848076,0.607037,0.52472687,0.4355576,0.29837412,0.3566771,0.3806842,0.34295875,0.2503599,0.15090185,0.106317215,0.14404267,0.14747226,0.10288762,0.08916927,0.16804978,0.1920569,0.17490897,0.15776102,0.23321195,0.14747226,0.0548734,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.116605975,0.25378948,0.34638834,0.18176813,0.12003556,0.15090185,0.23321195,0.28122616,0.22292319,0.19891608,0.16462019,0.17833854,0.37382504,0.65162164,0.75450927,0.805953,0.88826317,1.0631721,0.70649505,0.58302987,0.5555932,0.5727411,0.67219913,0.6893471,0.6241849,0.64476246,0.77851635,0.89169276,0.72707254,0.7510797,0.8779744,1.0288762,1.155771,1.0357354,0.7510797,0.5590228,0.59674823,0.89169276,0.6379033,0.4664239,0.4046913,0.45613512,0.6036074,0.47671264,0.37725464,0.32238123,0.32238123,0.36353627,0.38754338,0.37039545,0.34638834,0.3566771,0.4698535,0.4046913,0.1920569,0.07545093,0.09602845,0.09602845,0.0548734,0.044584636,0.072021335,0.13375391,0.20577525,0.28122616,0.5178677,0.51100856,0.22635277,0.0034295875,0.0,0.017147938,0.0274367,0.0274367,0.01371835,0.0034295875,0.0,0.0034295875,0.01371835,0.024007112,0.034295876,0.01371835,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.07545093,0.37725464,0.881404,1.2998136,1.097468,1.0940384,1.4678634,1.6770682,1.4815818,0.939707,0.90541106,0.86082643,1.1351935,1.5570327,1.4541451,1.2620882,1.2243627,1.2312219,1.1694894,0.9328478,1.1283343,1.5707511,1.7353712,1.6633499,1.9548649,1.8073926,1.9445761,2.2806756,2.6064866,2.5619018,2.2155135,2.0268862,1.978872,2.0337453,2.1194851,2.352697,2.386993,2.627064,3.000889,2.9631636,2.9048605,2.6785078,2.4007113,2.1572106,1.9891608,1.9720128,1.9274281,1.6599203,1.2312219,0.94999576,0.85739684,1.2860953,1.2826657,0.70649505,0.22978236,0.23321195,0.4115505,0.41498008,0.26064864,0.31895164,0.4629943,0.4972902,0.44927597,0.3806842,0.36353627,0.37039545,0.34981793,0.28122616,0.19548649,0.15433143,0.16119061,0.1371835,0.09602845,0.05144381,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.06516216,0.072021335,0.07888051,0.082310095,0.07545093,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.020577524,0.0034295875,0.01371835,0.024007112,0.034295876,0.020577524,0.01371835,0.010288762,0.0034295875,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.07888051,0.0,0.0,0.0548734,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.034295876,0.01371835,0.017147938,0.044584636,0.044584636,0.106317215,0.09602845,0.7922347,2.8739944,6.927767,3.9611735,4.931747,4.955754,2.8877127,1.313532,1.6770682,5.0929375,7.1061053,6.138962,3.4776018,2.6716487,1.8485477,1.7319417,2.0577524,1.5570327,0.9328478,1.1180456,1.0425946,0.6173257,0.70306545,0.8128122,0.9774324,0.939707,0.8025235,1.0220171,2.085189,2.952875,3.234101,2.651071,1.0528834,0.5144381,0.216064,0.06516216,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.082310095,0.082310095,0.030866288,0.15090185,0.4938606,0.7990939,0.82996017,0.58645946,0.30523327,0.26750782,0.38754338,0.48014224,0.45270553,0.30523327,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.106317215,0.17147937,0.24350071,0.23321195,0.18176813,0.1097468,0.037725464,0.0,0.0,0.037725464,0.0548734,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.048014224,0.0,0.048014224,0.024007112,0.061732575,0.19891608,0.3806842,0.45613512,0.59331864,0.7339317,0.9911508,1.6633499,3.117495,3.0317552,2.0303159,1.0494537,1.3443983,1.6736387,1.7353712,1.5398848,1.2175035,1.0220171,0.77851635,0.5418748,0.44584638,0.42869842,0.26064864,0.05144381,0.1920569,0.33952916,0.41498008,0.61046654,0.6824879,0.5178677,0.40126175,0.4081209,0.39783216,0.42183927,0.3806842,0.34638834,0.36010668,0.45613512,0.39783216,0.40126175,0.36353627,0.28465575,0.26064864,0.19891608,0.09259886,0.037725464,0.06516216,0.1371835,0.08916927,0.14061308,0.19548649,0.20920484,0.18176813,0.048014224,0.024007112,0.037725464,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.05144381,0.15090185,0.31895164,0.18519773,0.116605975,0.08573969,0.1097468,0.24350071,0.45270553,0.4389872,0.30523327,0.23664154,0.5178677,0.9328478,1.1008976,1.1797781,1.4027013,2.0749004,1.1351935,0.7613684,0.5727411,0.45270553,0.548734,0.64819205,0.67219913,0.6824879,0.67219913,0.548734,0.65848076,0.7613684,0.89512235,1.0460242,1.1454822,0.8265306,0.64819205,0.5693115,0.61046654,0.85396725,0.4629943,0.22978236,0.14404267,0.17833854,0.274367,0.32238123,0.35324752,0.30523327,0.20577525,0.16804978,0.14404267,0.1371835,0.18176813,0.28808534,0.45613512,0.4698535,0.26407823,0.18862732,0.26750782,0.18176813,0.072021335,0.037725464,0.030866288,0.044584636,0.106317215,0.09602845,0.16462019,0.17833854,0.09945804,0.01371835,0.0034295875,0.044584636,0.058302987,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.06859175,0.14747226,0.24350071,0.30523327,0.47671264,0.85739684,1.2003556,1.2312219,0.67219913,0.40126175,0.490431,0.83338976,1.2860953,1.6633499,1.3821237,1.1489118,0.9842916,0.9568549,1.1900668,1.371835,1.6016173,1.529596,1.2346514,1.2209331,1.8176813,2.5001693,2.3046827,1.6839274,2.503599,2.6716487,2.0097382,1.4369972,1.3238207,1.4953002,1.6907866,1.9857311,2.620205,3.5599117,4.4996185,3.2821152,2.8739944,2.8568463,2.952875,3.0523329,2.3801336,1.8554068,1.3546871,0.84024894,0.34981793,0.53501564,1.3684053,1.5673214,0.9842916,0.59674823,0.6207553,1.2860953,1.2860953,0.58645946,0.42869842,0.5624523,0.6962063,0.66533995,0.48357183,0.34981793,0.29151493,0.22978236,0.16804978,0.12003556,0.106317215,0.18176813,0.14404267,0.08916927,0.058302987,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08573969,0.14404267,0.09945804,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.024007112,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.15090185,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.006859175,0.0034295875,0.0034295875,0.010288762,0.010288762,0.020577524,0.0274367,0.33266997,1.2517995,3.1072063,1.4404267,2.5001693,4.125794,4.245829,0.8848336,1.3478279,3.1552205,5.007198,5.055212,0.89169276,1.0528834,1.0117283,1.3889829,2.0577524,2.153781,2.3424082,3.0420442,2.2463799,0.42526886,0.5178677,0.84367853,0.9294182,1.0254467,1.138623,1.0460242,0.9842916,1.3786942,1.961724,2.2326615,1.4438564,0.7407909,0.53844523,0.6756287,0.72364295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.061732575,0.12346515,0.17833854,0.29494452,0.28122616,0.22292319,0.20234565,0.29151493,0.5796003,0.82996017,1.0082988,1.0871792,1.039165,0.83338976,0.48014224,0.216064,0.09602845,0.0,0.058302987,0.072021335,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.034295876,0.048014224,0.106317215,0.1097468,0.06516216,0.006859175,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.010288762,0.048014224,0.1097468,0.18519773,0.26064864,0.274367,0.28808534,0.37725464,0.58988905,0.91912943,1.3066728,1.4164196,1.2209331,1.039165,1.5261664,2.0303159,2.1674993,2.0508933,1.8999915,2.0474637,1.8725548,1.3615463,0.9911508,0.86082643,0.69963586,0.70649505,0.5693115,0.5555932,0.70649505,0.84367853,0.8093826,0.4389872,0.31552204,0.4972902,0.5418748,0.17833854,0.20920484,0.33266997,0.4389872,0.6036074,0.6893471,0.6790583,0.58645946,0.4046913,0.07545093,0.15090185,0.1097468,0.116605975,0.16804978,0.07545093,0.24350071,0.17147937,0.1097468,0.12346515,0.1097468,0.024007112,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0,0.0,0.01371835,0.048014224,0.07545093,0.037725464,0.006859175,0.0,0.030866288,0.07888051,0.09602845,0.037725464,0.010288762,0.01371835,0.044584636,0.08916927,0.15776102,0.13375391,0.07888051,0.0548734,0.12346515,0.37725464,0.42183927,0.41498008,0.4355576,0.48357183,0.65162164,0.66533995,0.5727411,0.51100856,0.6824879,0.37725464,0.29494452,0.28465575,0.28808534,0.36696586,0.4938606,0.4972902,0.4698535,0.48014224,0.5727411,0.7133542,1.0563129,1.371835,1.5261664,1.4850113,1.1489118,1.1900668,1.371835,1.5364552,1.6359133,1.2826657,0.823101,0.432128,0.21263443,0.21263443,0.23321195,0.24007112,0.24007112,0.24007112,0.24007112,0.18862732,0.116605975,0.08573969,0.12003556,0.20234565,0.20234565,0.1097468,0.05144381,0.0548734,0.048014224,0.0274367,0.020577524,0.048014224,0.11317638,0.1920569,0.13032432,0.09259886,0.061732575,0.030866288,0.0034295875,0.0,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.034295876,0.041155048,0.030866288,0.01371835,0.024007112,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0274367,0.07888051,0.13032432,0.13375391,0.25721905,0.45613512,0.7510797,0.9602845,0.72021335,0.42183927,0.40126175,0.48357183,0.58302987,0.69963586,0.7990939,0.85739684,0.7888051,0.66533995,0.70306545,0.805953,0.94999576,0.9945804,0.96714365,1.0631721,1.6324836,2.1434922,2.527606,2.7813954,2.952875,3.0866287,2.8156912,2.2909644,1.7696671,1.6187652,1.5604624,1.6221949,1.8382589,2.1915064,2.633923,2.428148,2.2120838,2.1297739,2.1572106,2.0989075,1.8965619,1.5776103,1.1351935,0.6859175,0.45956472,0.8505377,2.5756202,4.3109913,4.681387,2.2806756,2.5001693,3.4192986,4.081209,3.9028704,2.6613598,1.6736387,1.5021594,1.2106444,0.64819205,0.48357183,0.3566771,0.2777966,0.20234565,0.13032432,0.12003556,0.14404267,0.14747226,0.14061308,0.1371835,0.14404267,0.12689474,0.09945804,0.07888051,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.09602845,0.13032432,0.1097468,0.020577524,0.0,0.0,0.0,0.0,0.13375391,0.15433143,0.15433143,0.17490897,0.18176813,0.09602845,0.030866288,0.0,0.0,0.0,0.0,0.030866288,0.030866288,0.0,0.0,0.037725464,0.020577524,0.020577524,0.048014224,0.048014224,0.010288762,0.0,0.0034295875,0.020577524,0.048014224,0.06859175,0.07888051,0.05144381,0.010288762,0.05144381,0.01371835,0.0034295875,0.0034295875,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.08573969,0.33952916,0.86082643,0.32238123,0.7579388,1.5673214,1.8348293,0.31209245,0.50757897,1.1111864,1.8725548,1.9925903,0.12346515,0.32924038,0.5521636,1.2792361,2.2806756,2.6064866,1.728512,1.6393428,1.138623,0.28465575,0.39097297,0.6962063,0.7956643,0.9774324,1.2312219,1.2346514,1.0768905,1.1763484,1.4815818,1.7730967,1.6427724,1.1900668,1.3821237,1.7182233,1.6667795,0.66876954,0.17147937,0.017147938,0.020577524,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.08916927,0.22978236,0.45270553,0.39097297,0.26750782,0.32238123,0.8128122,0.6001778,0.6893471,0.90884066,1.1420527,1.3306799,1.1283343,0.8128122,0.4664239,0.17490897,0.0,0.030866288,0.08573969,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.037725464,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.0548734,0.06516216,0.10288762,0.09259886,0.1371835,0.106317215,0.116605975,0.20234565,0.32924038,0.42869842,0.53844523,0.5693115,0.6036074,0.8745448,1.214074,1.2998136,1.4061309,1.6599203,2.037175,1.704505,1.4369972,1.2620882,1.1592005,1.0666018,0.7956643,0.78537554,0.9877212,1.1111864,0.5796003,0.51100856,0.6962063,0.864256,0.84367853,0.5521636,0.432128,0.38754338,0.44927597,0.5521636,0.53158605,0.70306545,0.65848076,0.5418748,0.39097297,0.11317638,0.16462019,0.1097468,0.1097468,0.17490897,0.17833854,0.18862732,0.18176813,0.15090185,0.09945804,0.037725464,0.006859175,0.0,0.0034295875,0.048014224,0.20234565,0.18519773,0.1371835,0.09259886,0.07545093,0.09259886,0.07545093,0.058302987,0.116605975,0.20577525,0.15433143,0.030866288,0.006859175,0.10288762,0.32924038,0.66191036,0.50757897,0.20920484,0.034295876,0.030866288,0.020577524,0.08573969,0.14747226,0.216064,0.25378948,0.20234565,0.25721905,0.28465575,0.30523327,0.37382504,0.58302987,0.7956643,0.7373613,0.7442205,0.9294182,1.2037852,0.97057325,0.864256,0.77851635,0.72707254,0.8162418,0.8676856,0.7888051,0.89855194,1.2312219,1.5227368,1.3546871,1.4987297,1.5707511,1.4644338,1.3341095,1.1523414,1.2415106,1.2003556,1.1146159,1.5570327,0.96714365,0.58988905,0.3566771,0.23664154,0.26407823,0.20234565,0.18519773,0.20920484,0.2503599,0.26750782,0.15776102,0.082310095,0.044584636,0.041155048,0.072021335,0.06516216,0.037725464,0.017147938,0.01371835,0.024007112,0.010288762,0.010288762,0.044584636,0.09945804,0.15090185,0.13375391,0.07888051,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.048014224,0.061732575,0.041155048,0.01371835,0.041155048,0.06859175,0.09259886,0.12003556,0.17833854,0.216064,0.15433143,0.082310095,0.041155048,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.072021335,0.12003556,0.14747226,0.26750782,0.48357183,0.65505123,0.5041494,0.29494452,0.25378948,0.274367,0.29151493,0.26407823,0.3806842,0.41840968,0.41840968,0.4355576,0.5624523,0.61046654,0.7613684,0.8025235,0.77851635,0.9945804,1.2346514,1.4850113,2.020027,2.6407824,2.6750782,2.452155,2.3972816,2.1160555,1.7079345,1.7765263,2.2909644,2.3904223,2.085189,1.611906,1.4164196,1.3924125,1.3169615,1.5673214,1.9857311,1.879414,2.020027,2.085189,1.6976458,1.0768905,1.0185875,1.488441,2.6167753,4.3007026,6.4304767,8.879202,7.8537555,6.6533995,6.7459984,8.196714,9.702303,6.9209075,4.5167665,3.4947495,3.6387923,3.5118976,2.6407824,1.3889829,0.607037,0.45956472,0.42526886,0.42183927,0.4424168,0.4698535,0.5007198,0.53501564,0.4698535,0.3841138,0.31209245,0.2469303,0.1371835,0.09259886,0.061732575,0.0274367,0.0,0.0,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.07888051,0.17490897,0.34638834,0.58645946,0.2503599,0.1097468,0.08573969,0.12689474,0.22978236,0.29494452,0.26064864,0.2194936,0.2194936,0.274367,0.14404267,0.06516216,0.020577524,0.006859175,0.037725464,0.037725464,0.058302987,0.058302987,0.037725464,0.037725464,0.0274367,0.01371835,0.030866288,0.061732575,0.061732575,0.041155048,0.01371835,0.0034295875,0.010288762,0.024007112,0.07888051,0.10288762,0.08573969,0.048014224,0.024007112,0.034295876,0.01371835,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.09602845,0.16462019,0.18519773,0.09259886,0.072021335,0.16119061,0.20577525,0.17833854,0.1920569,0.4115505,0.72021335,1.430138,2.2395205,2.253239,0.89855194,0.31209245,0.14404267,0.17833854,0.34295875,0.5624523,0.84024894,1.196926,1.5124481,1.5227368,1.4507155,1.2826657,1.3958421,1.7422304,1.8554068,1.4369972,1.6290541,2.1023371,2.369845,1.7902447,0.77165717,0.47328308,0.4938606,0.66876954,1.0734608,1.4644338,1.3101025,0.9945804,0.72021335,0.50757897,0.2777966,0.1920569,0.14747226,0.15433143,0.32581082,0.70649505,0.7510797,0.6344737,0.65162164,1.214074,1.1420527,1.2380811,1.2689474,1.2346514,1.371835,1.0768905,0.8471081,0.58645946,0.28808534,0.030866288,0.006859175,0.048014224,0.06516216,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.034295876,0.01371835,0.030866288,0.0,0.044584636,0.020577524,0.0,0.006859175,0.037725464,0.08916927,0.13375391,0.16462019,0.18862732,0.2469303,0.36353627,0.38754338,0.5658819,0.91912943,1.2380811,1.0666018,1.0151579,0.96714365,0.89169276,0.864256,0.5212973,0.58302987,0.84367853,0.9534253,0.41498008,0.31895164,0.5796003,0.823101,0.83338976,0.5453044,0.5453044,0.4698535,0.4664239,0.5144381,0.41498008,0.53844523,0.5693115,0.5590228,0.490431,0.26407823,0.26750782,0.1920569,0.15090185,0.17147937,0.18519773,0.16462019,0.2469303,0.24007112,0.13375391,0.08573969,0.13032432,0.16804978,0.23321195,0.39440256,0.7682276,0.72021335,0.59674823,0.48357183,0.37382504,0.14747226,0.14061308,0.1097468,0.14061308,0.20234565,0.16119061,0.030866288,0.010288762,0.116605975,0.39783216,0.89512235,0.7339317,0.35324752,0.116605975,0.09602845,0.058302987,0.058302987,0.11317638,0.20920484,0.2777966,0.18862732,0.12689474,0.13032432,0.17147937,0.39097297,1.0768905,1.7079345,1.8279701,1.9994495,2.318401,2.4212887,1.7593783,1.5330256,1.6736387,1.9582944,1.9994495,1.5776103,1.3375391,1.313532,1.430138,1.4918705,1.2929544,1.3101025,1.3341095,1.3032433,1.3101025,1.3203912,1.2860953,1.0528834,0.8196714,1.1592005,0.59674823,0.34638834,0.2709374,0.28465575,0.35324752,0.24007112,0.18176813,0.17833854,0.20920484,0.23321195,0.13032432,0.06859175,0.041155048,0.044584636,0.09259886,0.07545093,0.037725464,0.01371835,0.017147938,0.024007112,0.010288762,0.01371835,0.037725464,0.058302987,0.06516216,0.07888051,0.048014224,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.020577524,0.030866288,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.07888051,0.09259886,0.048014224,0.010288762,0.0274367,0.058302987,0.09945804,0.16119061,0.28808534,0.32581082,0.31552204,0.2469303,0.1371835,0.034295876,0.006859175,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.082310095,0.06859175,0.14061308,0.274367,0.38754338,0.33952916,0.25721905,0.24350071,0.2503599,0.23664154,0.1371835,0.20234565,0.18176813,0.16804978,0.216064,0.35324752,0.38754338,0.5590228,0.6859175,0.77851635,1.0254467,1.0597426,1.0871792,1.5741806,2.2360911,2.0508933,1.8691251,2.4555845,2.6887965,2.386993,2.318401,2.867135,3.093488,2.7402403,1.8725548,0.89169276,0.8779744,0.9431366,1.611906,2.5138876,2.3972816,2.5893385,2.7745364,2.4830213,1.8382589,1.5673214,1.7593783,2.1503513,3.1312134,5.2987127,9.465661,9.592556,7.98408,7.8503256,10.082987,13.265644,10.467101,7.9086285,7.531374,8.790032,8.663138,6.6876955,4.554492,3.0248961,2.2360911,1.7182233,1.646202,1.4438564,1.3821237,1.4781522,1.4987297,1.3512574,1.1934965,1.0357354,0.86082643,0.61389613,0.52472687,0.4972902,0.4664239,0.41498008,0.36010668,0.28808534,0.16462019,0.058302987,0.0,0.0,0.0,0.0,0.05144381,0.12689474,0.12346515,0.08916927,0.058302987,0.037725464,0.030866288,0.030866288,0.07545093,0.15090185,0.33609957,0.64476246,1.0323058,0.8025235,0.61046654,0.4389872,0.34981793,0.4664239,0.6344737,0.58645946,0.4664239,0.36696586,0.33609957,0.22292319,0.16462019,0.106317215,0.05144381,0.06859175,0.06859175,0.07545093,0.07888051,0.06859175,0.041155048,0.01371835,0.006859175,0.030866288,0.06516216,0.061732575,0.061732575,0.024007112,0.0,0.0034295875,0.024007112,0.07888051,0.09945804,0.09602845,0.072021335,0.0,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.034295876,0.12346515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.1920569,0.32581082,0.37382504,0.20920484,0.14747226,0.23664154,0.26407823,0.24007112,0.37725464,0.6893471,1.0357354,1.4918705,1.7902447,1.3032433,0.5453044,0.18519773,0.07888051,0.16119061,0.44584638,0.6241849,1.0220171,1.4575747,1.786815,1.9239986,1.7079345,1.2586586,1.2895249,1.728512,1.7319417,1.2346514,1.0700313,1.4815818,2.177788,2.3389788,1.3203912,1.0734608,1.255229,1.7490896,2.644212,3.532475,3.350707,2.8088322,2.311542,1.978872,1.546744,1.1317638,0.7682276,0.53501564,0.5555932,0.922559,1.0597426,1.0254467,0.9877212,1.2209331,1.7422304,1.8999915,1.6907866,1.3409687,1.2826657,0.9774324,0.8093826,0.6824879,0.5041494,0.216064,0.18519773,0.14061308,0.13032432,0.12346515,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.17490897,0.24350071,0.4389872,0.4355576,0.33952916,0.24350071,0.24350071,0.17147937,0.16119061,0.216064,0.31895164,0.42869842,0.35324752,0.19548649,0.2469303,0.48014224,0.52472687,0.3806842,0.34295875,0.34981793,0.34638834,0.28122616,0.35324752,0.48357183,0.59674823,0.6036074,0.39783216,0.39783216,0.33609957,0.2469303,0.15776102,0.06859175,0.18519773,0.31895164,0.33952916,0.28465575,0.32238123,0.38754338,0.4389872,0.53501564,0.7613684,1.2346514,1.1454822,0.9774324,0.823101,0.607037,0.1097468,0.14404267,0.15776102,0.14061308,0.09945804,0.06516216,0.020577524,0.010288762,0.061732575,0.2503599,0.7099246,0.66191036,0.4046913,0.2194936,0.17833854,0.15090185,0.14061308,0.09602845,0.08916927,0.11317638,0.09602845,0.09259886,0.10288762,0.18519773,0.5658819,1.6496316,2.644212,3.0146074,3.3026927,3.5599117,3.3541365,2.4967396,2.1880767,2.5413244,3.1723683,3.175798,2.218943,1.7182233,1.2860953,0.8128122,0.45613512,0.5624523,0.72021335,0.99801,1.3409687,1.5638919,1.5981878,1.4198492,1.2380811,1.1043272,0.939707,0.78537554,0.61046654,0.48014224,0.42526886,0.47328308,0.37382504,0.274367,0.21263443,0.19548649,0.1920569,0.1371835,0.082310095,0.0548734,0.07888051,0.15090185,0.14404267,0.06859175,0.020577524,0.01371835,0.01371835,0.01371835,0.020577524,0.024007112,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.044584636,0.06859175,0.0548734,0.0274367,0.006859175,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0034295875,0.017147938,0.041155048,0.09602845,0.09945804,0.044584636,0.010288762,0.020577524,0.024007112,0.041155048,0.09945804,0.2469303,0.24350071,0.34295875,0.33952916,0.18862732,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.09259886,0.18176813,0.26750782,0.28122616,0.31552204,0.31552204,0.2469303,0.12346515,0.17490897,0.18862732,0.13375391,0.048014224,0.048014224,0.08916927,0.23321195,0.5144381,0.8779744,1.1592005,1.2312219,1.1660597,1.488441,1.9342873,1.4507155,1.7216529,3.0146074,3.758828,3.5633414,3.2135234,3.100347,3.223812,3.0729103,2.369845,1.0666018,1.2003556,1.3958421,2.2738166,3.3781435,3.1860867,3.0866287,3.069481,2.9322972,2.5413244,1.8279701,1.5261664,1.5707511,1.9685832,2.7299516,3.882293,6.217842,6.3378778,6.790583,8.669997,11.602294,10.518545,10.0041065,11.039842,12.847235,12.895248,10.72432,8.7317295,6.8728933,5.3090014,4.389872,4.016047,3.309552,2.9940298,3.1072063,3.0111778,2.6304936,2.3629858,2.1091962,1.7971039,1.3889829,1.2312219,1.1832076,1.1317638,1.0254467,0.84367853,0.58988905,0.34295875,0.13032432,0.0,0.0,0.0,0.030866288,0.14061308,0.29494452,0.36010668,0.28808534,0.20577525,0.14404267,0.1097468,0.09945804,0.116605975,0.23321195,0.5007198,0.8745448,1.2037852,1.4369972,1.3821237,1.1111864,0.83681935,0.89855194,1.2689474,1.2277923,0.9842916,0.6790583,0.40126175,0.34295875,0.33609957,0.2709374,0.15433143,0.09945804,0.08916927,0.09259886,0.09602845,0.082310095,0.030866288,0.017147938,0.006859175,0.0274367,0.061732575,0.05144381,0.05144381,0.024007112,0.0034295875,0.010288762,0.048014224,0.058302987,0.06859175,0.072021335,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.13375391,0.47328308,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.024007112,0.12346515,0.024007112,0.0,0.06859175,0.18176813,0.24350071,0.048014224,0.274367,0.7510797,1.1214751,0.84024894,0.2777966,0.09259886,0.14747226,0.3841138,0.823101,1.0323058,0.9842916,0.90884066,1.2277923,2.534465,1.9480057,1.2895249,0.7510797,0.4355576,0.34981793,0.51100856,0.42183927,0.274367,0.23664154,0.45956472,0.59331864,0.8093826,1.5604624,2.5001693,2.486451,3.0111778,3.6559403,4.0880685,4.3452873,4.822,4.9694724,3.758828,2.3801336,1.4575747,1.0666018,1.0940384,1.1180456,1.1900668,1.2072148,0.91569984,0.6344737,0.22635277,0.29151493,0.805953,1.097468,1.2826657,1.2826657,1.1214751,0.89855194,0.77851635,0.864256,0.7099246,0.48014224,0.28122616,0.18176813,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14747226,0.14747226,0.0,0.0,0.12346515,0.15090185,0.09259886,0.037725464,0.18176813,0.35324752,0.45956472,0.48014224,0.42869842,0.36696586,0.32924038,0.23664154,0.2503599,0.28122616,0.0,0.35324752,0.31552204,0.25378948,0.29837412,0.33609957,0.3841138,0.41498008,0.274367,0.041155048,0.030866288,0.041155048,0.2194936,0.45613512,0.66533995,0.7613684,0.64133286,0.490431,0.36353627,0.33266997,0.5041494,0.39440256,0.26407823,0.12003556,0.0,0.0,0.072021335,0.18176813,0.2194936,0.16119061,0.07545093,0.05144381,0.017147938,0.024007112,0.19891608,0.7476501,0.84367853,0.5590228,0.26064864,0.15090185,0.274367,0.36010668,0.28122616,0.19548649,0.18176813,0.24350071,0.31895164,0.40126175,0.490431,0.7339317,1.4198492,1.7490896,1.9582944,2.277246,2.7573884,3.2821152,3.8308492,3.5290456,2.935727,2.5413244,2.760818,2.1743584,1.2963841,0.6241849,0.33609957,0.274367,0.50757897,0.9568549,1.4232788,1.7319417,1.7696671,1.4164196,1.3443983,1.3752645,1.3924125,1.3443983,1.646202,1.5947582,1.2243627,0.764798,0.65505123,0.64476246,0.5590228,0.48014224,0.4115505,0.29151493,0.16804978,0.09945804,0.06859175,0.0548734,0.030866288,0.09259886,0.06859175,0.034295876,0.01371835,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.024007112,0.030866288,0.017147938,0.006859175,0.030866288,0.10288762,0.17833854,0.18862732,0.13032432,0.044584636,0.044584636,0.0274367,0.010288762,0.0034295875,0.01371835,0.041155048,0.037725464,0.017147938,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.072021335,0.16804978,0.20577525,0.15090185,0.07545093,0.0274367,0.17833854,0.19891608,0.048014224,0.0,0.01371835,0.05144381,0.29151493,0.7682276,1.4027013,1.5741806,1.5913286,1.5638919,1.4850113,1.2037852,1.6804979,2.4041407,3.0283258,3.4947495,4.0434837,3.6285036,2.9665933,2.2841053,1.8382589,1.9239986,2.287535,2.534465,3.1415021,3.7725463,3.2958336,2.6476414,2.4247184,2.4967396,2.4761622,1.6942163,1.2037852,1.0014396,1.5673214,2.551613,2.7470996,1.8176813,2.5653315,3.7691166,5.5730796,9.489669,9.345626,9.263316,9.434795,9.962952,10.878652,11.646879,10.816919,9.345626,8.23444,8.515666,7.281014,5.9297566,5.2266912,5.1238036,4.746549,3.7211025,3.2272418,2.901431,2.5619018,2.1812177,1.8416885,1.5536032,1.2860953,0.9877212,0.61046654,0.36696586,0.19548649,0.072021335,0.0,0.0,0.0,0.14747226,0.34295875,0.50757897,0.5796003,0.5555932,0.45613512,0.34295875,0.2469303,0.19891608,0.17490897,0.22292319,0.42526886,0.7373613,1.0082988,1.5433143,1.9171394,2.0063086,1.9480057,2.1057668,2.3492675,2.2635276,1.7696671,1.0357354,0.47328308,0.4355576,0.52815646,0.4972902,0.31895164,0.19891608,0.1371835,0.11317638,0.106317215,0.10288762,0.09259886,0.030866288,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.058302987,0.32581082,1.1454822,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0034295875,0.024007112,0.0034295875,0.0,0.01371835,0.037725464,0.048014224,0.010288762,0.0548734,0.20234565,0.39783216,0.4972902,0.5693115,0.6756287,0.6962063,0.72707254,1.08032,1.0940384,0.90541106,0.90198153,1.0666018,1.0082988,1.1043272,0.77851635,0.37725464,0.13032432,0.13032432,0.2503599,0.34981793,0.42869842,0.44584638,0.32238123,0.4664239,0.6927767,0.89855194,1.2723769,2.3149714,2.9974594,3.210094,3.316411,3.6147852,4.3349986,4.9180284,4.866585,4.0880685,2.9220085,2.1434922,2.0406046,2.3458378,3.426158,4.5442033,3.8685746,2.7779658,2.3801336,1.7833855,1.1351935,1.6221949,1.6976458,1.313532,0.90198153,0.6893471,0.6927767,0.9259886,0.9568549,0.8779744,0.7442205,0.548734,0.19891608,0.044584636,0.0,0.0,0.0,0.0,0.020577524,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.030866288,0.0,0.0,0.024007112,0.030866288,0.017147938,0.006859175,0.037725464,0.072021335,0.09259886,0.12003556,0.16804978,0.24350071,0.5212973,0.37382504,0.274367,0.2709374,0.0,0.14061308,0.14747226,0.10288762,0.106317215,0.29837412,0.12346515,0.082310095,0.08916927,0.082310095,0.030866288,0.082310095,0.22292319,0.29494452,0.26064864,0.20234565,0.274367,0.18862732,0.1371835,0.16119061,0.1371835,0.08573969,0.05144381,0.024007112,0.0034295875,0.01371835,0.037725464,0.07545093,0.12346515,0.14747226,0.09945804,0.037725464,0.017147938,0.030866288,0.106317215,0.28465575,0.4115505,0.45270553,0.48700142,0.48357183,0.31209245,0.2709374,0.53158605,0.7990939,0.823101,0.41498008,0.29151493,0.29837412,0.33609957,0.39440256,0.5418748,0.7613684,0.922559,1.1146159,1.4335675,1.9857311,2.702515,2.9700227,3.0420442,3.3850029,4.6779575,4.355576,3.1552205,1.8108221,0.8471081,0.5796003,0.8025235,1.2586586,1.546744,1.6359133,1.8691251,1.7765263,1.8897027,2.020027,1.99602,1.6839274,1.5124481,1.4781522,1.2586586,0.8745448,0.71678376,0.6173257,0.48014224,0.42183927,0.42526886,0.34981793,0.2194936,0.17147937,0.1371835,0.08573969,0.041155048,0.044584636,0.030866288,0.020577524,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.006859175,0.017147938,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.024007112,0.020577524,0.0548734,0.19548649,0.31552204,0.30523327,0.16462019,0.020577524,0.030866288,0.082310095,0.13032432,0.13375391,0.0274367,0.01371835,0.044584636,0.058302987,0.041155048,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.034295876,0.041155048,0.030866288,0.0274367,0.006859175,0.044584636,0.048014224,0.010288762,0.0,0.01371835,0.030866288,0.14747226,0.4389872,0.9774324,1.0700313,1.0048691,1.0597426,1.3478279,1.8416885,2.335549,2.1915064,2.0303159,2.0063086,1.821111,1.7490896,1.8691251,2.4487255,3.2306714,3.4227283,3.8788633,4.4927597,4.8117113,4.5784993,3.724532,4.1120753,3.9097297,3.275256,2.49331,1.9754424,1.5741806,1.488441,1.6290541,1.9102802,2.2223728,2.651071,3.3061223,4.290414,5.6656785,7.466212,7.6685576,7.3393173,7.160979,7.596536,8.851766,10.696883,12.535142,12.898679,11.677745,10.113853,9.661148,7.1884155,5.3227196,5.099797,5.9400454,5.0140567,4.40359,4.40359,4.465323,3.2066643,2.4761622,1.937717,1.546744,1.1900668,0.6962063,0.3841138,0.216064,0.13375391,0.09602845,0.09602845,0.12689474,0.18519773,0.26750782,0.36353627,0.44584638,0.52815646,0.61046654,0.6036074,0.50757897,0.42869842,0.38754338,0.37039545,0.48014224,0.69963586,0.90884066,1.0460242,1.728512,2.3081124,2.5824795,2.7882545,3.9028704,4.32128,3.5221863,1.8897027,0.6927767,0.5693115,0.6824879,0.94999576,1.155771,0.9568549,0.58988905,0.32924038,0.18862732,0.14061308,0.12689474,0.09602845,0.058302987,0.034295876,0.024007112,0.01371835,0.0548734,0.0274367,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.041155048,0.32238123,1.2312219,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.14404267,0.2503599,0.3566771,0.4938606,0.6310441,0.61389613,0.4938606,0.5212973,0.6824879,0.58988905,0.5041494,0.48700142,0.41498008,0.4355576,0.3806842,0.31552204,0.2469303,0.13032432,0.13032432,0.4424168,0.6001778,0.48700142,0.35324752,0.35324752,0.5144381,0.65162164,0.7888051,1.1660597,1.6221949,1.6256244,1.6496316,1.9411465,2.5173173,2.6647894,2.7059445,2.3972816,1.8588364,1.5604624,1.2723769,1.5844694,2.510458,3.8342788,5.0929375,5.6005163,4.2698364,3.2375305,3.426158,4.554492,3.3609958,3.1037767,2.4315774,1.3375391,1.1763484,1.2826657,1.3032433,1.2586586,1.1763484,1.0906088,0.51100856,0.2503599,0.10288762,0.0,0.0,0.030866288,0.024007112,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.041155048,0.08573969,0.22635277,0.20920484,0.15776102,0.106317215,0.0,0.14404267,0.09602845,0.0548734,0.082310095,0.116605975,0.024007112,0.034295876,0.0548734,0.044584636,0.01371835,0.037725464,0.11317638,0.14061308,0.1097468,0.106317215,0.18519773,0.1097468,0.048014224,0.048014224,0.017147938,0.0034295875,0.0,0.0,0.0,0.006859175,0.017147938,0.034295876,0.09259886,0.23321195,0.48357183,0.6001778,0.29494452,0.08916927,0.14061308,0.24007112,0.33952916,0.34981793,0.4629943,0.6824879,0.84367853,0.980862,0.90884066,0.78537554,0.65505123,0.4664239,0.3018037,0.20234565,0.15776102,0.15090185,0.16462019,0.26407823,0.3566771,0.4698535,0.64133286,0.9294182,1.3375391,1.728512,2.2086544,2.952875,4.214963,4.40359,3.642222,2.5447538,1.6016173,1.1592005,1.3341095,1.6667795,1.7593783,1.605047,1.5638919,1.6187652,1.7696671,1.8485477,1.7662375,1.5124481,1.4610043,1.5158776,1.3786942,1.0288762,0.7339317,0.61046654,0.5041494,0.4424168,0.39783216,0.28465575,0.16462019,0.11317638,0.09259886,0.072021335,0.037725464,0.024007112,0.024007112,0.020577524,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0034295875,0.010288762,0.0274367,0.037725464,0.030866288,0.024007112,0.05144381,0.1371835,0.22978236,0.23321195,0.14061308,0.034295876,0.044584636,0.11317638,0.17147937,0.17490897,0.08573969,0.0548734,0.06859175,0.10288762,0.11317638,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.006859175,0.0,0.010288762,0.017147938,0.017147938,0.010288762,0.01371835,0.01371835,0.0548734,0.17490897,0.40126175,0.45270553,0.48014224,0.65162164,0.9945804,1.4232788,1.7833855,2.0646117,2.2841053,2.411,2.3835633,1.9720128,2.0646117,2.4555845,2.8945718,3.07634,3.5016088,3.9028704,4.016047,3.865145,3.7485392,6.0566516,5.8337283,4.671098,3.525616,2.6956558,2.7402403,2.5584722,2.4315774,2.417859,2.3664153,2.7985435,3.340418,4.331569,5.4187484,5.528495,5.2438393,5.48734,5.844017,6.200694,6.7459984,8.447074,9.952662,10.127572,9.626852,10.933525,12.370522,9.932085,6.7459984,4.98662,5.885172,5.586798,5.096367,5.086078,5.15467,3.8377085,2.5927682,1.9857311,1.7250825,1.5158776,1.0563129,0.77165717,0.53844523,0.40126175,0.31209245,0.15090185,0.15090185,0.15433143,0.16462019,0.17490897,0.16462019,0.33266997,0.5761707,0.6859175,0.6276145,0.53501564,0.6173257,0.84367853,0.91569984,0.8505377,0.9945804,1.0666018,1.4678634,1.961724,2.5653315,3.5564823,5.0106273,5.3878818,4.290414,2.386993,1.3992717,1.0082988,1.0906088,1.5090185,1.9445761,1.8862731,1.4027013,0.8848336,0.48357183,0.2709374,0.22978236,0.21263443,0.14747226,0.08573969,0.048014224,0.05144381,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.13032432,0.5007198,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.116605975,0.16462019,0.1920569,0.23664154,0.30523327,0.32924038,0.26750782,0.106317215,0.2469303,0.23321195,0.14404267,0.23664154,0.9568549,0.4389872,0.30523327,0.3841138,0.48700142,0.38754338,0.26407823,0.4629943,0.548734,0.42869842,0.31895164,0.20920484,0.26407823,0.37382504,0.41840968,0.26407823,0.4355576,0.39440256,0.40126175,0.5693115,0.84024894,0.70649505,0.65848076,0.6173257,0.58302987,0.65162164,0.42526886,0.6001778,1.0117283,1.8005334,3.3952916,4.3590055,3.175798,2.527606,3.2992632,4.5510626,3.5530527,3.8205605,3.4021509,2.253239,2.2429502,2.6887965,2.9734523,2.9322972,2.5927682,2.1812177,1.4164196,0.86082643,0.44927597,0.16804978,0.06859175,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.0548734,0.0,0.0,0.0,0.044584636,0.0548734,0.030866288,0.024007112,0.11317638,0.18176813,0.19548649,0.16119061,0.12689474,0.024007112,0.058302987,0.07545093,0.037725464,0.006859175,0.020577524,0.037725464,0.06516216,0.1097468,0.17833854,0.17147937,0.08573969,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.020577524,0.06516216,0.20577525,0.53844523,1.0494537,0.764798,0.37725464,0.23321195,0.33952916,0.44584638,0.34981793,0.37039545,0.6379033,1.097468,1.3924125,1.0837497,0.65848076,0.39440256,0.36353627,0.24007112,0.1371835,0.07545093,0.05144381,0.048014224,0.07888051,0.12003556,0.17490897,0.24350071,0.30866286,0.42869842,0.69963586,1.1626302,1.8176813,2.620205,3.100347,2.9871707,2.5173173,1.8965619,1.3169615,1.2415106,1.3752645,1.4232788,1.313532,1.2072148,1.2312219,1.3169615,1.313532,1.1934965,1.08032,1.2277923,1.2895249,1.1694894,0.90198153,0.6344737,0.4938606,0.41498008,0.37382504,0.31895164,0.19891608,0.106317215,0.07888051,0.082310095,0.07888051,0.037725464,0.01371835,0.017147938,0.024007112,0.020577524,0.010288762,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.006859175,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.01371835,0.030866288,0.034295876,0.0274367,0.024007112,0.041155048,0.072021335,0.12346515,0.14061308,0.106317215,0.0274367,0.06516216,0.15433143,0.18519773,0.13375391,0.09602845,0.09945804,0.07888051,0.08573969,0.10288762,0.061732575,0.0274367,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.010288762,0.024007112,0.034295876,0.034295876,0.034295876,0.0274367,0.034295876,0.0548734,0.06859175,0.08916927,0.16462019,0.33609957,0.5624523,0.7339317,0.91912943,1.5570327,2.2120838,2.5756202,2.4795918,1.9857311,1.9102802,1.845118,1.7250825,1.8485477,2.1332035,2.411,2.8911421,3.340418,3.083199,5.3330083,5.3981705,4.7431192,4.15666,3.7519686,3.3952916,3.069481,2.8911421,2.7985435,2.5619018,2.9048605,3.018037,3.7142432,4.57164,3.9371665,3.549623,3.981751,4.6436615,5.055212,4.822,6.1492505,7.3564653,7.5931067,7.8674736,11.067279,12.655178,10.326488,7.267296,5.874883,7.764586,8.532814,7.3873315,5.977771,4.8185706,3.2718265,2.1297739,1.6084765,1.4232788,1.313532,1.0563129,0.881404,0.6859175,0.5178677,0.36696586,0.16804978,0.09945804,0.07545093,0.06516216,0.06516216,0.1097468,0.20920484,0.44584638,0.61046654,0.64476246,0.6207553,0.85396725,1.3581166,1.5913286,1.5021594,1.5124481,1.8348293,2.287535,2.784825,3.2821152,3.7931237,5.4736214,5.744559,4.5956473,2.7470996,1.6530612,1.1489118,1.1592005,1.5776103,2.1023371,2.253239,2.0714707,1.9651536,1.6153357,1.0151579,0.48357183,0.3566771,0.25378948,0.15776102,0.082310095,0.06859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.1097468,0.23321195,0.13375391,0.0548734,0.09259886,0.18519773,0.53844523,1.6496316,0.8025235,0.4355576,0.41498008,0.53844523,0.5727411,0.4629943,0.39440256,0.3806842,0.3566771,0.20577525,0.13032432,0.09602845,0.09945804,0.09602845,0.0274367,0.0274367,0.017147938,0.006859175,0.0034295875,0.01371835,0.024007112,0.034295876,0.058302987,0.09602845,0.16804978,0.19548649,0.31209245,0.4629943,0.607037,0.72021335,0.65162164,0.53501564,0.5590228,0.85396725,1.4918705,1.9342873,2.6373527,2.819121,2.6373527,3.1620796,4.105216,4.791134,4.8905916,4.389872,3.5702004,2.6853669,1.8073926,1.1317638,0.6962063,0.4115505,0.20577525,0.106317215,0.0548734,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.034295876,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.020577524,0.020577524,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12003556,0.12003556,0.0,0.0,0.0,0.0,0.024007112,0.058302987,0.048014224,0.037725464,0.2709374,0.34638834,0.23321195,0.25721905,0.05144381,0.05144381,0.09602845,0.09945804,0.030866288,0.06859175,0.06516216,0.08916927,0.15090185,0.20920484,0.15090185,0.06859175,0.01371835,0.0,0.0,0.0,0.024007112,0.041155048,0.037725464,0.0274367,0.030866288,0.024007112,0.024007112,0.06516216,0.20920484,0.99801,1.0940384,0.8196714,0.53158605,0.64819205,0.69963586,0.5178677,0.3806842,0.4664239,0.8471081,1.1077567,0.91569984,0.59674823,0.33609957,0.20920484,0.15776102,0.12003556,0.08573969,0.058302987,0.041155048,0.08573969,0.11317638,0.116605975,0.09945804,0.09945804,0.15776102,0.26750782,0.44584638,0.70649505,1.0666018,1.5021594,1.9239986,2.1400626,1.961724,1.1832076,0.67219913,0.5727411,0.66191036,0.7922347,0.91569984,0.8265306,0.8093826,0.7442205,0.6310441,0.6036074,0.7613684,0.7476501,0.6344737,0.5007198,0.42183927,0.28465575,0.2194936,0.21263443,0.2194936,0.15776102,0.11317638,0.12346515,0.1371835,0.12003556,0.044584636,0.017147938,0.024007112,0.037725464,0.037725464,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.017147938,0.024007112,0.037725464,0.041155048,0.058302987,0.08573969,0.09945804,0.07545093,0.0034295875,0.058302987,0.16119061,0.15433143,0.061732575,0.072021335,0.12346515,0.082310095,0.041155048,0.0274367,0.017147938,0.037725464,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.037725464,0.048014224,0.048014224,0.05144381,0.05144381,0.05144381,0.030866288,0.034295876,0.06516216,0.13375391,0.20920484,0.23664154,0.29494452,0.75450927,1.3546871,1.6942163,1.2449403,1.097468,1.0117283,0.8093826,0.58302987,0.6756287,0.8196714,1.1660597,2.1674993,3.117495,2.1400626,2.5447538,3.0386145,3.4844608,3.8514268,4.2218223,2.9803114,2.6579304,2.6579304,2.6304936,2.4624438,2.9631636,2.6716487,3.059192,3.923448,3.415869,3.549623,3.4192986,3.5873485,3.875434,3.3678548,4.647091,5.960623,6.7391396,7.740579,11.039842,10.991828,8.745448,7.373613,8.364764,11.609154,12.881531,10.192734,6.660259,3.9063,2.0749004,1.5330256,1.1420527,0.8711152,0.71678376,0.6790583,0.66533995,0.6036074,0.4664239,0.29494452,0.20234565,0.07545093,0.041155048,0.044584636,0.106317215,0.31209245,0.30523327,0.42526886,0.5555932,0.64133286,0.6859175,0.96714365,1.5433143,2.1057668,2.4658735,2.5584722,3.1106358,4.0366244,4.791134,4.945465,4.1943855,5.6313825,5.830299,4.9008803,3.2306714,1.4644338,0.9945804,0.91569984,1.2037852,1.6942163,2.095478,2.4452958,3.0866287,3.0351849,2.1126258,0.939707,0.5453044,0.36353627,0.23664154,0.12346515,0.06859175,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.15776102,0.24350071,0.19548649,0.4664239,0.91912943,1.1111864,0.30523327,0.36696586,0.35324752,0.23664154,0.072021335,0.0,0.2194936,0.44927597,0.5212973,0.4115505,0.22978236,0.33952916,0.3018037,0.30866286,0.31895164,0.07545093,0.0274367,0.006859175,0.0,0.0034295875,0.01371835,0.05144381,0.041155048,0.030866288,0.082310095,0.29151493,0.32581082,0.78537554,1.371835,1.8691251,2.136633,2.428148,1.9720128,1.2586586,0.6756287,0.5041494,0.5144381,0.7305021,1.0151579,1.4781522,2.4418662,2.7230926,3.1586502,3.782835,4.3521466,4.3624353,3.3987212,2.7093742,2.1983654,1.7799559,1.3889829,0.88826317,0.52472687,0.26750782,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09259886,0.16462019,0.14747226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.09945804,0.082310095,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.10288762,0.10288762,0.1097468,0.1097468,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14747226,0.072021335,0.061732575,0.12346515,0.0,0.0,0.0,0.08573969,0.18862732,0.09259886,0.14061308,0.16119061,0.15433143,0.12346515,0.061732575,0.17147937,0.106317215,0.0274367,0.0,0.0,0.0,0.12689474,0.20920484,0.18519773,0.1371835,0.11317638,0.061732575,0.030866288,0.041155048,0.07545093,0.3566771,0.6927767,1.0666018,1.4027013,1.587899,1.2209331,0.881404,0.66191036,0.5418748,0.39783216,0.42183927,0.47328308,0.45613512,0.35324752,0.24350071,0.28122616,0.17147937,0.07888051,0.06859175,0.09259886,0.21263443,0.29151493,0.22292319,0.07545093,0.07545093,0.17490897,0.30866286,0.4115505,0.4938606,0.64133286,0.9568549,1.6770682,2.5756202,2.9665933,1.7079345,0.8162418,0.4389872,0.36010668,0.42869842,0.548734,0.53844523,0.45956472,0.37382504,0.31209245,0.274367,0.23664154,0.20920484,0.18519773,0.16462019,0.15090185,0.15090185,0.14404267,0.1371835,0.14747226,0.18176813,0.20920484,0.19548649,0.16462019,0.12003556,0.044584636,0.044584636,0.082310095,0.106317215,0.08916927,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.041155048,0.06516216,0.07545093,0.07545093,0.07545093,0.06516216,0.041155048,0.01371835,0.0034295875,0.0,0.017147938,0.061732575,0.12346515,0.13375391,0.12003556,0.07545093,0.030866288,0.030866288,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.030866288,0.030866288,0.041155048,0.06516216,0.08916927,0.09945804,0.07545093,0.12346515,0.28465575,0.37382504,0.32924038,0.18176813,0.23321195,0.20920484,0.20234565,0.2709374,0.4424168,0.6859175,0.8196714,1.1694894,1.7010754,2.0303159,2.054323,2.417859,2.8396983,2.9631636,2.3664153,1.6804979,1.7388009,2.1126258,2.352697,1.9994495,2.3046827,2.609916,3.806842,5.3330083,5.171818,5.6965446,4.722542,3.532475,2.819121,2.6853669,4.3933015,3.9165888,3.8857226,6.1561093,11.794352,11.074138,9.794902,10.288762,12.55915,14.280802,13.612033,9.259886,5.23698,3.1483612,2.1983654,1.7319417,1.3238207,0.9328478,0.6173257,0.5178677,0.65162164,0.65162164,0.5453044,0.4081209,0.33609957,0.2503599,0.20920484,0.22978236,0.31209245,0.45613512,0.6790583,0.8162418,0.83338976,0.7476501,0.6241849,0.7099246,0.9534253,1.7833855,3.059192,4.057202,4.1943855,5.271276,6.2041235,6.601956,6.759717,6.368744,6.23499,5.6245236,4.149801,1.7696671,1.1832076,1.0117283,1.0940384,1.4507155,2.2429502,2.719663,3.0866287,3.0489032,2.5138876,1.587899,0.84367853,0.48357183,0.29837412,0.17833854,0.09259886,0.06859175,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.030866288,0.048014224,0.037725464,0.09259886,0.18519773,0.22292319,0.061732575,0.11317638,0.17833854,0.16462019,0.07888051,0.024007112,0.048014224,0.08916927,0.11317638,0.12003556,0.14404267,0.17490897,0.12003556,0.07545093,0.06516216,0.0274367,0.006859175,0.0,0.0,0.0,0.0034295875,0.020577524,0.020577524,0.01371835,0.017147938,0.058302987,0.11317638,0.20920484,0.4629943,0.97400284,1.8176813,3.2443898,3.1860867,2.253239,1.1694894,0.78537554,0.66876954,0.5796003,0.5144381,0.48014224,0.48700142,0.96371406,1.4335675,1.646202,1.5433143,1.2517995,1.097468,0.99801,0.9602845,0.94656616,0.88826317,0.7305021,0.5178677,0.32581082,0.18176813,0.08573969,0.017147938,0.0,0.0,0.0,0.0,0.0,0.017147938,0.034295876,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.020577524,0.0,0.0,0.0,0.0,0.030866288,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.06859175,0.12346515,0.072021335,0.01371835,0.25721905,0.5007198,0.6001778,0.5624523,0.2777966,0.082310095,0.0,0.0,0.0,0.0,0.0,0.034295876,0.082310095,0.072021335,0.01371835,0.0,0.0,0.006859175,0.041155048,0.037725464,0.024007112,0.020577524,0.020577524,0.0,0.020577524,0.048014224,0.06516216,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.01371835,0.01371835,0.024007112,0.0,0.0,0.020577524,0.06516216,0.09259886,0.041155048,0.034295876,0.048014224,0.05144381,0.034295876,0.01371835,0.034295876,0.020577524,0.006859175,0.01371835,0.072021335,0.0548734,0.044584636,0.041155048,0.048014224,0.07545093,0.09945804,0.048014224,0.010288762,0.024007112,0.05144381,0.26407823,0.7579388,1.430138,2.0303159,2.1846473,2.318401,1.9548649,1.3615463,0.7888051,0.50757897,0.490431,0.70306545,1.0048691,1.0940384,0.47671264,0.2777966,0.30866286,0.33952916,0.28465575,0.20234565,0.14747226,0.26064864,0.3018037,0.21263443,0.12346515,0.15433143,0.28465575,0.36696586,0.3566771,0.34638834,0.4698535,0.75450927,1.1180456,1.3889829,1.2929544,0.84367853,0.4424168,0.2194936,0.18519773,0.2194936,0.2469303,0.22292319,0.17147937,0.12003556,0.10288762,0.116605975,0.1097468,0.09259886,0.07888051,0.06859175,0.058302987,0.061732575,0.07545093,0.08916927,0.09602845,0.09259886,0.09602845,0.08916927,0.07888051,0.082310095,0.05144381,0.061732575,0.08573969,0.10288762,0.08916927,0.037725464,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.058302987,0.06516216,0.06859175,0.07888051,0.09945804,0.082310095,0.06859175,0.048014224,0.017147938,0.0034295875,0.0,0.0,0.006859175,0.034295876,0.08573969,0.116605975,0.11317638,0.082310095,0.041155048,0.030866288,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.006859175,0.006859175,0.017147938,0.030866288,0.058302987,0.082310095,0.07545093,0.13375391,0.26750782,0.2469303,0.08916927,0.048014224,0.08916927,0.08916927,0.08573969,0.09259886,0.1371835,0.34295875,0.52472687,0.72364295,1.0768905,1.845118,2.3286898,2.9322972,3.3369887,3.5873485,4.0606318,3.3884325,2.7368107,2.3767042,2.3561265,2.510458,3.1963756,3.8617156,4.763697,5.576509,5.381023,4.938606,4.2046742,3.6593697,3.5633414,3.9543142,3.7005248,4.8768735,4.7088237,3.8034124,6.1321025,11.074138,10.429376,9.2153015,9.259886,9.205012,9.441654,6.4064693,4.081209,3.5770597,3.1620796,2.452155,1.728512,1.1180456,0.71678376,0.5796003,0.5761707,0.5693115,0.5144381,0.432128,0.39783216,0.4081209,0.48014224,0.5590228,0.6173257,0.66533995,0.7579388,0.83338976,0.8471081,0.78537554,0.6756287,0.66191036,0.6893471,0.9534253,1.4747226,2.1057668,2.884283,4.314421,5.6313825,6.5367937,7.174697,7.654839,7.874333,7.3050213,5.785714,3.5530527,1.9891608,1.3375391,1.0940384,1.1043272,1.546744,2.2395205,2.9803114,3.3438478,3.1380725,2.4041407,1.4747226,0.90541106,0.53501564,0.2777966,0.15090185,0.09945804,0.072021335,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.017147938,0.024007112,0.058302987,0.13032432,0.19548649,0.16804978,0.061732575,0.020577524,0.01371835,0.0274367,0.048014224,0.20920484,0.106317215,0.010288762,0.010288762,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.024007112,0.0274367,0.09945804,0.4115505,1.2072148,1.7593783,1.7593783,1.8485477,2.3492675,3.2718265,2.4658735,2.1812177,1.8005334,1.1214751,0.33952916,0.3566771,0.490431,0.52472687,0.39440256,0.18862732,0.20920484,0.22978236,0.26064864,0.29494452,0.30523327,0.31895164,0.26750782,0.19891608,0.13375391,0.041155048,0.05144381,0.020577524,0.01371835,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.044584636,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.030866288,0.05144381,0.08573969,0.1097468,0.072021335,0.09945804,0.082310095,0.037725464,0.0,0.0,0.15433143,0.09259886,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.061732575,0.037725464,0.09602845,0.26407823,0.432128,0.5418748,0.61046654,0.25721905,0.06859175,0.0,0.0,0.0,0.006859175,0.020577524,0.048014224,0.13032432,0.32924038,0.14061308,0.07545093,0.07545093,0.116605975,0.2194936,0.24007112,0.22978236,0.2194936,0.17490897,0.0,0.082310095,0.09945804,0.09602845,0.09259886,0.06516216,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.0274367,0.01371835,0.0034295875,0.006859175,0.010288762,0.0034295875,0.0,0.0,0.0,0.0034295875,0.017147938,0.044584636,0.0274367,0.010288762,0.0,0.0034295875,0.024007112,0.11317638,0.06516216,0.017147938,0.017147938,0.0274367,0.12689474,0.40126175,0.85396725,1.587899,2.8122618,3.2066643,3.07634,2.5413244,1.8725548,1.4953002,1.4575747,1.8519772,2.3732746,2.6545007,2.2566686,2.1023371,2.1263442,2.0165975,1.6427724,1.0357354,0.5041494,0.2777966,0.18176813,0.12346515,0.06516216,0.09259886,0.1920569,0.274367,0.29151493,0.25721905,0.24007112,0.30523327,0.432128,0.5796003,0.6962063,0.48700142,0.24350071,0.09602845,0.061732575,0.072021335,0.09602845,0.08916927,0.06516216,0.037725464,0.034295876,0.044584636,0.048014224,0.048014224,0.037725464,0.017147938,0.020577524,0.024007112,0.0274367,0.034295876,0.048014224,0.037725464,0.037725464,0.037725464,0.034295876,0.037725464,0.020577524,0.0274367,0.044584636,0.061732575,0.06859175,0.037725464,0.01371835,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.0548734,0.072021335,0.08573969,0.10288762,0.116605975,0.13375391,0.14747226,0.11317638,0.058302987,0.01371835,0.010288762,0.0034295875,0.006859175,0.010288762,0.024007112,0.058302987,0.08573969,0.10288762,0.09259886,0.06516216,0.030866288,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.044584636,0.058302987,0.10288762,0.16462019,0.13375391,0.034295876,0.006859175,0.034295876,0.0548734,0.0548734,0.05144381,0.07888051,0.17833854,0.4115505,0.7099246,1.0700313,1.5536032,2.3286898,3.2683969,3.782835,3.99204,4.7431192,4.7671266,4.091498,3.3061223,2.860276,3.059192,3.4844608,3.8685746,4.2423997,4.547633,4.616225,3.7794054,3.1449318,2.901431,3.0454736,3.3678548,3.1860867,4.0057583,4.108646,3.57363,4.2835546,9.582268,13.673765,13.203912,9.400499,8.080108,7.130112,5.1683884,3.7279615,3.309552,3.357566,2.983741,2.1846473,1.3958421,0.8779744,0.6859175,0.5624523,0.5212973,0.5007198,0.47671264,0.4664239,0.490431,0.58988905,0.6927767,0.7579388,0.78194594,0.83338976,0.89512235,0.9431366,0.9534253,0.8779744,0.864256,0.7888051,0.7476501,0.805953,0.9774324,1.2792361,2.1743584,3.2992632,4.461893,5.658819,6.8145905,7.654839,7.706283,6.742569,4.756838,3.4398763,2.3732746,1.646202,1.3306799,1.5090185,2.0714707,2.8808534,3.625074,4.180667,4.5853586,3.3609958,2.4830213,1.5913286,0.7339317,0.34295875,0.1920569,0.12346515,0.08573969,0.05144381,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.017147938,0.0034295875,0.006859175,0.072021335,0.16462019,0.15433143,0.061732575,0.024007112,0.024007112,0.0274367,0.006859175,0.16804978,0.106317215,0.034295876,0.030866288,0.01371835,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.072021335,0.13032432,0.1371835,0.22978236,0.7373613,0.8745448,1.2277923,1.9720128,3.1483612,4.633373,4.15323,3.7553983,3.865145,3.6936657,1.2415106,0.48014224,0.18519773,0.106317215,0.08916927,0.048014224,0.06516216,0.07545093,0.048014224,0.006859175,0.041155048,0.1097468,0.13032432,0.13032432,0.11317638,0.072021335,0.10288762,0.058302987,0.037725464,0.048014224,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.044584636,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.030866288,0.05144381,0.08573969,0.1097468,0.072021335,0.12003556,0.15090185,0.14747226,0.12689474,0.12346515,0.23664154,0.1371835,0.037725464,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08916927,0.1371835,0.19891608,0.29837412,0.44584638,0.23321195,0.07545093,0.0034295875,0.0,0.0,0.01371835,0.06859175,0.12689474,0.21263443,0.42869842,0.2469303,0.21263443,0.25721905,0.34981793,0.52472687,0.6036074,0.6276145,0.6207553,0.5590228,0.34638834,0.32238123,0.20920484,0.106317215,0.06516216,0.06516216,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.0274367,0.010288762,0.0034295875,0.0,0.0,0.0,0.08916927,0.07545093,0.041155048,0.020577524,0.010288762,0.037725464,0.11317638,0.30523327,0.8505377,2.1572106,3.0351849,3.4913201,3.234101,2.5619018,2.3389788,2.4315774,2.760818,3.2615378,3.7348208,3.8342788,3.2958336,3.0351849,2.9494452,2.8465576,2.4212887,1.3375391,0.5796003,0.16804978,0.048014224,0.11317638,0.061732575,0.08916927,0.15433143,0.22292319,0.25721905,0.15776102,0.13032432,0.15776102,0.216064,0.25721905,0.17490897,0.082310095,0.024007112,0.01371835,0.024007112,0.030866288,0.0274367,0.017147938,0.010288762,0.01371835,0.024007112,0.024007112,0.020577524,0.01371835,0.0,0.006859175,0.010288762,0.006859175,0.0034295875,0.017147938,0.010288762,0.01371835,0.01371835,0.006859175,0.006859175,0.0,0.006859175,0.01371835,0.0274367,0.034295876,0.0274367,0.01371835,0.01371835,0.020577524,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.041155048,0.0548734,0.072021335,0.09259886,0.106317215,0.1097468,0.16119061,0.11317638,0.048014224,0.01371835,0.01371835,0.006859175,0.010288762,0.020577524,0.030866288,0.05144381,0.061732575,0.072021335,0.07545093,0.06516216,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.048014224,0.061732575,0.05144381,0.0274367,0.006859175,0.017147938,0.034295876,0.037725464,0.034295876,0.06859175,0.1097468,0.28808534,0.5761707,0.8848336,1.0940384,1.728512,2.551613,3.1209247,3.474172,4.1429415,4.6093655,4.4756117,3.9508848,3.3987212,3.3301294,3.340418,3.2718265,3.1106358,2.952875,3.000889,2.3664153,1.961724,1.9342873,2.2292318,2.5790498,2.8911421,2.9974594,3.083199,3.3266997,3.9200184,8.947794,15.343974,16.019604,11.214751,8.501947,6.4304767,4.773986,3.4535947,2.651071,2.8019729,2.7779658,2.3046827,1.728512,1.2243627,0.78537554,0.6893471,0.64476246,0.61389613,0.5796003,0.53844523,0.58302987,0.66191036,0.764798,0.8505377,0.8779744,0.90198153,0.96371406,1.039165,1.097468,1.0940384,1.0940384,0.9945804,0.86082643,0.7407909,0.6824879,0.5727411,0.78194594,1.255229,1.9548649,2.8637056,3.8137012,4.7842746,5.425607,5.3707337,4.2389703,3.3712845,2.5241764,1.8965619,1.5810398,1.5638919,2.1263442,2.9906003,3.9371665,4.928317,6.0806584,5.3261495,4.506478,3.216953,1.7113642,0.922559,0.44584638,0.23321195,0.14747226,0.106317215,0.08916927,0.041155048,0.0274367,0.024007112,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.048014224,0.0,0.0034295875,0.07888051,0.106317215,0.06859175,0.017147938,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06516216,0.01371835,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.006859175,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.010288762,0.024007112,0.017147938,0.0034295875,0.010288762,0.030866288,0.041155048,0.01371835,0.030866288,0.061732575,0.06859175,0.044584636,0.01371835,0.024007112,0.024007112,0.017147938,0.0034295875,0.0,0.0,0.0,0.0034295875,0.020577524,0.048014224,0.14747226,0.26407823,0.28808534,0.29494452,0.5658819,1.1592005,2.061182,2.7573884,3.2272418,3.9474552,4.972902,4.756838,5.586798,6.3138704,2.352697,0.94656616,0.29151493,0.09602845,0.106317215,0.12346515,0.16462019,0.17833854,0.116605975,0.048014224,0.13375391,0.22292319,0.24350071,0.25378948,0.26750782,0.24350071,0.18176813,0.1371835,0.13375391,0.15090185,0.14404267,0.07545093,0.034295876,0.024007112,0.020577524,0.010288762,0.0034295875,0.0,0.0034295875,0.006859175,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07888051,0.15776102,0.2194936,0.25378948,0.24350071,0.18862732,0.17147937,0.1371835,0.07545093,0.0274367,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.030866288,0.0274367,0.048014224,0.11317638,0.23321195,0.23321195,0.14747226,0.05144381,0.0,0.0,0.010288762,0.09945804,0.1920569,0.2503599,0.26750782,0.23664154,0.28808534,0.37382504,0.48357183,0.65848076,0.7579388,0.8093826,0.8162418,0.78537554,0.72021335,0.5041494,0.28122616,0.1097468,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.017147938,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.08573969,0.017147938,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.01371835,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.037725464,0.017147938,0.0034295875,0.0,0.0,0.0,0.030866288,0.06516216,0.06516216,0.030866288,0.0,0.010288762,0.044584636,0.13032432,0.29837412,0.6001778,1.8073926,2.7402403,2.8088322,2.2909644,2.3286898,2.5619018,2.6236343,2.942586,3.5153272,3.923448,2.9117198,2.3458378,2.4144297,2.9391565,3.3472774,2.16064,1.0666018,0.33266997,0.072021335,0.22292319,0.07545093,0.024007112,0.048014224,0.12346515,0.2194936,0.116605975,0.06859175,0.058302987,0.06859175,0.07888051,0.058302987,0.030866288,0.010288762,0.0034295875,0.01371835,0.01371835,0.01371835,0.006859175,0.0034295875,0.01371835,0.030866288,0.0274367,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.01371835,0.0034295875,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.020577524,0.030866288,0.041155048,0.048014224,0.041155048,0.09945804,0.0548734,0.01371835,0.01371835,0.01371835,0.017147938,0.024007112,0.041155048,0.061732575,0.06516216,0.048014224,0.041155048,0.044584636,0.044584636,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.017147938,0.020577524,0.020577524,0.044584636,0.09602845,0.15433143,0.2709374,0.45613512,0.6790583,0.91569984,1.196926,1.6393428,2.2120838,2.74367,3.1552205,3.6044965,3.707384,3.4535947,3.2066643,3.0283258,2.6647894,2.1572106,1.6427724,1.3581166,1.1592005,1.1111864,1.2929544,1.7388009,2.428148,3.1209247,2.8739944,2.5207467,2.760818,4.1600895,8.738589,15.440002,17.439453,13.615462,8.549961,6.2727156,4.40702,2.9082901,1.937717,1.862266,1.9891608,2.054323,1.9925903,1.704505,1.0528834,0.939707,0.8711152,0.8162418,0.7476501,0.65505123,0.77165717,0.90198153,0.94999576,0.9431366,1.0082988,0.9945804,1.039165,1.0871792,1.1317638,1.2037852,1.2483698,1.2003556,1.097468,0.99801,0.980862,0.8711152,0.67219913,0.45613512,0.31209245,0.31209245,0.4355576,0.939707,1.670209,2.2738166,2.2223728,1.6736387,1.5158776,1.488441,1.4507155,1.3992717,2.1091962,3.0283258,3.957744,4.9180284,6.1458206,6.6876955,6.2967224,4.897451,3.0043187,1.7319417,0.8265306,0.41498008,0.24007112,0.15090185,0.116605975,0.08916927,0.07545093,0.06859175,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.38754338,0.53844523,0.34638834,0.09259886,0.09259886,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.07545093,0.31895164,0.06516216,0.0,0.0,0.0,0.0,0.01371835,0.06859175,0.082310095,0.037725464,0.0,0.0,0.017147938,0.030866288,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.072021335,0.037725464,0.048014224,0.116605975,0.09259886,0.017147938,0.017147938,0.017147938,0.0,0.0,0.0,0.017147938,0.024007112,0.01371835,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.034295876,0.12003556,0.29494452,0.5658819,0.85739684,1.6907866,2.527606,2.959734,2.7162333,5.1580997,5.857735,5.7308407,4.90431,2.7299516,1.4129901,0.52472687,0.19548649,0.23321195,0.12346515,0.19548649,0.15090185,0.11317638,0.14747226,0.24350071,0.45270553,0.5212973,0.6241849,0.70649505,0.48700142,0.32924038,0.32581082,0.4424168,0.5590228,0.47328308,0.32581082,0.17833854,0.11317638,0.106317215,0.044584636,0.020577524,0.006859175,0.01371835,0.034295876,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.082310095,0.082310095,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1097468,0.274367,0.29837412,0.18519773,0.1371835,0.08916927,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.044584636,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.15090185,0.1371835,0.06516216,0.0,0.0,0.0,0.22978236,0.22978236,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.0548734,0.061732575,0.061732575,0.061732575,0.061732575,0.061732575,0.072021335,0.09602845,0.12346515,0.024007112,0.0548734,0.10288762,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.08573969,0.08916927,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041155048,0.08573969,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.058302987,0.061732575,0.0,0.0,0.017147938,0.048014224,0.09945804,0.19891608,0.37039545,0.66876954,0.96714365,1.1454822,1.0837497,1.0357354,1.0048691,1.2655178,1.6770682,1.6770682,1.4953002,1.2758065,1.1420527,1.2860953,1.9685832,1.9445761,1.2792361,0.5453044,0.09945804,0.07545093,0.07545093,0.030866288,0.0,0.0,0.0,0.024007112,0.030866288,0.030866288,0.030866288,0.030866288,0.030866288,0.020577524,0.010288762,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0274367,0.05144381,0.05144381,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.024007112,0.06859175,0.10288762,0.11317638,0.07545093,0.05144381,0.06516216,0.06859175,0.061732575,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.030866288,0.030866288,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.05144381,0.06859175,0.06859175,0.106317215,0.16804978,0.1920569,0.26064864,0.432128,0.7613684,0.97057325,0.9294182,0.96714365,1.2415106,1.7559488,2.095478,2.2360911,2.3149714,2.4624438,2.7916842,2.877424,2.5893385,2.0989075,1.5913286,1.2346514,0.9294182,1.0837497,1.3821237,1.8691251,2.9288676,4.4447455,3.9611735,3.192946,3.4398763,5.6005163,5.73427,18.135658,23.256033,16.21852,6.8043017,4.791134,3.1895163,2.1160555,1.5330256,1.2517995,1.4472859,1.7319417,1.9891608,2.0920484,1.9068506,1.1866373,0.9328478,0.9294182,0.97400284,0.89855194,1.1454822,1.5913286,1.4987297,1.0185875,1.1900668,1.1763484,1.155771,1.0837497,1.0220171,1.1454822,1.3649758,1.4472859,1.3992717,1.3101025,1.3581166,1.2106444,1.0014396,0.7613684,0.5418748,0.39783216,0.28808534,0.2503599,0.274367,0.31895164,0.30523327,0.29151493,0.41840968,0.5453044,0.6790583,0.94656616,1.5193073,2.2326615,3.000889,3.9371665,5.3398676,7.2707253,7.174697,5.857735,4.0023284,2.1983654,1.1832076,0.66533995,0.39783216,0.23664154,0.15090185,0.116605975,0.106317215,0.09602845,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.07888051,0.1097468,0.07545093,0.0548734,0.07545093,0.09602845,0.17833854,0.24007112,0.072021335,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.082310095,0.2469303,0.09945804,0.024007112,0.0,0.0,0.0,0.45270553,1.6221949,1.5776103,0.37725464,0.08573969,0.31895164,0.2709374,0.21263443,0.21263443,0.16119061,0.1097468,0.082310095,0.08916927,0.17147937,0.41498008,0.5658819,0.41840968,0.2777966,0.25378948,0.23664154,0.26407823,0.26407823,0.16119061,0.010288762,0.0,0.010288762,0.017147938,0.01371835,0.0034295875,0.0034295875,0.020577524,0.0548734,0.058302987,0.058302987,0.13375391,0.4081209,0.3806842,0.25721905,0.1920569,0.26750782,0.2503599,0.18519773,0.18862732,0.37725464,0.8711152,0.6241849,0.6207553,0.90541106,1.5158776,2.4727325,4.201245,5.15467,5.857735,6.636252,7.6274023,6.0737996,3.8514268,2.1023371,1.0871792,0.20920484,0.07545093,0.16804978,0.40126175,0.77165717,1.3684053,1.2620882,0.94656616,0.6824879,0.65162164,0.939707,0.7510797,0.59674823,0.53158605,0.53844523,0.5212973,0.3566771,0.1371835,0.15090185,0.33266997,0.29151493,0.061732575,0.058302987,0.106317215,0.1097468,0.082310095,0.09602845,0.06859175,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.017147938,0.0,0.0,0.0,0.0,0.020577524,0.0548734,0.072021335,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.0548734,0.058302987,0.07888051,0.23664154,0.22635277,0.23664154,0.20920484,0.14404267,0.08573969,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.030866288,0.0274367,0.01371835,0.0,0.0,0.0,0.12689474,0.32581082,0.48357183,0.41498008,0.13032432,0.024007112,0.09602845,0.26064864,0.32924038,0.30866286,0.216064,0.106317215,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.020577524,0.024007112,0.0034295875,0.010288762,0.020577524,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.017147938,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.082310095,0.024007112,0.034295876,0.01371835,0.0,0.0034295875,0.0,0.010288762,0.0548734,0.0548734,0.010288762,0.0,0.0,0.006859175,0.010288762,0.01371835,0.0,0.0,0.010288762,0.020577524,0.037725464,0.07545093,0.15090185,0.25721905,0.3806842,0.48700142,0.53501564,0.5144381,0.490431,0.5796003,0.7613684,0.90884066,0.91227025,0.8128122,0.7613684,0.91227025,1.4198492,1.8039631,1.7902447,1.3649758,0.72364295,0.26064864,0.11317638,0.08916927,0.082310095,0.0548734,0.024007112,0.020577524,0.010288762,0.010288762,0.017147938,0.006859175,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.024007112,0.044584636,0.058302987,0.058302987,0.05144381,0.058302987,0.048014224,0.037725464,0.037725464,0.037725464,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.034295876,0.072021335,0.08573969,0.07888051,0.07545093,0.082310095,0.08573969,0.07545093,0.05144381,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.01371835,0.024007112,0.0274367,0.030866288,0.037725464,0.044584636,0.06859175,0.12003556,0.30866286,0.5521636,0.5693115,0.5693115,0.53844523,0.6036074,0.823101,1.1694894,1.1900668,1.255229,1.4850113,1.8999915,2.4247184,3.0386145,3.4604537,3.4055803,2.9391565,2.4555845,2.767677,3.525616,3.5633414,3.0454736,3.5050385,4.2938433,4.355576,4.0229063,3.8034124,4.389872,4.0949273,7.888051,13.516005,15.995596,7.599966,4.108646,2.2120838,1.3443983,1.0185875,0.83681935,0.9911508,1.1592005,1.2415106,1.2449403,1.2860953,1.1008976,0.91569984,0.8711152,0.94999576,0.9842916,1.1626302,1.4507155,1.862266,2.2155135,2.1434922,1.4953002,1.2209331,1.1077567,1.0837497,1.2037852,1.3272504,1.5090185,1.646202,1.6599203,1.5055889,1.2689474,0.9945804,0.72707254,0.490431,0.274367,0.21263443,0.18176813,0.22635277,0.32924038,0.41498008,0.3841138,0.3806842,0.5212973,0.8162418,1.1523414,1.5124481,2.1194851,2.585909,2.9391565,3.6319332,5.0414934,6.0566516,6.245279,5.8200097,5.6142344,2.7470996,1.3546871,0.7442205,0.45613512,0.274367,0.17833854,0.13375391,0.11317638,0.09259886,0.061732575,0.05144381,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.0274367,0.044584636,0.08916927,0.14747226,0.18176813,0.072021335,0.017147938,0.0,0.0,0.0,0.0,0.0,0.16119061,0.34638834,0.12003556,0.024007112,0.0,0.006859175,0.034295876,0.09259886,0.041155048,0.01371835,0.0,0.0,0.0,0.22292319,0.805953,0.77851635,0.18519773,0.041155048,0.16119061,0.13375391,0.106317215,0.116605975,0.106317215,0.15433143,0.17147937,0.28465575,0.5658819,1.0323058,1.1592005,0.9877212,0.8128122,0.7339317,0.64133286,1.4369972,1.3341095,0.805953,0.29494452,0.2469303,0.26064864,0.31209245,0.38754338,0.4389872,0.39440256,0.16804978,0.116605975,0.07888051,0.030866288,0.08573969,0.23664154,0.24350071,0.20577525,0.20920484,0.34638834,0.3806842,0.36010668,0.29494452,0.53844523,1.8073926,1.587899,1.7113642,1.8176813,1.8519772,2.0646117,2.7059445,3.0523329,3.426158,4.091498,5.2506986,4.7842746,4.7328305,4.3658648,3.1415021,0.7133542,0.5521636,1.9651536,4.149801,5.871454,5.456474,5.3227196,4.0846386,2.5413244,1.646202,2.5001693,1.5501735,1.2037852,1.0768905,0.9259886,0.67219913,0.4424168,0.26407823,0.25378948,0.37725464,0.45270553,0.18519773,0.07545093,0.05144381,0.05144381,0.037725464,0.048014224,0.034295876,0.044584636,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.037725464,0.044584636,0.12689474,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.10288762,0.13375391,0.20577525,0.25721905,0.26750782,0.25378948,0.2194936,0.17147937,0.08916927,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12689474,0.32238123,0.45613512,0.32581082,0.08916927,0.01371835,0.1097468,0.30866286,0.4389872,0.20577525,0.10288762,0.048014224,0.010288762,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.006859175,0.0274367,0.048014224,0.072021335,0.14404267,0.13032432,0.05144381,0.017147938,0.037725464,0.0,0.0,0.0,0.034295876,0.08573969,0.09945804,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.072021335,0.12346515,0.048014224,0.017147938,0.0274367,0.06516216,0.09945804,0.07545093,0.13032432,0.12003556,0.034295876,0.010288762,0.010288762,0.010288762,0.006859175,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.0274367,0.0548734,0.08573969,0.12346515,0.17147937,0.22292319,0.24007112,0.23664154,0.26064864,0.33952916,0.48014224,0.5555932,0.48357183,0.42869842,0.5418748,0.9602845,1.5227368,1.5707511,1.2895249,0.823101,0.2777966,0.09602845,0.0548734,0.05144381,0.034295876,0.01371835,0.006859175,0.0034295875,0.0034295875,0.006859175,0.010288762,0.01371835,0.006859175,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0274367,0.041155048,0.037725464,0.034295876,0.0548734,0.082310095,0.048014224,0.0274367,0.034295876,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0034295875,0.010288762,0.030866288,0.061732575,0.116605975,0.17490897,0.17490897,0.20920484,0.22635277,0.19548649,0.14404267,0.15090185,0.116605975,0.07545093,0.048014224,0.0274367,0.010288762,0.0034295875,0.010288762,0.017147938,0.020577524,0.024007112,0.037725464,0.034295876,0.030866288,0.0274367,0.020577524,0.020577524,0.044584636,0.18519773,0.4629943,0.8471081,0.5658819,0.38754338,0.32924038,0.4046913,0.6379033,0.7682276,0.72707254,0.922559,1.430138,1.99602,2.8637056,3.566771,3.82399,3.7862647,3.998899,4.629943,5.2609873,5.178677,4.557922,4.4516044,6.1321025,7.623973,8.48137,8.05953,5.5079174,4.856296,4.9488945,8.2481575,12.490558,10.700313,4.681387,1.8691251,0.83338976,0.5555932,0.4115505,0.45613512,0.5007198,0.548734,0.6036074,0.67219913,0.71678376,0.66191036,0.6790583,0.84367853,1.1249046,1.2277923,1.3855534,1.8142518,2.428148,2.8294096,2.6167753,2.1640697,1.7559488,1.5501735,1.5776103,1.6667795,1.8862731,2.1674993,2.3458378,2.153781,1.9651536,1.4747226,0.9842916,0.6276145,0.3806842,0.2503599,0.2194936,0.32581082,0.52472687,0.67219913,0.64133286,0.5521636,0.5418748,0.6927767,1.039165,1.3889829,1.8828435,2.5961976,3.5633414,4.7774153,5.576509,6.0875177,6.6739774,7.5279446,8.666568,6.783724,3.998899,1.8416885,0.8471081,0.5418748,0.37382504,0.2503599,0.17147937,0.12689474,0.10288762,0.09259886,0.061732575,0.041155048,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.14747226,0.20234565,0.32581082,0.25721905,0.037725464,0.0,0.0,0.01371835,0.2503599,0.4972902,0.12346515,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.06516216,0.048014224,0.01371835,0.0274367,0.09945804,0.13375391,0.26064864,0.64476246,1.4781522,2.0131679,1.4987297,0.9842916,0.90198153,1.0666018,2.7711067,2.3424082,1.3992717,0.85739684,0.91227025,0.6379033,0.4698535,0.44584638,0.5144381,0.5418748,0.48014224,0.5693115,0.8162418,1.1043272,1.2037852,0.8471081,0.64819205,0.5453044,0.5453044,0.7305021,0.7990939,0.61389613,0.42183927,0.6859175,2.0989075,2.170929,2.877424,3.6627994,3.9165888,2.976882,2.9906003,2.6167753,2.7093742,3.3061223,3.6353626,3.0283258,3.4776018,3.8274195,3.199805,0.9877212,1.2655178,3.6627994,6.1801167,7.1541195,5.219832,5.223262,4.7602673,4.125794,3.7519686,4.214963,3.2786856,2.6647894,2.1469216,1.7456601,1.7559488,1.2689474,1.1763484,1.1283343,0.97400284,0.7682276,0.35324752,0.12689474,0.058302987,0.058302987,0.0,0.106317215,0.1097468,0.08573969,0.08573969,0.14061308,0.16119061,0.16804978,0.17147937,0.15090185,0.07888051,0.06516216,0.0548734,0.044584636,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.0274367,0.017147938,0.09259886,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.09259886,0.15433143,0.20234565,0.2469303,0.30523327,0.31552204,0.2469303,0.14747226,0.12689474,0.08916927,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.037725464,0.030866288,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072021335,0.072021335,0.01371835,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08916927,0.18176813,0.21263443,0.12003556,0.06859175,0.020577524,0.061732575,0.17833854,0.274367,0.07545093,0.010288762,0.037725464,0.09259886,0.09602845,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.020577524,0.01371835,0.061732575,0.14747226,0.12003556,0.07545093,0.072021335,0.1371835,0.14061308,0.0548734,0.017147938,0.041155048,0.024007112,0.0034295875,0.0,0.034295876,0.08573969,0.09945804,0.020577524,0.0,0.0,0.0,0.0,0.020577524,0.048014224,0.10288762,0.16462019,0.17147937,0.072021335,0.09602845,0.15090185,0.18519773,0.1920569,0.15433143,0.17147937,0.15090185,0.082310095,0.044584636,0.017147938,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.017147938,0.0274367,0.034295876,0.044584636,0.07545093,0.09945804,0.10288762,0.11317638,0.15090185,0.24007112,0.31895164,0.26750782,0.21263443,0.2709374,0.53501564,0.9534253,0.97400284,0.82996017,0.607037,0.22978236,0.06859175,0.017147938,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.020577524,0.034295876,0.030866288,0.024007112,0.061732575,0.082310095,0.05144381,0.037725464,0.044584636,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.01371835,0.01371835,0.0274367,0.041155048,0.061732575,0.116605975,0.18519773,0.20920484,0.25378948,0.30866286,0.34638834,0.34638834,0.28808534,0.2503599,0.19891608,0.14747226,0.09602845,0.034295876,0.017147938,0.017147938,0.020577524,0.020577524,0.024007112,0.06516216,0.06516216,0.048014224,0.034295876,0.034295876,0.020577524,0.017147938,0.061732575,0.2709374,0.823101,0.70306545,0.5007198,0.34638834,0.32924038,0.490431,0.8779744,0.94999576,1.0082988,1.2312219,1.6599203,2.417859,3.0557625,3.4844608,3.7382503,3.9783216,4.3933015,5.07236,5.4907694,5.518206,5.446185,7.5382333,9.966381,11.427385,10.679735,6.5710897,5.504488,4.90431,6.060081,8.769455,11.351934,6.4407654,2.6750782,0.7682276,0.39440256,0.18519773,0.15776102,0.16462019,0.22978236,0.32238123,0.37382504,0.47671264,0.51100856,0.58988905,0.75450927,0.9911508,1.1351935,1.2860953,1.6256244,2.1915064,2.8911421,3.1860867,2.9288676,2.503599,2.1640697,2.0303159,1.978872,2.1674993,2.6133456,3.1449318,3.3747141,3.2683969,2.7573884,1.9411465,1.1043272,0.7305021,0.52815646,0.42526886,0.53501564,0.8265306,1.1214751,1.4267083,1.3581166,1.1489118,1.0082988,1.1214751,1.4507155,1.6976458,2.4418662,3.8617156,5.7308407,6.619104,6.90033,7.5519514,8.992378,11.108434,11.4033785,8.611694,4.976331,2.1263442,1.0563129,0.7305021,0.48357183,0.31209245,0.21263443,0.15090185,0.1371835,0.1097468,0.08573969,0.06516216,0.030866288,0.024007112,0.01371835,0.006859175,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28122616,0.6276145,0.53844523,0.106317215,0.01371835,0.041155048,0.09945804,0.26064864,0.36696586,0.037725464,0.006859175,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.06859175,0.2194936,0.24007112,0.14404267,0.020577524,0.020577524,0.01371835,0.01371835,0.048014224,0.34638834,1.3238207,2.2806756,1.471293,0.7510797,0.96714365,1.9548649,4.033195,2.9871707,1.7936742,1.6324836,1.8691251,1.1729189,0.5727411,0.36010668,0.607037,1.1626302,1.7010754,2.469303,4.2698364,6.1492505,5.377593,3.426158,2.5790498,2.5241764,2.942586,3.4981792,2.9288676,1.8725548,1.214074,1.3512574,2.2052248,2.510458,3.2821152,4.715683,5.871454,4.681387,4.650521,4.1155047,4.413879,5.3501563,5.206114,3.0489032,2.061182,1.8005334,1.7216529,1.1797781,1.9102802,3.9954693,4.880303,3.6868064,1.2277923,1.3375391,2.901431,4.8322887,6.077229,5.597087,5.6348124,5.0929375,4.1292233,3.292404,3.5461934,3.175798,3.3472774,3.1380725,2.2909644,1.2175035,0.64476246,0.37725464,0.42869842,0.5796003,0.37382504,0.61046654,0.64819205,0.53501564,0.42526886,0.6036074,0.59674823,0.6036074,0.61046654,0.5796003,0.42869842,0.33266997,0.23664154,0.22978236,0.25721905,0.14747226,0.12346515,0.116605975,0.07888051,0.017147938,0.017147938,0.0034295875,0.0,0.072021335,0.16804978,0.10288762,0.18519773,0.1097468,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.05144381,0.07888051,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.061732575,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.072021335,0.1920569,0.28465575,0.32581082,0.31209245,0.28808534,0.2194936,0.10288762,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.06516216,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15433143,0.17147937,0.061732575,0.15090185,0.030866288,0.006859175,0.017147938,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08916927,0.044584636,0.0,0.006859175,0.034295876,0.044584636,0.020577524,0.07888051,0.18862732,0.13375391,0.0274367,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.01371835,0.017147938,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.044584636,0.037725464,0.19548649,0.3566771,0.20920484,0.05144381,0.01371835,0.05144381,0.17490897,0.2194936,0.2469303,0.2503599,0.18862732,0.06859175,0.0548734,0.082310095,0.08916927,0.0,0.0,0.006859175,0.01371835,0.020577524,0.024007112,0.06516216,0.10288762,0.21263443,0.31209245,0.17833854,0.11317638,0.20577525,0.29151493,0.29494452,0.23664154,0.20577525,0.16462019,0.13375391,0.13032432,0.14404267,0.037725464,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.006859175,0.0274367,0.0274367,0.0274367,0.030866288,0.05144381,0.106317215,0.14747226,0.1371835,0.116605975,0.12346515,0.18176813,0.29837412,0.36696586,0.37382504,0.3018037,0.16119061,0.0548734,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.024007112,0.024007112,0.0548734,0.0548734,0.048014224,0.048014224,0.05144381,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.030866288,0.030866288,0.041155048,0.05144381,0.07545093,0.09602845,0.12689474,0.19548649,0.2469303,0.32924038,0.45956472,0.53844523,0.36696586,0.38754338,0.37039545,0.32924038,0.26064864,0.15090185,0.12003556,0.08573969,0.044584636,0.010288762,0.017147938,0.09602845,0.08916927,0.061732575,0.058302987,0.08916927,0.082310095,0.048014224,0.020577524,0.08573969,0.37382504,0.65848076,0.59674823,0.48357183,0.48014224,0.59674823,1.0871792,1.3615463,1.3272504,1.2003556,1.4815818,1.9548649,2.3664153,2.7779658,3.0283258,2.7402403,2.5790498,4.1292233,5.813151,6.9209075,7.623973,8.14527,9.626852,10.316199,9.273604,6.375603,5.284994,5.2747054,5.5147767,6.217842,8.632272,7.9189177,4.0949273,1.2312219,0.50757897,0.19891608,0.14404267,0.17147937,0.24007112,0.31552204,0.37382504,0.5041494,0.6207553,0.69963586,0.72364295,0.66191036,0.90541106,1.155771,1.488441,1.9342873,2.4795918,2.8705647,2.9906003,2.8534167,2.5824795,2.3972816,2.1674993,2.3732746,2.952875,3.7348208,4.4584637,4.870014,4.8768735,3.875434,2.2498093,1.371835,1.1317638,0.9945804,1.0494537,1.2689474,1.5021594,2.2360911,2.4007113,2.294394,2.1572106,2.1400626,2.218943,1.9308578,2.0680413,3.0660512,5.0003386,6.526505,7.449064,8.2310095,9.47938,11.917816,14.352823,13.516005,9.997248,5.518206,2.9254382,1.6736387,0.99801,0.6036074,0.34638834,0.22292319,0.18519773,0.14747226,0.12003556,0.10288762,0.07888051,0.06859175,0.041155048,0.024007112,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.072021335,0.116605975,0.1371835,0.07545093,0.19891608,0.3566771,0.4046913,0.30523327,0.12346515,0.024007112,0.0,0.0,0.0034295875,0.01371835,0.041155048,0.017147938,0.0,0.0,0.0,0.0,0.0,0.017147938,0.09259886,0.274367,0.70306545,0.5624523,0.274367,0.09602845,0.106317215,0.06859175,0.034295876,0.041155048,0.07888051,0.09259886,0.09259886,0.18176813,0.70649505,2.0063086,4.4104495,5.521636,3.5633414,2.2223728,2.49331,2.6990852,2.0406046,1.2072148,1.1489118,2.2498093,4.3487167,5.288424,7.5450926,13.697772,19.730417,15.0456,9.002667,6.9346256,7.9086285,10.405369,12.298501,9.208443,5.919468,3.9680326,3.707384,4.3178506,4.465323,3.3369887,3.1312134,4.108646,4.6093655,4.547633,5.007198,5.693115,6.355026,6.8043017,3.8274195,4.1429415,4.108646,2.8396983,2.2429502,2.2292318,2.3286898,2.2052248,1.9239986,1.9239986,1.8485477,3.532475,5.528495,6.7802944,6.6225333,7.4524937,8.200144,7.7371492,6.1458206,4.729401,6.1458206,7.0958166,6.3207297,3.9508848,1.5090185,1.2792361,1.0734608,1.5570327,2.311542,1.862266,1.9823016,2.16064,2.1194851,1.8485477,1.6187652,1.3855534,1.3272504,1.3443983,1.371835,1.3581166,1.0151579,0.64819205,0.70306545,1.0014396,0.7339317,0.61046654,0.58988905,0.38754338,0.07888051,0.09259886,0.017147938,0.0,0.36696586,0.83681935,0.5178677,0.922559,0.5555932,0.14747226,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.25378948,0.39440256,0.29151493,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12689474,0.30523327,0.24350071,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.09259886,0.15090185,0.21263443,0.20234565,0.14747226,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.12346515,0.18519773,0.1371835,0.041155048,0.034295876,0.08916927,0.12346515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.16804978,0.034295876,0.0,0.037725464,0.072021335,0.0,0.0,0.0,0.037725464,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.017147938,0.0,0.0,0.0,0.061732575,0.08573969,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14747226,0.7339317,0.36696586,0.1097468,0.006859175,0.06516216,0.26064864,0.77165717,1.0563129,1.2277923,1.2037852,0.70306545,0.29837412,0.2709374,0.41840968,0.45270553,0.0,0.0,0.037725464,0.072021335,0.09602845,0.12346515,0.12346515,0.048014224,0.07888051,0.216064,0.29151493,0.15433143,0.15090185,0.20920484,0.274367,0.274367,0.21263443,0.13375391,0.08573969,0.13032432,0.34981793,0.12003556,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.020577524,0.044584636,0.058302987,0.061732575,0.0548734,0.048014224,0.061732575,0.09602845,0.13375391,0.15090185,0.1371835,0.07545093,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.030866288,0.030866288,0.030866288,0.030866288,0.030866288,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.024007112,0.01371835,0.01371835,0.0274367,0.058302987,0.09602845,0.14747226,0.24350071,0.35324752,0.40126175,0.4115505,0.41498008,0.42869842,0.53844523,0.6001778,0.607037,0.5658819,0.5041494,0.45613512,0.31552204,0.15433143,0.041155048,0.030866288,0.07888051,0.06516216,0.05144381,0.08916927,0.19891608,0.22292319,0.1371835,0.044584636,0.006859175,0.030866288,0.041155048,0.1097468,0.20920484,0.30523327,0.36696586,0.4629943,0.5144381,0.65162164,0.94656616,1.4335675,1.9342873,2.2155135,2.369845,2.5207467,2.8396983,2.3732746,5.9571934,9.513676,11.640019,13.581166,9.650859,6.883182,5.223262,4.5922174,4.897451,5.2164025,5.5422134,5.1580997,4.557922,5.446185,6.217842,4.513337,2.2120838,0.58988905,0.31895164,0.19891608,0.15090185,0.17490897,0.2503599,0.33609957,0.6036074,0.9362774,0.97400284,0.7339317,0.6241849,0.7613684,1.0940384,1.5398848,1.978872,2.2566686,2.369845,2.3595562,2.335549,2.386993,2.5927682,2.4590142,2.9494452,3.4433057,3.7142432,3.9200184,6.166398,7.5725293,6.941485,4.605936,2.393852,2.1400626,2.2292318,2.2841053,2.0131679,1.2209331,1.7216529,2.4795918,3.350707,4.2389703,5.0826488,4.4447455,3.1140654,1.9308578,1.5947582,2.6545007,4.290414,6.001778,7.0203657,7.658269,9.294182,13.029003,15.333686,15.29939,12.754636,8.285883,4.0263357,2.0886188,1.1214751,0.490431,0.31895164,0.22292319,0.17833854,0.16804978,0.15090185,0.09259886,0.07888051,0.07545093,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.072021335,0.20577525,0.28465575,0.09602845,0.037725464,0.15090185,0.6276145,1.0837497,0.5658819,0.4115505,0.30523327,0.23321195,0.2777966,0.6241849,1.1900668,1.704505,1.704505,1.214074,0.7476501,1.2689474,1.3066728,0.90198153,0.34981793,0.18176813,0.36010668,0.5796003,0.7099246,0.6241849,0.20234565,0.29494452,0.7099246,1.786815,2.983741,2.877424,1.2586586,0.6276145,0.34638834,0.274367,0.77508676,0.61046654,0.72364295,1.8931323,3.426158,3.1655092,1.961724,1.138623,1.0631721,1.7079345,2.6750782,3.9783216,4.297273,3.450165,2.2429502,2.4555845,3.3952916,5.919468,9.132992,11.622872,11.454823,7.0752387,7.4044795,9.870353,12.569438,14.277372,9.9869585,9.14328,9.386781,9.211872,7.966932,6.142391,4.880303,4.413879,4.5339146,4.5956473,5.267846,7.5725293,9.4862385,9.054111,4.389872,3.4021509,3.3815732,3.5359046,4.0949273,6.307011,5.4667625,4.3590055,3.5633414,3.069481,2.287535,2.3424082,2.3081124,2.6647894,3.4192986,4.1189346,4.383013,4.1189346,3.8102717,4.1360826,5.950334,6.5950966,5.147811,3.415869,2.318401,1.8897027,2.0474637,1.488441,1.704505,2.5996273,2.4590142,2.4830213,2.7093742,2.8328393,2.74367,2.534465,2.9940298,3.5187566,3.6696587,3.3884325,3.0043187,2.5070283,2.318401,2.5996273,3.1106358,3.223812,2.942586,2.74367,2.3389788,1.6873571,0.9945804,0.8128122,0.9945804,1.4747226,1.845118,1.3615463,1.313532,0.9534253,0.5693115,0.45956472,0.9259886,1.2483698,1.3101025,1.8931323,3.2032347,4.8322887,6.975781,5.4187484,2.74367,0.65505123,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.037725464,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.061732575,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.041155048,0.041155048,0.030866288,0.037725464,0.1097468,0.1097468,0.07888051,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.048014224,0.08916927,0.020577524,0.006859175,0.09602845,0.20577525,0.12346515,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.006859175,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.01371835,0.017147938,0.010288762,0.01371835,0.072021335,0.072021335,0.030866288,0.030866288,0.06859175,0.048014224,0.010288762,0.0,0.0,0.030866288,0.14747226,0.072021335,0.058302987,0.59331864,1.6599203,2.726522,3.649081,4.0709205,3.923448,3.2443898,2.1674993,1.1866373,1.0151579,0.97057325,0.69963586,0.15776102,0.25721905,0.48700142,0.7613684,1.0220171,1.2312219,0.9877212,0.6859175,0.47671264,0.3841138,0.29151493,0.20577525,0.16804978,0.20234565,0.32238123,0.5178677,0.42869842,0.31209245,0.20920484,0.16119061,0.20577525,0.1097468,0.072021335,0.048014224,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.020577524,0.024007112,0.030866288,0.030866288,0.020577524,0.024007112,0.041155048,0.058302987,0.06859175,0.061732575,0.041155048,0.010288762,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.010288762,0.017147938,0.020577524,0.030866288,0.020577524,0.017147938,0.017147938,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.017147938,0.020577524,0.0274367,0.0274367,0.048014224,0.12003556,0.13032432,0.106317215,0.19548649,0.3841138,0.5453044,0.6241849,0.5796003,0.37725464,0.42869842,0.53844523,0.58645946,0.5418748,0.42869842,0.42183927,0.45270553,0.45956472,0.4046913,0.274367,0.12689474,0.07888051,0.07545093,0.116605975,0.2469303,0.39783216,0.37382504,0.24007112,0.09259886,0.06859175,0.06859175,0.08916927,0.13375391,0.19891608,0.28122616,0.37725464,0.42183927,0.48014224,0.5658819,0.65162164,0.9774324,1.214074,1.4644338,1.7730967,2.1297739,2.3389788,3.4844608,4.5819287,5.137522,5.144381,3.841138,3.1517909,2.7059445,2.5824795,3.2992632,3.9303071,3.9371665,4.0023284,4.1326528,3.6765177,3.5564823,3.806842,4.105216,3.8445675,2.1503513,0.7990939,0.34638834,0.2503599,0.2469303,0.36010668,0.5418748,0.83681935,1.1043272,1.214074,1.0666018,1.3546871,1.4953002,1.7525192,2.194936,2.7093742,2.8088322,2.6236343,2.386993,2.2841053,2.4247184,2.2292318,2.2052248,2.1880767,2.1640697,2.2738166,4.99005,7.864044,8.621983,6.8557453,4.029765,2.9048605,3.0077481,3.9303071,5.1580997,6.0532217,5.6656785,4.2081037,3.6559403,4.5647807,6.0703697,7.4353456,7.881192,7.4696417,6.574519,5.888602,5.4839106,5.4016004,5.254128,5.3707337,6.800872,9.942374,12.826657,15.121051,16.13621,14.791811,10.854645,6.917478,4.0503426,2.3629858,1.039165,0.53158605,0.29151493,0.21263443,0.19548649,0.16462019,0.10288762,0.07545093,0.048014224,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0274367,0.07888051,0.13032432,0.06516216,0.048014224,0.34638834,0.7510797,0.94999576,0.50757897,0.26064864,0.4698535,0.9602845,1.2106444,0.3566771,0.22635277,0.16119061,0.1920569,0.48014224,1.3169615,1.937717,3.2958336,3.1655092,1.6084765,0.9945804,2.0063086,2.0577524,1.5536032,0.9534253,0.7613684,0.8025235,0.8745448,0.85396725,0.65505123,0.22978236,0.2709374,0.5624523,1.2929544,2.1743584,2.435007,1.5844694,1.1317638,1.039165,1.6667795,3.7759757,2.0440342,1.3855534,1.5227368,1.8039631,1.2072148,0.65505123,0.36353627,0.35324752,0.607037,1.0871792,1.9068506,2.503599,2.6922262,2.74367,3.4021509,5.4839106,8.522525,9.39707,8.162418,8.049242,6.711703,8.251588,10.100135,10.590566,8.947794,8.351046,11.88352,13.985858,13.200482,12.195613,9.047252,7.3050213,6.420188,5.960623,5.627953,5.65539,6.1046658,6.550512,6.293293,4.3624353,4.40702,3.9303071,3.4535947,3.590778,5.0826488,4.938606,4.32128,3.7931237,3.5187566,3.2683969,3.2958336,3.0248961,3.2649672,3.882293,3.82399,4.0709205,3.5153272,2.9734523,3.1072063,4.4447455,4.4687524,3.4707425,2.5310357,2.1297739,2.1194851,2.0989075,1.7353712,1.9445761,2.6167753,2.627064,2.4898806,2.5001693,2.4590142,2.311542,2.1400626,2.9288676,4.105216,4.420738,3.9646032,4.166949,3.8308492,3.4124396,4.1429415,5.874883,7.0752387,6.7802944,6.4819202,6.1561093,5.7274113,5.0655007,6.608815,7.7680154,8.495089,8.601405,7.723431,7.6171136,6.8728933,6.3790326,6.9723516,9.462232,9.674867,8.48137,7.0375133,6.0737996,5.878313,8.1487,5.6348124,2.2978237,0.29837412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.006859175,0.0034295875,0.010288762,0.020577524,0.0,0.0034295875,0.0034295875,0.010288762,0.020577524,0.0,0.08916927,0.082310095,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0548734,0.0548734,0.041155048,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041155048,0.21263443,0.15090185,0.09945804,0.082310095,0.10288762,0.116605975,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.14061308,0.18176813,0.13032432,0.034295876,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.12689474,0.8779744,2.3286898,4.139512,6.1904054,7.3598948,7.5519514,6.831738,5.435896,3.8137012,2.5824795,1.5981878,0.91569984,0.7579388,1.039165,1.4129901,1.8485477,2.294394,2.6922262,2.3732746,2.1400626,2.085189,1.9651536,1.2243627,0.8711152,0.5041494,0.30523327,0.36010668,0.66191036,0.5144381,0.30523327,0.15090185,0.09602845,0.09602845,0.09945804,0.09602845,0.061732575,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.006859175,0.01371835,0.020577524,0.01371835,0.006859175,0.010288762,0.020577524,0.0274367,0.0274367,0.020577524,0.010288762,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.0034295875,0.01371835,0.020577524,0.01371835,0.01371835,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.041155048,0.048014224,0.05144381,0.082310095,0.082310095,0.06516216,0.09945804,0.2503599,0.45613512,0.59674823,0.61046654,0.5212973,0.6379033,0.64476246,0.6036074,0.5418748,0.44927597,0.4698535,0.5590228,0.6310441,0.6241849,0.51100856,0.3566771,0.274367,0.21263443,0.17490897,0.18519773,0.32581082,0.38754338,0.41840968,0.4046913,0.28808534,0.13375391,0.12689474,0.19891608,0.29494452,0.36010668,0.5007198,0.6859175,0.7579388,0.66191036,0.4664239,0.5727411,0.67219913,0.83338976,1.0254467,1.1283343,1.3375391,1.6496316,1.9582944,2.0714707,1.6804979,1.2380811,1.1146159,1.1111864,1.2860953,1.9548649,3.1346428,3.2581081,3.4192986,3.841138,3.865145,2.4555845,2.4555845,2.9906003,3.3609958,3.0386145,1.6153357,0.7888051,0.4938606,0.5418748,0.65162164,0.6756287,0.6893471,0.78537554,0.97400284,1.1763484,1.4164196,1.3924125,1.4472859,1.7490896,2.301253,2.867135,3.1826572,3.3541365,3.4981792,3.707384,3.450165,3.2546785,3.0146074,2.7093742,2.428148,3.9508848,6.6122446,7.747438,6.5196457,3.9371665,3.4947495,3.940596,5.953764,9.15014,12.079007,11.489118,9.071259,6.5710897,5.394741,6.619104,8.347616,10.158438,11.928105,13.179905,13.05301,11.177026,10.247607,10.076128,10.494537,11.362224,12.329367,13.138749,13.978998,14.7197895,14.898128,14.63062,14.634049,14.417986,12.895248,8.399059,2.976882,0.9945804,0.4664239,0.28465575,0.20920484,0.13032432,0.08573969,0.061732575,0.044584636,0.034295876,0.01371835,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.058302987,0.14747226,0.21263443,0.082310095,0.05144381,0.30866286,0.65162164,0.8093826,0.45613512,0.2469303,0.40126175,0.65848076,0.6824879,0.082310095,0.037725464,0.044584636,0.116605975,0.37382504,1.0220171,1.4267083,2.644212,2.568761,1.2312219,0.805953,1.99602,2.4761622,2.1091962,1.3924125,1.4747226,1.7525192,1.605047,1.2689474,0.9602845,0.864256,0.96371406,0.77508676,0.6927767,0.86082643,1.1592005,1.155771,1.097468,1.4335675,2.5447538,4.7534084,3.175798,2.8019729,2.2292318,1.2826657,0.99801,2.07833,1.8862731,1.0666018,0.24350071,0.017147938,0.50757897,2.3149714,3.474172,4.040054,6.118384,9.407358,12.3911,12.908967,11.183885,9.818909,8.97523,10.010965,11.039842,11.019264,9.753747,12.260776,15.354263,16.901007,16.362562,14.802099,11.135871,8.601405,7.455923,7.291303,7.0203657,6.2727156,5.693115,5.209543,4.9420357,5.195825,5.2918534,4.5167665,3.673088,3.2306714,3.3301294,3.8274195,4.2423997,4.184097,3.899441,4.2869844,4.9523244,4.9180284,4.822,4.729401,4.1120753,4.3281393,3.7348208,3.1380725,2.8637056,2.7539587,2.8122618,2.5721905,2.2395205,1.9411465,1.7319417,1.5021594,1.3958421,1.9651536,2.9803114,3.457024,2.5756202,2.311542,2.3321195,2.277246,1.7319417,2.4418662,3.3747141,3.9303071,4.1635194,4.7979927,4.5784993,3.7965534,4.2835546,6.3138704,8.601405,8.255017,7.864044,8.038953,8.553391,8.354475,9.97667,11.290202,11.952112,11.852654,11.122152,11.201033,10.789482,10.244178,10.302481,12.096155,12.024134,10.63858,8.501947,6.2692857,4.681387,5.501058,3.4364467,1.1523414,0.0,0.0,0.0,0.0548734,0.0548734,0.0,0.0,0.0,0.010288762,0.017147938,0.010288762,0.0,0.01371835,0.037725464,0.058302987,0.061732575,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.0,0.11317638,0.10288762,0.044584636,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05144381,0.2503599,0.3018037,0.16804978,0.044584636,0.010288762,0.0548734,0.14747226,0.18176813,0.11317638,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16119061,0.19548649,0.15090185,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.5521636,0.8025235,1.3649758,2.4761622,3.99204,6.6053853,8.690575,9.952662,10.254466,9.633711,7.8091707,5.874883,4.0263357,2.5756202,1.9480057,2.1812177,2.4247184,2.8054025,3.3026927,3.74168,3.6353626,4.029765,4.5956473,4.887162,4.3349986,3.6970954,2.6133456,1.5227368,0.7682276,0.5761707,0.37382504,0.18519773,0.07545093,0.05144381,0.05144381,0.07545093,0.07545093,0.041155048,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0034295875,0.01371835,0.006859175,0.01371835,0.020577524,0.01371835,0.0,0.0,0.010288762,0.01371835,0.01371835,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.006859175,0.017147938,0.020577524,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.010288762,0.024007112,0.048014224,0.072021335,0.048014224,0.041155048,0.041155048,0.041155048,0.041155048,0.14061308,0.33609957,0.48014224,0.5212973,0.4972902,0.6893471,0.70306545,0.6207553,0.5453044,0.59674823,0.6756287,0.72364295,0.7510797,0.7373613,0.65505123,0.5693115,0.48357183,0.39440256,0.29837412,0.20577525,0.23664154,0.29837412,0.41840968,0.5178677,0.3841138,0.16119061,0.15090185,0.23321195,0.32924038,0.40126175,0.548734,0.7990939,1.0940384,1.1900668,0.66876954,0.548734,0.52472687,0.53501564,0.51100856,0.41498008,0.5761707,0.8745448,1.0185875,0.89512235,0.5693115,0.33952916,0.26407823,0.31552204,0.53844523,1.0288762,2.2258022,2.5173173,2.5653315,2.7059445,2.9563043,1.6324836,1.4095604,1.6393428,1.9685832,2.3252604,1.4472859,0.89855194,0.6036074,0.5144381,0.6001778,0.66876954,0.5761707,0.52472687,0.64476246,1.0220171,1.2003556,1.1832076,1.1694894,1.2929544,1.6359133,2.3286898,2.9734523,3.6216443,4.290414,4.976331,5.192395,5.3261495,5.329579,5.15467,4.746549,5.439326,7.1232533,8.069819,7.723431,6.684266,7.040943,7.905199,11.012405,16.095055,20.886189,19.54179,16.04018,12.144169,9.338767,8.820899,9.39707,11.108434,13.920695,17.072487,19.044498,18.423744,18.03963,18.492336,19.737276,21.085104,20.76958,19.356592,17.566347,16.04361,15.337115,17.916164,22.669573,26.047716,25.44068,19.174824,10.851214,5.9983487,2.7745364,0.65505123,0.42526886,0.216064,0.13032432,0.09259886,0.06859175,0.05144381,0.0274367,0.017147938,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.06516216,0.1371835,0.16462019,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.15776102,0.40126175,0.5178677,0.4698535,0.38754338,1.2826657,2.2292318,2.1640697,1.4644338,1.9548649,2.7093742,2.6785078,2.2498093,1.8862731,2.1503513,2.352697,1.9925903,1.6530612,1.546744,1.5330256,1.6942163,1.6804979,2.1400626,3.0660512,3.8308492,3.9440255,4.715683,4.4275975,3.1963756,3.000889,4.722542,4.1326528,2.3835633,0.6344737,0.030866288,0.86082643,4.4413157,5.6210938,4.9248877,8.556821,10.89237,12.507706,13.958421,14.740367,13.2862215,12.277924,12.88839,13.605173,14.085316,15.151917,17.28512,16.269962,15.937293,16.300829,13.588025,10.813489,8.333898,7.3873315,7.750868,7.7577267,6.9792104,7.06838,6.8728933,6.193835,5.785714,5.8337283,5.147811,4.437886,3.8891523,3.1552205,3.858286,5.336438,5.7068334,5.0312047,5.3432975,7.085528,6.944915,5.7239814,4.482471,4.540774,4.5030484,3.5873485,2.9048605,2.6064866,1.8931323,2.633923,2.318401,1.7353712,1.2689474,0.89512235,0.6756287,0.66876954,1.9514352,3.99204,4.636802,2.5173173,1.9754424,2.2120838,2.3492675,1.4061309,1.7593783,1.8245405,2.4727325,3.590778,4.098357,3.9097297,3.0386145,2.8054025,3.875434,6.2692857,5.9571934,5.6245236,6.3447366,7.740579,7.9600725,7.956643,8.522525,8.848335,8.742019,8.632272,8.958082,9.3593445,8.923786,7.7028537,6.708273,6.509357,6.2898636,5.56965,4.40359,3.350707,2.6716487,2.1229146,1.4815818,0.83338976,0.5453044,0.45613512,0.6001778,0.70306545,0.7888051,1.2037852,1.371835,1.097468,0.65162164,0.28465575,0.20577525,0.29151493,0.32924038,0.274367,0.14747226,0.024007112,0.0034295875,0.020577524,0.048014224,0.061732575,0.041155048,0.048014224,0.12346515,0.18862732,0.20234565,0.14404267,0.12003556,0.07888051,0.041155048,0.010288762,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.13375391,0.30866286,0.14061308,0.0274367,0.07888051,0.12346515,0.48014224,0.5658819,0.33952916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.116605975,0.058302987,0.072021335,0.14747226,0.0,0.0,0.0,0.0,0.0,0.0,1.1043272,1.6221949,2.0749004,2.5584722,2.7230926,4.746549,7.2021337,9.496528,11.283342,12.46312,11.324498,9.616563,7.5519514,5.4976287,3.974892,3.9303071,3.9543142,4.249259,4.746549,5.120374,5.2609873,6.0669403,6.9689217,7.630832,7.963502,7.205563,5.456474,3.3987212,1.605047,0.53844523,0.22292319,0.09945804,0.09259886,0.11317638,0.061732575,0.082310095,0.0548734,0.020577524,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.01371835,0.020577524,0.020577524,0.010288762,0.0034295875,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.017147938,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.017147938,0.0274367,0.05144381,0.082310095,0.041155048,0.041155048,0.037725464,0.024007112,0.024007112,0.09945804,0.22978236,0.35324752,0.4081209,0.32581082,0.51100856,0.6344737,0.61389613,0.5555932,0.7613684,0.9259886,0.89855194,0.805953,0.7305021,0.70649505,0.64819205,0.58302987,0.52472687,0.4664239,0.37382504,0.29494452,0.28122616,0.32924038,0.39783216,0.37382504,0.20577525,0.17147937,0.18519773,0.22292319,0.31895164,0.4389872,0.65505123,1.1900668,1.6393428,0.9774324,0.7510797,0.65162164,0.5144381,0.31895164,0.1920569,0.3566771,0.7510797,0.8025235,0.4698535,0.2194936,0.14061308,0.09602845,0.08916927,0.17833854,0.48014224,1.1214751,1.4747226,1.4747226,1.2312219,1.0117283,0.7990939,0.864256,0.97400284,0.9534253,0.6824879,0.4355576,0.5555932,0.4664239,0.17490897,0.28465575,0.48014224,0.50757897,0.47671264,0.5007198,0.70649505,0.90541106,1.0185875,1.0425946,1.0220171,1.0494537,1.4164196,1.937717,2.6887965,3.683377,4.846007,5.830299,6.5950966,7.226141,7.6616983,7.689135,8.718011,9.856634,10.878652,11.835506,13.056439,13.96871,15.247946,18.87302,24.696459,30.451307,28.222075,23.739605,19.53836,16.592344,14.280802,13.210771,13.320518,14.826107,17.61779,21.253153,23.664154,24.43581,25.474976,27.464136,29.85113,30.122066,28.458717,25.756203,22.875349,20.635828,23.211449,29.305824,34.055805,34.4262,29.230373,22.158566,15.282242,8.488229,2.8877127,0.82996017,0.39097297,0.21263443,0.14061308,0.09602845,0.06859175,0.048014224,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.030866288,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.034295876,0.06859175,0.106317215,0.22978236,0.432128,0.7442205,1.1763484,1.7250825,2.2738166,3.216953,3.5770597,3.3850029,3.6765177,4.0434837,4.839148,5.6039457,6.060081,6.1321025,6.5470824,5.627953,5.0277753,5.2472687,5.6005163,5.442755,5.967482,6.2727156,6.0635104,5.662249,5.086078,3.2855449,1.6804979,0.77508676,0.15090185,0.44584638,3.7965534,4.173808,2.7093742,7.689135,3.5393343,1.8073926,2.7162333,5.120374,6.4990683,12.394529,16.743246,17.178804,13.687484,8.621983,6.584808,6.842027,7.531374,7.507367,6.3481665,6.9346256,7.6376915,7.606825,6.9037595,6.4990683,6.9037595,6.601956,6.0395036,5.5662203,5.4324665,7.130112,7.1129646,6.39961,5.4153185,3.998899,5.3158607,7.9875093,8.995808,7.932636,7.0032177,8.968371,7.8023114,5.24041,3.6147852,5.857735,5.470192,3.3678548,1.5673214,0.96371406,1.3443983,2.9048605,1.9308578,0.8471081,0.5521636,0.4424168,0.37039545,0.37039545,2.5893385,5.610805,4.4413157,1.2655178,0.37382504,0.274367,0.19891608,0.07545093,0.07545093,0.15090185,0.26064864,0.38754338,0.53501564,0.5212973,0.39097297,0.31895164,0.4081209,0.70306545,0.9602845,1.1694894,1.6016173,2.0886188,2.0131679,2.0508933,2.4075704,2.6956558,2.7985435,2.884283,3.2855449,3.4055803,3.2581081,2.935727,2.5927682,2.8259802,3.340418,3.7553983,4.046913,4.547633,4.962613,5.761707,5.5422134,4.1600895,2.7299516,2.2806756,2.4590142,2.9665933,3.9508848,6.025785,6.8557453,5.3707337,3.100347,1.3169615,1.039165,1.3066728,1.2723769,0.864256,0.28122616,0.0,0.0,0.09945804,0.23664154,0.30866286,0.19891608,0.2469303,0.6173257,0.94656616,1.0117283,0.71678376,0.34981793,0.20577525,0.12346515,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13375391,0.39097297,0.61046654,1.039165,1.0151579,0.5590228,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1729189,2.5447538,3.0866287,1.7079345,2.1126258,3.3850029,5.06893,7.1781263,10.192734,11.036412,10.319629,9.033533,7.8537555,7.1712675,6.9517736,7.2638664,7.9292064,8.659708,9.0644,8.831187,8.05953,7.4113383,7.2295704,7.5210853,6.910619,5.5147767,3.9954693,2.6133456,1.2209331,0.5727411,0.26407823,0.25378948,0.31895164,0.061732575,0.2194936,0.16804978,0.06859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.030866288,0.0548734,0.082310095,0.044584636,0.034295876,0.07545093,0.06516216,0.0,0.0,0.037725464,0.0548734,0.20920484,0.42526886,0.4115505,0.44927597,0.53158605,0.5727411,0.59331864,0.70306545,0.9328478,0.90884066,0.7133542,0.548734,0.7339317,0.58645946,0.4664239,0.4972902,0.6276145,0.64133286,0.6036074,0.5693115,0.47671264,0.4081209,0.5796003,0.432128,0.24007112,0.11317638,0.08916927,0.1371835,0.28465575,0.5693115,0.85396725,1.039165,1.039165,1.039165,0.85396725,0.6036074,0.38754338,0.29151493,0.082310095,0.041155048,0.041155048,0.037725464,0.061732575,0.14747226,0.12346515,0.06859175,0.041155048,0.07545093,0.26064864,0.607037,1.0528834,1.3786942,1.2209331,0.6344737,0.2503599,0.06859175,0.048014224,0.12346515,0.048014224,0.10288762,0.14061308,0.18519773,0.4424168,0.4046913,0.432128,0.4698535,0.45956472,0.34981793,0.66876954,0.8025235,0.77851635,0.67219913,0.61046654,0.78194594,0.9877212,1.1900668,1.4644338,2.0131679,3.0283258,4.197815,5.4736214,6.7391396,7.8126,9.925226,12.439114,14.990726,17.473747,20.049368,21.976797,23.760181,26.380386,30.228384,35.125835,33.990643,30.447878,27.01143,24.912523,24.106571,22.813616,20.814167,18.800999,17.87158,19.5315,22.703869,23.242313,23.948809,25.67732,27.313234,29.535606,31.325851,32.58794,33.218983,33.109238,32.951477,33.69227,34.851467,35.34533,33.476204,29.569902,25.10458,18.495766,9.911508,1.2826657,0.64819205,0.33266997,0.19891608,0.14404267,0.106317215,0.09602845,0.072021335,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.16462019,0.17147937,0.037725464,0.034295876,0.19548649,0.48357183,0.6276145,0.6036074,0.6241849,0.70649505,0.881404,0.85396725,0.6756287,0.7339317,0.96371406,1.4129901,1.9308578,2.4144297,2.7882545,3.0866287,2.9803114,2.6785078,2.2669573,1.6942163,1.4472859,1.6393428,1.7422304,1.6187652,1.4987297,1.5124481,1.0357354,0.5178677,0.28122616,0.50757897,1.2277923,1.8897027,1.5947582,1.2998136,3.8102717,5.195825,7.006647,8.858624,9.304471,5.8405876,8.056101,7.4353456,6.3138704,5.65539,5.0312047,7.9737906,8.39563,6.9620624,4.7362604,3.1860867,3.4776018,3.5530527,3.5564823,3.7519686,4.5099077,4.434457,3.6970954,3.234101,3.474172,4.3452873,5.3090014,7.39762,8.855195,8.652849,6.475061,8.107545,9.23245,8.608265,6.509357,4.722542,4.8905916,4.870014,4.184097,3.2478194,3.3952916,3.6559403,2.633923,1.6187652,1.255229,1.5261664,1.9171394,1.4335675,0.78194594,0.35324752,0.23664154,0.26064864,0.40126175,2.5824795,5.164959,2.9391565,0.88826317,0.33952916,0.28808534,0.24350071,0.26064864,0.29837412,0.2777966,0.26064864,0.25721905,0.22978236,0.29494452,0.2777966,0.22292319,0.19548649,0.26407823,0.31209245,0.34981793,0.42526886,0.5212973,0.53844523,0.66191036,0.85739684,1.0185875,1.1111864,1.1866373,1.2963841,1.313532,1.3101025,1.3649758,1.5673214,1.9171394,2.352697,2.9940298,3.8034124,4.5956473,5.099797,5.7822843,6.0737996,5.754848,4.9420357,4.9180284,4.6573796,4.386442,4.6127954,6.101236,7.7885933,8.093826,7.130112,5.535354,4.4447455,4.341858,3.5976372,2.620205,1.7388009,1.2312219,1.4953002,2.0508933,1.8588364,0.91227025,0.23664154,0.12689474,0.14404267,0.18862732,0.20234565,0.14404267,0.06859175,0.041155048,0.024007112,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06859175,0.034295876,0.0,0.0,0.0,0.07888051,0.12689474,0.08916927,0.01371835,0.072021335,0.0548734,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.061732575,0.048014224,0.0,0.0,0.0,0.2503599,0.6036074,0.5007198,0.89855194,0.7373613,0.33952916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19548649,0.6036074,1.1008976,1.646202,2.2841053,1.961724,1.6393428,2.4452958,3.5359046,2.0886188,1.5433143,1.8759843,3.6010668,6.276145,8.508806,10.367643,11.516555,12.123591,12.548861,13.347955,14.946142,15.9750185,15.741806,13.9309845,10.6145735,7.9120584,5.744559,4.180667,3.2203827,2.8122618,2.8465576,2.627064,2.170929,1.5604624,0.939707,0.607037,0.37382504,0.22635277,0.12346515,0.024007112,0.0548734,0.037725464,0.01371835,0.0034295875,0.01371835,0.030866288,0.037725464,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.020577524,0.020577524,0.024007112,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.030866288,0.05144381,0.08573969,0.12003556,0.106317215,0.07545093,0.044584636,0.020577524,0.01371835,0.010288762,0.010288762,0.072021335,0.18862732,0.31552204,0.26407823,0.39097297,0.52815646,0.6344737,0.7613684,0.9842916,0.90541106,0.6790583,0.4972902,0.61046654,0.6207553,0.4972902,0.4698535,0.5693115,0.64133286,0.50757897,0.548734,0.77508676,1.0220171,0.9568549,0.6859175,0.61389613,0.51100856,0.33266997,0.23664154,0.23664154,0.29837412,0.41498008,0.53158605,0.5624523,0.5727411,0.5453044,0.4938606,0.4629943,0.5212973,0.29494452,0.23321195,0.17490897,0.08916927,0.08573969,0.11317638,0.072021335,0.0274367,0.006859175,0.01371835,0.061732575,0.17833854,0.37039545,0.52815646,0.42869842,0.20234565,0.06859175,0.017147938,0.020577524,0.024007112,0.058302987,0.22978236,0.5144381,0.90541106,1.4061309,1.0666018,0.58645946,0.28122616,0.20920484,0.16804978,0.26064864,0.32581082,0.36353627,0.40126175,0.47671264,0.91227025,1.1694894,1.2620882,1.2723769,1.3443983,1.5158776,1.9548649,2.5824795,3.2786856,3.8925817,5.0483527,6.4098988,8.110974,10.179015,12.531713,15.9921665,19.675543,23.077694,26.00999,28.571894,31.624226,30.26268,26.02714,21.36633,19.641247,19.850452,19.181683,17.240536,14.4145565,11.866373,12.538571,12.284782,11.410237,11.087856,13.347955,16.595774,18.914175,20.635828,22.072824,23.516682,25.156025,26.767931,28.2598,29.374416,29.693369,28.424421,26.003132,22.12084,16.698662,9.873782,4.417309,1.5261664,0.4046913,0.23664154,0.17833854,0.274367,0.1920569,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.13375391,0.17147937,0.19548649,0.26064864,0.45613512,0.490431,0.274367,0.082310095,0.010288762,0.006859175,0.07545093,0.19891608,0.24007112,0.18519773,0.14061308,0.12689474,0.12003556,0.06859175,0.0,0.0,0.07888051,0.22292319,0.4046913,0.6001778,0.78194594,0.88826317,0.9259886,0.83681935,0.61046654,0.28808534,0.17833854,0.22292319,0.2469303,0.20920484,0.18176813,0.274367,0.20920484,0.09602845,0.061732575,0.23664154,0.59331864,0.7339317,0.9259886,1.4610043,2.6716487,4.4104495,5.8337283,7.0889573,8.018375,8.176137,9.0369625,8.81061,7.8263187,6.210983,3.8891523,5.1683884,5.7239814,5.5079174,4.6916757,3.6970954,3.6799474,3.309552,2.976882,2.976882,3.5016088,3.7965534,3.57363,3.2546785,3.1209247,3.3129816,3.3850029,4.3521466,5.439326,5.970912,5.3844523,6.1561093,6.6533995,6.2247014,4.9660425,3.7108135,3.1963756,3.625074,3.758828,3.5359046,4.0949273,4.07435,3.666229,3.1312134,2.6545007,2.3492675,2.8568463,1.978872,1.2415106,1.0666018,0.7613684,0.881404,1.1317638,2.3732746,3.542764,1.6290541,0.70306545,0.7305021,0.8745448,0.85396725,0.94656616,0.864256,0.6276145,0.42526886,0.31895164,0.25378948,0.21263443,0.15776102,0.1097468,0.082310095,0.08916927,0.09602845,0.09259886,0.09259886,0.10288762,0.13032432,0.18862732,0.25721905,0.31552204,0.36353627,0.4046913,0.42869842,0.432128,0.4698535,0.5727411,0.75450927,0.91912943,1.0906088,1.3752645,1.7662375,2.136633,2.411,2.7779658,3.175798,3.4467354,3.3232703,4.4927597,5.2918534,4.9180284,3.99204,4.57164,5.950334,6.4373355,6.327589,5.936616,5.579939,5.1855364,4.4756117,4.0229063,4.2286816,5.329579,5.1340923,4.770556,3.6147852,1.879414,0.59331864,0.1371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034295876,0.061732575,0.044584636,0.0,0.0,0.037725464,0.06516216,0.044584636,0.006859175,0.037725464,0.0274367,0.010288762,0.024007112,0.05144381,0.0,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.030866288,0.024007112,0.0,0.22635277,0.33266997,0.5007198,0.6790583,0.59331864,0.6893471,0.45270553,0.4629943,0.58645946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.082310095,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.25721905,0.7407909,1.4541451,3.0420442,6.7700057,8.237869,6.228131,4.149801,3.0900583,1.8073926,1.2826657,1.6359133,3.4055803,6.276145,9.074688,10.864933,12.096155,13.306799,14.627191,15.772673,16.979887,16.45516,14.023583,10.319629,6.7802944,4.8288593,3.5530527,2.6613598,2.0097382,1.6153357,1.9925903,2.3664153,2.3321195,1.8005334,1.0082988,0.5521636,0.44584638,0.30523327,0.072021335,0.034295876,0.0274367,0.01371835,0.006859175,0.0,0.006859175,0.058302987,0.05144381,0.037725464,0.030866288,0.010288762,0.0034295875,0.0,0.0,0.0,0.006859175,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.030866288,0.017147938,0.041155048,0.044584636,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.041155048,0.06516216,0.06516216,0.024007112,0.010288762,0.024007112,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.020577524,0.041155048,0.08573969,0.16462019,0.116605975,0.05144381,0.020577524,0.020577524,0.01371835,0.010288762,0.010288762,0.024007112,0.06859175,0.16119061,0.18519773,0.2503599,0.34638834,0.47671264,0.66876954,0.70649505,0.65505123,0.5418748,0.4629943,0.58988905,0.5796003,0.44584638,0.48014224,0.69963586,0.8505377,0.64819205,0.6173257,0.8505377,1.1934965,1.2277923,0.96714365,0.99801,0.96714365,0.72021335,0.32238123,0.4389872,0.5590228,0.6207553,0.64819205,0.7442205,0.70649505,0.6790583,0.6276145,0.5761707,0.607037,0.45613512,0.45956472,0.4664239,0.4081209,0.3018037,0.23321195,0.13375391,0.058302987,0.048014224,0.12689474,0.044584636,0.058302987,0.11317638,0.15090185,0.09945804,0.048014224,0.01371835,0.0034295875,0.0034295875,0.0,0.024007112,0.12689474,0.3806842,0.7922347,1.2826657,1.0425946,0.7579388,0.6344737,0.6344737,0.48014224,0.33266997,0.23321195,0.18176813,0.18862732,0.26750782,0.6241849,0.78537554,0.90541106,1.0528834,1.2312219,1.2586586,1.3066728,1.4267083,1.6393428,1.9342873,2.5413244,3.3266997,4.5613513,6.217842,7.9875093,10.257896,13.327377,16.317978,18.849012,21.04395,23.821915,23.69845,20.399187,15.402277,11.931535,11.993267,12.668896,11.900668,9.239308,5.857735,5.5113473,5.31929,4.746549,4.1463714,4.7774153,6.684266,7.956643,8.951223,10.237319,12.603734,15.035312,16.986746,18.893597,21.081675,23.749893,24.69303,23.986534,22.216867,19.589804,15.940722,11.173596,6.5299344,2.767677,0.50757897,0.2709374,0.37039545,0.37382504,0.28465575,0.16804978,0.1371835,0.058302987,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.13375391,0.17147937,0.19548649,0.26064864,0.45613512,0.48014224,0.19548649,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.034295876,0.037725464,0.058302987,0.09259886,0.09259886,0.274367,0.7305021,1.5021594,2.3424082,2.7230926,3.0969174,3.426158,3.8342788,4.6848164,6.5710897,6.931196,8.124693,9.047252,8.724871,6.293293,4.245829,4.887162,6.9037595,8.827758,9.040393,8.872343,8.704293,7.6342616,5.9914894,5.3673043,5.096367,4.4447455,3.6285036,2.860276,2.318401,1.9548649,1.8176813,2.0817597,2.627064,3.0626216,3.2306714,3.4707425,3.5016088,3.3541365,3.3644254,2.8054025,3.508468,3.9680326,3.9783216,4.6265135,4.3624353,4.623084,4.9420357,4.897451,4.1326528,3.8102717,2.8499873,2.2600982,2.0131679,1.039165,1.2758065,1.4404267,1.646202,1.6633499,0.90884066,1.0014396,1.2517995,1.2586586,1.1249046,1.4472859,1.3101025,0.980862,0.6893471,0.52815646,0.47328308,0.36696586,0.2194936,0.09602845,0.034295876,0.034295876,0.041155048,0.05144381,0.072021335,0.09602845,0.106317215,0.08573969,0.09259886,0.1097468,0.13032432,0.15433143,0.16462019,0.18176813,0.2194936,0.26750782,0.30866286,0.30866286,0.3018037,0.30866286,0.33609957,0.36696586,0.45613512,0.58988905,0.84367853,1.155771,1.3101025,2.4898806,3.4433057,3.333559,2.5584722,2.7642474,3.4295874,3.7451096,4.180667,4.863155,5.597087,5.305572,4.722542,4.48933,4.962613,6.193835,6.2384195,5.528495,3.858286,1.7902447,0.65848076,0.2194936,0.044584636,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07545093,0.09602845,0.048014224,0.048014224,0.07888051,0.06859175,0.034295876,0.0,0.0,0.0,0.0,0.024007112,0.061732575,0.048014224,0.030866288,0.058302987,0.048014224,0.0034295875,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.0548734,0.0548734,0.044584636,0.048014224,0.048014224,0.037725464,0.020577524,0.0034295875,0.0,0.0,0.0,0.09602845,0.20234565,0.06859175,0.24007112,0.33266997,0.4046913,0.47671264,0.52472687,0.65162164,0.48700142,0.6824879,0.9431366,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.024007112,0.037725464,0.15433143,0.4115505,0.082310095,0.0,0.0,0.010288762,0.0548734,0.2709374,0.7133542,1.6633499,4.2938433,10.666017,13.522863,10.693454,6.3824625,3.1449318,1.8725548,1.5741806,1.879414,3.333559,5.90575,9.009526,10.847785,12.05157,13.289652,14.54831,15.13134,15.854982,14.332246,10.943813,6.783724,3.6627994,2.4624438,2.0749004,2.1194851,2.301253,2.4212887,2.9700227,3.4433057,3.2855449,2.4247184,1.2689474,0.58988905,0.4938606,0.47328308,0.34981793,0.26407823,0.2469303,0.18862732,0.1097468,0.041155048,0.006859175,0.09945804,0.12346515,0.1371835,0.14061308,0.06516216,0.01371835,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.006859175,0.0,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.017147938,0.05144381,0.09259886,0.14747226,0.16119061,0.15433143,0.12689474,0.06859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.020577524,0.034295876,0.061732575,0.09602845,0.13375391,0.09259886,0.05144381,0.037725464,0.034295876,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.020577524,0.030866288,0.06859175,0.14061308,0.106317215,0.048014224,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.010288762,0.024007112,0.05144381,0.13375391,0.16462019,0.216064,0.33952916,0.5693115,0.5727411,0.5590228,0.52815646,0.53158605,0.6756287,0.7510797,0.6001778,0.5555932,0.72707254,0.9842916,0.8711152,0.84024894,0.9602845,1.1694894,1.2758065,1.0666018,1.0666018,1.0220171,0.8162418,0.45613512,0.59331864,0.66876954,0.6824879,0.69963586,0.8162418,0.71678376,0.6344737,0.58988905,0.5658819,0.5041494,0.39783216,0.42526886,0.48357183,0.48357183,0.3566771,0.24350071,0.1371835,0.07545093,0.082310095,0.15090185,0.0548734,0.05144381,0.058302987,0.041155048,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.024007112,0.15433143,0.39783216,0.6893471,0.6344737,0.64819205,0.7407909,0.7956643,0.5761707,0.33266997,0.18519773,0.09945804,0.072021335,0.1097468,0.274367,0.34981793,0.5041494,0.77508676,1.0666018,1.3684053,1.4850113,1.3786942,1.1832076,1.1832076,1.5364552,2.2738166,3.2306714,4.2081037,4.996909,5.9126086,7.857185,10.268185,12.672326,14.647768,15.745236,16.37285,14.760944,11.129011,7.6788464,6.40304,6.691125,6.6739774,5.528495,3.4638834,2.702515,2.6750782,2.8568463,2.8122618,2.1812177,2.428148,2.5138876,2.5653315,3.0351849,4.681387,6.5813785,8.532814,10.672876,13.306799,16.914726,19.46291,20.330595,20.21056,19.521212,18.427174,15.810398,11.550851,6.927767,3.1963756,1.5707511,0.9294182,0.6859175,0.5590228,0.42869842,0.34638834,0.1920569,0.12003556,0.06516216,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.01371835,0.06516216,0.15776102,0.23664154,0.19891608,0.51100856,1.1351935,1.9685832,2.6167753,2.4075704,1.9308578,1.9857311,2.194936,2.2395205,1.8554068,1.9754424,3.216953,5.73427,8.484799,9.211872,6.2041235,6.7700057,9.709162,13.087306,14.246507,13.906977,14.246507,12.740917,9.633711,7.939495,6.23156,4.461893,2.983741,1.9651536,1.3615463,1.1077567,0.980862,0.9294182,0.9534253,1.1249046,1.3066728,1.3958421,1.5707511,2.1126258,3.391862,3.0523329,4.0229063,4.804852,4.9008803,4.8322887,4.187526,4.605936,5.4496145,5.9331865,5.1580997,3.566771,3.1072063,2.9665933,2.4452958,0.9534253,1.1008976,1.0082988,0.66191036,0.34638834,0.65505123,1.3066728,1.5741806,1.4129901,1.2037852,1.7799559,1.5193073,1.1523414,0.83338976,0.64133286,0.5693115,0.4972902,0.32238123,0.1371835,0.01371835,0.01371835,0.017147938,0.08573969,0.22635277,0.33609957,0.20920484,0.09602845,0.061732575,0.072021335,0.10288762,0.12003556,0.12003556,0.14404267,0.16804978,0.18176813,0.17833854,0.15090185,0.13032432,0.1371835,0.16462019,0.1920569,0.2469303,0.30866286,0.3566771,0.39097297,0.42183927,0.5144381,0.5453044,0.72707254,1.0837497,1.4781522,1.6221949,1.9171394,2.5241764,3.4673128,4.636802,4.8014226,4.4275975,4.0434837,3.8308492,3.6319332,4.2595477,3.9474552,2.6236343,0.980862,0.5041494,0.31209245,0.18176813,0.07545093,0.0,0.0,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.106317215,0.09602845,0.09602845,0.15776102,0.13375391,0.06516216,0.0,0.0,0.0,0.017147938,0.024007112,0.034295876,0.09602845,0.020577524,0.116605975,0.14404267,0.072021335,0.07888051,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.01371835,0.020577524,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072021335,0.19548649,0.34981793,0.51100856,0.70649505,0.72707254,0.67219913,0.6379033,0.70649505,0.78537554,0.6379033,0.37725464,0.13375391,0.041155048,0.024007112,0.037725464,0.25721905,0.4938606,0.21263443,0.1371835,0.048014224,0.034295876,0.18862732,0.59331864,0.83681935,0.78194594,0.823101,0.8093826,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09602845,0.06859175,0.030866288,0.17147937,0.7476501,0.33952916,0.14747226,0.09259886,0.12346515,0.2194936,0.30523327,0.6756287,1.862266,4.979761,11.72233,14.925565,12.994707,8.923786,5.0826488,3.2066643,2.7711067,3.0969174,3.9783216,5.3330083,7.2158523,9.256456,11.002116,12.662037,13.941273,14.04759,14.2190695,12.751206,10.189304,7.181556,4.4996185,3.0729103,2.4418662,2.6236343,3.3266997,3.9646032,4.5030484,4.6402316,4.07435,2.901431,1.5776103,0.84367853,0.65162164,0.72707254,0.823101,0.70649505,0.6790583,0.53844523,0.34295875,0.16119061,0.0548734,0.15090185,0.25378948,0.35324752,0.37039545,0.14404267,0.05144381,0.01371835,0.0,0.0034295875,0.010288762,0.044584636,0.024007112,0.0034295875,0.006859175,0.024007112,0.030866288,0.020577524,0.006859175,0.0034295875,0.0,0.0,0.0,0.010288762,0.058302987,0.18176813,0.22292319,0.23321195,0.24007112,0.22292319,0.13375391,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.037725464,0.05144381,0.058302987,0.061732575,0.06859175,0.14404267,0.15090185,0.1097468,0.061732575,0.058302987,0.044584636,0.030866288,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.0274367,0.034295876,0.06859175,0.09259886,0.061732575,0.030866288,0.020577524,0.024007112,0.020577524,0.010288762,0.006859175,0.01371835,0.01371835,0.07545093,0.12346515,0.1920569,0.31209245,0.53844523,0.70306545,0.7305021,0.7133542,0.7339317,0.8676856,1.1317638,1.0014396,0.7990939,0.7476501,0.9602845,1.0014396,1.0871792,1.1214751,1.1146159,1.1797781,1.0871792,0.96714365,0.8162418,0.67219913,0.6310441,0.6790583,0.58302987,0.50757897,0.52472687,0.6173257,0.48700142,0.34981793,0.33609957,0.40126175,0.31552204,0.24350071,0.2194936,0.24007112,0.25721905,0.20920484,0.12346515,0.06516216,0.0548734,0.072021335,0.05144381,0.030866288,0.048014224,0.0548734,0.041155048,0.024007112,0.020577524,0.006859175,0.0,0.0,0.0,0.0034295875,0.01371835,0.048014224,0.10288762,0.14747226,0.18176813,0.29494452,0.41840968,0.45956472,0.31552204,0.15090185,0.09945804,0.082310095,0.058302987,0.044584636,0.061732575,0.106317215,0.24007112,0.44927597,0.65162164,1.2072148,1.6290541,1.611906,1.2586586,1.0837497,1.3409687,2.1469216,2.8328393,3.0900583,2.9494452,3.2889743,4.4241676,6.3378778,8.546532,10.124143,10.100135,10.854645,10.604284,9.132992,7.8023114,5.3330083,3.9337368,3.7005248,4.0777793,3.8479972,2.9048605,2.8122618,3.4364467,4.1189346,3.6627994,3.0351849,2.6545007,2.2738166,1.862266,1.6187652,2.1400626,3.4776018,5.2026844,7.4456344,10.906088,14.044161,16.273392,17.648657,18.310568,18.45461,17.178804,14.79524,11.626302,8.093826,4.7019644,2.6476414,1.5501735,1.0151579,0.7510797,0.5693115,0.40126175,0.34295875,0.25378948,0.11317638,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0274367,0.15776102,0.274367,0.2709374,0.07545093,0.0274367,0.07888051,0.30523327,0.5041494,0.19891608,0.3566771,0.78194594,1.9274281,3.1380725,2.6236343,3.07634,2.5481834,2.07833,2.7059445,5.4770513,6.931196,7.082098,7.298162,7.8983397,8.179566,7.164408,7.133542,6.9552035,6.166398,4.9591837,2.8705647,1.7079345,1.0425946,0.64133286,0.45613512,0.4081209,0.37725464,0.35324752,0.3566771,0.4424168,0.5658819,0.6310441,1.0460242,2.0714707,3.8308492,3.6970954,4.7431192,6.23156,7.459353,7.750868,5.2472687,3.6525106,2.609916,1.9480057,1.6770682,1.6290541,1.5981878,1.5810398,1.5021594,1.2209331,0.64819205,0.32924038,0.2503599,0.29151493,0.22978236,0.34981793,1.3512574,2.07833,2.2909644,2.6716487,1.7182233,0.9842916,0.490431,0.20577525,0.044584636,0.020577524,0.006859175,0.0,0.0,0.0,0.024007112,0.29494452,0.8265306,1.2072148,0.61046654,0.25721905,0.08573969,0.041155048,0.058302987,0.044584636,0.058302987,0.061732575,0.061732575,0.06859175,0.09259886,0.10288762,0.116605975,0.14747226,0.1920569,0.22978236,0.25378948,0.2777966,0.28465575,0.274367,0.274367,0.29837412,0.38754338,0.48014224,0.6241849,0.9774324,1.2209331,1.3992717,1.5536032,1.6942163,1.8176813,2.4007113,2.959734,3.3026927,3.3987212,3.3884325,2.7642474,1.99602,1.6359133,1.5398848,0.8711152,0.34638834,0.4698535,0.3841138,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09259886,0.12689474,0.072021335,0.0,0.0,0.1097468,0.2503599,0.31209245,0.15090185,0.09259886,0.030866288,0.0,0.0,0.0,0.0,0.06516216,0.09602845,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36696586,0.9842916,1.7456601,2.5619018,3.1483612,3.0660512,2.8225505,2.7539587,3.0351849,3.4398763,2.8088322,1.6770682,0.6173257,0.21263443,0.116605975,0.1920569,0.33266997,0.432128,0.39783216,0.5555932,0.23664154,0.0,0.34981793,1.7559488,1.1077567,0.91912943,0.7613684,0.47671264,0.18176813,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09945804,0.15433143,0.12346515,0.07545093,0.96714365,0.7407909,0.45956472,0.5007198,0.548734,0.4389872,0.61389613,1.6873571,4.1292233,8.255017,11.965831,13.296511,12.600305,10.251037,6.636252,5.3432975,7.0443726,7.6788464,6.1629686,4.3933015,5.6656785,8.169277,11.880091,15.621771,17.075916,14.5585985,12.394529,10.978109,10.251037,9.688584,8.309891,6.3447366,5.051782,4.8322887,5.2335505,5.442755,4.8322887,3.998899,3.0797696,1.786815,1.3958421,1.1694894,1.0666018,1.0597426,1.1454822,1.1077567,0.9431366,0.6790583,0.39783216,0.21263443,0.20234565,0.37382504,0.65848076,0.764798,0.16804978,0.15433143,0.061732575,0.0,0.010288762,0.044584636,0.082310095,0.0548734,0.024007112,0.024007112,0.061732575,0.08573969,0.072021335,0.041155048,0.01371835,0.0,0.0,0.0,0.006859175,0.048014224,0.18176813,0.037725464,0.010288762,0.010288762,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.017147938,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.10288762,0.14061308,0.10288762,0.030866288,0.030866288,0.07545093,0.1371835,0.15433143,0.044584636,0.034295876,0.041155048,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.017147938,0.030866288,0.0548734,0.061732575,0.0548734,0.048014224,0.061732575,0.037725464,0.020577524,0.010288762,0.0034295875,0.01371835,0.01371835,0.08916927,0.20577525,0.3566771,0.5658819,0.84367853,0.9877212,1.0185875,1.0254467,1.1592005,1.4027013,1.4472859,1.3924125,1.2415106,0.90198153,0.864256,1.0460242,1.1454822,1.1214751,1.2037852,1.4129901,1.3169615,1.0734608,0.84024894,0.77851635,0.9602845,0.91569984,0.70649505,0.50757897,0.5796003,0.5178677,0.31209245,0.17147937,0.18176813,0.29151493,0.42526886,0.31895164,0.1920569,0.13375391,0.12346515,0.08573969,0.048014224,0.024007112,0.01371835,0.01371835,0.01371835,0.006859175,0.017147938,0.048014224,0.061732575,0.048014224,0.017147938,0.0,0.0,0.0,0.01371835,0.024007112,0.07888051,0.13375391,0.061732575,0.037725464,0.08573969,0.116605975,0.106317215,0.106317215,0.12003556,0.18519773,0.18519773,0.106317215,0.044584636,0.034295876,0.041155048,0.06859175,0.12346515,0.19891608,0.39440256,0.7990939,1.1043272,1.2175035,1.2655178,1.4267083,1.6564908,1.9274281,2.1194851,2.061182,1.8897027,2.2395205,3.1552205,4.6779575,6.852316,7.133542,6.6431108,6.2658563,6.495639,7.4627824,6.094377,4.3692946,3.3815732,3.2992632,3.3712845,2.6167753,2.3252604,2.959734,4.173808,4.822,4.273266,4.4447455,4.6093655,4.2046742,2.8396983,2.4247184,1.7593783,1.762808,3.4364467,7.905199,9.966381,13.011855,16.21509,18.660385,19.332584,18.087645,16.492886,14.692352,12.562579,9.719451,6.375603,3.7176728,1.99602,1.1454822,0.77851635,0.66876954,0.66876954,0.6379033,0.4629943,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.041155048,0.041155048,0.01371835,0.0034295875,0.006859175,0.030866288,0.0548734,0.0548734,0.01371835,0.006859175,0.017147938,0.061732575,0.09945804,0.041155048,0.072021335,0.16462019,0.39783216,0.64133286,0.548734,0.64819205,0.85396725,2.170929,5.0003386,9.139851,9.55826,7.3118806,4.8734436,3.5290456,3.3678548,3.4021509,3.0866287,2.2909644,1.3443983,1.0528834,0.6173257,0.39440256,0.2469303,0.12689474,0.09259886,0.082310095,0.082310095,0.08916927,0.15776102,0.41840968,1.8176813,2.294394,2.0063086,1.4438564,1.4267083,2.0234566,3.07634,3.8445675,3.974892,3.5153272,4.1292233,3.5804894,3.415869,3.5359046,2.201795,1.9994495,1.6633499,1.4232788,1.4438564,1.8554068,1.2929544,0.6310441,0.2469303,0.16462019,0.09602845,0.07888051,0.2709374,0.42183927,0.4698535,0.5453044,0.36696586,0.22292319,0.20234565,0.26064864,0.22978236,0.08573969,0.020577524,0.0,0.0,0.0,0.0034295875,0.38754338,0.89512235,1.0837497,0.32924038,0.09259886,0.017147938,0.006859175,0.010288762,0.010288762,0.010288762,0.01371835,0.0274367,0.06516216,0.12689474,0.16804978,0.18176813,0.20234565,0.25721905,0.36353627,0.45613512,0.47671264,0.4389872,0.39783216,0.44584638,0.4698535,1.2998136,1.4438564,0.84367853,0.85396725,0.84367853,0.9328478,1.1180456,1.3615463,1.5707511,1.6496316,1.6633499,1.6633499,1.7113642,1.8862731,2.153781,2.1400626,1.7456601,1.0666018,0.39440256,0.24007112,0.20920484,0.16119061,0.22292319,0.7682276,0.69963586,0.53844523,0.36010668,0.22292319,0.13375391,0.08573969,0.12346515,0.216064,0.29151493,0.24350071,0.07888051,0.044584636,0.037725464,0.024007112,0.024007112,0.0548734,0.048014224,0.048014224,0.09602845,0.23321195,0.12346515,0.037725464,0.0,0.0,0.0,0.010288762,0.024007112,0.034295876,0.0548734,0.09602845,0.16462019,0.09602845,0.05144381,0.061732575,0.030866288,0.08573969,0.08573969,0.09259886,0.12689474,0.14747226,0.25378948,0.45613512,0.5727411,0.51100856,0.25721905,0.08916927,0.020577524,0.0,0.044584636,0.2194936,0.7373613,1.7662375,3.093488,4.396731,5.2747054,5.809721,6.1629686,5.953764,4.897451,2.8156912,1.3924125,0.7579388,0.5178677,0.45956472,0.5555932,0.14404267,0.048014224,0.06516216,0.08573969,0.07888051,0.22978236,0.106317215,0.0,0.06859175,0.34981793,0.32924038,0.42869842,0.490431,0.432128,0.25721905,0.36353627,0.50757897,0.34981793,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20577525,0.4389872,0.5555932,0.48700142,0.23321195,0.07545093,0.01371835,0.0034295875,0.01371835,0.01371835,0.25721905,0.58645946,0.7682276,0.70649505,0.4424168,0.7373613,0.6927767,0.8676856,1.3306799,1.6736387,1.2209331,0.9568549,1.4164196,3.0523329,6.2418494,12.199042,19.027351,22.899355,21.887627,15.951012,14.568888,15.820687,16.37971,14.160767,8.351046,5.3707337,5.2987127,6.6465406,8.361334,9.822338,9.856634,8.913498,9.338767,11.063849,11.605724,12.229909,13.649758,12.843805,9.685155,6.9552035,5.305572,4.962613,4.6608095,3.8514268,2.6647894,2.2360911,1.9239986,1.6256244,1.371835,1.3409687,1.2826657,1.1489118,1.0185875,1.0425946,1.4472859,1.4815818,1.9445761,2.1469216,1.8931323,1.4610043,0.9911508,0.53158605,0.24007112,0.16462019,0.22978236,0.20577525,0.09945804,0.037725464,0.08916927,0.23321195,0.31552204,0.2503599,0.12346515,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.010288762,0.037725464,0.006859175,0.017147938,0.034295876,0.0548734,0.072021335,0.08573969,0.034295876,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.037725464,0.10288762,0.18519773,0.26750782,0.31209245,0.08573969,0.041155048,0.058302987,0.07888051,0.106317215,0.0548734,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.020577524,0.017147938,0.017147938,0.024007112,0.037725464,0.030866288,0.020577524,0.010288762,0.0,0.0034295875,0.01371835,0.030866288,0.06859175,0.15776102,0.3566771,0.70649505,1.0357354,1.1934965,1.155771,1.039165,1.1660597,1.3101025,1.4267083,1.4438564,1.2792361,1.1351935,1.2689474,1.5227368,1.6976458,1.5604624,1.6016173,1.4507155,1.2655178,1.1420527,1.1214751,1.3821237,1.6907866,1.8313997,1.7353712,1.5090185,1.2106444,0.9842916,0.78194594,0.59674823,0.4115505,0.45956472,0.44927597,0.44927597,0.41498008,0.20920484,0.14061308,0.17147937,0.1371835,0.030866288,0.0034295875,0.01371835,0.01371835,0.024007112,0.048014224,0.061732575,0.048014224,0.017147938,0.0,0.0,0.0,0.030866288,0.11317638,0.14061308,0.106317215,0.12346515,0.23321195,0.29494452,0.2777966,0.29837412,0.6310441,0.72364295,0.8745448,0.89855194,0.7099246,0.32581082,0.20577525,0.12003556,0.072021335,0.06859175,0.11317638,0.18176813,0.29151493,0.5144381,0.83338976,1.1454822,1.7422304,2.318401,3.7005248,5.15467,4.389872,2.551613,2.0749004,2.702515,4.3109913,6.924337,8.357904,6.341307,4.8254294,5.5833683,8.217292,5.9640527,5.65539,4.8940215,3.6079261,4.091498,4.1155047,3.9268777,4.122364,4.8494368,5.7994323,5.9914894,5.641671,5.0174866,4.540774,4.7534084,3.9474552,2.428148,1.6221949,2.335549,4.7431192,5.0174866,8.032094,12.096155,15.913286,18.574646,19.263992,18.660385,17.243965,15.391989,13.358243,10.871792,8.032094,5.212973,2.8980014,1.6804979,0.91569984,0.67219913,0.65848076,0.6207553,0.35324752,0.28465575,0.15090185,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.01371835,0.017147938,0.18176813,0.99801,2.585909,4.698535,5.1238036,3.9097297,2.4075704,1.5193073,1.6907866,2.3046827,1.8142518,0.89855194,0.15090185,0.06859175,0.05144381,0.041155048,0.0274367,0.010288762,0.010288762,0.0034295875,0.0034295875,0.006859175,0.048014224,0.1920569,1.2312219,2.0337453,2.287535,2.0097382,1.546744,1.6324836,2.0131679,2.352697,2.469303,2.3561265,3.4467354,4.314421,4.3007026,3.4295874,2.369845,2.1846473,1.6942163,1.3272504,1.2072148,1.1249046,0.72707254,0.33952916,0.14404267,0.12346515,0.08916927,0.024007112,0.0034295875,0.0034295875,0.006859175,0.006859175,0.010288762,0.01371835,0.072021335,0.15776102,0.12689474,0.058302987,0.09259886,0.14404267,0.14404267,0.0548734,0.010288762,0.18176813,0.39783216,0.44927597,0.10288762,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.06516216,0.1097468,0.1371835,0.1371835,0.15776102,0.20577525,0.26750782,0.31895164,0.42183927,0.5212973,0.5693115,0.53501564,0.6379033,1.0357354,1.0734608,0.8128122,1.0151579,0.9362774,0.85396725,0.83681935,0.88826317,0.9431366,0.91569984,0.8505377,0.78194594,0.7510797,0.7888051,0.939707,0.980862,0.805953,0.45956472,0.15433143,0.10288762,0.06516216,0.07888051,0.18176813,0.44927597,0.4081209,0.5007198,0.6927767,1.097468,1.961724,2.7368107,2.8396983,2.3664153,1.6084765,1.0666018,1.4507155,1.6770682,1.3169615,0.548734,0.16804978,0.14747226,0.17147937,0.1920569,0.20577525,0.24350071,0.14061308,0.09602845,0.082310095,0.07888051,0.06516216,0.06859175,0.09259886,0.16119061,0.3018037,0.5418748,0.51100856,0.42526886,0.25378948,0.061732575,0.017147938,0.12003556,0.28808534,0.44584638,0.5007198,0.3566771,0.31552204,0.3841138,0.4424168,0.4081209,0.25721905,0.072021335,0.010288762,0.0,0.50757897,2.534465,4.338428,5.5559316,7.023795,8.570539,9.009526,7.7542973,6.138962,4.417309,2.7573884,1.2346514,0.51100856,0.16462019,0.1097468,0.22978236,0.3841138,0.14404267,0.034295876,0.0,0.0,0.0,0.058302987,0.030866288,0.0,0.0,0.0,0.274367,0.6893471,0.96371406,0.980862,0.7682276,1.0357354,0.91912943,0.52472687,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10288762,0.5555932,0.9259886,0.96714365,0.6207553,0.5796003,0.53844523,0.4115505,0.20577525,0.05144381,0.17490897,0.37382504,0.6756287,0.9774324,1.0563129,1.0940384,1.3238207,1.862266,2.534465,2.867135,2.6167753,3.309552,4.90431,7.4353456,11.008976,16.516893,20.728426,21.829325,19.442331,14.599753,12.339656,11.72233,12.236768,12.850664,12.010415,9.678296,7.6616983,6.1766872,5.518206,6.060081,5.610805,4.962613,5.6793966,7.613684,8.9100685,9.716022,10.851214,10.371073,8.22758,6.2487082,5.3158607,5.096367,4.698535,3.8857226,3.0386145,2.6819375,2.6613598,2.4658735,1.9857311,1.5364552,1.5913286,1.488441,1.6187652,2.0508933,2.5413244,2.74367,3.3438478,3.9474552,4.3109913,4.338428,3.4913201,2.3458378,1.5021594,1.0220171,0.45613512,0.39097297,0.39440256,0.274367,0.08916927,0.12689474,0.26407823,0.26064864,0.19891608,0.13032432,0.06859175,0.020577524,0.0034295875,0.0,0.0,0.0,0.006859175,0.0274367,0.07545093,0.13375391,0.16462019,0.14061308,0.25721905,0.2777966,0.15776102,0.06516216,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.09602845,0.17490897,0.22635277,0.2709374,0.17490897,0.15433143,0.17833854,0.2194936,0.26064864,0.16119061,0.06516216,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.006859175,0.017147938,0.020577524,0.020577524,0.017147938,0.01371835,0.010288762,0.010288762,0.006859175,0.006859175,0.034295876,0.14404267,0.39783216,0.66876954,0.83338976,0.9294182,1.0117283,1.1351935,1.0425946,1.0323058,1.0631721,1.0837497,1.0357354,1.1043272,1.3649758,1.646202,1.7971039,1.6667795,1.6153357,1.5433143,1.430138,1.2689474,1.0597426,1.1489118,1.529596,1.8073926,1.8416885,1.7490896,1.5055889,1.2860953,1.2175035,1.2346514,1.0666018,0.8128122,0.6241849,0.5624523,0.52472687,0.23664154,0.16462019,0.16804978,0.13375391,0.05144381,0.010288762,0.0274367,0.044584636,0.058302987,0.072021335,0.106317215,0.06516216,0.0274367,0.017147938,0.030866288,0.037725464,0.09602845,0.24007112,0.33266997,0.32924038,0.28465575,0.32924038,0.28465575,0.20234565,0.20234565,0.48014224,1.3958421,1.7902447,1.670209,1.1900668,0.6790583,0.3566771,0.17833854,0.08573969,0.05144381,0.082310095,0.11317638,0.16804978,0.31552204,0.5693115,0.90198153,1.4575747,2.0817597,3.1483612,4.2423997,4.1600895,2.9254382,2.1263442,1.8999915,2.5824795,4.681387,6.944915,5.90232,4.4996185,4.763697,7.795452,5.161529,4.57507,4.417309,4.2595477,4.8322887,4.866585,4.5099077,4.4584637,4.962613,5.813151,6.0806584,5.9469047,5.439326,4.7774153,4.355576,3.6936657,2.49331,1.6427724,1.6290541,2.5619018,2.719663,4.7259717,8.004657,11.89038,15.63206,18.193962,19.79901,19.95334,18.608942,16.170506,13.900118,11.664027,9.273604,6.8557453,4.863155,3.2786856,2.2155135,1.587899,1.2312219,0.90198153,0.6893471,0.38754338,0.15433143,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.12003556,0.3566771,0.6790583,1.0357354,0.9602845,0.70306545,0.5590228,0.89855194,1.4061309,1.0906088,0.5693115,0.20920484,0.1097468,0.106317215,0.09259886,0.06516216,0.034295876,0.010288762,0.0034295875,0.0,0.0,0.006859175,0.0274367,0.3806842,0.94999576,1.3958421,1.5227368,1.2723769,1.0323058,0.97400284,1.0906088,1.3306799,1.605047,2.2292318,3.2306714,3.2546785,2.411,2.2600982,2.3458378,2.1229146,1.8519772,1.5844694,1.155771,0.70649505,0.3806842,0.22978236,0.19891608,0.12003556,0.030866288,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.020577524,0.048014224,0.017147938,0.017147938,0.08573969,0.14404267,0.14747226,0.061732575,0.01371835,0.017147938,0.030866288,0.030866288,0.006859175,0.006859175,0.037725464,0.08916927,0.13375391,0.13375391,0.17490897,0.16119061,0.12003556,0.07545093,0.061732575,0.06859175,0.06516216,0.08916927,0.16804978,0.30523327,0.6379033,0.77851635,0.71678376,0.548734,0.48357183,0.71678376,0.881404,0.91227025,0.9259886,1.2243627,1.0906088,0.7888051,0.5521636,0.45270553,0.4046913,0.39783216,0.37382504,0.32924038,0.274367,0.20920484,0.15433143,0.12003556,0.10288762,0.08573969,0.044584636,0.017147938,0.010288762,0.034295876,0.072021335,0.06859175,0.072021335,0.2503599,0.53501564,1.0631721,2.1469216,3.1449318,3.4810312,3.3438478,3.0420442,3.0043187,3.758828,4.437886,4.0366244,2.7813954,2.1503513,2.1434922,2.136633,2.0920484,1.9925903,1.8313997,1.3581166,0.90198153,0.6344737,0.6173257,0.8093826,0.7956643,0.64476246,0.65505123,0.881404,1.1420527,0.8848336,0.70649505,0.5727411,0.432128,0.20577525,0.23321195,0.64476246,1.0048691,1.3821237,2.352697,1.7559488,1.3752645,1.0323058,0.8265306,1.1214751,0.7922347,1.3786942,2.9974594,5.6828265,9.369633,8.491658,8.800322,10.199594,11.677745,11.327928,8.333898,5.0003386,2.277246,0.65848076,0.15776102,0.16462019,0.07888051,0.034295876,0.061732575,0.12689474,0.33952916,0.23321195,0.07545093,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24350071,0.7099246,1.1489118,1.3752645,1.2826657,1.5981878,1.4027013,1.0494537,0.66191036,0.17833854,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33609957,0.8745448,1.2758065,0.97400284,1.0528834,1.1351935,0.9294182,0.48014224,0.16119061,0.09259886,0.10288762,0.30523327,0.66876954,1.0014396,1.0185875,1.3066728,1.9514352,2.719663,3.059192,3.566771,5.144381,8.011517,11.396519,13.543441,15.450292,15.45715,13.910407,11.547421,9.510246,7.438775,5.9160385,6.3893213,8.954653,12.3533745,12.22648,9.3079,6.4236174,5.055212,5.360445,5.164959,4.602506,4.479041,4.98662,5.7102633,5.9434752,5.8165803,5.2918534,4.5819287,4.1326528,4.273266,4.064061,3.6970954,3.391862,3.3815732,3.223812,3.508468,3.6353626,3.3541365,2.7745364,2.5619018,2.2223728,2.3218307,2.884283,3.3781435,3.8308492,5.1100855,6.6636887,7.7680154,7.5245147,6.392751,4.7534084,3.4295874,2.469303,1.1592005,0.8505377,0.8162418,0.6790583,0.39097297,0.24350071,0.2709374,0.34638834,0.4115505,0.44584638,0.45613512,0.32924038,0.12346515,0.0034295875,0.0034295875,0.017147938,0.16119061,0.36696586,0.6036074,0.7922347,0.7922347,0.66191036,0.7682276,0.78194594,0.5658819,0.1920569,0.16119061,0.061732575,0.01371835,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.10288762,0.17490897,0.20234565,0.216064,0.28122616,0.29151493,0.29151493,0.28122616,0.216064,0.16804978,0.07888051,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.01371835,0.0274367,0.030866288,0.024007112,0.010288762,0.0034295875,0.0,0.030866288,0.12689474,0.33609957,0.5144381,0.5555932,0.59674823,0.72021335,0.9534253,0.86082643,0.8093826,0.8196714,0.85739684,0.85739684,1.1146159,1.5330256,1.8656956,1.9480057,1.7147937,1.5844694,1.605047,1.587899,1.4335675,1.1249046,1.0837497,1.3409687,1.6084765,1.8005334,2.0063086,2.1126258,1.9068506,1.7696671,1.7525192,1.6153357,1.2037852,0.9431366,0.89512235,0.90541106,0.6173257,0.42183927,0.32238123,0.29151493,0.26407823,0.16119061,0.12689474,0.12689474,0.12689474,0.12003556,0.12346515,0.09259886,0.07545093,0.08916927,0.13032432,0.17147937,0.24007112,0.36010668,0.45956472,0.47328308,0.34981793,0.274367,0.17147937,0.09945804,0.09945804,0.20577525,1.1214751,1.6084765,1.7113642,1.5261664,1.2037852,0.65848076,0.36696586,0.19891608,0.106317215,0.106317215,0.14061308,0.23321195,0.32238123,0.432128,0.65162164,1.1351935,1.6084765,2.1023371,2.609916,3.0969174,2.836269,2.270387,1.6907866,1.5501735,2.4830213,4.3281393,4.256118,3.5702004,3.6559403,5.9812007,3.8342788,3.1277838,3.350707,3.974892,4.4584637,4.955754,4.979761,4.8905916,4.9934793,5.56965,5.9160385,6.118384,6.0737996,5.6965446,4.8905916,4.0537724,2.8122618,1.7971039,1.3306799,1.4267083,1.6907866,2.627064,4.5442033,7.3873315,10.741467,13.756075,17.353712,19.929333,20.522652,18.825006,16.417435,14.2533655,12.319078,10.64201,9.290752,7.366754,5.4736214,3.8617156,2.633923,1.7388009,1.1694894,0.66533995,0.31209245,0.13032432,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.14747226,0.16462019,0.20920484,0.23664154,0.22292319,0.14747226,0.15776102,0.15433143,0.12003556,0.058302987,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.05144381,0.1097468,0.07888051,0.044584636,0.072021335,0.20920484,0.4629943,0.64133286,0.6824879,0.8025235,1.1111864,1.6496316,1.99602,2.2326615,2.1983654,1.9445761,1.7113642,1.1420527,0.64819205,0.36696586,0.25721905,0.1097468,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0034295875,0.01371835,0.044584636,0.09945804,0.19891608,0.29494452,0.35324752,0.35324752,0.30866286,0.36696586,0.32924038,0.21263443,0.072021335,0.01371835,0.01371835,0.024007112,0.12003556,0.36353627,0.8128122,1.4061309,1.3615463,0.89855194,0.42526886,0.53844523,0.9911508,1.4095604,1.4541451,1.2175035,1.2346514,1.0906088,0.6207553,0.2709374,0.17147937,0.14747226,0.14061308,0.12346515,0.09945804,0.07888051,0.048014224,0.030866288,0.017147938,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.034295876,0.044584636,0.058302987,0.16462019,0.53844523,0.96371406,1.5193073,2.3904223,3.549623,4.722542,5.353586,6.327589,6.4579134,5.6005163,4.6436615,5.127233,5.192395,5.188966,5.24041,5.2747054,4.6676683,3.690236,2.901431,2.620205,2.8945718,2.6750782,1.9651536,1.5433143,1.6599203,2.0406046,1.3684053,1.0425946,1.0425946,1.1283343,0.8505377,0.980862,1.7147937,2.3492675,3.2821152,6.029215,5.593657,4.8734436,3.8342788,3.223812,4.5647807,4.705394,5.9812007,8.447074,11.571428,14.222499,9.318189,8.577398,9.935514,11.413667,11.122152,7.9292064,4.664239,2.2052248,0.8676856,0.39440256,0.31552204,0.14747226,0.030866288,0.0,0.0,0.50757897,0.4081209,0.15433143,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.28808534,0.7133542,1.155771,1.3066728,1.4918705,1.5604624,1.5604624,1.2998136,0.35324752,0.22292319,0.07545093,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4664239,1.1214751,0.939707,1.0460242,1.214074,1.0425946,0.5727411,0.2777966,0.116605975,0.030866288,0.0,0.06516216,0.31895164,0.4355576,0.5761707,1.0563129,1.7765263,2.2223728,3.3712845,4.9420357,7.905199,10.971251,10.597425,8.707723,6.975781,5.751418,5.284994,5.744559,5.0655007,3.8171308,3.957744,6.125243,9.616563,11.026124,8.539673,6.0566516,5.3501563,6.0395036,7.239859,6.948344,6.036074,5.1821065,4.8597255,3.9954693,2.8705647,1.9925903,1.6393428,1.8416885,2.2909644,2.0989075,2.0646117,2.5721905,3.566771,3.6970954,4.0023284,4.338428,4.513337,4.280125,3.6696587,3.0729103,2.9974594,3.4707425,4.0503426,4.955754,7.390761,9.897789,11.101575,9.736599,8.008087,6.138962,4.6436615,3.457024,1.9239986,1.3169615,1.1249046,1.0837497,0.9945804,0.7099246,0.45613512,0.52472687,0.6927767,0.83681935,0.9259886,0.6824879,0.31895164,0.17833854,0.33266997,0.59331864,1.1797781,1.7559488,2.335549,2.8396983,3.0729103,2.9734523,2.8054025,2.5173173,1.9239986,0.72364295,0.41498008,0.15090185,0.0548734,0.09259886,0.05144381,0.0274367,0.020577524,0.017147938,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.1097468,0.18862732,0.23321195,0.23321195,0.33609957,0.33952916,0.29151493,0.19548649,0.020577524,0.061732575,0.044584636,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.037725464,0.048014224,0.030866288,0.0034295875,0.0,0.0,0.017147938,0.058302987,0.13375391,0.28465575,0.36353627,0.41498008,0.47671264,0.5590228,0.65505123,0.72364295,0.8128122,0.90541106,0.9294182,1.2758065,1.7936742,2.1400626,2.1160555,1.6599203,1.611906,1.6804979,1.6393428,1.4335675,1.1797781,1.1626302,1.2792361,1.4987297,1.8142518,2.2395205,2.7299516,2.5584722,2.1743584,1.8313997,1.6084765,1.3032433,1.2003556,1.3066728,1.430138,1.1866373,0.9602845,0.805953,0.75450927,0.7373613,0.5693115,0.4046913,0.29837412,0.24007112,0.20234565,0.1371835,0.16462019,0.21263443,0.2709374,0.32581082,0.36353627,0.4081209,0.41840968,0.42183927,0.39097297,0.26407823,0.1371835,0.072021335,0.06516216,0.08916927,0.08573969,0.17490897,0.5007198,1.0014396,1.546744,1.9411465,1.2929544,0.8265306,0.4972902,0.28122616,0.19891608,0.22978236,0.41840968,0.53844523,0.5418748,0.5590228,1.0494537,1.3752645,1.7730967,2.301253,2.8225505,2.620205,2.4624438,2.16064,1.762808,1.5638919,2.07833,2.0920484,2.1503513,2.6545007,3.858286,2.9940298,2.8088322,2.9220085,3.1346428,3.391862,4.3590055,5.0483527,5.1683884,5.038064,5.56965,5.936616,6.3173003,6.824879,7.2467184,7.0478024,5.8543057,4.2355404,2.8568463,1.937717,1.2586586,1.1832076,1.4061309,2.1263442,3.4124396,5.195825,7.160979,11.410237,16.184223,19.86417,20.982216,18.893597,16.235666,14.054449,12.919256,12.919256,11.684605,9.6817255,7.438775,5.329579,3.5839188,2.417859,1.5536032,0.9362774,0.53158605,0.31552204,0.17833854,0.07545093,0.017147938,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.034295876,0.0548734,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.12689474,0.20920484,0.23664154,0.19891608,0.08916927,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.06859175,0.20920484,0.4424168,0.9294182,1.0906088,0.864256,0.42869842,0.19891608,0.09945804,0.041155048,0.010288762,0.0034295875,0.01371835,0.0034295875,0.0548734,0.3841138,1.08032,2.1057668,1.8005334,1.1283343,0.6241849,0.61046654,1.2209331,2.1229146,2.4795918,2.136633,1.3546871,0.7922347,0.91569984,0.4972902,0.15433143,0.08573969,0.061732575,0.037725464,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.034295876,0.05144381,0.08573969,0.18176813,0.31895164,0.5693115,1.1077567,1.9548649,2.9906003,3.309552,3.799983,4.8905916,5.5490727,3.2649672,5.377593,6.0806584,6.715132,7.8606143,9.338767,10.508256,10.179015,9.009526,7.706283,7.034084,6.0703697,4.280125,2.7299516,2.311542,3.7382503,2.2738166,2.0440342,2.0131679,1.937717,2.3664153,3.4021509,4.605936,5.672538,6.958633,9.458802,12.315649,12.281353,10.497967,9.434795,12.878101,15.87899,16.11906,12.236768,5.871454,1.6496316,1.3924125,1.9582944,3.4535947,5.7754254,8.604835,7.936065,6.9689217,5.4941993,3.590778,1.6633499,1.5158776,0.59331864,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041155048,0.14747226,0.30523327,0.061732575,0.4115505,0.8196714,0.8162418,0.0,0.7682276,0.3841138,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.072021335,0.0,0.09602845,0.048014224,0.0,0.044584636,0.22978236,0.106317215,0.030866288,0.0,0.0,0.0,0.19548649,0.32581082,0.52815646,0.8779744,1.4027013,1.6839274,2.2052248,3.069481,4.0777793,4.698535,5.212973,5.751418,6.046363,6.159539,6.4990683,6.8283086,5.099797,4.07435,4.9420357,7.3084507,8.457363,7.9086285,6.4887795,5.1855364,5.171818,5.9434752,6.15268,6.4579134,7.1026754,7.932636,4.8837323,2.8019729,1.5913286,1.0494537,0.85396725,0.805953,0.82996017,1.0323058,1.6153357,2.884283,3.2855449,3.1037767,2.9322972,3.059192,3.450165,3.3369887,3.2478194,3.5461934,4.2218223,4.866585,6.711703,9.945804,12.240198,12.260776,9.674867,6.2075534,4.012617,2.726522,1.99602,1.4953002,1.0563129,0.96371406,1.2277923,1.5398848,1.2963841,0.69963586,0.59674823,0.78537554,0.9602845,0.71678376,0.33952916,0.41840968,0.85739684,1.6324836,2.7916842,4.341858,5.305572,6.217842,7.346176,8.711152,9.235879,8.735159,7.534804,5.5559316,2.335549,0.7476501,0.21263443,0.15776102,0.19891608,0.1371835,0.11317638,0.106317215,0.08916927,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06859175,0.14404267,0.19548649,0.18176813,0.20920484,0.21263443,0.19548649,0.14404267,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.024007112,0.01371835,0.01371835,0.0034295875,0.0,0.006859175,0.024007112,0.061732575,0.28122616,0.3806842,0.45613512,0.53501564,0.59674823,0.6927767,0.75450927,0.77851635,0.8093826,0.9294182,1.4815818,1.9823016,2.0646117,1.6976458,1.2209331,1.7593783,1.8176813,1.3478279,0.65505123,0.4115505,0.51100856,0.7442205,1.0185875,1.313532,1.6770682,2.020027,1.9685832,1.6324836,1.1694894,0.77851635,0.71678376,0.89512235,1.1797781,1.3821237,1.2346514,1.6153357,1.6530612,1.5501735,1.4267083,1.3272504,0.9842916,0.6173257,0.40126175,0.34638834,0.26064864,0.34638834,0.4938606,0.6173257,0.6310441,0.47328308,0.45956472,0.33952916,0.19891608,0.106317215,0.106317215,0.09602845,0.072021335,0.06859175,0.08573969,0.12346515,0.12346515,0.14061308,0.25721905,0.90198153,2.867135,2.4658735,1.6873571,1.0288762,0.65162164,0.3806842,0.34638834,0.8025235,1.155771,1.1454822,0.84024894,1.1934965,1.6770682,2.767677,4.1772375,4.835718,3.1415021,2.7333813,2.5619018,2.2360911,2.0303159,1.9068506,1.8485477,2.1915064,2.942586,3.782835,4.554492,4.588788,4.2183924,3.7725463,3.6010668,2.952875,3.2032347,3.8891523,4.8254294,6.118384,5.65539,6.1149545,7.2878733,8.56025,8.927217,8.340756,7.6274023,6.368744,4.40702,1.8313997,1.0631721,0.8711152,0.9842916,1.1934965,1.3272504,1.961724,4.722542,9.647429,15.803539,21.287449,21.297739,18.818146,15.731518,13.406258,12.710052,13.625751,13.104454,11.773774,9.993818,7.857185,5.8817425,4.2423997,2.867135,1.7799559,1.0837497,0.7888051,0.37725464,0.09259886,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.041155048,0.048014224,0.041155048,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.030866288,0.010288762,0.0034295875,0.020577524,0.048014224,0.09602845,0.09602845,0.1097468,0.116605975,0.0,0.06859175,0.19548649,0.25378948,0.20920484,0.15090185,0.26750782,0.28808534,0.2194936,0.106317215,0.041155048,0.020577524,0.006859175,0.006859175,0.01371835,0.01371835,0.072021335,0.77165717,1.2380811,1.1729189,0.86082643,0.58645946,0.42526886,0.51100856,0.7990939,1.097468,1.2003556,1.2312219,1.1660597,1.0460242,0.96371406,0.52815646,0.22292319,0.061732575,0.017147938,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0034295875,0.01371835,0.09259886,0.33609957,0.90198153,1.0185875,0.980862,0.9945804,1.0631721,0.9877212,0.77851635,0.823101,1.08032,1.2895249,0.97057325,1.4918705,2.393852,3.2066643,3.865145,4.7362604,5.0586414,5.3673043,5.576509,5.7308407,5.9983487,6.869464,7.010077,6.3310184,5.1238036,4.081209,3.0454736,3.1517909,3.0523329,2.9220085,4.4516044,5.051782,5.754848,6.018926,5.8165803,5.6656785,5.9126086,5.1752477,4.2423997,4.0606318,5.7239814,4.996909,5.336438,4.1429415,1.5810398,0.5624523,0.51100856,0.7990939,1.728512,3.2889743,5.164959,7.099246,9.469091,10.710602,9.602845,5.2506986,1.8725548,0.4698535,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.08573969,0.34295875,0.15776102,0.274367,0.432128,0.4424168,0.17147937,0.52815646,0.6962063,0.64819205,0.40126175,0.0,0.0,0.0,0.048014224,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.07888051,0.13375391,0.17490897,0.2709374,0.41840968,0.48014224,0.20577525,0.19891608,0.08573969,0.048014224,0.16462019,0.4389872,0.40126175,0.42183927,0.4972902,0.7476501,1.4267083,2.0406046,2.4007113,2.9220085,3.7965534,5.003768,5.576509,5.778855,5.0757895,4.0434837,4.3624353,4.897451,4.722542,4.232111,4.314421,6.3207297,10.88551,12.034423,9.414218,4.773986,1.9857311,1.8965619,1.9582944,2.0680413,2.428148,3.5393343,3.7108135,3.1380725,2.3252604,1.605047,1.1351935,0.939707,0.8265306,0.881404,1.2346514,2.0646117,2.9391565,3.223812,3.1552205,2.8877127,2.4967396,2.6304936,2.7539587,2.9803114,3.333559,3.7553983,5.305572,7.363324,8.769455,8.838047,7.3427467,5.5833683,4.513337,3.542764,2.633923,2.287535,1.5673214,1.1249046,1.2209331,1.5844694,1.4198492,1.0357354,0.8093826,0.7305021,0.77851635,0.9259886,0.9568549,0.8093826,0.72021335,0.85739684,1.3169615,2.054323,3.2855449,5.2987127,7.98065,10.813489,11.670886,12.099585,11.036412,8.241299,4.32471,1.8485477,0.6962063,0.30523327,0.2503599,0.26064864,0.25378948,0.1371835,0.07545093,0.082310095,0.024007112,0.01371835,0.0034295875,0.0034295875,0.017147938,0.037725464,0.048014224,0.061732575,0.09259886,0.13032432,0.15776102,0.14404267,0.23664154,0.274367,0.22292319,0.14404267,0.037725464,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.0274367,0.0274367,0.024007112,0.017147938,0.01371835,0.020577524,0.037725464,0.12003556,0.29494452,0.432128,0.4698535,0.42526886,0.45270553,0.58645946,0.7579388,0.88826317,0.89512235,1.1694894,1.611906,1.8828435,1.8416885,1.5501735,1.7559488,1.99602,1.7079345,1.0048691,0.6927767,1.1214751,1.4335675,1.3821237,1.1008976,1.1043272,1.4164196,1.5570327,1.5261664,1.3752645,1.1694894,1.0700313,1.1934965,1.3238207,1.3203912,1.1249046,1.6804979,2.194936,2.218943,1.8245405,1.6084765,1.0597426,0.58988905,0.29151493,0.18519773,0.18519773,0.24350071,0.28808534,0.37382504,0.47328308,0.51100856,0.9362774,0.6241849,0.22978236,0.0548734,0.044584636,0.18862732,0.18519773,0.13032432,0.08573969,0.072021335,0.06516216,0.058302987,0.08916927,0.37039545,1.2826657,2.9391565,2.5070283,1.9857311,1.9411465,1.5158776,0.980862,0.9945804,1.2037852,1.3272504,1.1214751,1.0631721,1.3992717,2.3424082,3.642222,4.5922174,3.6970954,4.214963,3.8857226,2.5721905,2.2978237,2.311542,2.668219,3.0077481,3.316411,3.9543142,4.166949,3.625074,3.8308492,5.4016004,8.093826,6.8591747,4.057202,3.0454736,4.57507,6.776865,6.2658563,5.967482,6.660259,8.217292,9.609704,9.249598,8.577398,7.689135,6.351596,3.9783216,1.5398848,0.75450927,0.6790583,0.78194594,0.9259886,1.2277923,2.1880767,4.722542,9.297611,15.940722,20.670124,22.12427,20.982216,18.190533,14.942713,13.478279,13.450842,13.666906,13.032433,10.556271,7.034084,4.184097,2.2909644,1.2655178,0.6207553,0.33609957,0.13032432,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.01371835,0.0034295875,0.0034295875,0.010288762,0.024007112,0.048014224,0.048014224,0.0548734,0.058302987,0.0,0.048014224,0.1920569,0.2194936,0.106317215,0.030866288,0.041155048,0.041155048,0.037725464,0.0274367,0.010288762,0.11317638,0.29151493,0.50757897,0.7579388,1.0940384,1.4987297,1.5193073,1.4232788,1.3306799,1.2277923,1.1694894,0.94999576,0.72707254,0.61389613,0.6927767,0.82996017,0.85396725,0.7510797,0.5727411,0.4115505,0.17490897,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.044584636,0.082310095,0.12003556,0.116605975,0.20920484,0.42869842,0.6790583,0.6001778,0.4698535,0.38754338,0.33609957,0.19548649,0.058302987,0.030866288,0.05144381,0.08916927,0.15776102,0.216064,0.61046654,0.9774324,1.2209331,1.5158776,1.7079345,2.3492675,2.9906003,3.3781435,3.4398763,4.190956,4.770556,4.90431,4.9180284,5.7479887,5.994919,6.3481665,6.509357,6.5813785,7.1061053,7.191845,6.824879,6.701414,7.0443726,7.6171136,6.6293926,5.4941993,4.6436615,4.125794,3.625074,2.1126258,2.884283,2.9665933,1.920569,1.845118,2.1400626,2.0817597,1.8999915,1.821111,2.0406046,3.1140654,4.5510626,5.470192,5.15467,3.0557625,1.2792361,0.66876954,0.4081209,0.14061308,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.14061308,0.116605975,0.23664154,0.37382504,0.432128,0.37725464,0.40126175,0.5007198,0.53844523,0.39783216,0.0,0.072021335,0.037725464,0.06516216,0.13032432,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.034295876,0.06859175,0.07545093,0.2777966,0.4698535,0.490431,0.216064,0.18176813,0.072021335,0.14061308,0.36353627,0.45613512,0.28122616,0.20234565,0.20577525,0.33609957,0.72021335,1.2415106,1.5673214,1.8588364,2.5207467,4.173808,4.3281393,4.6265135,4.8597255,5.24041,6.392751,7.514226,8.296172,8.512236,8.546532,9.414218,11.598865,10.244178,6.6465406,2.6579304,0.6962063,0.4629943,0.45613512,0.5453044,0.7888051,1.4541451,2.2326615,2.3321195,2.0406046,1.6221949,1.3341095,1.1008976,1.0460242,1.1832076,1.4678634,1.7799559,1.9994495,2.3904223,2.9288676,3.3472774,3.1277838,3.0969174,3.2889743,3.5187566,3.666229,3.6799474,4.314421,5.5079174,7.0272245,7.8091707,5.970912,5.3432975,5.223262,4.846007,4.108646,3.5770597,3.069481,2.651071,2.3149714,2.0474637,1.8416885,1.8142518,1.3306799,0.82996017,0.5590228,0.59331864,0.5727411,0.8745448,1.138623,1.3238207,1.704505,1.9342873,2.668219,4.273266,6.7322803,9.606275,11.046701,11.369082,10.024684,7.1987042,3.7965534,1.9342873,0.7990939,0.274367,0.16119061,0.17147937,0.26750782,0.24350071,0.17833854,0.116605975,0.041155048,0.034295876,0.030866288,0.034295876,0.05144381,0.082310095,0.13032432,0.18176813,0.23664154,0.3018037,0.39097297,0.2777966,0.32581082,0.32924038,0.22978236,0.10288762,0.024007112,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.041155048,0.041155048,0.024007112,0.01371835,0.006859175,0.006859175,0.01371835,0.061732575,0.18519773,0.30523327,0.3806842,0.41840968,0.44584638,0.5144381,0.7510797,1.0666018,1.1592005,1.4610043,1.6427724,1.646202,1.5090185,1.3684053,1.4953002,1.7182233,1.704505,1.5021594,1.5227368,1.9548649,2.0508933,1.7388009,1.2312219,0.99801,1.0906088,1.08032,1.0460242,1.0014396,0.90884066,0.7476501,0.7339317,0.7990939,0.8711152,0.89855194,1.255229,1.6907866,1.7971039,1.529596,1.2106444,0.7510797,0.44927597,0.26750782,0.17833854,0.15776102,0.22292319,0.274367,0.29151493,0.28122616,0.26407823,0.490431,0.33609957,0.12346515,0.017147938,0.01371835,0.09945804,0.1371835,0.14061308,0.12346515,0.09602845,0.09259886,0.072021335,0.061732575,0.21263443,0.7922347,2.4830213,2.7162333,2.5207467,2.2978237,1.8279701,1.2346514,1.0014396,0.96371406,0.9602845,0.8505377,0.8162418,1.097468,1.8862731,3.018037,3.9646032,3.6936657,4.3452873,4.266407,3.2135234,2.3561265,3.1072063,3.1826572,3.1380725,3.2683969,3.6044965,4.8494368,4.479041,4.5099077,5.994919,9.006097,6.958633,4.5339146,4.314421,5.7239814,5.0106273,5.5422134,6.293293,8.124693,10.100135,9.506817,8.755736,8.40249,8.158989,7.531374,5.8337283,2.9700227,1.3855534,0.7888051,0.7373613,0.65162164,0.7373613,1.0357354,2.1469216,4.8082814,9.887501,16.654078,22.391777,25.94826,26.925692,25.711617,24.363789,23.664154,22.566685,20.484926,17.29198,12.792361,8.889491,5.878313,3.6593697,1.7113642,0.90541106,0.4046913,0.12689474,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.010288762,0.006859175,0.020577524,0.1097468,0.15090185,0.16804978,0.31209245,0.32581082,0.29151493,0.32581082,0.432128,0.5041494,0.5555932,0.75450927,1.0528834,1.430138,1.8965619,2.253239,1.6667795,1.1694894,1.155771,1.3684053,1.2723769,0.94656616,0.5624523,0.2777966,0.26407823,0.44584638,0.48700142,0.3841138,0.18519773,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.034295876,0.09259886,0.20920484,0.21263443,0.16119061,0.18862732,0.274367,0.2469303,0.12346515,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.044584636,0.07545093,0.082310095,0.22978236,0.6824879,1.1077567,1.3272504,1.3409687,1.8828435,2.3801336,2.726522,3.292404,4.945465,5.9400454,6.759717,7.548522,8.261876,8.669997,9.088407,8.700864,8.457363,8.680285,9.071259,7.720001,6.667118,5.857735,5.07236,3.9371665,3.2683969,3.8857226,4.201245,3.8685746,3.799983,4.033195,3.5461934,2.5001693,1.2689474,0.4355576,0.45270553,0.5727411,0.6859175,0.7133542,0.59674823,0.4938606,0.53844523,0.45613512,0.22978236,0.1097468,0.09945804,0.08573969,0.07545093,0.061732575,0.037725464,0.006859175,0.048014224,0.116605975,0.17147937,0.17147937,0.034295876,0.0,0.0,0.0,0.0,0.044584636,0.14404267,0.23664154,0.29151493,0.29151493,0.21263443,0.26407823,0.39097297,0.45613512,0.274367,0.30866286,0.12689474,0.041155048,0.07888051,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14747226,0.26064864,0.25378948,0.1371835,0.09259886,0.034295876,0.116605975,0.29494452,0.30523327,0.16462019,0.09602845,0.0548734,0.05144381,0.14747226,0.38754338,0.8025235,1.097468,1.4747226,2.620205,2.6785078,3.1380725,4.180667,5.6793966,7.222711,8.416207,9.249598,9.595985,9.417647,8.748878,8.697433,6.1972647,3.1792276,0.9602845,0.24350071,0.12003556,0.106317215,0.216064,0.42869842,0.70649505,1.1934965,1.4061309,1.430138,1.3615463,1.3101025,1.2003556,1.138623,1.2312219,1.4095604,1.4267083,1.2449403,1.5158776,2.2120838,3.0386145,3.415869,3.8377085,4.197815,4.3178506,4.2595477,4.3041325,4.8734436,5.5490727,6.6705475,7.2775846,5.1238036,4.671098,4.8117113,4.887162,4.65395,4.273266,4.057202,3.9680326,3.673088,3.1140654,2.5138876,2.8945718,2.2841053,1.313532,0.4972902,0.23321195,0.29151493,1.0288762,1.7250825,2.07833,2.1812177,2.1194851,2.527606,3.4776018,5.099797,7.5862474,8.752307,8.333898,6.8591747,4.8254294,2.6853669,1.6770682,0.939707,0.5144381,0.34638834,0.26750782,0.31895164,0.31895164,0.2709374,0.19548649,0.13032432,0.1371835,0.14747226,0.16804978,0.20577525,0.26407823,0.34981793,0.41840968,0.45956472,0.48357183,0.5418748,0.4081209,0.36353627,0.34638834,0.2709374,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.037725464,0.044584636,0.0274367,0.006859175,0.0,0.0,0.0,0.030866288,0.07545093,0.14061308,0.22292319,0.3018037,0.32581082,0.34638834,0.5453044,0.8745448,1.08032,1.3821237,1.3649758,1.1660597,0.9431366,0.86082643,0.9945804,1.1934965,1.3375391,1.4335675,1.6221949,1.9342873,1.9891608,1.7456601,1.313532,0.94999576,0.89169276,0.7956643,0.69963586,0.6173257,0.53158605,0.39783216,0.42869842,0.6001778,0.84367853,1.0631721,1.2415106,1.3341095,1.2895249,1.1008976,0.8093826,0.6859175,0.64476246,0.6241849,0.6001778,0.58645946,0.5658819,0.6173257,0.59674823,0.50757897,0.5007198,0.45613512,0.31552204,0.16804978,0.061732575,0.017147938,0.0274367,0.07545093,0.1097468,0.11317638,0.09602845,0.11317638,0.09259886,0.07888051,0.19891608,0.64819205,1.6290541,1.99602,2.0234566,1.9102802,1.7593783,1.2758065,1.0768905,0.9328478,0.75450927,0.607037,0.6310441,0.8162418,1.5673214,2.6990852,3.4467354,3.5050385,3.9680326,3.9680326,3.3850029,2.843128,4.166949,3.789694,3.2135234,3.0866287,3.2135234,4.389872,4.40702,4.9008803,6.3653145,8.1384115,5.8988905,4.4241676,4.6916757,5.785714,4.931747,4.7499785,5.453044,7.5245147,9.791472,9.407358,8.519095,8.529384,8.80718,8.752307,7.7885933,5.2987127,3.2066643,1.961724,1.3615463,0.5212973,0.5007198,0.59331864,0.980862,2.1434922,4.870014,10.6317215,17.88873,24.641586,29.76539,32.99949,36.24388,39.73863,42.708652,44.92074,46.70755,46.55665,41.446564,32.18668,20.848463,10.7757635,5.5730796,2.5207467,0.9259886,0.23321195,0.030866288,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.0274367,0.044584636,0.09602845,0.07888051,0.12003556,0.1920569,0.26064864,0.25378948,0.15090185,0.12003556,0.22292319,0.5041494,0.9842916,1.2380811,1.097468,0.96714365,0.9911508,1.0528834,0.9294182,0.94999576,1.1111864,1.3684053,1.6221949,1.5947582,1.0631721,0.65848076,0.607037,0.72021335,0.42869842,0.1920569,0.0548734,0.010288762,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.1097468,0.25721905,0.18862732,0.09602845,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.08916927,0.39097297,1.0460242,1.4335675,1.6153357,1.7113642,1.9068506,2.6853669,3.9097297,5.23698,6.5367937,7.891481,9.160428,9.887501,9.993818,9.493098,8.467651,7.3873315,6.680836,5.9914894,5.284994,4.8425775,5.288424,5.271276,5.120374,4.945465,4.6402316,4.465323,3.6936657,2.4967396,1.2380811,0.45613512,0.42869842,0.274367,0.106317215,0.0,0.0,0.0,0.08916927,0.15776102,0.18519773,0.24350071,0.2503599,0.25378948,0.26064864,0.26407823,0.23664154,0.17833854,0.22292319,0.32238123,0.4081209,0.3841138,0.07545093,0.0,0.01371835,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17147937,0.37382504,0.5453044,0.6756287,0.6173257,0.30866286,0.14747226,0.15776102,0.0,0.0,0.034295876,0.061732575,0.061732575,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.18862732,0.15433143,0.14747226,0.08916927,0.0,0.0,0.030866288,0.52815646,0.9362774,1.0768905,1.1283343,1.371835,1.7765263,2.651071,3.9097297,5.0757895,5.7136927,6.012067,6.012067,5.5147767,4.057202,3.8102717,2.6373527,1.3409687,0.41840968,0.082310095,0.0274367,0.0274367,0.12346515,0.29494452,0.47328308,0.67219913,0.7442205,0.823101,0.9328478,0.99801,1.0700313,0.9534253,0.8779744,0.91569984,0.9602845,1.0014396,1.1111864,1.4061309,1.9342873,2.6819375,3.6593697,4.173808,4.197815,4.081209,4.5442033,5.8200097,6.2967224,6.451054,6.125243,4.530485,3.9371665,3.9714622,4.3041325,4.6436615,4.7328305,4.6265135,4.846007,4.8905916,4.431027,3.3026927,3.8034124,3.2512488,2.0406046,0.77165717,0.22635277,0.5555932,1.4164196,2.253239,2.627064,2.218943,1.9685832,2.3458378,2.9322972,3.841138,5.7136927,5.7925735,4.6882463,3.5118976,2.6819375,1.9480057,1.4918705,1.2929544,1.1660597,0.99801,0.7339317,0.5521636,0.4115505,0.33952916,0.31552204,0.2709374,0.3018037,0.34295875,0.39097297,0.44584638,0.51100856,0.58645946,0.6207553,0.61389613,0.5658819,0.48357183,0.4046913,0.32581082,0.33952916,0.34295875,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.041155048,0.034295876,0.01371835,0.0,0.0,0.0034295875,0.0,0.0,0.01371835,0.044584636,0.072021335,0.072021335,0.09602845,0.18862732,0.35324752,0.5624523,0.7407909,0.6927767,0.548734,0.40126175,0.31209245,0.4355576,0.64476246,0.78537554,0.83681935,0.91912943,1.1317638,1.3341095,1.3581166,1.1626302,0.8196714,0.7579388,0.7407909,0.67219913,0.53501564,0.4046913,0.36696586,0.6173257,1.0185875,1.3992717,1.5638919,1.6427724,1.4575747,1.1866373,0.94999576,0.8025235,1.039165,1.1283343,1.1592005,1.1797781,1.2003556,1.0460242,1.0357354,0.9911508,0.922559,1.0528834,0.94656616,0.66191036,0.37725464,0.18176813,0.058302987,0.034295876,0.05144381,0.061732575,0.0548734,0.0548734,0.09259886,0.08573969,0.09259886,0.18862732,0.45956472,0.8505377,0.88826317,0.9945804,1.2792361,1.5501735,1.155771,1.0940384,1.0151579,0.7990939,0.5590228,0.53501564,0.5796003,1.2689474,2.3972816,2.9734523,3.2478194,3.7313912,3.8342788,3.6079261,3.74168,5.0174866,4.540774,3.7039545,3.2032347,3.059192,3.1380725,3.457024,4.8322887,6.557371,6.39961,4.9488945,4.1772375,4.040054,4.7259717,6.6636887,5.051782,4.4241676,5.099797,6.81802,8.7317295,8.210432,8.604835,9.366203,9.918367,9.650859,8.117833,6.108095,4.40702,3.0489032,1.3341095,0.6756287,0.47671264,0.548734,0.91227025,1.7833855,4.619654,10.062409,16.739817,23.825344,31.003471,40.201626,50.747604,61.715427,72.86159,84.614784,93.161316,87.25556,68.893555,44.351425,24.17859,13.018714,6.3653145,2.7128036,0.922559,0.23664154,0.09259886,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.08916927,0.14404267,0.2194936,0.48700142,0.40126175,0.5178677,0.84367853,1.1934965,1.2037852,0.6927767,0.4629943,0.59331864,1.0666018,1.8005334,2.9220085,2.627064,1.7113642,0.7956643,0.31895164,0.19891608,0.13032432,0.082310095,0.048014224,0.061732575,0.061732575,0.034295876,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.29837412,0.939707,1.5158776,0.9294182,1.0151579,1.7525192,2.551613,3.216953,3.9371665,5.0003386,6.509357,7.98065,8.944365,8.958082,8.772884,8.086967,7.1095347,6.101236,5.3570156,5.7822843,5.7891436,4.787704,3.210094,2.503599,2.2223728,1.7662375,1.3101025,1.0288762,1.1146159,1.1763484,0.7888051,0.31209245,0.0,0.0,0.0,0.0,0.0,0.024007112,0.12346515,0.24350071,0.40126175,0.5624523,0.70306545,0.823101,0.823101,0.64133286,0.45270553,0.32238123,0.21263443,0.041155048,0.0,0.06859175,0.13375391,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12003556,0.12003556,0.12346515,0.6241849,0.72364295,0.64819205,0.7442205,0.7922347,0.0,0.0,0.17490897,0.30866286,0.31209245,0.21263443,0.041155048,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.274367,0.10288762,0.024007112,0.0,0.0,0.0,0.15776102,0.47328308,0.764798,0.922559,0.8848336,0.6893471,0.59674823,0.7099246,1.097468,1.7559488,1.8656956,2.037175,2.1229146,2.2120838,2.6407824,2.0920484,1.3855534,0.78194594,0.38754338,0.16804978,0.034295876,0.0,0.01371835,0.034295876,0.044584636,0.06859175,0.11317638,0.18176813,0.2777966,0.4115505,0.48357183,0.548734,0.5693115,0.6207553,0.90198153,1.155771,1.3032433,1.3581166,1.3889829,1.5090185,1.0700313,1.2449403,1.6187652,2.0303159,2.5790498,3.690236,4.197815,4.2081037,4.0194764,4.105216,4.6916757,5.422178,6.118384,6.6122446,6.759717,6.478491,6.3893213,5.9743414,5.096367,3.998899,3.7279615,3.2581081,2.4830213,1.5433143,0.823101,1.1523414,1.903421,2.6236343,2.9391565,2.5481834,2.085189,2.0063086,2.3458378,2.942586,3.4192986,2.7951138,2.037175,1.5604624,1.471293,1.5570327,1.5330256,1.7833855,2.0508933,2.0646117,1.5398848,1.0666018,0.72707254,0.51100856,0.39440256,0.31895164,0.41840968,0.50757897,0.5727411,0.59674823,0.548734,0.52472687,0.490431,0.52815646,0.5453044,0.29151493,0.22978236,0.28808534,0.35324752,0.32924038,0.12346515,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.030866288,0.01371835,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.037725464,0.061732575,0.13375391,0.19891608,0.20577525,0.15090185,0.09259886,0.17833854,0.32581082,0.4424168,0.5041494,0.5658819,0.7613684,0.84367853,0.84367853,0.7956643,0.7476501,0.72364295,0.75450927,0.7956643,0.8093826,0.7476501,0.69963586,1.0700313,1.6324836,2.0268862,1.7696671,1.5364552,1.5090185,1.4472859,1.3272504,1.3272504,1.5364552,1.3684053,1.1763484,1.1008976,1.0528834,0.91912943,0.8128122,0.6790583,0.6001778,0.8093826,0.8711152,0.72021335,0.4938606,0.2777966,0.106317215,0.044584636,0.020577524,0.020577524,0.030866288,0.030866288,0.06859175,0.07545093,0.08916927,0.13032432,0.22978236,0.5590228,0.7956643,1.0357354,1.2312219,1.2209331,0.8162418,0.5693115,0.5144381,0.5590228,0.47328308,0.40126175,0.3806842,0.61389613,1.1523414,1.9239986,2.7642474,4.091498,5.312431,5.693115,4.3624353,4.8288593,5.15467,4.945465,4.180667,3.2032347,3.998899,4.4447455,5.3090014,5.8508763,3.799983,4.0194764,4.880303,5.0929375,4.955754,6.3481665,7.5210853,6.824879,5.470192,4.6402316,5.5079174,5.4839106,6.495639,8.258447,10.041832,10.6488695,10.6488695,9.451943,7.870903,6.2898636,4.65395,1.5536032,0.5761707,0.45613512,0.51100856,0.67219913,1.2826657,3.5599117,7.5690994,13.193623,20.128248,28.475864,38.82293,50.579556,64.75404,83.97002,98.81327,93.96041,72.7587,45.260265,28.242653,17.511473,10.39165,5.552502,2.3595562,0.8711152,0.34638834,0.10288762,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.0274367,0.010288762,0.0,0.0,0.0,0.0034295875,0.017147938,0.0274367,0.061732575,0.18176813,0.16462019,0.29151493,0.41840968,0.5761707,0.94999576,0.77851635,0.4355576,0.53501564,1.2998136,2.568761,2.901431,1.5673214,0.4629943,0.20234565,0.07545093,0.041155048,0.0274367,0.017147938,0.010288762,0.01371835,0.01371835,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.058302987,0.18862732,0.3018037,0.18519773,0.20234565,0.70306545,1.1317638,1.3512574,1.6427724,2.627064,3.765687,4.722542,5.4599032,6.23499,7.6445503,7.7131424,7.466212,7.298162,6.992929,6.7048435,6.3961806,5.579939,4.3178506,3.199805,3.1895163,3.2443898,2.819121,1.9445761,1.2003556,0.66533995,0.39097297,0.2777966,0.22978236,0.17147937,0.26750782,0.116605975,0.09259886,0.22978236,0.2194936,0.08916927,0.16804978,0.37725464,0.66533995,1.0323058,1.371835,1.5261664,1.5158776,1.1592005,0.041155048,0.106317215,0.048014224,0.01371835,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.024007112,0.082310095,0.4046913,0.6001778,0.67219913,0.89855194,1.1660597,0.9774324,0.5658819,0.8779744,1.0837497,0.78537554,0.041155048,0.006859175,0.0,0.13032432,0.33609957,0.36696586,0.072021335,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.19548649,0.3018037,0.28808534,0.1920569,0.13375391,0.0274367,0.0,0.020577524,0.06859175,0.15090185,0.17833854,0.072021335,0.020577524,0.06859175,0.14747226,0.061732575,0.09602845,0.25721905,0.4424168,0.44584638,0.33952916,0.31552204,0.39440256,0.53501564,0.65505123,0.5521636,0.5453044,0.607037,0.6927767,0.7476501,0.6962063,0.8196714,0.9362774,0.8848336,0.51100856,0.2777966,0.09602845,0.010288762,0.010288762,0.020577524,0.017147938,0.024007112,0.037725464,0.058302987,0.09602845,0.13032432,0.12346515,0.17833854,0.30866286,0.45956472,0.6790583,1.5536032,1.9857311,1.8073926,1.7902447,1.4198492,1.0837497,0.83681935,0.7442205,0.89512235,1.4198492,1.8897027,2.194936,2.369845,2.5893385,3.7039545,4.7945633,5.501058,5.6793966,5.40503,5.3501563,5.0586414,4.5030484,3.7039545,2.7539587,2.0749004,1.7593783,1.5398848,1.255229,0.83681935,1.2346514,1.8691251,2.253239,2.2360911,2.0097382,1.8416885,1.8108221,1.8862731,2.0337453,2.2463799,2.4624438,2.352697,2.0680413,1.9548649,2.5584722,2.4830213,2.627064,2.7916842,2.7402403,2.1743584,1.7765263,1.4164196,1.0494537,0.764798,0.7613684,0.7305021,0.764798,0.7990939,0.8265306,0.91569984,0.83338976,0.75450927,0.6310441,0.44584638,0.22978236,0.22635277,0.34981793,0.4355576,0.36353627,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.030866288,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.024007112,0.037725464,0.05144381,0.05144381,0.048014224,0.0548734,0.1097468,0.20234565,0.29837412,0.38754338,0.48014224,0.5761707,0.6001778,0.58645946,0.5624523,0.5521636,0.6756287,0.83681935,1.0494537,1.2860953,1.4815818,1.196926,1.1077567,1.3855534,1.7079345,1.2586586,1.2415106,1.0151579,0.7305021,0.4972902,0.40126175,0.51100856,0.5212973,0.4664239,0.39783216,0.41840968,0.39097297,0.274367,0.21263443,0.2709374,0.42869842,0.4424168,0.33266997,0.2194936,0.16119061,0.15433143,0.11317638,0.05144381,0.010288762,0.006859175,0.006859175,0.024007112,0.048014224,0.072021335,0.17147937,0.5212973,0.764798,0.8471081,0.8505377,0.8265306,0.7922347,0.65505123,0.59674823,0.65848076,0.7990939,0.88826317,0.8745448,0.69963586,0.6241849,0.78194594,1.1900668,1.7696671,3.000889,4.763697,6.3001523,6.217842,5.3741636,5.219832,5.267846,5.2026844,4.887162,5.5662203,5.2644167,4.5784993,3.9200184,3.5187566,3.9337368,4.8494368,5.3707337,5.2815647,5.055212,5.3570156,5.4187484,4.73969,3.5976372,3.0317552,4.3933015,5.295283,6.385892,7.888051,9.599416,11.321068,11.567999,10.816919,9.56512,8.327039,5.8234396,2.9220085,1.1454822,0.764798,0.805953,0.9945804,1.7971039,3.7965534,7.06838,11.190743,17.70696,24.970827,31.061773,35.962654,41.56317,49.632988,52.088573,46.834446,36.72745,29.573332,22.906214,17.758404,12.898679,8.090397,4.091498,1.9651536,0.8128122,0.2709374,0.072021335,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.041155048,0.09259886,0.14061308,0.30866286,0.91227025,0.71678376,0.33609957,0.22978236,0.5418748,1.1043272,1.1592005,0.5212973,0.061732575,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17490897,0.32238123,0.40126175,0.5453044,0.9911508,1.4027013,1.7079345,2.0508933,2.7813954,4.3521466,5.2472687,5.7377,6.0223556,6.193835,6.1972647,7.006647,7.0718093,5.953764,4.314421,3.7039545,3.2581081,2.836269,2.2909644,1.4781522,0.8676856,0.59674823,0.4389872,0.32238123,0.31552204,0.26064864,0.2194936,0.24007112,0.25721905,0.09602845,0.020577524,0.044584636,0.13032432,0.31895164,0.70649505,1.1729189,1.5193073,1.6770682,1.5501735,1.0254467,1.0528834,0.96714365,0.72021335,0.34981793,0.0,0.06516216,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.10288762,0.5144381,0.82996017,0.86082643,0.84024894,0.86082643,0.85396725,0.48014224,0.78537554,1.1420527,1.0768905,0.28465575,0.1371835,0.15090185,0.39440256,0.72707254,0.77851635,0.41840968,0.25721905,0.23664154,0.26407823,0.22978236,0.19891608,0.116605975,0.106317215,0.16119061,0.1371835,0.08573969,0.08916927,0.1920569,0.32581082,0.31209245,0.30523327,0.22292319,0.14404267,0.09602845,0.06859175,0.01371835,0.0,0.010288762,0.0548734,0.17833854,0.18519773,0.12003556,0.11317638,0.19891608,0.31209245,0.28122616,0.18519773,0.17490897,0.23664154,0.18862732,0.3018037,0.35324752,0.4081209,0.4389872,0.31895164,0.12346515,0.06859175,0.09259886,0.12346515,0.1097468,0.14061308,0.2709374,0.4938606,0.7682276,1.0357354,1.2037852,1.155771,0.9534253,0.6756287,0.41840968,0.20920484,0.061732575,0.0,0.0,0.006859175,0.06859175,0.12689474,0.12346515,0.09259886,0.14061308,0.31895164,0.8265306,1.1249046,1.1694894,1.4129901,1.4918705,1.3101025,0.9911508,0.71678376,0.72021335,0.7407909,0.8025235,0.8676856,0.9259886,1.0220171,1.5570327,2.0337453,2.3835633,2.5481834,2.4830213,2.352697,2.3149714,2.0646117,1.5570327,1.0117283,0.8779744,0.7442205,0.6824879,0.6790583,0.6276145,0.88826317,1.2346514,1.4232788,1.4027013,1.2998136,1.1934965,1.0940384,0.97400284,1.1420527,2.2566686,2.9082901,2.9700227,2.5413244,2.0131679,2.0577524,2.2120838,2.4624438,2.5207467,2.2463799,1.6221949,1.5193073,1.3512574,1.2346514,1.1934965,1.1626302,0.9774324,0.922559,0.922559,0.9259886,0.9259886,0.7682276,0.6379033,0.5144381,0.37725464,0.21263443,0.20234565,0.29494452,0.31209245,0.20234565,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.020577524,0.020577524,0.017147938,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.017147938,0.044584636,0.09259886,0.16119061,0.24007112,0.32924038,0.39440256,0.41498008,0.42526886,0.4698535,0.58645946,0.66533995,0.7613684,0.9534253,1.2792361,1.762808,1.5398848,1.1008976,0.922559,1.0494537,1.0940384,1.2826657,1.0460242,0.64133286,0.28808534,0.15776102,0.20920484,0.274367,0.29494452,0.29151493,0.34981793,0.45270553,0.48700142,0.48014224,0.44927597,0.39097297,0.45613512,0.4698535,0.45613512,0.4115505,0.32238123,0.31552204,0.26064864,0.18519773,0.12003556,0.082310095,0.09602845,0.07545093,0.0548734,0.09259886,0.26407823,0.36010668,0.4081209,0.4115505,0.41498008,0.4938606,0.53158605,0.5761707,0.64476246,0.7305021,0.7888051,0.8848336,0.85739684,0.75450927,0.6824879,0.83338976,1.2860953,1.9548649,3.4604537,5.2301207,5.4839106,5.051782,5.5387836,5.9469047,5.717122,4.7499785,6.262427,6.3035817,5.4153185,4.201245,3.3198407,3.3232703,3.6010668,3.940596,4.187526,4.2183924,4.3109913,4.5030484,4.3281393,3.5770597,2.2841053,3.7485392,5.267846,6.090947,6.5367937,7.98408,10.820349,12.55229,13.039291,12.47341,11.38966,9.544542,7.010077,4.588788,2.5996273,0.8745448,0.823101,1.0117283,1.8039631,3.316411,5.422178,10.532263,16.770683,22.299177,26.236343,28.654203,30.880005,31.740831,31.66881,30.897154,29.43272,25.073713,20.954779,17.322845,13.786942,9.290752,5.360445,2.7470996,1.2072148,0.45270553,0.15090185,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.034295876,0.048014224,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.106317215,0.33952916,0.64476246,0.42869842,0.17147937,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.12003556,0.17833854,0.1920569,0.19891608,0.28808534,0.61389613,1.5741806,2.3904223,3.018037,3.4433057,3.6765177,4.1600895,5.4599032,6.1321025,5.7136927,4.698535,4.057202,3.426158,2.8980014,2.486451,2.136633,1.6667795,1.1832076,0.7922347,0.5796003,0.6241849,0.490431,0.4664239,0.44584638,0.34295875,0.13375391,0.09602845,0.18176813,0.22292319,0.274367,0.59674823,0.8676856,1.0528834,1.2209331,1.3615463,1.3924125,1.3924125,1.3615463,1.1180456,0.65162164,0.1097468,0.116605975,0.048014224,0.0,0.0034295875,0.024007112,0.07888051,0.23321195,0.4115505,0.6001778,0.8711152,0.9259886,0.7579388,0.5555932,0.4664239,0.58645946,0.34295875,0.4629943,0.85739684,1.1523414,0.6859175,0.5144381,0.5590228,0.82996017,1.2517995,1.6393428,1.6942163,1.1454822,0.7373613,0.72707254,0.881404,1.0151579,1.0288762,1.097468,1.1660597,0.96714365,0.6241849,0.48014224,0.53501564,0.64476246,0.5418748,0.31209245,0.16462019,0.08916927,0.0548734,0.0,0.0,0.0,0.0,0.024007112,0.12689474,0.106317215,0.08573969,0.10288762,0.17833854,0.31209245,0.28122616,0.18519773,0.17833854,0.274367,0.36010668,0.4046913,0.4355576,0.47671264,0.4664239,0.26407823,0.061732575,0.017147938,0.010288762,0.0,0.0,0.0,0.030866288,0.20920484,0.5144381,0.7956643,1.0666018,1.1489118,1.0357354,0.823101,0.6927767,0.39440256,0.1920569,0.061732575,0.0,0.0,0.05144381,0.12003556,0.09259886,0.0,0.0,0.09602845,0.17833854,0.26750782,0.4355576,0.8265306,1.1008976,1.1832076,1.0906088,0.9602845,1.039165,0.83338976,0.6379033,0.5007198,0.42869842,0.38754338,0.3841138,0.34638834,0.36696586,0.44927597,0.4938606,0.35324752,0.4389872,0.41498008,0.216064,0.037725464,0.216064,0.1920569,0.16804978,0.22978236,0.33609957,0.4424168,0.5453044,0.65848076,0.7373613,0.6893471,0.5761707,0.4355576,0.29494452,0.48357183,1.646202,2.2498093,2.4418662,2.2326615,1.8142518,1.5193073,1.4644338,1.6667795,1.6770682,1.4129901,1.1249046,1.255229,1.2312219,1.2586586,1.3684053,1.4267083,1.255229,1.0563129,0.88826317,0.8128122,0.91912943,0.6344737,0.41498008,0.29151493,0.23664154,0.15090185,0.1371835,0.17147937,0.15090185,0.06859175,0.030866288,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.01371835,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.017147938,0.0274367,0.0548734,0.09602845,0.15776102,0.20577525,0.23664154,0.28465575,0.37382504,0.53158605,0.5555932,0.58988905,0.7613684,1.1763484,1.9342873,1.8862731,1.3101025,0.85739684,0.8128122,1.1214751,1.2792361,1.0734608,0.75450927,0.4664239,0.274367,0.2469303,0.30523327,0.36010668,0.3806842,0.4046913,0.58302987,0.8025235,0.864256,0.71678376,0.4629943,0.5007198,0.5590228,0.5761707,0.52815646,0.42183927,0.4081209,0.37382504,0.29494452,0.1920569,0.12346515,0.116605975,0.082310095,0.048014224,0.030866288,0.0274367,0.041155048,0.07888051,0.09945804,0.12689474,0.23321195,0.35324752,0.41840968,0.4424168,0.44584638,0.45613512,0.5796003,0.70649505,0.7682276,0.8162418,1.0220171,1.1351935,1.5227368,2.5893385,3.8514268,3.940596,3.9851806,4.955754,5.7925735,5.7925735,4.5819287,5.7891436,6.012067,5.288424,4.064061,3.1723683,2.7333813,2.4761622,2.6853669,3.2821152,3.8514268,3.6799474,3.6765177,3.7279615,3.4844608,2.3732746,2.9734523,4.1635194,4.852866,5.113515,6.1904054,8.796892,11.358793,13.296511,14.239647,14.020154,12.6757555,10.909517,8.752307,6.2864337,3.6353626,1.5638919,0.91569984,1.039165,1.5810398,2.4795918,6.029215,11.183885,16.71238,21.489796,24.504402,24.367218,22.786179,22.820475,24.53184,24.981115,23.341772,21.102251,19.171394,17.20624,13.649758,9.012956,5.346727,2.8054025,1.3066728,0.5178677,0.19548649,0.06516216,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.07888051,0.116605975,0.1097468,0.058302987,0.0034295875,0.0,0.0,0.006859175,0.034295876,0.07545093,0.09945804,0.041155048,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18176813,0.39440256,0.17147937,0.06516216,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.106317215,0.14747226,0.1097468,0.33609957,0.39440256,0.61046654,0.9259886,0.90541106,1.5021594,2.1880767,2.8259802,3.3438478,3.7211025,3.8171308,3.6216443,3.0797696,2.5173173,2.644212,2.5138876,1.8725548,1.3341095,1.1489118,1.1832076,1.0768905,0.94999576,0.83338976,0.7133542,0.5453044,0.34295875,0.51100856,0.65505123,0.7373613,1.0940384,0.8745448,0.6001778,0.5727411,0.7613684,0.805953,0.86082643,0.9431366,0.90198153,0.66191036,0.2194936,0.13032432,0.07545093,0.06859175,0.12689474,0.274367,0.61389613,1.1077567,1.4987297,1.605047,1.3272504,0.881404,0.4938606,0.29837412,0.34981793,0.6001778,0.45956472,0.35324752,0.65162164,1.1420527,1.0528834,0.922559,1.0563129,1.4747226,2.2086544,3.3232703,4.091498,3.1140654,2.095478,1.8965619,2.5310357,2.9734523,3.069481,3.0386145,2.8739944,2.335549,1.6221949,1.1797781,0.922559,0.7579388,0.59674823,0.39440256,0.32581082,0.25721905,0.14061308,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.010288762,0.05144381,0.044584636,0.05144381,0.26407823,0.20577525,0.1920569,0.29837412,0.51100856,0.7339317,0.47671264,0.41840968,0.42869842,0.39097297,0.22635277,0.116605975,0.08573969,0.048014224,0.0,0.0,0.0,0.058302987,0.22978236,0.34295875,0.0034295875,0.0,0.082310095,0.17490897,0.3018037,0.5727411,0.37725464,0.25721905,0.12346515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06859175,0.34638834,0.45613512,0.607037,0.7613684,0.91912943,1.1420527,1.0082988,0.8745448,0.78537554,0.7339317,0.65848076,0.5555932,0.44927597,0.33952916,0.22978236,0.12003556,0.08573969,0.048014224,0.024007112,0.01371835,0.0,0.010288762,0.0034295875,0.01371835,0.048014224,0.08573969,0.106317215,0.12003556,0.22978236,0.36696586,0.31552204,0.19548649,0.09602845,0.061732575,0.13375391,0.34638834,0.58988905,0.89512235,1.1660597,1.3101025,1.2380811,0.7133542,0.69963586,0.72364295,0.6962063,0.9259886,1.138623,1.1934965,1.196926,1.2586586,1.4781522,1.4164196,1.1146159,0.77508676,0.6207553,0.90198153,0.5212973,0.23321195,0.08916927,0.061732575,0.05144381,0.05144381,0.05144381,0.041155048,0.0274367,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.041155048,0.017147938,0.0034295875,0.0,0.0034295875,0.024007112,0.044584636,0.07888051,0.14404267,0.23321195,0.32924038,0.3806842,0.44927597,0.6824879,1.1900668,2.0474637,2.2498093,1.7662375,1.2586586,1.0563129,1.1420527,1.08032,0.91227025,0.8162418,0.7682276,0.52472687,0.37725464,0.39440256,0.45270553,0.47328308,0.42183927,0.548734,0.8265306,0.9294182,0.764798,0.4698535,0.39440256,0.4046913,0.41840968,0.4046913,0.4046913,0.34638834,0.31552204,0.26064864,0.17833854,0.11317638,0.07545093,0.06516216,0.05144381,0.030866288,0.010288762,0.010288762,0.0274367,0.020577524,0.006859175,0.041155048,0.1920569,0.26750782,0.26407823,0.20577525,0.15433143,0.21263443,0.37382504,0.61389613,0.94999576,1.4164196,1.1900668,1.7388009,2.6373527,3.391862,3.426158,2.9082901,3.5118976,4.5510626,5.1821065,4.420738,4.434457,4.5990767,4.2869844,3.590778,3.3369887,2.8088322,2.3835633,2.4590142,3.117495,4.125794,3.6079261,3.2786856,3.2375305,3.2478194,2.7299516,2.1640697,2.1263442,2.6545007,3.6387923,4.822,6.3207297,8.669997,11.266195,13.526293,14.911846,14.534592,13.395968,12.085866,10.738038,9.047252,4.6745276,2.609916,1.862266,1.7765263,2.0406046,3.782835,7.2604365,11.646879,16.098484,19.764713,20.502073,19.137098,18.28656,18.674105,19.13024,20.018501,19.709839,18.890167,17.724108,15.827546,11.9040985,8.049242,4.856296,2.5824795,1.1489118,0.53844523,0.22292319,0.07545093,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041155048,0.16462019,0.39783216,0.5796003,0.5418748,0.29837412,0.01371835,0.0,0.0,0.0,0.01371835,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.061732575,0.0274367,0.07545093,0.12689474,0.2194936,0.41498008,0.75450927,1.2655178,1.8039631,1.9754424,1.9925903,1.9342873,1.7388009,2.411,2.311542,2.0989075,2.0268862,1.9514352,1.7593783,1.6907866,1.6667795,1.5947582,1.3889829,0.764798,0.7579388,1.0254467,1.4747226,2.2429502,1.3889829,0.69963586,0.31552204,0.24350071,0.36696586,0.40126175,0.53158605,0.5178677,0.30523327,0.0,0.13375391,0.23321195,0.34638834,0.59331864,1.1283343,2.287535,3.192946,3.3884325,2.7916842,1.6942163,1.1694894,0.75450927,0.59674823,0.6756287,0.8093826,0.83338976,0.78537554,0.9911508,1.3341095,1.2346514,0.8196714,1.1934965,2.352697,4.1292233,6.1801167,7.3393173,6.6876955,5.446185,4.8494368,6.118384,6.728851,6.2212715,5.164959,4.0674906,3.3712845,2.7368107,1.9925903,1.1866373,0.58645946,0.67219913,0.9259886,0.70649505,0.39097297,0.17490897,0.07545093,0.01371835,0.0,0.0,0.0,0.0,0.048014224,0.25378948,0.22978236,0.12003556,0.59674823,0.8745448,0.96371406,0.9568549,0.8676856,0.61046654,0.35324752,0.29151493,0.20920484,0.10288762,0.15090185,0.28808534,0.26407823,0.1371835,0.0,0.0,0.0,0.0,0.09602845,0.19891608,0.01371835,0.0034295875,0.010288762,0.010288762,0.01371835,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.15090185,0.15090185,0.16119061,0.26407823,0.45613512,0.64133286,0.7133542,0.7682276,0.8128122,0.82996017,0.7922347,0.67219913,0.5590228,0.44927597,0.33952916,0.22978236,0.15433143,0.1097468,0.06859175,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.15090185,0.22978236,0.16804978,0.058302987,0.01371835,0.01371835,0.0274367,0.01371835,0.01371835,0.024007112,0.1097468,0.2503599,0.33609957,0.14061308,0.09945804,0.12003556,0.15433143,0.22978236,0.5212973,0.8162418,1.0117283,1.1214751,1.2826657,1.0734608,0.91227025,0.7956643,0.6962063,0.548734,0.30523327,0.116605975,0.024007112,0.01371835,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.034295876,0.08573969,0.18176813,0.34295875,0.5555932,0.89169276,1.3512574,1.8759843,2.5001693,2.253239,1.6736387,1.1420527,0.8848336,0.77508676,0.7099246,0.77165717,0.8779744,0.7922347,0.48700142,0.39440256,0.4664239,0.5796003,0.5178677,0.42183927,0.42526886,0.42869842,0.3841138,0.274367,0.18862732,0.20577525,0.26407823,0.33266997,0.3806842,0.28465575,0.20577525,0.17490897,0.17490897,0.1371835,0.09945804,0.082310095,0.06859175,0.058302987,0.044584636,0.010288762,0.0,0.0,0.01371835,0.07545093,0.30866286,0.51100856,0.5555932,0.4115505,0.16804978,0.15433143,0.26407823,0.42869842,0.6824879,1.1592005,1.4027013,2.095478,3.3952916,4.9420357,5.844017,3.1449318,2.452155,2.8808534,3.3438478,2.5653315,3.07634,4.057202,5.1238036,5.5730796,4.3624353,4.3041325,3.7759757,3.1037767,3.1620796,5.3707337,5.079219,4.3624353,3.9611735,3.8171308,3.0969174,2.1194851,1.704505,1.99602,3.0283258,4.698535,5.895461,6.917478,7.534804,8.440215,11.262765,13.824667,13.972139,13.512574,13.516005,14.29795,12.257345,8.570539,5.5387836,4.091498,3.799983,3.9097297,6.142391,9.373062,12.902108,16.479168,18.324286,18.766703,18.509483,18.61923,20.522652,20.426622,18.653526,17.051908,16.314548,15.9613,13.495427,10.295622,6.9517736,4.016047,2.0131679,1.0254467,0.47671264,0.19548649,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.072021335,0.34638834,0.40126175,0.34295875,0.29494452,0.40126175,0.823101,1.0220171,1.0768905,1.1111864,1.3238207,1.6633499,1.4747226,0.94999576,0.34295875,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.006859175,0.01371835,0.2194936,0.23664154,0.17833854,0.15090185,0.25378948,0.44927597,0.65162164,0.96371406,1.3203912,1.5090185,1.8485477,2.5824795,3.1586502,3.2889743,2.942586,2.6579304,2.7368107,2.884283,2.9322972,2.8534167,2.1126258,2.3767042,2.9665933,3.6113555,4.4413157,3.2135234,1.9548649,1.0014396,0.4629943,0.23321195,0.24007112,0.36696586,0.3566771,0.16804978,0.0,0.14404267,0.4424168,0.70306545,1.0460242,1.8862731,2.8877127,3.542764,3.566771,2.976882,2.085189,1.8245405,1.7388009,1.5776103,1.2517995,0.8093826,0.980862,1.2826657,1.8759843,2.5824795,2.8945718,3.2032347,4.187526,5.1855364,6.0497923,7.143831,7.7851634,7.3255987,6.6568294,6.5642304,7.706283,7.6616983,6.5230756,5.144381,4.040054,3.3850029,2.4761622,2.0646117,1.6770682,1.2620882,1.2209331,0.99801,1.1934965,1.5021594,1.6942163,1.6256244,1.605047,1.3924125,1.0220171,0.5727411,0.18176813,0.048014224,0.2777966,0.3566771,0.2469303,0.40126175,0.4938606,0.44927597,0.36353627,0.31209245,0.32924038,0.26750782,0.31895164,0.24350071,0.058302987,0.030866288,0.1371835,0.16462019,0.09945804,0.0,0.0,0.0,0.0,0.020577524,0.041155048,0.0034295875,0.0,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.030866288,0.030866288,0.05144381,0.1097468,0.22635277,0.2503599,0.35324752,0.48357183,0.6001778,0.67219913,0.66533995,0.6344737,0.58302987,0.5212973,0.45956472,0.4081209,0.28465575,0.15433143,0.0548734,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.030866288,0.044584636,0.034295876,0.010288762,0.0034295875,0.0034295875,0.006859175,0.0034295875,0.0034295875,0.01371835,0.037725464,0.072021335,0.07888051,0.041155048,0.061732575,0.13375391,0.20234565,0.16804978,0.1371835,0.23321195,0.3806842,0.548734,0.7579388,0.75450927,0.6276145,0.42869842,0.274367,0.35324752,0.4698535,0.23321195,0.034295876,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.044584636,0.12346515,0.31895164,0.6756287,1.1317638,1.6256244,2.0714707,2.3732746,2.3595562,2.1297739,1.7799559,1.3992717,0.97400284,0.6344737,0.47328308,0.4698535,0.51100856,0.4629943,0.4664239,0.5796003,0.805953,1.1043272,0.94999576,0.805953,0.6824879,0.61046654,0.6276145,0.45613512,0.33266997,0.274367,0.29494452,0.3806842,0.4389872,0.47328308,0.4115505,0.28465575,0.19891608,0.13375391,0.12003556,0.13032432,0.13375391,0.13032432,0.07545093,0.06859175,0.072021335,0.082310095,0.12346515,0.3566771,0.71678376,1.0425946,1.039165,0.2777966,0.16804978,0.16804978,0.26750782,0.4355576,0.65848076,0.7682276,1.1180456,1.8073926,2.6887965,3.3678548,3.1380725,2.8225505,3.069481,3.5873485,3.1380725,4.187526,4.9351764,5.178677,4.962613,4.5853586,4.07435,3.9371665,4.15666,4.6882463,5.4941993,5.9228973,5.0895076,4.314421,4.0846386,4.0366244,3.7622573,2.819121,2.510458,3.2478194,4.540774,4.866585,4.9488945,5.223262,5.8645945,6.7802944,9.551401,11.080997,12.106443,13.241637,14.970149,14.874121,12.758065,9.585697,6.447624,4.5442033,4.537344,5.086078,6.557371,9.3764925,14.027013,17.147938,17.720678,17.21996,17.339994,19.987637,22.103691,22.666143,21.27716,18.331144,15.0078745,12.9809885,10.604284,7.9772205,5.336438,3.0523329,1.6633499,0.823101,0.3566771,0.12003556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.20920484,0.33266997,0.45270553,0.7579388,1.611906,0.8265306,0.69963586,0.7099246,0.77165717,1.2277923,1.7353712,1.6804979,1.1934965,0.5144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09602845,0.09602845,0.048014224,0.0,0.0,0.044584636,0.13375391,0.33609957,0.6173257,0.85396725,1.097468,1.646202,2.1812177,2.5241764,2.6304936,2.860276,3.3747141,3.7862647,3.9474552,3.9440255,4.65395,4.852866,4.9214582,5.0449233,5.23698,3.9783216,2.5310357,1.3684053,0.6824879,0.37382504,0.39440256,0.31209245,0.18519773,0.06516216,0.0274367,0.116605975,0.31552204,0.48357183,0.6379033,0.96714365,1.3752645,1.7525192,2.0165975,2.1126258,2.0268862,2.0646117,2.253239,2.3664153,2.3252604,2.2086544,2.270387,2.6887965,3.7279615,5.312431,7.0478024,8.80718,9.815479,10.628291,10.655728,8.162418,7.3050213,6.783724,6.8454566,7.6033955,9.0369625,9.414218,8.834618,8.2310095,7.747438,6.756287,2.9082901,1.6187652,1.2895249,1.1832076,1.4027013,2.5207467,3.82399,4.8597255,5.4976287,5.950334,5.5422134,3.899441,2.0131679,0.64133286,0.29151493,0.1920569,0.274367,0.29151493,0.20920484,0.18519773,0.16804978,0.2503599,0.38754338,0.52815646,0.607037,0.5144381,0.5727411,0.48014224,0.20234565,0.0,0.037725464,0.09602845,0.09945804,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.0548734,0.10288762,0.18862732,0.28808534,0.39440256,0.47671264,0.53501564,0.5658819,0.5796003,0.5727411,0.48014224,0.32924038,0.18519773,0.07888051,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.006859175,0.006859175,0.020577524,0.0548734,0.08573969,0.061732575,0.017147938,0.041155048,0.09602845,0.16462019,0.26064864,0.32238123,0.29151493,0.18176813,0.07888051,0.14061308,0.26064864,0.15776102,0.044584636,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.061732575,0.26064864,0.65162164,1.138623,1.6324836,2.037175,2.294394,2.3321195,2.1469216,1.7971039,1.4335675,0.9774324,0.66876954,0.44584638,0.30523327,0.30523327,0.41840968,0.42526886,0.44584638,0.5796003,0.90198153,0.97400284,0.8711152,0.72707254,0.66876954,0.83681935,0.91227025,0.6893471,0.4938606,0.45956472,0.52815646,0.6173257,0.7613684,0.805953,0.67219913,0.34295875,0.26750782,0.23664154,0.20920484,0.17490897,0.16119061,0.13032432,0.14061308,0.1920569,0.23321195,0.18176813,0.23321195,0.5761707,1.1900668,1.6290541,1.0460242,0.40126175,0.15433143,0.12689474,0.18176813,0.23321195,0.26064864,0.37382504,0.61389613,0.9602845,1.3169615,1.6564908,1.8519772,2.1743584,2.5310357,2.4555845,3.625074,5.1580997,5.7822843,5.288424,4.537344,4.389872,3.8377085,4.0503426,5.0449233,5.689686,5.5079174,4.99005,4.2252517,3.566771,3.6319332,4.506478,4.5270553,4.0434837,3.5016088,3.4295874,3.5976372,3.858286,4.3452873,4.8905916,5.038064,7.7920227,10.302481,12.171606,13.437123,14.568888,15.151917,14.46257,12.836946,10.518545,7.6685576,5.9126086,4.6573796,4.434457,5.7068334,8.899779,12.123591,13.347955,13.186764,13.025573,15.0078745,19.586374,23.34863,24.85422,23.485815,19.44919,15.7966795,12.3911,9.417647,6.944915,4.9420357,3.4433057,2.3252604,1.5021594,0.84367853,0.18176813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.13375391,0.29151493,0.65162164,1.5090185,0.5007198,0.59674823,0.59674823,0.35324752,0.78194594,1.1729189,1.1626302,0.8505377,0.40126175,0.048014224,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06516216,0.16462019,0.29837412,0.4664239,0.6962063,1.0323058,1.4918705,2.0268862,2.7745364,3.7451096,4.5030484,5.0414934,5.802862,7.06495,6.7631464,6.186976,5.861165,5.5250654,4.201245,2.7402403,1.6599203,1.0768905,0.7373613,0.805953,0.5727411,0.29837412,0.14061308,0.17490897,0.15776102,0.15776102,0.17147937,0.18862732,0.18519773,0.3018037,0.4115505,0.6962063,1.138623,1.5501735,1.99602,2.7093742,3.649081,4.605936,5.1752477,4.9591837,5.3227196,6.4544835,8.165848,9.914937,11.458252,11.97269,12.596875,12.55229,9.177576,7.205563,6.526505,7.058091,8.460793,10.134431,10.88551,10.508256,10.696883,11.005547,8.855195,4.996909,3.8960114,4.170378,5.0586414,6.3961806,8.186425,9.709162,10.566559,10.5597,9.678296,7.891481,5.5730796,3.542764,2.5721905,3.3678548,3.9063,3.1312134,1.5947582,0.17147937,0.044584636,0.010288762,0.29494452,0.72707254,1.0666018,1.0220171,0.86082643,0.7922347,0.6001778,0.2709374,0.0,0.09259886,0.12346515,0.10288762,0.05144381,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.07545093,0.15090185,0.23321195,0.31209245,0.3841138,0.4389872,0.4629943,0.3841138,0.274367,0.17147937,0.09259886,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.024007112,0.024007112,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.017147938,0.01371835,0.058302987,0.072021335,0.048014224,0.010288762,0.017147938,0.058302987,0.061732575,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.15433143,0.45270553,0.85739684,1.2929544,1.6290541,1.862266,1.9171394,1.7799559,1.5124481,1.2277923,0.91569984,0.78537554,0.59331864,0.34295875,0.26750782,0.35324752,0.34638834,0.32924038,0.37725464,0.5624523,0.7099246,0.6962063,0.6241849,0.6173257,0.823101,0.9568549,0.78194594,0.61046654,0.5796003,0.66876954,0.78194594,1.0185875,1.1626302,1.0563129,0.59674823,0.42869842,0.35324752,0.31895164,0.2777966,0.20577525,0.15433143,0.15090185,0.2194936,0.31209245,0.30523327,0.274367,0.47328308,1.0288762,1.5364552,1.0700313,0.45956472,0.20577525,0.12689474,0.106317215,0.09602845,0.08916927,0.07545093,0.082310095,0.13032432,0.24350071,0.4664239,0.8505377,1.196926,1.4335675,1.6084765,2.3835633,3.7211025,4.773986,5.2644167,5.501058,5.9160385,5.284994,4.99005,5.394741,5.871454,4.8082814,4.249259,3.9543142,3.8205605,3.875434,4.6402316,5.079219,4.8322887,4.07435,3.508468,2.8637056,2.884283,3.3884325,4.029765,4.3178506,5.6313825,7.7714453,10.052121,12.044711,13.560589,14.627191,14.740367,14.695783,14.390549,12.812939,10.72775,8.436785,6.944915,6.831738,8.268735,10.861504,12.500846,12.5145645,11.283342,10.216741,13.214201,18.173384,22.748453,25.121729,24.02083,20.821026,16.767254,12.624311,8.999237,6.327589,4.616225,3.3987212,2.551613,1.8519772,0.9877212,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.06859175,0.082310095,0.082310095,0.11317638,0.14747226,0.19548649,0.26407823,0.37382504,0.35324752,1.0220171,1.0288762,0.36010668,0.3566771,0.490431,0.39097297,0.23664154,0.14747226,0.14404267,0.06859175,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.030866288,0.048014224,0.106317215,0.22292319,0.4629943,0.8745448,1.471293,2.3801336,3.542764,4.5956473,5.6519604,7.2775846,7.8777623,7.2707253,6.540223,6.0635104,5.4941993,4.266407,3.0077481,2.0989075,1.5707511,1.1077567,1.155771,0.96371406,0.64819205,0.3841138,0.4115505,0.30866286,0.14061308,0.030866288,0.037725464,0.14404267,0.4115505,0.3566771,0.52815646,1.0288762,1.5364552,2.1812177,3.192946,4.7328305,6.468202,7.579388,7.4284863,7.9257765,8.958082,10.028113,10.244178,9.72288,9.4862385,9.945804,10.511685,9.626852,7.8366075,7.0546613,7.4284863,8.766026,10.521975,12.490558,13.588025,15.326826,16.640358,13.862392,13.656617,14.400838,15.223939,15.268523,13.704632,13.745787,14.109323,14.201921,13.22106,10.14129,7.0615206,5.2301207,4.40702,4.756838,6.831738,7.915488,6.142391,2.9391565,0.14747226,0.0,0.0274367,0.39440256,0.9328478,1.3409687,1.1797781,1.0117283,0.78194594,0.48014224,0.18862732,0.058302987,0.2469303,0.216064,0.09602845,0.0,0.0034295875,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.044584636,0.07888051,0.13032432,0.18176813,0.20577525,0.19548649,0.16462019,0.12689474,0.08573969,0.041155048,0.010288762,0.0,0.0,0.0,0.0,0.0,0.020577524,0.058302987,0.09602845,0.116605975,0.1371835,0.106317215,0.061732575,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.01371835,0.030866288,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.01371835,0.024007112,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.037725464,0.17147937,0.4115505,0.7099246,0.9534253,1.1214751,1.2106444,1.214074,1.1214751,0.9362774,0.82996017,0.8676856,0.75450927,0.490431,0.3566771,0.2777966,0.25378948,0.26750782,0.3018037,0.34295875,0.36353627,0.4046913,0.44584638,0.5041494,0.65505123,0.64819205,0.6859175,0.75450927,0.84367853,0.939707,0.9911508,1.2963841,1.4747226,1.3512574,0.9568549,0.6790583,0.52815646,0.44584638,0.37725464,0.28808534,0.22292319,0.17833854,0.20920484,0.31209245,0.42183927,0.42526886,0.45956472,0.6824879,0.85396725,0.36696586,0.31209245,0.26750782,0.22635277,0.1920569,0.18862732,0.16804978,0.14061308,0.09602845,0.05144381,0.058302987,0.14747226,0.36353627,0.58988905,0.7922347,1.0014396,1.2003556,1.4027013,2.3595562,4.2183924,6.550512,7.795452,7.5107965,6.560801,5.641671,5.302142,4.033195,3.3369887,3.7965534,4.8734436,4.8905916,4.5990767,4.616225,4.557922,4.3761535,4.355576,3.2203827,2.6922262,2.750529,3.210094,3.7142432,3.0900583,3.7862647,5.9914894,9.139851,11.928105,13.687484,14.1299,14.898128,16.359133,17.607502,17.20967,15.241087,13.306799,12.271064,12.247057,13.790371,15.817257,16.61292,15.138199,11.005547,8.7283,11.417097,16.47231,21.685282,25.234905,25.289778,22.275171,17.484037,12.243628,7.9086285,5.3913116,3.858286,3.0111778,2.510458,1.9582944,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.20234565,0.34638834,0.4115505,0.4115505,0.5590228,0.7407909,0.881404,0.9362774,0.89855194,0.88826317,1.0048691,0.9294182,0.5658819,0.01371835,0.34638834,0.29837412,0.17833854,0.14404267,0.22978236,0.20577525,0.09602845,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.11317638,0.29837412,0.64133286,1.2380811,1.9823016,3.059192,4.2389703,4.897451,5.446185,6.125243,6.217842,5.579939,4.6402316,4.417309,3.8514268,2.9117198,1.8279701,1.0837497,0.8745448,0.90541106,0.84367853,0.65505123,0.59674823,0.5212973,0.29151493,0.09259886,0.044584636,0.22978236,0.64476246,0.6927767,1.4198492,2.7951138,3.724532,3.673088,3.4776018,3.5050385,3.9783216,5.003768,6.1904054,7.6651278,9.15014,10.014396,9.294182,6.924337,6.1046658,6.4579134,7.466212,8.453933,8.587687,7.8983397,7.160979,7.2638664,9.2153015,16.173935,24.823355,31.42874,34.49136,34.772587,37.73918,40.887543,40.119312,31.881445,13.169616,7.9943686,6.451054,6.824879,7.174697,5.3570156,3.8308492,2.452155,1.6324836,1.6221949,2.486451,2.2429502,0.9911508,0.12003556,0.0,0.0,0.13375391,0.21263443,0.39783216,0.64476246,0.71678376,0.607037,0.4046913,0.17490897,0.058302987,0.29151493,0.31552204,0.20920484,0.082310095,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.034295876,0.044584636,0.044584636,0.0548734,0.0548734,0.041155048,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0274367,0.11317638,0.23664154,0.33609957,0.48357183,0.42869842,0.274367,0.1097468,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.024007112,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0274367,0.082310095,0.18176813,0.36696586,0.5727411,0.6893471,0.72021335,0.6927767,0.65505123,0.65505123,0.6927767,0.6927767,0.6001778,0.3806842,0.23664154,0.13375391,0.07888051,0.072021335,0.12346515,0.13375391,0.17490897,0.2469303,0.36353627,0.53501564,0.6927767,1.0357354,1.5055889,1.879414,1.7696671,1.3924125,1.728512,1.9102802,1.6770682,1.371835,1.2380811,0.9568549,0.5693115,0.26407823,0.39783216,0.5178677,0.47671264,0.4081209,0.37382504,0.33609957,0.20234565,0.2777966,0.3806842,0.41498008,0.36696586,0.29151493,0.22978236,0.20920484,0.21263443,0.15090185,0.15090185,0.17833854,0.15090185,0.06859175,0.044584636,0.106317215,0.16804978,0.25378948,0.34295875,0.36696586,0.5727411,0.78194594,1.1180456,2.0817597,4.547633,7.64798,7.140401,5.7239814,4.420738,2.5790498,2.6407824,3.0214665,4.0846386,5.2301207,4.914599,4.972902,5.144381,4.314421,2.9254382,2.976882,5.0277753,5.3741636,4.7328305,3.7759757,3.1277838,3.1415021,2.8225505,4.122364,6.944915,9.156999,11.561139,12.655178,13.491997,14.935853,17.669235,19.085653,19.109661,18.015623,16.139639,13.869251,14.112752,17.689812,22.196291,25.056566,23.544119,17.28169,14.160767,14.092175,16.715809,21.37662,24.7822,24.912523,22.415783,18.005335,12.449403,7.970361,4.9180284,2.983741,1.9582944,1.7388009,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.06859175,0.082310095,0.082310095,0.11317638,0.15433143,0.22292319,0.32581082,0.47328308,0.53844523,0.5796003,0.6344737,0.6859175,0.6756287,0.48700142,0.31895164,0.4389872,0.90884066,1.5604624,1.4850113,1.0871792,0.64819205,0.36010668,0.32924038,0.32924038,0.3018037,0.23321195,0.13032432,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.061732575,0.14061308,0.3566771,0.7305021,1.2758065,1.9925903,2.8465576,3.532475,3.666229,3.4810312,3.2409601,3.2581081,3.4295874,3.3061223,2.9734523,2.5413244,2.1091962,1.8828435,1.4369972,1.0048691,0.805953,1.0597426,1.5433143,1.7833855,1.6496316,1.3478279,1.4129901,1.2517995,1.3101025,1.8759843,2.784825,3.4295874,3.292404,2.9665933,2.9631636,3.6147852,5.079219,6.036074,7.6925645,8.676856,8.220721,6.142391,5.446185,6.543653,8.05953,8.985519,8.683716,7.658269,6.927767,7.267296,9.537683,14.685493,20.70442,25.080574,26.593021,24.703318,19.552078,14.640909,12.507706,11.129011,8.64256,3.3678548,2.07833,1.7936742,2.4041407,3.3747141,3.7451096,3.3129816,2.585909,1.7456601,0.9774324,0.4972902,0.58645946,0.31209245,0.06859175,0.061732575,0.30523327,0.5453044,0.64476246,0.6173257,0.4938606,0.31552204,0.3018037,0.35324752,0.38754338,0.37382504,0.3018037,0.37382504,0.17490897,0.017147938,0.0,0.0034295875,0.18862732,0.09259886,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.010288762,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.01371835,0.044584636,0.08573969,0.116605975,0.21263443,0.22635277,0.17147937,0.07888051,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.037725464,0.08573969,0.14747226,0.18862732,0.216064,0.22635277,0.22978236,0.24007112,0.31552204,0.4081209,0.45613512,0.39440256,0.2469303,0.12346515,0.0548734,0.058302987,0.14747226,0.31552204,0.39440256,0.41840968,0.45613512,0.607037,0.823101,1.1797781,1.5398848,1.7422304,1.611906,1.4095604,1.5021594,1.5330256,1.3649758,1.08032,0.89855194,0.8093826,0.7133542,0.6241849,0.6893471,0.64476246,0.67219913,0.70649505,0.6344737,0.274367,0.16119061,0.16119061,0.20234565,0.22978236,0.2194936,0.16462019,0.11317638,0.12003556,0.15090185,0.09259886,0.061732575,0.07545093,0.09259886,0.10288762,0.106317215,0.08916927,0.12346515,0.16462019,0.18519773,0.17147937,0.29151493,0.4698535,0.85396725,1.6187652,2.9734523,4.8425775,5.7479887,5.7102633,5.23698,5.336438,4.605936,4.307562,5.7754254,7.956643,7.414768,6.5196457,5.3158607,3.957744,2.7128036,1.961724,2.9494452,4.173808,5.0414934,4.955754,3.309552,2.054323,1.9994495,2.527606,3.5118976,5.3227196,7.531374,9.942374,12.106443,13.9138365,15.594335,17.899017,19.500635,20.316875,20.131678,18.595222,17.686382,17.87501,19.720127,22.648996,24.970827,22.751883,18.560926,15.285671,14.308239,15.505165,20.436913,22.988525,23.094843,20.94792,17.003895,12.524854,8.694004,5.7274113,3.532475,1.7388009,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.06859175,0.14747226,0.18176813,0.19548649,0.23321195,0.3018037,0.3806842,0.41498008,0.7099246,1.1626302,1.5261664,1.4267083,1.0700313,0.7510797,0.52815646,0.42183927,0.42183927,0.42183927,0.40126175,0.34638834,0.23664154,0.05144381,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0548734,0.16462019,0.34981793,0.66533995,1.2072148,1.7902447,2.136633,2.5001693,3.0283258,3.782835,3.7965534,3.690236,3.5770597,3.5564823,3.7005248,3.4467354,2.9151495,2.369845,2.0749004,2.2738166,3.2546785,4.180667,4.602506,4.4859004,4.2081037,3.4192986,2.8156912,2.5756202,2.7779658,3.4124396,4.0880685,4.3487167,4.434457,4.65395,5.3707337,7.6205435,7.301592,5.9571934,4.6127954,3.7622573,5.693115,8.625413,10.316199,9.743458,7.1232533,5.6210938,5.147811,5.4804807,6.5333643,8.361334,10.545981,12.082437,12.329367,10.906088,7.671987,4.4927597,2.9185789,2.5481834,2.393852,0.88826317,0.61389613,0.97057325,1.9514352,3.1415021,3.690236,3.0111778,2.8259802,2.253239,1.2620882,0.65162164,0.72707254,0.7579388,0.7373613,0.70306545,0.764798,0.8505377,0.881404,0.8676856,0.7579388,0.432128,0.40126175,0.6310441,0.78537554,0.75450927,0.65162164,0.6344737,0.4389872,0.25721905,0.16462019,0.12003556,0.23321195,0.12689474,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.024007112,0.058302987,0.07545093,0.06859175,0.037725464,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.024007112,0.037725464,0.05144381,0.058302987,0.061732575,0.1097468,0.19548649,0.2777966,0.26750782,0.16462019,0.082310095,0.041155048,0.061732575,0.14404267,0.28465575,0.37382504,0.47328308,0.6344737,0.881404,1.1660597,1.3169615,1.3649758,1.3101025,1.1214751,1.0151579,1.0837497,1.1146159,1.0014396,0.7407909,0.6927767,0.67219913,0.6927767,0.7407909,0.7888051,0.7476501,0.7133542,0.66876954,0.5693115,0.34981793,0.2194936,0.17490897,0.15776102,0.14061308,0.12003556,0.07888051,0.048014224,0.06516216,0.12003556,0.14061308,0.10288762,0.06859175,0.09602845,0.19548649,0.32238123,0.22978236,0.15776102,0.12689474,0.116605975,0.08573969,0.17490897,0.37725464,0.7442205,1.3169615,2.1126258,4.5030484,5.4907694,5.552502,5.2918534,5.4599032,4.846007,4.314421,4.7431192,6.0566516,7.208993,6.5059276,5.23698,4.5819287,4.5270553,3.8617156,2.9631636,3.1826572,3.8891523,4.3795834,3.8891523,2.0406046,1.5981878,1.6084765,1.9102802,3.1380725,4.5956473,6.619104,8.755736,10.768905,12.63117,14.997586,17.463459,19.764713,21.43835,21.836184,21.150267,19.925903,19.510923,20.382038,22.144846,22.340332,20.135109,17.051908,14.568888,14.085316,16.156786,19.12681,21.153696,21.287449,19.459478,16.283682,13.05301,9.897789,6.9209075,4.201245,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.017147938,0.044584636,0.20577525,0.58302987,0.96371406,1.0906088,0.66876954,0.34638834,0.216064,0.20920484,0.2503599,0.274367,0.47328308,0.5453044,0.432128,0.20577525,0.05144381,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.09945804,0.29151493,0.6310441,1.0768905,1.7113642,2.5378947,3.4913201,3.7622573,3.9097297,4.108646,4.4413157,4.928317,4.698535,4.3658648,4.1429415,4.125794,4.2698364,5.6348124,6.574519,6.958633,6.866034,6.5642304,6.101236,5.3570156,4.4687524,3.765687,3.7519686,4.605936,5.0312047,5.079219,4.8185706,4.338428,6.0840883,5.0174866,3.3472774,2.4315774,2.7916842,5.055212,7.3050213,7.9772205,6.6739774,4.170378,3.5599117,3.8960114,4.57164,5.0003386,4.6093655,4.0606318,3.782835,3.5530527,3.2546785,2.8637056,2.1434922,1.6359133,1.5844694,1.6153357,0.72364295,0.4972902,0.89855194,1.8725548,3.083199,3.9200184,3.758828,3.9680326,3.8342788,3.309552,3.000889,2.767677,2.4384367,2.0268862,1.605047,1.2963841,1.2415106,1.2037852,1.1763484,1.08032,0.7682276,0.66876954,0.77508676,0.8128122,0.7373613,0.72707254,0.78194594,0.6962063,0.5041494,0.31552204,0.32581082,0.30523327,0.22292319,0.15776102,0.12689474,0.07888051,0.017147938,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.0274367,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.034295876,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0034295875,0.006859175,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.024007112,0.06516216,0.116605975,0.12346515,0.07888051,0.037725464,0.020577524,0.041155048,0.09602845,0.16804978,0.2503599,0.39097297,0.61046654,0.91227025,1.1660597,1.1523414,1.0288762,0.89169276,0.7510797,0.7133542,0.805953,0.89169276,0.89169276,0.78537554,0.7990939,0.7510797,0.7133542,0.70306545,0.69963586,0.6927767,0.65848076,0.6241849,0.6036074,0.61389613,0.53158605,0.6173257,0.5453044,0.29837412,0.17490897,0.15776102,0.19891608,0.26750782,0.33266997,0.34295875,0.274367,0.274367,0.35324752,0.50757897,0.7133542,0.5658819,0.34981793,0.18519773,0.1097468,0.072021335,0.14061308,0.34295875,0.6310441,1.0323058,1.6496316,3.6044965,4.2938433,4.482471,4.6608095,5.0620713,5.1683884,4.8905916,4.605936,4.852866,6.355026,5.7377,4.6916757,4.2698364,4.636802,5.099797,4.3041325,3.7176728,3.3987212,3.350707,3.5461934,3.1792276,2.7368107,2.1400626,1.7422304,2.3424082,3.1140654,4.3041325,5.645101,7.1026754,8.882631,11.231899,13.989287,16.722668,19.250275,21.623549,22.422644,22.093403,21.506943,21.218857,21.496655,22.179142,22.007662,20.584383,18.434032,17.017612,16.005884,17.329706,19.21255,20.460918,20.481497,18.897026,16.736387,14.212211,11.461681,8.567109,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0034295875,0.017147938,0.037725464,0.4355576,0.58988905,0.4081209,0.072021335,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.037725464,0.13032432,0.33266997,0.6824879,1.1866373,1.8313997,2.6236343,3.2272418,3.8617156,4.557922,5.144381,5.127233,5.1512403,5.422178,5.830299,5.9743414,7.239859,7.6171136,7.596536,7.514226,7.56224,7.747438,7.2021337,6.060081,4.6848164,3.673088,3.9165888,4.091498,4.190956,3.9371665,2.8122618,2.4075704,2.1846473,2.1846473,2.452155,3.0557625,3.4707425,3.1415021,2.3424082,1.5055889,1.2277923,1.9994495,3.0797696,4.3349986,5.425607,5.796003,5.007198,3.9543142,3.093488,2.8019729,3.3644254,2.8122618,2.153781,1.4850113,0.90884066,0.5212973,0.33952916,0.4389872,1.0151579,2.1915064,4.0194764,5.2609873,5.7377,6.0806584,6.495639,6.756287,6.447624,5.6348124,4.465323,3.1517909,1.9685832,1.7250825,1.6221949,1.5193073,1.3409687,1.0734608,0.82996017,0.6173257,0.44584638,0.36010668,0.42869842,0.64133286,0.6824879,0.5453044,0.38754338,0.53844523,0.4664239,0.432128,0.38754338,0.31552204,0.22978236,0.05144381,0.020577524,0.034295876,0.041155048,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.058302987,0.058302987,0.01371835,0.017147938,0.010288762,0.0034295875,0.0,0.006859175,0.01371835,0.037725464,0.058302987,0.0548734,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.006859175,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.024007112,0.024007112,0.010288762,0.0,0.006859175,0.0274367,0.082310095,0.16462019,0.26407823,0.39440256,0.61046654,0.7305021,0.66876954,0.58988905,0.5590228,0.5453044,0.6036074,0.7373613,0.90541106,1.0631721,1.1523414,1.0940384,0.96371406,0.8025235,0.65848076,0.607037,0.58988905,0.6241849,0.69963586,0.805953,0.90884066,0.91569984,1.1763484,1.0837497,0.64819205,0.490431,0.48700142,0.58988905,0.69963586,0.7442205,0.6790583,0.6379033,0.6756287,0.7682276,0.89855194,1.0563129,0.89169276,0.65162164,0.4046913,0.2194936,0.12346515,0.14404267,0.29151493,0.4629943,0.71678376,1.2792361,1.7730967,2.277246,2.8294096,3.5187566,4.5030484,5.4633327,5.895461,5.994919,6.0395036,6.3790326,5.593657,4.633373,3.8137012,3.6285036,4.7499785,5.2747054,4.8117113,3.7485392,2.6853669,2.4418662,4.262977,4.523626,3.690236,2.6236343,2.551613,3.0283258,3.57363,3.940596,4.32471,5.360445,7.582818,10.1481495,12.456262,14.730078,18.025911,20.587814,22.463799,23.592133,24.010542,23.86307,23.852781,24.43238,24.497543,23.413794,21.0268,18.787281,17.929884,18.28999,19.394318,20.45063,20.28944,19.29143,17.775553,15.8138275,13.203912,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.058302987,0.12003556,0.23321195,0.42869842,0.72021335,1.2517995,2.0646117,3.059192,3.998899,4.5853586,4.9591837,5.178677,5.267846,5.219832,5.195825,5.535354,6.262427,7.085528,7.414768,6.293293,4.73969,3.3952916,2.4247184,1.5124481,1.6084765,2.2841053,3.210094,3.957744,3.981751,3.433017,2.983741,2.8019729,2.9803114,3.5564823,3.433017,2.3046827,1.2620882,0.77508676,0.70306545,0.90884066,1.1729189,1.5673214,2.0234566,2.3046827,2.510458,2.170929,1.704505,1.5090185,1.9239986,2.1057668,1.9514352,1.5398848,1.0220171,0.59674823,0.47328308,0.39783216,0.6824879,1.8108221,4.4104495,6.0806584,6.783724,7.5210853,8.735159,10.285333,11.125582,10.813489,9.1981535,6.4373355,3.0043187,2.1263442,1.8897027,1.8416885,1.6599203,1.1592005,0.5727411,0.29151493,0.1920569,0.18176813,0.18176813,0.18176813,0.1920569,0.26064864,0.4046913,0.6241849,0.69963586,0.7442205,0.6173257,0.38754338,0.34981793,0.09602845,0.09602845,0.17490897,0.20577525,0.106317215,0.034295876,0.006859175,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.05144381,0.07545093,0.08916927,0.0548734,0.017147938,0.006859175,0.030866288,0.06859175,0.08573969,0.0548734,0.006859175,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.1371835,0.26064864,0.31552204,0.29151493,0.24350071,0.20920484,0.15433143,0.12346515,0.13032432,0.16804978,0.40126175,0.6962063,1.0082988,1.2517995,1.313532,1.1660597,0.9568549,0.8196714,0.8162418,0.89855194,0.8162418,0.7922347,0.83681935,0.89855194,0.8848336,0.8711152,0.91569984,0.91569984,0.9294182,1.1763484,1.1008976,1.0940384,1.08032,1.0597426,1.0837497,1.3032433,1.138623,0.96714365,0.922559,0.8848336,0.7510797,0.881404,0.85739684,0.5761707,0.26064864,0.20920484,0.24350071,0.29151493,0.40126175,0.71678376,1.2792361,1.7490896,2.0165975,2.1469216,2.3664153,3.707384,5.178677,6.5642304,7.658269,8.268735,8.014946,7.1712675,6.7322803,6.385892,4.5167665,3.2478194,3.2135234,3.1895163,2.7333813,2.1983654,2.8088322,4.0674906,4.647091,4.173808,3.234101,3.8685746,3.9543142,3.758828,3.6285036,3.981751,5.1683884,7.0923867,9.112414,11.043272,13.169616,15.916716,18.938183,21.592682,23.485815,24.473536,24.415234,24.7822,24.837072,23.554407,19.6241,18.04649,17.600643,17.837284,18.495766,19.486916,20.69413,21.061096,20.107672,17.977898,15.426285,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.12346515,0.37725464,0.4664239,0.26064864,0.06516216,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.020577524,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.048014224,0.09602845,0.216064,0.42526886,0.8676856,1.5844694,2.4967396,3.2786856,3.899441,4.461893,4.931747,5.144381,5.9297566,6.159539,6.252138,6.3035817,6.0978065,4.9248877,3.566771,2.651071,2.2360911,1.7799559,1.5536032,1.5330256,1.762808,2.1126258,2.2738166,2.3286898,2.3561265,2.352697,2.2841053,2.0646117,1.5913286,1.3512574,1.1180456,0.7956643,0.42183927,0.4424168,0.432128,0.490431,0.65505123,0.8745448,1.2998136,1.5947582,1.7147937,1.6976458,1.704505,1.9137098,2.0749004,1.99602,1.6427724,1.1077567,0.8093826,0.5521636,0.59674823,1.2449403,2.7985435,4.372724,5.686256,7.1781263,9.115844,11.616013,12.583157,11.746337,8.992378,5.2781353,2.6407824,1.7799559,1.6564908,2.061182,2.6613598,2.9906003,1.8759843,1.0425946,0.6001778,0.50757897,0.58645946,0.45956472,0.33952916,0.31895164,0.37382504,0.37039545,0.5693115,0.4115505,0.274367,0.29837412,0.38754338,0.36696586,0.38754338,0.41840968,0.3806842,0.15433143,0.034295876,0.0,0.0,0.0,0.0,0.061732575,0.044584636,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.034295876,0.08573969,0.09945804,0.07545093,0.044584636,0.037725464,0.05144381,0.06859175,0.12346515,0.13032432,0.09259886,0.041155048,0.0548734,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.020577524,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.037725464,0.08573969,0.116605975,0.116605975,0.09602845,0.08916927,0.072021335,0.05144381,0.041155048,0.058302987,0.14404267,0.3018037,0.45956472,0.5693115,0.5796003,0.5212973,0.44927597,0.4046913,0.4081209,0.48357183,0.45956472,0.42183927,0.39097297,0.37725464,0.3841138,0.39097297,0.41840968,0.4424168,0.48700142,0.61389613,0.6859175,0.8093826,0.9294182,1.0357354,1.155771,1.2792361,1.3238207,1.4747226,1.6599203,1.5570327,1.2072148,1.0494537,0.91227025,0.78194594,0.7956643,0.6207553,0.3806842,0.24007112,0.26750782,0.44927597,0.8848336,1.3889829,1.6942163,1.8142518,2.037175,3.57363,4.955754,6.3447366,7.517656,7.8537555,6.574519,5.796003,5.9400454,6.478491,5.967482,4.8151407,3.6627994,2.7333813,2.0817597,1.5741806,1.9514352,2.8156912,3.8102717,4.3281393,3.5153272,3.292404,3.426158,3.2786856,2.8877127,2.9563043,3.4192986,4.636802,6.2418494,7.8434668,9.030104,10.333347,12.442543,15.391989,18.691252,21.349182,22.813616,23.900795,24.511261,24.147726,21.904776,20.018501,19.46291,19.377169,19.239986,18.862732,19.476627,20.755863,20.79016,19.085653,16.561478,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.18862732,0.23321195,0.13032432,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.020577524,0.034295876,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.09602845,0.26407823,0.5693115,1.0048691,1.5638919,2.1469216,2.8259802,3.542764,4.1017866,4.7602673,4.972902,5.06893,5.1169443,4.945465,3.957744,2.877424,2.3629858,2.452155,2.5413244,2.311542,1.8519772,1.4369972,1.2243627,1.2895249,1.7216529,2.0989075,2.2738166,2.0714707,1.2826657,0.8093826,0.66191036,0.61046654,0.5178677,0.32238123,0.30523327,0.36010668,0.3806842,0.36353627,0.4081209,0.6962063,1.0597426,1.3478279,1.5604624,1.8588364,2.393852,2.8156912,2.9220085,2.5653315,1.6290541,1.5947582,1.1077567,0.7990939,1.0494537,1.9823016,3.5942078,5.24041,6.447624,7.6342616,10.134431,11.832077,12.010415,9.767465,5.844017,2.603057,1.9480057,2.5996273,3.6079261,4.3007026,4.280125,3.1826572,1.8931323,1.0768905,0.85739684,0.8162418,0.64133286,0.4938606,0.35324752,0.23664154,0.20577525,0.31209245,0.2503599,0.19548649,0.2709374,0.52472687,0.7442205,0.7407909,0.53501564,0.24350071,0.07545093,0.01371835,0.0,0.0,0.0,0.0,0.030866288,0.034295876,0.024007112,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.041155048,0.05144381,0.058302987,0.058302987,0.07545093,0.09259886,0.07545093,0.44584638,0.6001778,0.51100856,0.274367,0.08916927,0.09259886,0.07545093,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.017147938,0.017147938,0.01371835,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.0274367,0.030866288,0.024007112,0.030866288,0.030866288,0.020577524,0.010288762,0.030866288,0.06516216,0.15090185,0.216064,0.23664154,0.22292319,0.17833854,0.15090185,0.13032432,0.12346515,0.16119061,0.16462019,0.14404267,0.116605975,0.09945804,0.10288762,0.12346515,0.14061308,0.17147937,0.22635277,0.31895164,0.48014224,0.7442205,1.0117283,1.2346514,1.4404267,1.529596,1.5604624,1.6359133,1.7559488,1.8245405,2.0063086,1.9582944,1.5947582,1.1454822,1.1420527,0.939707,0.607037,0.36010668,0.28465575,0.34638834,0.5555932,0.91912943,1.1866373,1.3238207,1.4850113,2.5378947,3.4398763,4.57507,5.703404,5.9571934,5.0620713,4.605936,4.7534084,5.254128,5.470192,4.8768735,4.166949,3.758828,3.673088,3.5153272,3.093488,2.9048605,3.234101,3.9611735,4.5647807,2.750529,2.5241764,2.6579304,2.5756202,2.369845,2.6887965,3.1963756,3.9954693,4.9831905,5.826869,6.5024977,7.9463544,10.542552,14.143619,18.060207,20.834743,22.590693,23.334913,22.94051,21.167414,19.480057,20.12139,21.167414,21.565247,21.11597,20.567236,20.724997,20.220848,18.362011,15.107333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.017147938,0.0034295875,0.0,0.0034295875,0.010288762,0.010288762,0.024007112,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.037725464,0.082310095,0.15433143,0.3841138,0.69963586,1.1489118,1.7147937,2.318401,2.8088322,3.333559,3.8445675,4.122364,3.7725463,3.3232703,2.983741,2.8945718,3.1140654,3.6147852,3.724532,3.2581081,2.4761622,1.6976458,1.3066728,1.6427724,2.0028791,2.2909644,2.2429502,1.4095604,1.0940384,0.823101,0.5761707,0.3841138,0.32924038,0.51100856,0.7888051,1.0082988,1.0425946,0.78194594,0.69963586,0.85739684,1.1797781,1.6599203,2.352697,2.959734,3.3232703,3.5599117,3.6627994,3.5016088,3.2409601,2.4041407,1.7216529,1.6187652,2.2155135,4.125794,5.7377,6.5950966,7.332458,9.647429,11.461681,12.3533745,11.026124,7.5382333,3.316411,2.1091962,3.4776018,5.1409516,5.885172,5.56965,4.57164,2.983741,1.6907866,1.0494537,0.8745448,0.65505123,0.50757897,0.35324752,0.19548649,0.15433143,0.19548649,0.2709374,0.31895164,0.36010668,0.52472687,0.8848336,0.94999576,0.6790583,0.2469303,0.058302987,0.017147938,0.010288762,0.017147938,0.024007112,0.024007112,0.024007112,0.07888051,0.07888051,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.030866288,0.044584636,0.07888051,0.12003556,0.13032432,0.70649505,1.3101025,1.3615463,0.8128122,0.15090185,0.11317638,0.12003556,0.106317215,0.058302987,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0274367,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.01371835,0.01371835,0.024007112,0.034295876,0.06859175,0.08916927,0.07888051,0.06859175,0.044584636,0.034295876,0.020577524,0.010288762,0.0274367,0.0548734,0.07545093,0.06516216,0.037725464,0.024007112,0.024007112,0.030866288,0.0548734,0.1097468,0.18862732,0.37039545,0.66533995,0.97057325,1.2312219,1.4472859,1.5330256,1.5536032,1.5604624,1.6153357,1.7833855,2.311542,2.5721905,2.311542,1.7765263,1.7319417,1.4095604,1.0528834,0.78537554,0.6310441,0.51100856,0.4355576,0.5555932,0.72707254,0.881404,1.0220171,1.6153357,2.1263442,2.7916842,3.4535947,3.5633414,3.333559,3.3369887,3.5564823,3.9303071,4.3624353,4.523626,4.8151407,4.7774153,4.372724,3.998899,3.673088,3.7794054,4.3624353,4.887162,4.2595477,2.318401,2.0406046,3.1620796,4.465323,3.7862647,3.0969174,3.0523329,3.1483612,3.3198407,3.9268777,4.173808,5.2438393,7.507367,11.012405,15.470869,18.931322,20.793589,21.157125,20.388897,19.11652,18.488907,19.898466,21.633839,22.717587,22.926792,22.165424,21.311457,19.70298,16.698662,11.7086115,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.072021335,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.07545093,0.22978236,0.5453044,1.0117283,1.8313997,2.6785078,3.1243541,2.6476414,3.0626216,3.6147852,3.8445675,3.865145,4.3487167,4.7191124,4.48933,3.7622573,2.8705647,2.3904223,2.0680413,2.0063086,2.2395205,2.49331,2.201795,2.1057668,1.7559488,1.1832076,0.6310441,0.5212973,1.0220171,1.3889829,1.6770682,1.7525192,1.2895249,1.0048691,1.0014396,1.3272504,1.9720128,2.860276,3.223812,3.3198407,3.6456516,4.434457,5.672538,4.9591837,3.9268777,3.0043187,2.534465,2.7539587,5.353586,7.0375133,7.9257765,8.690575,10.569988,11.808069,12.583157,12.048141,9.630281,5.0277753,2.486451,3.6182148,5.5902276,6.852316,7.143831,6.3207297,4.650521,2.877424,1.5673214,1.0700313,0.69963586,0.490431,0.36353627,0.2777966,0.22292319,0.28465575,0.39097297,0.4698535,0.48357183,0.42526886,0.823101,1.0734608,0.9602845,0.5590228,0.25378948,0.08573969,0.034295876,0.034295876,0.05144381,0.058302987,0.05144381,0.1371835,0.12346515,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05144381,0.18862732,0.33266997,0.29837412,0.97400284,2.2326615,2.668219,1.8965619,0.58645946,0.216064,0.14747226,0.16119061,0.14061308,0.072021335,0.034295876,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.048014224,0.030866288,0.006859175,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.017147938,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.030866288,0.034295876,0.0274367,0.020577524,0.037725464,0.08916927,0.14747226,0.14747226,0.10288762,0.09602845,0.041155048,0.024007112,0.037725464,0.072021335,0.13032432,0.28122616,0.4938606,0.7373613,0.9842916,1.2003556,1.2963841,1.3752645,1.4164196,1.4369972,1.5090185,1.8931323,2.3595562,2.4727325,2.311542,2.4727325,1.9308578,1.5947582,1.430138,1.3238207,1.0734608,0.77851635,0.69963586,0.7373613,0.8162418,0.8711152,1.2415106,1.5947582,1.8039631,1.8313997,1.7319417,1.8073926,2.2052248,2.7539587,3.2581081,3.4844608,4.0263357,4.9694724,4.928317,3.882293,3.1689389,3.7279615,5.0140567,6.3653145,6.3790326,2.9117198,1.961724,1.8554068,3.74168,6.217842,5.3261495,3.6525106,3.4913201,3.3026927,2.8534167,3.2272418,3.1586502,3.9440255,5.826869,8.865483,12.932974,16.352274,18.139088,18.605513,18.30028,17.995045,18.663815,19.840164,21.102251,22.158566,22.847912,22.86163,22.035099,19.723558,15.37827,8.536243,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.044584636,0.12003556,0.3018037,0.6310441,1.1489118,1.8931323,3.333559,3.9131594,4.040054,3.9337368,3.6147852,3.275256,3.0077481,2.8054025,3.0248961,4.3795834,2.9151495,2.2086544,2.0508933,2.311542,2.9460156,3.1655092,2.7059445,1.9548649,1.3032433,1.1454822,1.7422304,1.6736387,1.2072148,0.71678376,0.65505123,0.9842916,1.2243627,1.4678634,1.8965619,2.760818,2.9700227,3.093488,3.4227283,4.012617,4.6848164,4.7808447,4.331569,3.5050385,2.568761,1.862266,5.6348124,8.570539,9.764035,9.626852,9.932085,10.957532,11.55428,11.907528,11.2421875,7.8126,4.0263357,2.9185789,4.1635194,6.7665763,9.047252,8.889491,7.4113383,5.446185,3.549623,1.9994495,1.2655178,0.7888051,0.48014224,0.31895164,0.3806842,0.4424168,0.40126175,0.3841138,0.4355576,0.53501564,0.9602845,1.4267083,1.4610043,1.0837497,0.77851635,0.29151493,0.06859175,0.006859175,0.020577524,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2194936,0.7339317,1.1523414,0.64133286,1.7147937,3.4947495,4.4413157,3.8925817,2.0749004,0.65848076,0.21263443,0.15776102,0.17147937,0.18176813,0.13375391,0.06859175,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.072021335,0.072021335,0.041155048,0.01371835,0.0034295875,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.044584636,0.034295876,0.01371835,0.0,0.061732575,0.12346515,0.12689474,0.12346515,0.24350071,0.1097468,0.06859175,0.0548734,0.044584636,0.044584636,0.15433143,0.32924038,0.5555932,0.84367853,1.2346514,1.3821237,1.4747226,1.3992717,1.2037852,1.0666018,1.1420527,1.2895249,1.5090185,1.9102802,2.7162333,2.0680413,1.8416885,1.9720128,2.2223728,2.1983654,1.9891608,1.9480057,1.8485477,1.5913286,1.1763484,1.2723769,1.5090185,1.704505,1.7422304,1.5707511,1.4747226,1.9068506,2.7745364,3.532475,3.2032347,2.8396983,3.2581081,3.9851806,4.7191124,5.3398676,5.888602,6.310441,6.159539,5.1683884,3.2649672,1.5433143,0.9294182,1.0117283,1.3821237,1.6633499,2.2360911,2.784825,2.8877127,2.7368107,3.1277838,3.3232703,3.4638834,4.1155047,5.658819,8.272165,11.153018,13.96871,17.093063,19.86417,20.584383,21.181131,21.699,21.815605,21.554956,21.287449,21.650986,21.568676,19.977346,16.067617,9.294182,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.034295876,0.08573969,0.216064,0.5178677,1.1351935,1.7662375,2.1503513,2.3904223,2.5584722,2.6887965,2.8156912,2.6064866,2.4418662,2.510458,2.7916842,2.5790498,2.4624438,2.4075704,2.428148,2.603057,2.959734,3.1209247,2.819121,2.2463799,2.061182,2.1297739,2.2669573,2.07833,1.6187652,1.3649758,2.4830213,3.3232703,2.9391565,1.937717,2.4795918,2.4041407,2.8122618,3.415869,3.9851806,4.355576,4.8151407,4.8494368,4.461893,4.341858,5.8405876,8.488229,10.964391,12.960411,14.2533655,14.692352,12.264205,10.741467,10.405369,10.593996,9.692014,6.3378778,4.0537724,3.649081,5.178677,7.949784,10.113853,9.716022,8.028665,5.8988905,3.7451096,2.270387,1.2792361,0.7442205,0.5658819,0.5761707,0.75450927,0.6859175,0.58302987,0.53844523,0.51100856,1.0734608,1.2792361,1.0906088,0.6893471,0.45956472,0.23664154,0.07888051,0.01371835,0.020577524,0.044584636,0.037725464,0.058302987,0.08916927,0.08916927,0.0,0.0,0.0,0.048014224,0.1097468,0.061732575,0.020577524,0.0548734,0.106317215,0.106317215,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05144381,0.19891608,0.3566771,0.32238123,0.6173257,1.6359133,2.6887965,3.1963756,2.6853669,1.8759843,1.3546871,0.8676856,0.4389872,0.35324752,0.29494452,0.17490897,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.0274367,0.0274367,0.01371835,0.01371835,0.034295876,0.0548734,0.061732575,0.06516216,0.09602845,0.05144381,0.06859175,0.09259886,0.11317638,0.13032432,0.18176813,0.20234565,0.23664154,0.3018037,0.37039545,0.42869842,0.5178677,0.58302987,0.6207553,0.70306545,0.78537554,0.881404,0.980862,1.1523414,1.5673214,1.8691251,1.8931323,1.8073926,1.7319417,1.7456601,1.8108221,1.9754424,2.0440342,1.9068506,1.5398848,2.1091962,2.4452958,2.4555845,2.2326615,2.0714707,2.1503513,2.3424082,2.4555845,2.4590142,2.4590142,2.6304936,3.5221863,4.448175,4.9488945,4.791134,5.1066556,4.8837323,4.5647807,4.232111,3.6079261,2.3732746,1.6187652,1.3375391,1.4129901,1.6256244,1.6942163,1.8999915,2.301253,2.8396983,3.3472774,3.7965534,4.1017866,4.712253,5.7411294,6.975781,8.128122,10.103564,13.214201,16.684942,18.656956,19.233126,19.277712,19.065077,18.811287,18.650097,19.023922,19.473198,18.996485,16.732958,11.941824,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.044584636,0.15433143,0.432128,0.69963586,0.9294182,1.1660597,1.4335675,1.7422304,1.9514352,2.0989075,2.1846473,2.311542,2.651071,2.6407824,2.5619018,2.568761,2.726522,3.0317552,3.7142432,3.8205605,3.6319332,3.340418,3.0214665,2.8225505,2.6750782,2.3286898,1.845118,1.605047,2.8808534,3.566771,3.525616,3.3198407,4.2218223,4.245829,4.170378,4.184097,4.1943855,3.8514268,4.482471,4.722542,5.1100855,6.0052075,7.596536,8.89635,10.172156,12.298501,15.704081,20.399187,14.757515,11.05699,9.451943,9.537683,10.347065,8.467651,5.813151,4.314421,4.705394,6.5299344,9.935514,11.396519,11.132441,9.362774,6.2967224,3.5153272,1.9891608,1.1866373,0.84367853,0.94656616,1.2860953,1.0940384,0.86082643,0.84024894,1.0425946,1.3032433,1.2003556,1.2106444,1.2860953,0.8676856,0.5693115,0.274367,0.09259886,0.048014224,0.072021335,0.08916927,0.13032432,0.14404267,0.10288762,0.010288762,0.0034295875,0.12689474,0.20234565,0.15776102,0.041155048,0.020577524,0.030866288,0.05144381,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.017147938,0.010288762,0.030866288,0.07545093,0.12346515,0.26750782,0.71678376,1.5707511,2.417859,2.3424082,1.7799559,1.5227368,1.155771,0.6344737,0.26750782,0.29494452,0.16804978,0.072021335,0.0548734,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.034295876,0.041155048,0.034295876,0.030866288,0.05144381,0.058302987,0.044584636,0.034295876,0.037725464,0.06516216,0.09945804,0.116605975,0.09602845,0.106317215,0.09602845,0.10288762,0.12003556,0.106317215,0.09945804,0.13032432,0.1920569,0.2777966,0.3806842,0.45956472,0.5212973,0.59674823,0.71678376,0.91569984,1.3272504,1.605047,1.7353712,1.7765263,1.8416885,1.8588364,2.0989075,2.2498093,2.201795,2.0165975,2.7093742,3.2375305,3.1689389,2.6407824,2.3801336,2.486451,2.5927682,2.6373527,2.5927682,2.4658735,2.3972816,2.983741,3.9165888,4.712253,4.7191124,4.396731,4.3624353,4.465323,4.479041,4.0777793,4.4241676,3.957744,2.836269,1.7422304,1.8999915,1.8039631,1.5913286,1.5810398,1.9582944,2.7882545,3.4638834,4.262977,5.586798,7.3839016,9.160428,9.201583,9.438225,10.731179,12.843805,14.438563,14.30138,14.339106,14.723219,15.364552,15.913286,16.582056,17.391438,17.751545,16.928444,14.023583,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.048014224,0.072021335,0.01371835,0.0034295875,0.017147938,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0548734,0.15090185,0.25721905,0.4081209,0.61389613,0.8745448,1.0597426,1.4678634,1.7182233,1.821111,2.1880767,2.3286898,2.4452958,2.627064,2.8980014,3.2272418,3.9783216,4.57164,4.746549,4.523626,4.2046742,4.0846386,3.6970954,3.1620796,2.7093742,2.6922262,3.3884325,3.82399,3.9646032,4.1326528,4.9934793,5.7411294,5.7377,5.06893,4.1292233,3.6182148,4.2046742,4.523626,5.3913116,7.051232,9.187865,10.508256,10.271614,11.146159,14.466,20.21056,15.285671,11.657167,9.647429,9.283894,10.302481,9.661148,7.473071,5.7308407,5.4084597,6.444195,10.432805,12.902108,13.598314,12.500846,9.815479,5.861165,3.4981792,2.2600982,1.7525192,1.6359133,1.5741806,1.2037852,0.9877212,1.1111864,1.471293,1.2826657,1.0048691,1.1111864,1.4335675,1.1523414,0.77851635,0.45613512,0.26750782,0.1920569,0.10288762,0.13375391,0.17490897,0.20577525,0.19548649,0.09602845,0.06859175,0.21263443,0.28465575,0.22292319,0.1371835,0.11317638,0.12346515,0.07888051,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09259886,0.31209245,0.64133286,1.0323058,1.3752645,1.6633499,1.9068506,2.1194851,2.1023371,1.9514352,2.1400626,2.5001693,2.253239,1.546744,1.2037852,0.939707,0.607037,0.20920484,0.3841138,0.33266997,0.22978236,0.15776102,0.072021335,0.058302987,0.024007112,0.0034295875,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.006859175,0.020577524,0.0548734,0.09259886,0.08916927,0.048014224,0.044584636,0.044584636,0.030866288,0.01371835,0.030866288,0.048014224,0.06516216,0.072021335,0.041155048,0.034295876,0.034295876,0.044584636,0.061732575,0.058302987,0.030866288,0.0274367,0.0548734,0.116605975,0.20920484,0.2777966,0.3018037,0.36010668,0.47671264,0.6276145,0.881404,1.1523414,1.3855534,1.587899,1.8382589,1.8039631,2.0577524,2.3629858,2.5721905,2.6167753,2.959734,3.4021509,3.5873485,3.3644254,2.8019729,3.0214665,2.8945718,2.7470996,2.6785078,2.568761,2.428148,2.6887965,3.4021509,4.280125,4.698535,3.957744,4.0880685,4.413879,4.479041,4.064061,4.6402316,4.2081037,3.0043187,1.7936742,1.8588364,1.5981878,1.2826657,1.0906088,1.2380811,1.9720128,2.7128036,3.5050385,4.955754,7.1952744,9.877212,10.477389,10.233889,10.14472,10.587136,11.30735,10.912948,10.494537,10.532263,11.201033,12.401388,13.581166,14.445422,15.155347,15.518884,15.011304,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.024007112,0.07888051,0.1371835,0.15433143,0.030866288,0.006859175,0.030866288,0.05144381,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.048014224,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.06516216,0.1371835,0.23664154,0.4081209,0.7888051,1.0082988,1.0288762,1.1489118,1.6256244,2.1263442,2.5070283,2.7642474,3.018037,3.5153272,4.791134,5.422178,5.2164025,5.1992545,5.5079174,5.353586,4.98662,4.6882463,4.770556,4.523626,4.6848164,4.5270553,4.122364,4.341858,5.593657,6.1801167,5.5662203,4.4516044,4.7774153,4.996909,4.9934793,5.528495,7.15069,10.182446,13.094165,12.603734,11.808069,12.428825,14.808959,13.865822,12.511135,11.204462,10.323058,10.127572,9.750318,8.309891,6.941485,6.4544835,7.31531,11.14273,13.612033,14.678635,14.644339,14.188204,9.5205345,6.0395036,4.0229063,3.1620796,2.5550427,1.786815,1.1763484,0.97057325,1.1351935,1.371835,0.9774324,0.7922347,0.9534253,1.3169615,1.4575747,0.85396725,0.6276145,0.52815646,0.39783216,0.16462019,0.18176813,0.20234565,0.26407823,0.31552204,0.20920484,0.16462019,0.20920484,0.25378948,0.28465575,0.35324752,0.32238123,0.32581082,0.20234565,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18519773,0.6790583,1.5364552,2.469303,3.3232703,4.0263357,4.5819287,5.079219,4.822,4.201245,3.6113555,3.0900583,2.3321195,1.3581166,0.7099246,0.432128,0.45270553,0.5727411,1.0185875,1.039165,0.8471081,0.5521636,0.15776102,0.12689474,0.058302987,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.0274367,0.06859175,0.12003556,0.12689474,0.0548734,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.020577524,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.017147938,0.030866288,0.020577524,0.024007112,0.037725464,0.06859175,0.15776102,0.2194936,0.22292319,0.2503599,0.34295875,0.48357183,0.58645946,0.67219913,0.8093826,1.0528834,1.4507155,1.5330256,1.7559488,2.1572106,2.5996273,2.7882545,2.668219,2.860276,3.450165,3.957744,3.3266997,3.6010668,3.1723683,2.6853669,2.4795918,2.6167753,2.702515,2.784825,3.059192,3.6113555,4.389872,3.9646032,3.9714622,3.9851806,3.8034124,3.433017,2.9940298,2.417859,1.9342873,1.6564908,1.5741806,1.0871792,0.89855194,0.89855194,1.0220171,1.2620882,1.7765263,2.0886188,2.9494452,4.746549,7.507367,9.647429,10.4705305,10.422516,10.086417,10.203023,10.30591,9.294182,8.080108,7.613684,8.89635,10.556271,11.38623,12.157887,13.375391,15.29253,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.12689474,0.22635277,0.20577525,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.23664154,0.2194936,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.15090185,0.2194936,0.31209245,0.490431,0.8093826,1.2723769,1.6907866,1.9720128,2.2841053,3.0660512,3.309552,3.5187566,3.8171308,4.297273,5.003768,6.0052075,6.8969,7.4044795,7.380472,6.8214493,6.077229,5.470192,5.0243454,4.695105,4.3795834,3.9508848,4.256118,5.305572,6.9963584,9.108984,8.450503,7.040943,6.0326443,6.142391,7.6445503,12.528283,15.789821,15.501736,12.902108,12.3911,13.697772,14.38026,13.934414,12.411677,10.422516,9.163857,7.6033955,6.4579134,6.1321025,6.728851,9.06097,11.842365,14.037301,15.909856,18.996485,14.078457,9.513676,6.1458206,4.214963,3.3712845,2.6990852,1.762808,1.0494537,0.7133542,0.5796003,0.70306545,0.9602845,1.7662375,2.7779658,2.8980014,1.2860953,0.9842916,0.83338976,0.4698535,0.33609957,0.274367,0.26064864,0.25378948,0.23321195,0.18176813,0.17147937,0.17833854,0.18176813,0.24350071,0.48700142,0.5727411,0.4389872,0.20920484,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29151493,1.4644338,2.2223728,2.942586,3.5221863,3.9783216,4.4550343,4.3933015,3.974892,3.3644254,2.527606,1.2209331,0.40126175,0.15433143,0.14061308,0.51100856,1.8931323,2.843128,2.7333813,2.3389788,1.7216529,0.24350071,0.08573969,0.037725464,0.024007112,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.034295876,0.044584636,0.041155048,0.030866288,0.006859175,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.030866288,0.030866288,0.037725464,0.048014224,0.061732575,0.12346515,0.18176813,0.23321195,0.24007112,0.16804978,0.13032432,0.2503599,0.47671264,0.70649505,0.77851635,1.1454822,1.2277923,1.2689474,1.3615463,1.4335675,1.5673214,1.9411465,2.4967396,3.117495,3.6319332,3.3884325,3.0523329,2.8259802,2.8019729,2.959734,2.8980014,2.5173173,2.1880767,2.352697,3.525616,4.5613513,4.4721823,3.7965534,3.0077481,2.5173173,2.469303,2.4384367,2.3149714,2.0886188,1.8313997,1.2449403,0.88826317,0.78537554,0.8471081,0.8848336,0.7133542,0.96371406,1.605047,2.5756202,3.782835,5.994919,7.8366075,8.97866,9.445084,9.626852,10.446524,10.220171,8.803751,7.2124224,7.613684,9.321619,10.583707,11.749766,13.365103,16.160215,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.13375391,0.06516216,0.041155048,0.030866288,0.020577524,0.0,0.048014224,0.1920569,0.4081209,0.52472687,0.2194936,0.082310095,0.044584636,0.044584636,0.041155048,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.048014224,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.06516216,0.11317638,0.18862732,0.31895164,0.5418748,0.77851635,1.0117283,1.2963841,1.786815,2.294394,2.7059445,3.018037,3.350707,3.9440255,4.73969,5.8337283,6.931196,7.764586,8.090397,7.939495,7.490219,6.869464,6.159539,5.3913116,4.787704,4.383013,4.7499785,6.15268,8.546532,9.918367,9.640571,7.9875093,6.258997,6.7528577,9.167287,10.851214,11.897239,12.648318,13.708061,14.349394,15.234227,15.676644,15.590904,15.488017,13.430264,10.840926,8.7317295,7.7577267,8.217292,10.031544,12.456262,14.856973,16.983316,18.948471,15.542891,11.372512,7.822889,5.7136927,5.302142,6.025785,4.9180284,3.2272418,1.7559488,0.86082643,0.8265306,1.1043272,1.4369972,1.6427724,1.6187652,1.8519772,1.8588364,1.5055889,0.94999576,0.6276145,0.53844523,0.48014224,0.5624523,0.64819205,0.36696586,0.26750782,0.6379033,0.9877212,1.0734608,0.9294182,0.85739684,0.66191036,0.40126175,0.15090185,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.29151493,0.51100856,0.6276145,0.939707,1.1008976,1.3512574,1.6873571,2.2155135,3.1483612,4.729401,5.144381,4.5784993,3.3952916,2.1469216,1.3889829,0.99801,0.9328478,1.2929544,2.318401,3.6627994,3.649081,3.0523329,2.2155135,1.0631721,0.4629943,0.15776102,0.034295876,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.0,0.01371835,0.020577524,0.020577524,0.020577524,0.017147938,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.017147938,0.0274367,0.06859175,0.106317215,0.13032432,0.13375391,0.12689474,0.14061308,0.16462019,0.18862732,0.20577525,0.15776102,0.1371835,0.16119061,0.24007112,0.36353627,0.67219913,0.97400284,1.2175035,1.3821237,1.4815818,1.5981878,1.8999915,2.2360911,2.5996273,3.1449318,2.860276,2.726522,2.6613598,2.5756202,2.3732746,2.2052248,2.1332035,1.903421,1.6084765,1.704505,1.8656956,1.762808,1.5638919,1.4129901,1.430138,1.5981878,1.5261664,1.8142518,2.2155135,1.6496316,1.0323058,0.72707254,0.8025235,1.1351935,1.3855534,0.91227025,1.0871792,1.5844694,2.0714707,2.1846473,3.340418,4.9694724,6.6293926,8.038953,9.091836,10.045261,10.477389,10.261326,9.671436,9.373062,9.764035,10.621432,11.753197,13.066729,14.572317,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.14747226,0.20234565,0.09602845,0.044584636,0.06859175,0.08573969,0.061732575,0.0,0.030866288,0.1097468,0.29151493,0.42526886,0.16462019,0.058302987,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.06859175,0.09259886,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.048014224,0.09602845,0.18176813,0.31552204,0.5212973,0.8025235,1.1351935,1.4610043,1.8519772,2.3595562,2.867135,3.0900583,3.6765177,4.5030484,5.593657,6.8283086,7.939495,8.549961,8.525954,8.117833,7.5862474,7.174697,6.9380555,6.341307,5.871454,5.8508763,6.447624,7.1849856,8.035523,7.64798,6.420188,6.5024977,7.082098,7.7680154,9.139851,11.252477,13.63604,13.773223,13.828096,13.865822,13.910407,13.917266,12.435684,11.228469,10.823778,10.796341,9.781183,10.206452,12.044711,14.623761,17.1205,18.578075,16.736387,13.7938,10.158438,7.040943,6.451054,8.381912,7.8674736,5.8645945,3.3644254,1.3992717,0.91569984,0.86082643,0.94999576,1.0494537,1.1763484,1.4129901,1.704505,1.7662375,1.4507155,0.7476501,0.607037,0.4629943,0.45613512,0.53158605,0.4664239,0.52815646,0.86082643,1.1351935,1.1043272,0.6344737,0.9877212,0.8128122,0.47671264,0.18862732,0.034295876,0.048014224,0.0548734,0.034295876,0.0034295875,0.010288762,0.0034295875,0.17490897,0.4081209,0.64133286,0.85396725,0.7922347,0.5590228,0.490431,0.75450927,1.3581166,2.417859,3.0626216,3.0969174,2.6236343,2.0406046,1.6256244,1.3958421,1.3992717,1.6633499,2.170929,2.6579304,2.5207467,2.085189,1.5227368,0.84367853,0.3806842,0.14747226,0.058302987,0.034295876,0.017147938,0.010288762,0.01371835,0.01371835,0.010288762,0.017147938,0.010288762,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0034295875,0.010288762,0.0,0.0034295875,0.006859175,0.010288762,0.01371835,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.006859175,0.024007112,0.06516216,0.11317638,0.15776102,0.17833854,0.18519773,0.18519773,0.16804978,0.14747226,0.14061308,0.12689474,0.11317638,0.106317215,0.11317638,0.13032432,0.2709374,0.5624523,0.90198153,1.2277923,1.5055889,1.5913286,1.8485477,2.3629858,3.0077481,3.433017,3.0146074,3.0077481,3.1037767,3.199805,3.391862,3.333559,3.2032347,2.9151495,2.5927682,2.568761,1.9754424,1.4850113,1.1626302,1.0151579,1.0220171,1.0288762,1.0220171,1.2346514,1.4678634,1.0631721,0.7613684,0.7373613,0.9911508,1.4267083,1.8485477,1.7765263,1.704505,1.7490896,1.8691251,1.8965619,2.0028791,3.0043187,4.4584637,6.029215,7.5210853,8.7145815,9.770895,10.401938,10.4705305,9.993818,9.856634,9.863494,10.065839,10.576848,11.55771,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.09259886,0.19548649,0.24007112,0.18862732,0.0274367,0.01371835,0.048014224,0.06859175,0.05144381,0.0,0.006859175,0.01371835,0.08916927,0.16462019,0.0548734,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.06859175,0.09259886,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.041155048,0.10288762,0.23321195,0.42869842,0.67219913,0.91227025,1.255229,1.7353712,2.1915064,2.2600982,2.5996273,3.069481,3.865145,5.0277753,6.4579134,7.8434668,8.56368,8.796892,8.7145815,8.505377,8.543102,8.001227,6.9071894,5.552502,4.496189,4.554492,5.761707,6.5162163,6.5127864,6.7185616,6.776865,7.099246,7.9429245,9.373062,11.266195,12.178465,12.3911,12.466551,12.4802685,12.017275,10.545981,9.983529,10.556271,11.427385,10.690024,9.990388,10.943813,13.29994,16.245956,18.420315,17.754974,15.649208,12.127021,8.47451,7.2158523,9.277034,9.6645775,8.193284,5.456474,2.8019729,1.6942163,1.3272504,1.1797781,1.0563129,1.0871792,1.0631721,1.3272504,1.5604624,1.5330256,1.1146159,0.7476501,0.48357183,0.39440256,0.4698535,0.6001778,0.75450927,1.0014396,1.3101025,1.3889829,0.6893471,1.0906088,0.96371406,0.6276145,0.3018037,0.11317638,0.07545093,0.061732575,0.041155048,0.020577524,0.05144381,0.030866288,0.037725464,0.15090185,0.3566771,0.53158605,0.4698535,0.29494452,0.15776102,0.15433143,0.33952916,0.58645946,0.96714365,1.2037852,1.2483698,1.2963841,1.1797781,1.08032,1.1214751,1.2826657,1.4267083,1.2826657,1.1214751,0.90884066,0.64476246,0.3566771,0.15776102,0.07888051,0.05144381,0.037725464,0.024007112,0.020577524,0.0274367,0.024007112,0.017147938,0.017147938,0.010288762,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.006859175,0.024007112,0.0548734,0.09945804,0.16119061,0.216064,0.2503599,0.2469303,0.20234565,0.1371835,0.08573969,0.08916927,0.09602845,0.10288762,0.09602845,0.058302987,0.08916927,0.32581082,0.6859175,1.0631721,1.3032433,1.4095604,1.6873571,2.4898806,3.5564823,4.0023284,3.3061223,3.2786856,3.5804894,4.0503426,4.722542,4.7979927,4.7499785,4.7328305,4.6676683,4.266407,2.8739944,2.0131679,1.5570327,1.3306799,1.1214751,0.85739684,0.8848336,1.0357354,1.1111864,0.86082643,0.77165717,0.939707,1.2243627,1.5330256,1.8382589,2.1400626,2.2909644,2.4898806,2.836269,3.3369887,2.201795,2.3046827,3.0900583,4.256118,5.7479887,7.3530354,8.992378,10.209882,10.755186,10.563129,10.124143,9.424506,8.995808,9.167287,10.093276,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.034295876,0.09945804,0.19548649,0.29494452,0.31895164,0.1920569,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.037725464,0.09945804,0.2469303,0.548734,0.84367853,1.0666018,1.2346514,1.4232788,1.6084765,1.8897027,2.3664153,3.1415021,4.3349986,6.3618846,7.7748747,8.745448,9.23245,9.012956,8.954653,8.495089,6.9826403,4.8288593,3.5187566,3.590778,4.2526884,5.144381,6.029215,6.8111606,7.5245147,7.9189177,8.052671,8.004657,7.8537555,9.860064,11.2421875,12.21962,12.672326,12.147599,10.254466,9.153569,9.177576,10.124143,11.2421875,10.408798,10.484249,12.13731,15.148488,18.392878,18.025911,16.101913,13.114742,10.000677,8.128122,9.263316,10.600855,10.031544,7.490219,4.9248877,3.333559,2.8122618,2.4075704,1.7971039,1.3032433,1.3478279,1.2415106,1.1592005,1.2243627,1.488441,0.91227025,0.5727411,0.48357183,0.58988905,0.7476501,0.7956643,1.0254467,1.5090185,1.8519772,1.1832076,1.1660597,1.097468,0.8676856,0.5418748,0.34981793,0.14061308,0.048014224,0.020577524,0.037725464,0.08573969,0.0548734,0.020577524,0.0,0.0034295875,0.0,0.010288762,0.23321195,0.31552204,0.22635277,0.25721905,0.33952916,0.2777966,0.16804978,0.15433143,0.41498008,0.41498008,0.34295875,0.34638834,0.432128,0.45270553,0.34295875,0.3018037,0.22978236,0.11317638,0.037725464,0.010288762,0.017147938,0.020577524,0.01371835,0.01371835,0.020577524,0.024007112,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.020577524,0.048014224,0.09602845,0.17490897,0.26750782,0.31209245,0.29494452,0.23321195,0.15090185,0.07545093,0.06516216,0.06859175,0.072021335,0.072021335,0.072021335,0.10288762,0.29494452,0.6001778,0.8676856,0.84024894,1.0082988,1.3169615,2.1812177,3.3644254,3.9611735,3.2443898,3.1277838,3.5290456,4.3109913,5.302142,5.4016004,5.5490727,5.9400454,6.186976,5.3330083,3.4776018,2.503599,2.0714707,1.8313997,1.3924125,0.9534253,0.9431366,1.155771,1.3169615,1.1008976,1.0631721,1.1694894,1.2929544,1.371835,1.4232788,1.8039631,2.5138876,3.4398763,4.4721823,5.4941993,3.799983,3.0900583,2.959734,3.3026927,4.3041325,6.0497923,7.8023114,9.153569,9.97667,10.408798,10.055551,9.421077,9.283894,9.952662,11.283342,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.0034295875,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.17147937,0.4629943,0.7922347,0.70649505,0.274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.06516216,0.17833854,0.29837412,0.44584638,0.70306545,1.0940384,1.4918705,1.8656956,2.2738166,2.884283,5.24041,6.495639,7.6274023,8.755736,9.170717,8.742019,8.241299,6.111525,3.3472774,3.4947495,3.117495,2.8465576,3.0969174,4.0777793,5.7994323,7.3598948,7.805741,8.2653055,8.477941,6.8043017,7.208993,8.783174,10.63858,12.096155,12.696333,12.181894,11.616013,11.345076,11.657167,12.754636,13.087306,12.96727,13.670336,15.498305,17.806417,16.317978,14.610043,12.912396,11.338216,9.873782,9.945804,12.21619,11.770344,8.453933,6.866034,5.4496145,4.8117113,4.2938433,3.4878905,2.2429502,2.2806756,1.6496316,1.1489118,1.0254467,0.9774324,0.7339317,0.52472687,0.45613512,0.5521636,0.7476501,0.5521636,0.70649505,1.0288762,1.2929544,1.2209331,1.0871792,1.1249046,1.0288762,0.8265306,0.89855194,0.38754338,0.12346515,0.017147938,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.037725464,0.18176813,0.7442205,0.58302987,0.26064864,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.12346515,0.24350071,0.36696586,0.39097297,0.33266997,0.24007112,0.15090185,0.07545093,0.06516216,0.061732575,0.061732575,0.061732575,0.061732575,0.1097468,0.20577525,0.33952916,0.4115505,0.22978236,0.4355576,0.64476246,0.96714365,1.4472859,2.0440342,2.411,2.3458378,2.3972816,2.9563043,4.2869844,4.2526884,4.1326528,4.2286816,4.5270553,4.6848164,3.6216443,2.9185789,2.4041407,1.9274281,1.3443983,0.9534253,0.881404,1.0117283,1.1626302,1.1146159,1.3101025,1.0666018,0.89512235,0.9842916,1.1900668,1.5433143,2.2360911,3.450165,4.9180284,5.919468,6.3001523,5.422178,4.280125,3.508468,3.3884325,4.0709205,4.65395,5.1855364,5.8817425,7.1266828,8.1384115,8.961512,10.124143,11.917816,14.359683,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25721905,0.33952916,0.29494452,0.22292319,0.28122616,0.6344737,0.8025235,0.5624523,0.09945804,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25378948,0.52472687,0.7373613,0.83681935,0.805953,0.58302987,0.24007112,0.058302987,0.061732575,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.041155048,0.09259886,0.18176813,0.36010668,0.7613684,1.3375391,1.862266,2.2841053,2.7368107,3.3541365,4.184097,5.422178,6.927767,8.241299,8.05953,7.6925645,6.5779486,4.979761,3.981751,3.3781435,3.0489032,2.8637056,2.8122618,2.9906003,4.90431,6.7700057,8.766026,10.535692,11.187314,10.446524,9.033533,9.15014,10.933525,12.452832,11.653738,11.516555,12.394529,14.164196,16.19794,16.431154,14.918706,14.033872,14.846684,17.12393,16.619781,15.391989,14.057879,12.7272,11.008976,9.997248,12.185325,12.452832,10.021255,8.453933,8.824328,8.961512,7.7611566,5.381023,3.2546785,2.8156912,2.369845,1.9823016,1.6496316,1.3169615,1.0837497,0.9431366,0.85739684,0.78537554,0.69963586,0.72707254,0.83338976,0.9877212,1.1832076,1.4404267,1.5501735,1.1317638,0.8779744,0.9431366,0.9362774,0.64819205,0.39440256,0.17833854,0.030866288,0.01371835,0.020577524,0.017147938,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.14747226,0.116605975,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.037725464,0.116605975,0.2194936,0.29151493,0.2777966,0.23321195,0.17147937,0.1097468,0.06516216,0.05144381,0.0548734,0.061732575,0.061732575,0.061732575,0.072021335,0.12003556,0.18519773,0.22978236,0.20577525,0.274367,0.44927597,0.77851635,1.2346514,1.7147937,2.4247184,3.2066643,3.7691166,3.957744,3.7759757,4.6265135,5.4770513,6.3310184,7.1061053,7.6274023,6.81802,6.060081,5.1512403,4.1120753,3.1723683,2.294394,1.6633499,1.3409687,1.3101025,1.4541451,1.0837497,0.9842916,1.0048691,1.1180456,1.4335675,2.6373527,4.715683,7.2467184,9.06097,8.213862,8.134981,6.4716315,4.856296,3.865145,3.0214665,3.5393343,4.4104495,5.1409516,5.662249,6.3207297,7.6959944,9.571979,11.674315,13.505715,14.345964,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12689474,0.16804978,0.14747226,0.1097468,0.14061308,0.31552204,0.40126175,0.28122616,0.05144381,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.59674823,0.9362774,0.9842916,0.7956643,0.50757897,0.28122616,0.10288762,0.030866288,0.030866288,0.006859175,0.044584636,0.0548734,0.044584636,0.0274367,0.0274367,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.08916927,0.061732575,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.06516216,0.16462019,0.41498008,0.86082643,1.3375391,1.8142518,2.3904223,2.7642474,3.309552,4.0537724,4.880303,5.5490727,5.9743414,6.252138,6.307011,6.036074,5.295283,4.245829,3.7142432,3.3678548,3.1277838,3.1689389,3.9165888,5.171818,6.708273,8.292743,9.702303,10.676306,9.630281,9.266746,10.288762,11.4205265,10.100135,9.033533,9.362774,11.266195,13.982429,14.791811,13.903547,13.289652,13.934414,15.844694,16.503176,15.844694,14.870691,13.680624,11.465111,10.05898,11.46854,12.476839,11.914387,10.652299,10.220171,9.836057,8.443645,6.276145,4.8905916,4.57164,4.197815,3.6627994,2.860276,1.6873571,1.3169615,1.0871792,0.9568549,0.8745448,0.7956643,0.881404,0.9877212,0.9877212,0.9534253,1.1489118,1.2963841,1.0357354,0.8676856,0.89512235,0.8265306,0.6893471,0.47328308,0.26407823,0.12346515,0.09602845,0.09602845,0.058302987,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.010288762,0.024007112,0.034295876,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.006859175,0.034295876,0.08573969,0.14061308,0.17490897,0.16462019,0.1371835,0.10288762,0.07545093,0.05144381,0.048014224,0.048014224,0.06516216,0.08916927,0.09602845,0.106317215,0.12689474,0.16119061,0.20577525,0.26407823,0.29151493,0.36010668,0.5144381,0.7613684,1.0666018,1.5364552,2.2052248,2.7402403,3.0214665,3.1346428,3.9371665,4.870014,5.960623,7.140401,8.241299,8.940934,8.035523,6.5230756,5.0106273,3.7142432,2.6407824,1.8931323,1.4438564,1.255229,1.2655178,0.90884066,0.71678376,0.64476246,0.7407909,1.1489118,2.7470996,4.763697,6.560801,7.421627,6.5539417,7.8674736,8.522525,7.4627824,5.1752477,3.6799474,3.210094,3.3644254,3.9303071,4.73969,5.662249,6.9860697,8.920357,11.122152,13.107883,14.243076,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.0548734,0.048014224,0.06859175,0.1371835,0.26750782,0.64133286,0.91569984,0.9259886,0.66876954,0.29837412,0.08573969,0.030866288,0.07545093,0.16119061,0.21263443,0.16119061,0.09945804,0.058302987,0.044584636,0.044584636,0.06859175,0.044584636,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.030866288,0.12346515,0.23321195,0.12689474,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.030866288,0.037725464,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.06859175,0.17833854,0.4389872,0.78194594,1.214074,1.8142518,2.335549,2.7882545,3.199805,3.4776018,3.4295874,3.8377085,4.3521466,4.99005,5.521636,5.4667625,4.3658648,3.7622573,3.6079261,3.74168,3.9063,3.5633414,3.673088,4.1292233,4.9420357,6.228131,8.48137,8.522525,8.289313,8.635701,9.321619,8.423067,7.0546613,6.667118,7.723431,9.705732,10.878652,11.262765,11.7086115,12.682614,14.2533655,15.556609,15.306249,14.651197,13.735497,11.71547,10.329918,10.967821,12.562579,13.821238,13.248496,11.581717,10.086417,8.501947,7.1095347,6.7357097,6.7185616,6.2212715,5.188966,3.7691166,2.2978237,1.605047,1.1454822,0.9362774,0.90541106,0.90541106,1.0254467,1.1043272,1.0940384,1.0425946,1.08032,1.2209331,1.2689474,1.2312219,1.1283343,1.0117283,2.085189,2.1332035,1.6804979,1.0494537,0.39783216,0.26407823,0.116605975,0.0274367,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.006859175,0.020577524,0.030866288,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.020577524,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.017147938,0.034295876,0.058302987,0.07545093,0.08916927,0.08916927,0.07888051,0.06516216,0.061732575,0.058302987,0.058302987,0.058302987,0.07888051,0.12003556,0.14061308,0.15090185,0.16119061,0.18176813,0.23664154,0.34295875,0.42526886,0.44927597,0.4664239,0.52815646,0.6790583,0.8779744,1.1763484,1.5055889,1.9411465,2.7059445,3.5393343,4.214963,4.9831905,6.018926,7.4181976,8.755736,8.464222,7.517656,6.375603,4.9694724,3.6044965,2.9974594,2.702515,2.4761622,2.2669573,2.1572106,1.704505,1.3375391,1.3375391,1.8416885,3.2409601,4.3178506,4.773986,4.5853586,3.998899,5.48734,7.6033955,7.9257765,6.1766872,4.2423997,3.192946,2.6785078,2.7813954,3.4604537,4.57507,5.874883,7.623973,9.585697,11.417097,12.655178,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.116605975,0.12689474,0.13375391,0.21263443,0.40126175,0.6824879,0.58302987,0.7339317,0.7888051,0.61389613,0.28808534,0.06859175,0.048014224,0.22635277,0.4664239,0.5144381,0.31209245,0.14747226,0.058302987,0.037725464,0.041155048,0.06516216,0.058302987,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.041155048,0.15776102,0.28465575,0.12689474,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.034295876,0.072021335,0.09602845,0.06859175,0.034295876,0.01371835,0.0034295875,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.07888051,0.216064,0.42183927,0.7305021,1.2072148,1.7833855,2.16064,2.49331,2.719663,2.5824795,2.4075704,2.5619018,3.0111778,3.57363,3.9165888,3.3747141,3.0248961,3.2066643,3.7039545,3.7725463,3.1860867,2.6716487,2.510458,2.836269,3.649081,5.4907694,5.861165,5.768566,5.9331865,6.7871537,7.366754,6.9826403,6.427047,6.135532,6.1766872,7.0306544,8.292743,9.836057,11.4376745,12.785502,13.996146,13.934414,13.471419,12.854094,11.701753,10.744898,11.005547,12.8197975,15.155347,15.62863,13.680624,11.293632,9.253027,8.069819,7.997798,8.128122,7.548522,6.094377,4.2183924,3.0043187,2.0714707,1.4850113,1.2106444,1.1317638,1.039165,1.1900668,1.2175035,1.2792361,1.3855534,1.371835,1.5741806,1.7319417,1.762808,1.7250825,1.8073926,4.3761535,4.979761,4.3590055,3.0146074,1.2072148,0.607037,0.22978236,0.061732575,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.034295876,0.034295876,0.020577524,0.006859175,0.0,0.0034295875,0.0034295875,0.024007112,0.037725464,0.044584636,0.05144381,0.06859175,0.072021335,0.072021335,0.072021335,0.07545093,0.08916927,0.08573969,0.08573969,0.10288762,0.1371835,0.17833854,0.18862732,0.18862732,0.19891608,0.2503599,0.37725464,0.548734,0.6173257,0.61389613,0.59674823,0.65848076,0.7579388,0.8265306,0.9774324,1.3992717,2.3389788,3.3987212,3.9783216,4.650521,5.5387836,6.3138704,6.9826403,7.905199,8.525954,8.3922,7.15069,5.23698,4.8014226,4.8185706,4.7191124,4.389872,4.461893,3.899441,3.3609958,3.2889743,3.9028704,4.7191124,4.664239,4.0263357,3.1380725,2.3664153,2.486451,4.0503426,5.641671,6.101236,4.537344,3.6353626,2.9117198,2.5207467,2.5961976,3.2375305,4.7671266,6.40304,8.179566,9.770895,10.491108,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.09259886,0.10288762,0.18862732,0.39097297,0.6344737,0.7339317,1.2072148,1.2449403,1.0082988,0.64133286,0.274367,0.0548734,0.037725464,0.36010668,0.7339317,0.4424168,0.39440256,0.29151493,0.1371835,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.01371835,0.048014224,0.12346515,0.2194936,0.15090185,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.09945804,0.22978236,0.48700142,0.9774324,1.6496316,1.5673214,1.5193073,1.762808,2.0440342,1.862266,1.5947582,1.4507155,1.4507155,1.4507155,1.9137098,2.2498093,2.3904223,2.369845,2.318401,2.318401,2.311542,2.74367,3.4913201,3.8445675,4.3590055,4.0023284,3.4878905,3.6387923,5.3707337,7.48336,8.735159,8.453933,6.9346256,5.4324665,5.212973,6.2658563,8.488229,10.981539,12.055,12.6757555,12.703192,12.199042,11.4205265,10.834066,10.981539,11.290202,12.744347,15.079896,16.80155,16.091625,13.965281,11.149589,8.608265,7.5210853,7.3873315,7.298162,6.420188,4.7842746,3.2958336,2.7951138,2.651071,2.4247184,1.9514352,1.3443983,1.4267083,1.4575747,1.4335675,1.4198492,1.5398848,1.9823016,1.8142518,1.845118,2.417859,3.4192986,5.079219,6.4373355,6.7528577,5.627953,2.9906003,1.2449403,0.48700142,0.20920484,0.09259886,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.044584636,0.044584636,0.020577524,0.006859175,0.006859175,0.01371835,0.01371835,0.01371835,0.024007112,0.041155048,0.06859175,0.09259886,0.116605975,0.11317638,0.11317638,0.12346515,0.1371835,0.12346515,0.12346515,0.12689474,0.15433143,0.22978236,0.22978236,0.20920484,0.1920569,0.20920484,0.30523327,0.47671264,0.61046654,0.6344737,0.58645946,0.61046654,0.67219913,0.7133542,0.7922347,0.9842916,1.371835,2.0920484,3.1792276,5.5902276,7.9120584,6.3618846,6.2898636,7.857185,9.321619,9.678296,8.652849,6.025785,5.545643,5.8200097,6.001778,5.7822843,5.6965446,5.7754254,5.7754254,5.857735,6.5779486,6.992929,6.464772,5.2301207,3.6593697,2.2429502,1.8656956,2.49331,3.5873485,4.671098,5.3570156,4.756838,4.012617,3.57363,3.3232703,2.5790498,4.616225,6.0806584,7.9943686,10.124143,10.9541025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.16804978,0.31895164,0.21263443,0.09945804,0.10288762,0.19891608,0.42526886,0.85396725,1.0082988,1.0528834,1.1420527,1.2037852,0.9328478,0.18519773,0.006859175,0.072021335,0.14747226,0.08916927,0.116605975,0.29837412,0.6173257,0.980862,1.2003556,0.37725464,0.06859175,0.0,0.0,0.0,0.0,0.0,0.0,0.08916927,0.4389872,3.1037767,1.5090185,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.006859175,0.024007112,0.048014224,0.116605975,0.10288762,0.06516216,0.034295876,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.037725464,0.106317215,0.24007112,0.47671264,0.8676856,0.9328478,0.7888051,0.7613684,1.0254467,1.6290541,1.8965619,1.4267083,1.0768905,1.0871792,1.0940384,1.2380811,1.762808,2.3321195,2.633923,2.3801336,1.9891608,2.1469216,2.2635276,2.2566686,2.551613,3.4535947,3.82399,3.234101,2.3972816,3.1723683,4.2698364,5.809721,7.0752387,7.689135,7.5931067,6.893471,6.1732574,6.869464,8.769455,9.990388,11.30735,11.948683,11.749766,10.991828,10.405369,10.357354,10.840926,12.116733,14.020154,15.944152,16.839275,16.348843,13.4474125,9.448513,8.011517,7.5245147,7.5382333,7.4765005,6.9380555,5.7136927,4.2355404,3.841138,3.3129816,2.4041407,1.8416885,1.8416885,1.8039631,1.7182233,1.6016173,1.529596,1.6667795,1.6359133,1.7936742,2.318401,3.210094,4.314421,5.0414934,5.1580997,4.5167665,3.0523329,1.7662375,0.91912943,0.41840968,0.16119061,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.0274367,0.037725464,0.037725464,0.037725464,0.030866288,0.024007112,0.034295876,0.058302987,0.07545093,0.07545093,0.058302987,0.041155048,0.030866288,0.044584636,0.072021335,0.106317215,0.14061308,0.18519773,0.23664154,0.28465575,0.32238123,0.34638834,0.28465575,0.22292319,0.21263443,0.274367,0.42526886,0.5007198,0.36353627,0.22292319,0.17490897,0.19548649,0.2503599,0.31895164,0.37725464,0.4355576,0.53844523,0.6379033,0.6310441,0.5693115,0.52472687,0.59331864,0.84367853,1.2723769,2.2841053,3.4673128,3.566771,4.413879,5.936616,7.2021337,7.4181976,5.9434752,5.0277753,4.7431192,4.8494368,5.144381,5.4907694,5.6793966,5.2918534,4.8014226,4.5339146,4.6608095,4.479041,3.7382503,2.6887965,1.6873571,1.1797781,1.3478279,1.6016173,2.0886188,2.8294096,3.707384,4.1463714,4.530485,4.773986,4.715683,4.1155047,4.5819287,5.2266912,6.464772,8.186425,9.746887,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.010288762,0.006859175,0.0034295875,0.0034295875,0.006859175,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.044584636,0.044584636,0.034295876,0.017147938,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.01371835,0.017147938,0.01371835,0.01371835,0.024007112,0.0034295875,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.06516216,0.09945804,0.08573969,0.07545093,0.18519773,0.34638834,0.30866286,0.2503599,0.23664154,0.2777966,0.42526886,0.78537554,0.90884066,0.9328478,0.9602845,0.939707,0.6859175,0.1371835,0.0,0.0034295875,0.058302987,0.25721905,0.216064,0.216064,0.33266997,0.5453044,0.71678376,0.2777966,0.23664154,0.2194936,0.09602845,0.0,0.0,0.0,0.0,0.12689474,0.6310441,2.1400626,1.2037852,0.19891608,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0034295875,0.006859175,0.0,0.006859175,0.01371835,0.037725464,0.072021335,0.07545093,0.12346515,0.12003556,0.106317215,0.12346515,0.216064,0.42526886,0.4424168,0.31895164,0.15776102,0.1371835,0.17490897,0.15776102,0.22292319,0.41498008,0.70306545,0.5590228,0.4081209,0.36353627,0.5007198,0.8471081,1.0666018,0.89512235,0.7579388,0.78537554,0.83338976,0.9877212,1.2998136,1.5810398,1.8759843,2.4795918,2.6647894,2.7059445,2.4624438,2.1057668,2.1469216,2.6853669,2.9117198,2.4075704,1.5981878,1.7559488,2.4144297,3.5942078,4.880303,5.892031,6.310441,6.138962,5.675967,5.9400454,7.058091,8.285883,9.928656,11.118723,11.355364,10.768905,10.117283,9.602845,10.0041065,11.231899,13.090735,15.302819,17.364002,17.559488,15.354263,11.852654,9.798331,8.786603,8.447074,8.467651,8.323608,7.298162,5.8234396,4.962613,4.0846386,3.083199,2.3801336,2.4452958,2.2806756,2.07833,1.9102802,1.7353712,1.6221949,1.5021594,1.4918705,1.8005334,2.7093742,3.6010668,3.9714622,4.15666,4.139512,3.5530527,1.8759843,0.9328478,0.432128,0.17490897,0.048014224,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.024007112,0.037725464,0.044584636,0.061732575,0.06516216,0.048014224,0.041155048,0.0548734,0.072021335,0.07888051,0.07545093,0.072021335,0.08916927,0.11317638,0.15433143,0.216064,0.28122616,0.32924038,0.41840968,0.5007198,0.548734,0.5521636,0.4938606,0.41840968,0.3841138,0.42869842,0.5555932,0.6310441,0.4972902,0.34295875,0.26064864,0.23321195,0.2194936,0.2469303,0.31209245,0.41498008,0.53844523,0.6241849,0.6241849,0.5624523,0.48700142,0.45270553,0.47671264,0.5624523,0.82996017,1.2620882,1.7250825,2.4967396,3.6079261,4.5922174,4.9694724,4.2389703,3.7862647,3.5702004,3.5187566,3.6696587,4.180667,4.6265135,4.588788,4.383013,4.249259,4.3624353,4.173808,3.4295874,2.417859,1.5055889,1.1351935,1.2415106,1.2586586,1.3821237,1.7559488,2.4727325,3.2032347,3.8617156,4.290414,4.4275975,4.290414,4.3624353,4.928317,5.8337283,6.931196,8.090397,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.01371835,0.006859175,0.006859175,0.006859175,0.0,0.0,0.010288762,0.020577524,0.024007112,0.006859175,0.0,0.0034295875,0.006859175,0.006859175,0.01371835,0.030866288,0.0274367,0.024007112,0.024007112,0.017147938,0.030866288,0.017147938,0.0034295875,0.0,0.006859175,0.0,0.0034295875,0.017147938,0.037725464,0.058302987,0.058302987,0.048014224,0.0274367,0.006859175,0.006859175,0.006859175,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.017147938,0.020577524,0.017147938,0.024007112,0.01371835,0.020577524,0.030866288,0.037725464,0.024007112,0.020577524,0.010288762,0.0034295875,0.0,0.006859175,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.0034295875,0.0,0.0034295875,0.006859175,0.01371835,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.006859175,0.017147938,0.01371835,0.006859175,0.006859175,0.01371835,0.017147938,0.017147938,0.017147938,0.017147938,0.017147938,0.01371835,0.01371835,0.010288762,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.07888051,0.072021335,0.061732575,0.07888051,0.12003556,0.12346515,0.09259886,0.116605975,0.19548649,0.22292319,0.22292319,0.22292319,0.28122616,0.45613512,0.8196714,0.8471081,0.88826317,0.8093826,0.5727411,0.2469303,0.0548734,0.0034295875,0.034295876,0.20577525,0.6962063,0.52472687,0.23321195,0.0548734,0.05144381,0.12003556,0.08916927,0.20234565,0.2194936,0.09602845,0.0,0.0,0.0,0.0,0.082310095,0.4115505,0.58645946,0.44927597,0.19891608,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.006859175,0.017147938,0.024007112,0.017147938,0.020577524,0.0274367,0.07888051,0.20234565,0.3806842,0.4424168,0.4389872,0.45956472,0.5212973,0.5658819,0.8128122,0.8711152,0.7613684,0.58302987,0.5144381,0.48357183,0.39783216,0.33609957,0.35324752,0.48357183,0.4115505,0.39097297,0.45270553,0.5761707,0.70306545,0.58302987,0.5178677,0.52472687,0.58645946,0.66876954,0.7990939,0.91569984,0.9362774,1.0700313,1.8005334,2.4487255,2.6647894,2.6613598,2.651071,2.8396983,2.983741,2.8259802,2.3252604,1.6839274,1.3272504,1.5604624,2.2806756,3.0866287,3.7725463,4.314421,4.65395,4.9420357,5.377593,6.042933,6.90033,8.388771,9.757176,10.288762,9.928656,9.287323,8.457363,8.515666,9.56512,11.47197,13.831526,16.331696,16.743246,15.481158,13.37882,11.698323,10.31277,9.366203,8.886061,8.604835,7.936065,6.9620624,5.953764,4.897451,3.9303071,3.350707,3.2443898,2.836269,2.417859,2.1263442,1.9685832,1.7765263,1.6256244,1.4198492,1.4267083,2.2635276,3.0043187,3.3987212,3.8720043,4.2698364,3.865145,1.9068506,0.91227025,0.4389872,0.21263443,0.10288762,0.048014224,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.010288762,0.020577524,0.030866288,0.037725464,0.048014224,0.048014224,0.06516216,0.07888051,0.07888051,0.058302987,0.048014224,0.058302987,0.07545093,0.09602845,0.12689474,0.15433143,0.21263443,0.3018037,0.4115505,0.5007198,0.5727411,0.6859175,0.7579388,0.7510797,0.6859175,0.607037,0.53158605,0.48700142,0.48700142,0.53844523,0.59331864,0.51100856,0.39440256,0.29837412,0.24350071,0.22292319,0.2469303,0.31209245,0.41498008,0.53158605,0.58988905,0.6001778,0.5761707,0.5418748,0.50757897,0.45270553,0.42869842,0.4389872,0.52472687,0.764798,1.1694894,1.7662375,2.386993,2.8122618,2.7813954,2.503599,2.5001693,2.760818,3.1072063,3.1689389,3.4535947,3.6970954,3.8308492,3.9268777,4.187526,4.3692946,4.0057583,3.2272418,2.393852,2.0989075,2.0063086,1.8108221,1.7010754,1.8039631,2.177788,2.5447538,3.199805,3.724532,4.0091877,4.2423997,4.32471,4.8082814,5.442755,6.125243,6.90033,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.0274367,0.034295876,0.048014224,0.034295876,0.024007112,0.020577524,0.01371835,0.006859175,0.010288762,0.024007112,0.034295876,0.01371835,0.010288762,0.01371835,0.017147938,0.020577524,0.020577524,0.0548734,0.061732575,0.058302987,0.0548734,0.048014224,0.058302987,0.041155048,0.024007112,0.017147938,0.017147938,0.006859175,0.010288762,0.024007112,0.037725464,0.037725464,0.030866288,0.030866288,0.030866288,0.0274367,0.024007112,0.020577524,0.006859175,0.0,0.0,0.0034295875,0.0034295875,0.010288762,0.017147938,0.017147938,0.017147938,0.030866288,0.041155048,0.0548734,0.06516216,0.06516216,0.048014224,0.0274367,0.010288762,0.0034295875,0.01371835,0.0034295875,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0034295875,0.006859175,0.017147938,0.0274367,0.020577524,0.020577524,0.020577524,0.01371835,0.01371835,0.020577524,0.024007112,0.020577524,0.01371835,0.024007112,0.030866288,0.024007112,0.020577524,0.024007112,0.0274367,0.041155048,0.048014224,0.0548734,0.061732575,0.061732575,0.048014224,0.037725464,0.0274367,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.041155048,0.07545093,0.08573969,0.16804978,0.13375391,0.06859175,0.0274367,0.044584636,0.106317215,0.106317215,0.072021335,0.034295876,0.030866288,0.024007112,0.037725464,0.13032432,0.36010668,0.78194594,0.69963586,0.7922347,0.7133542,0.39097297,0.017147938,0.01371835,0.006859175,0.11317638,0.5212973,1.4815818,1.1111864,0.4698535,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.01371835,0.030866288,0.041155048,0.041155048,0.030866288,0.037725464,0.116605975,0.32924038,0.7305021,0.82996017,0.8196714,0.8779744,0.97400284,0.8711152,0.91569984,0.9842916,1.0117283,0.96714365,0.864256,0.7133542,0.64476246,0.5212973,0.36696586,0.34981793,0.42526886,0.5624523,0.7510797,0.9328478,0.9842916,0.6207553,0.42869842,0.40126175,0.4698535,0.52472687,0.5727411,0.71678376,0.7956643,0.78537554,0.77165717,1.2929544,1.8348293,2.486451,3.1826572,3.6970954,3.8548563,3.542764,3.0489032,2.5138876,1.9137098,1.6221949,1.9720128,2.287535,2.452155,2.9151495,3.4467354,4.262977,5.1512403,5.844017,6.0497923,7.040943,8.080108,8.611694,8.491658,8.018375,7.06495,6.697984,7.4970784,9.403929,11.729189,14.054449,14.613472,14.109323,13.293081,12.96727,11.646879,10.172156,8.999237,8.31332,8.042382,7.5759587,6.783724,5.7754254,4.870014,4.5853586,4.0846386,3.3678548,2.6647894,2.1812177,2.095478,2.0440342,2.0165975,1.7730967,1.5604624,2.1091962,2.5961976,3.059192,3.765687,4.3109913,3.5804894,1.879414,0.9294182,0.47328308,0.29151493,0.20920484,0.11317638,0.061732575,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.006859175,0.030866288,0.041155048,0.0548734,0.06859175,0.082310095,0.06859175,0.06859175,0.07888051,0.09259886,0.08916927,0.07545093,0.08916927,0.116605975,0.15776102,0.2194936,0.2469303,0.33952916,0.48357183,0.64133286,0.764798,0.8848336,1.0014396,1.0151579,0.90541106,0.7476501,0.6241849,0.5453044,0.5007198,0.47671264,0.4389872,0.4629943,0.42526886,0.34981793,0.2709374,0.23321195,0.22978236,0.26407823,0.31209245,0.37382504,0.4698535,0.52815646,0.5521636,0.5624523,0.5658819,0.53844523,0.4629943,0.4355576,0.45956472,0.490431,0.4698535,0.58302987,0.77851635,1.0323058,1.2792361,1.4232788,1.4095604,1.6770682,2.393852,3.069481,2.5447538,2.411,2.5927682,2.8499873,3.1312134,3.5461934,4.2081037,4.383013,4.07435,3.6285036,3.7313912,3.7142432,3.3850029,3.07634,2.9117198,2.836269,2.5550427,3.0454736,3.6353626,4.064061,4.4721823,4.5613513,4.756838,5.0826488,5.5902276,6.3824625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.024007112,0.041155048,0.06859175,0.106317215,0.13032432,0.09259886,0.07888051,0.09602845,0.061732575,0.037725464,0.01371835,0.006859175,0.01371835,0.01371835,0.041155048,0.037725464,0.030866288,0.034295876,0.044584636,0.06859175,0.06859175,0.0548734,0.048014224,0.061732575,0.061732575,0.07888051,0.09259886,0.07888051,0.030866288,0.017147938,0.01371835,0.034295876,0.061732575,0.061732575,0.037725464,0.041155048,0.058302987,0.072021335,0.061732575,0.037725464,0.01371835,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.020577524,0.030866288,0.030866288,0.041155048,0.0548734,0.048014224,0.041155048,0.07545093,0.05144381,0.0274367,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.010288762,0.01371835,0.01371835,0.01371835,0.0274367,0.048014224,0.06859175,0.07545093,0.07545093,0.05144381,0.06516216,0.06859175,0.061732575,0.061732575,0.048014224,0.037725464,0.037725464,0.041155048,0.01371835,0.041155048,0.06516216,0.09602845,0.12346515,0.12346515,0.09602845,0.072021335,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06516216,0.18519773,0.28122616,0.18176813,0.061732575,0.01371835,0.0,0.010288762,0.044584636,0.15433143,0.20920484,0.18519773,0.10288762,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.26750782,0.39097297,0.37382504,0.2503599,0.09259886,0.017147938,0.010288762,0.2777966,1.1420527,3.0214665,2.277246,0.96371406,0.12689474,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.01371835,0.0274367,0.06859175,0.14747226,0.2777966,0.47328308,0.58302987,0.58302987,0.6310441,0.7510797,0.823101,0.6893471,0.6207553,0.61389613,0.6207553,0.53501564,0.31552204,0.39783216,0.5178677,0.5693115,0.59674823,0.58302987,0.5693115,0.58988905,0.5590228,0.29151493,0.31552204,0.37382504,0.4046913,0.36696586,0.24350071,0.48700142,0.8711152,1.1249046,1.1626302,1.0528834,0.96714365,1.1763484,1.8691251,2.6750782,2.6236343,3.357566,3.4673128,3.3987212,3.3644254,3.340418,2.767677,2.6887965,2.4315774,1.9857311,1.9994495,2.8054025,4.0846386,5.5079174,6.4887795,6.193835,6.756287,6.9792104,7.160979,7.3221693,7.1884155,5.9434752,5.501058,6.2967224,8.176137,10.422516,12.483699,13.440554,13.183334,12.55229,13.320518,12.723769,11.283342,9.836057,8.872343,8.529384,8.114404,7.442205,6.601956,5.7925735,5.3398676,4.6436615,3.7211025,2.7916842,2.1332035,2.061182,2.3389788,2.4761622,2.452155,2.352697,2.3664153,2.4624438,2.2395205,2.6373527,3.2855449,2.5173173,1.4815818,0.77165717,0.41840968,0.34638834,0.3806842,0.23664154,0.14404267,0.082310095,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.0548734,0.05144381,0.06516216,0.09602845,0.106317215,0.13032432,0.12689474,0.1097468,0.09945804,0.1371835,0.17490897,0.18176813,0.22635277,0.30523327,0.36696586,0.45270553,0.51100856,0.61389613,0.7888051,1.0220171,1.1694894,1.2415106,1.1866373,1.0151579,0.8093826,0.6756287,0.58645946,0.5693115,0.5727411,0.48700142,0.40126175,0.35324752,0.32238123,0.31895164,0.36696586,0.35324752,0.34295875,0.31209245,0.28808534,0.33609957,0.48357183,0.5555932,0.6173257,0.65162164,0.5658819,0.41840968,0.35324752,0.36696586,0.42183927,0.45613512,0.44584638,0.4698535,0.5144381,0.5693115,0.64133286,0.77508676,0.90884066,1.1043272,1.2758065,1.1900668,1.1043272,1.2037852,1.5261664,2.0680413,2.7779658,3.6936657,3.9303071,4.046913,4.4413157,5.3570156,6.0497923,5.885172,5.305572,4.605936,3.9200184,3.40901,3.1792276,3.5221863,4.2766957,4.835718,4.897451,4.9420357,4.972902,5.195825,6.025785,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.0034295875,0.0,0.01371835,0.024007112,0.024007112,0.024007112,0.048014224,0.044584636,0.0274367,0.01371835,0.01371835,0.0034295875,0.010288762,0.01371835,0.017147938,0.0274367,0.0274367,0.020577524,0.020577524,0.034295876,0.06859175,0.07545093,0.082310095,0.08916927,0.08916927,0.072021335,0.058302987,0.030866288,0.017147938,0.030866288,0.041155048,0.06516216,0.061732575,0.05144381,0.044584636,0.058302987,0.09259886,0.12003556,0.12346515,0.11317638,0.13375391,0.106317215,0.07888051,0.06859175,0.06516216,0.0548734,0.024007112,0.024007112,0.030866288,0.048014224,0.09602845,0.10288762,0.082310095,0.05144381,0.030866288,0.037725464,0.041155048,0.024007112,0.006859175,0.006859175,0.0274367,0.048014224,0.05144381,0.05144381,0.05144381,0.030866288,0.05144381,0.06859175,0.07888051,0.08916927,0.07545093,0.12003556,0.09259886,0.041155048,0.0034295875,0.0,0.0,0.006859175,0.006859175,0.0,0.0034295875,0.010288762,0.01371835,0.020577524,0.030866288,0.05144381,0.15090185,0.19548649,0.22292319,0.2469303,0.2469303,0.22292319,0.23664154,0.20577525,0.1371835,0.09602845,0.12346515,0.15090185,0.15090185,0.116605975,0.06516216,0.058302987,0.061732575,0.06859175,0.072021335,0.072021335,0.06859175,0.06516216,0.05144381,0.037725464,0.024007112,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.048014224,0.08573969,0.037725464,0.26064864,0.4972902,0.58302987,0.42869842,0.037725464,0.01371835,0.0034295875,0.0,0.0034295875,0.010288762,0.05144381,0.16804978,0.20234565,0.12689474,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.44584638,0.4046913,0.21263443,0.058302987,0.017147938,0.034295876,0.15433143,0.3841138,0.7099246,1.1043272,0.7888051,0.34638834,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.006859175,0.017147938,0.0274367,0.041155048,0.14404267,0.23321195,0.29494452,0.4115505,0.764798,1.0597426,1.3924125,1.6736387,1.6290541,1.1729189,0.6927767,0.37382504,0.2503599,0.20577525,0.17147937,0.31209245,0.4698535,0.5521636,0.5590228,0.50757897,0.4938606,0.41840968,0.26750782,0.106317215,0.17147937,0.25721905,0.2777966,0.216064,0.12346515,0.25721905,0.45270553,0.6344737,0.8093826,1.039165,1.3649758,1.529596,1.9308578,2.4418662,2.393852,2.3629858,2.2978237,2.3218307,2.435007,2.5001693,2.8225505,3.0557625,2.860276,2.2738166,1.7319417,2.2052248,2.976882,4.57164,6.632822,7.939495,8.872343,9.205012,8.971801,8.289313,7.332458,6.3824625,5.802862,5.813151,6.6053853,8.333898,10.991828,12.579727,12.891819,12.620882,13.368532,13.612033,13.025573,11.880091,10.5597,9.554831,8.738589,7.857185,7.1198235,6.64997,6.4990683,6.1766872,5.103226,3.9200184,3.0626216,2.7573884,2.6167753,2.551613,2.6956558,3.2135234,4.2698364,3.2135234,3.2683969,3.8891523,4.386442,3.9200184,2.386993,1.0768905,0.41498008,0.34638834,0.34638834,0.2777966,0.2194936,0.15433143,0.07888051,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0,0.010288762,0.0034295875,0.0034295875,0.017147938,0.030866288,0.06516216,0.08573969,0.07888051,0.058302987,0.06859175,0.15433143,0.15776102,0.13375391,0.13032432,0.18519773,0.22292319,0.19548649,0.19548649,0.2503599,0.32924038,0.39440256,0.50757897,0.6310441,0.77508676,0.99801,1.1729189,1.313532,1.3375391,1.2277923,1.039165,0.8779744,0.6859175,0.5418748,0.48357183,0.52472687,0.4972902,0.4424168,0.37382504,0.34638834,0.4629943,0.64819205,0.6036074,0.52472687,0.5007198,0.5178677,0.53844523,0.58645946,0.6173257,0.58988905,0.4664239,0.36010668,0.31895164,0.34295875,0.3806842,0.36010668,0.34638834,0.32924038,0.32238123,0.36010668,0.48357183,0.7339317,0.96371406,0.94999576,0.72364295,0.5796003,0.52472687,0.59331864,0.85739684,1.4404267,2.5207467,3.1620796,3.216953,3.1277838,3.316411,4.170378,5.579939,5.7479887,5.470192,4.9934793,4.0057583,3.4947495,3.2272418,3.2032347,3.4810312,4.190956,5.7274113,6.2898636,6.159539,5.717122,5.453044,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.017147938,0.024007112,0.030866288,0.048014224,0.058302987,0.061732575,0.061732575,0.06859175,0.06516216,0.06859175,0.07545093,0.07888051,0.08573969,0.08573969,0.06516216,0.044584636,0.034295876,0.041155048,0.05144381,0.06859175,0.082310095,0.07888051,0.06859175,0.0548734,0.05144381,0.06516216,0.07888051,0.0548734,0.05144381,0.044584636,0.037725464,0.0274367,0.034295876,0.06859175,0.10288762,0.1097468,0.1097468,0.13375391,0.18519773,0.16119061,0.106317215,0.06516216,0.07888051,0.06516216,0.041155048,0.0274367,0.024007112,0.041155048,0.07545093,0.09259886,0.08916927,0.07545093,0.06859175,0.058302987,0.06859175,0.06859175,0.0548734,0.058302987,0.082310095,0.106317215,0.1097468,0.082310095,0.020577524,0.061732575,0.08916927,0.11317638,0.12346515,0.11317638,0.13032432,0.1371835,0.10288762,0.037725464,0.010288762,0.010288762,0.017147938,0.01371835,0.0,0.0,0.01371835,0.01371835,0.037725464,0.082310095,0.14404267,0.274367,0.34981793,0.40126175,0.42526886,0.4081209,0.37725464,0.34981793,0.28465575,0.19548649,0.15090185,0.14404267,0.14404267,0.1371835,0.12003556,0.09602845,0.061732575,0.05144381,0.058302987,0.06859175,0.06859175,0.061732575,0.05144381,0.037725464,0.024007112,0.01371835,0.006859175,0.006859175,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.11317638,0.14061308,0.09602845,0.037725464,0.13375391,0.24350071,0.2709374,0.18862732,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.030866288,0.14747226,0.16119061,0.06859175,0.017147938,0.0034295875,0.0,0.0034295875,0.020577524,0.072021335,0.26064864,0.19891608,0.07888051,0.006859175,0.010288762,0.08916927,0.33266997,0.58988905,0.70649505,0.53501564,0.29151493,0.13032432,0.07888051,0.08916927,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.017147938,0.06516216,0.1097468,0.14404267,0.21263443,0.4664239,0.7099246,0.881404,0.9774324,1.0357354,1.2003556,1.4747226,1.4541451,1.1317638,0.89169276,0.6036074,0.764798,1.1146159,1.3478279,1.097468,0.64133286,0.41840968,0.26750782,0.13375391,0.05144381,0.06516216,0.09945804,0.1097468,0.08916927,0.0548734,0.12003556,0.21263443,0.32924038,0.48700142,0.70649505,0.96714365,1.1866373,1.4472859,1.7662375,2.095478,2.4247184,2.4041407,2.3561265,2.4247184,2.5447538,3.0729103,3.3712845,3.2306714,2.7779658,2.5070283,2.5447538,2.860276,3.9508848,5.6348124,7.051232,8.052671,9.191295,9.424506,8.656279,7.7097125,7.233,6.9346256,6.759717,6.800872,7.3084507,9.091836,11.091286,12.109874,12.332796,13.327377,15.244516,14.925565,13.54687,11.96926,10.717461,9.582268,8.577398,7.888051,7.5039372,7.2021337,7.250148,6.416758,5.31929,4.3795834,3.799983,3.40901,3.1689389,3.2066643,3.5599117,4.1600895,3.3061223,3.1415021,3.532475,4.232111,4.866585,3.5016088,1.9102802,0.82996017,0.4698535,0.5453044,0.65162164,0.4664239,0.2709374,0.16462019,0.06859175,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.030866288,0.0548734,0.082310095,0.08573969,0.07888051,0.06859175,0.058302987,0.06516216,0.06859175,0.06516216,0.058302987,0.07888051,0.18519773,0.20234565,0.18862732,0.1920569,0.24350071,0.28808534,0.2709374,0.25378948,0.28465575,0.39440256,0.48357183,0.5796003,0.6962063,0.8745448,1.1763484,1.255229,1.313532,1.3101025,1.2312219,1.097468,0.9431366,0.7990939,0.83681935,0.96714365,0.8711152,0.7956643,0.8848336,1.1008976,1.3992717,1.7250825,1.6907866,1.3992717,1.0425946,0.7579388,0.6001778,0.6344737,0.72021335,0.72364295,0.6379033,0.607037,0.61046654,0.6036074,0.5796003,0.5658819,0.6001778,0.53844523,0.41840968,0.32581082,0.32238123,0.432128,0.6859175,1.0734608,1.2003556,1.0082988,0.78537554,0.6241849,0.5555932,0.6001778,0.84024894,1.4027013,1.7662375,1.8725548,1.9514352,2.1880767,2.7299516,3.5633414,3.9611735,4.105216,4.091498,3.9474552,3.7691166,3.5839188,3.8479972,4.2115335,3.542764,4.5030484,5.768566,6.4544835,6.368744,6.0052075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0034295875,0.010288762,0.017147938,0.030866288,0.05144381,0.07545093,0.09259886,0.09945804,0.106317215,0.116605975,0.13032432,0.1371835,0.12689474,0.1371835,0.12346515,0.10288762,0.082310095,0.061732575,0.048014224,0.061732575,0.07545093,0.07888051,0.06859175,0.07545093,0.09945804,0.12003556,0.12003556,0.07888051,0.07545093,0.06859175,0.058302987,0.044584636,0.034295876,0.0548734,0.072021335,0.07545093,0.072021335,0.09602845,0.19891608,0.20920484,0.16804978,0.11317638,0.1097468,0.106317215,0.082310095,0.061732575,0.048014224,0.037725464,0.07545093,0.11317638,0.13032432,0.12346515,0.09602845,0.09259886,0.12003556,0.12003556,0.07888051,0.05144381,0.07545093,0.106317215,0.12346515,0.11317638,0.082310095,0.12689474,0.15433143,0.17147937,0.17833854,0.17833854,0.15776102,0.17490897,0.15776102,0.09945804,0.07545093,0.058302987,0.048014224,0.034295876,0.017147938,0.01371835,0.01371835,0.024007112,0.058302987,0.12689474,0.22292319,0.34638834,0.44584638,0.48700142,0.47328308,0.4389872,0.42869842,0.37725464,0.29151493,0.20577525,0.18176813,0.1371835,0.12003556,0.11317638,0.106317215,0.09945804,0.058302987,0.044584636,0.061732575,0.07888051,0.06859175,0.05144381,0.034295876,0.020577524,0.01371835,0.006859175,0.006859175,0.0034295875,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0034295875,0.006859175,0.030866288,0.08916927,0.16804978,0.15776102,0.06516216,0.017147938,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0274367,0.09602845,0.08916927,0.01371835,0.0,0.0,0.0034295875,0.017147938,0.048014224,0.1097468,0.07888051,0.037725464,0.010288762,0.010288762,0.05144381,0.20234565,0.42183927,0.5693115,0.5521636,0.31552204,0.13032432,0.0548734,0.08573969,0.13375391,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.010288762,0.020577524,0.024007112,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.006859175,0.024007112,0.0548734,0.15776102,0.29494452,0.4115505,0.5007198,0.58302987,0.86082643,1.5124481,1.7833855,1.605047,1.5741806,1.5604624,1.6839274,1.6873571,1.5604624,1.5330256,1.0425946,0.77851635,0.607037,0.45270553,0.32581082,0.25721905,0.14061308,0.08916927,0.106317215,0.08573969,0.08916927,0.12346515,0.1920569,0.274367,0.34295875,0.41498008,0.61046654,0.8162418,1.0700313,1.5604624,2.1229146,2.4041407,2.4898806,2.534465,2.784825,3.3781435,3.799983,3.9646032,3.8720043,3.57363,3.6799474,3.799983,4.170378,4.839148,5.6348124,6.5539417,7.881192,8.573969,8.4264965,8.093826,8.028665,7.932636,7.6925645,7.349606,7.1266828,8.110974,9.914937,11.235329,11.80464,12.363663,14.503725,14.822677,14.078457,12.88839,11.742908,10.563129,9.626852,9.033533,8.683716,8.30646,8.39563,7.9120584,7.116394,6.2658563,5.6176643,4.9591837,4.372724,4.012617,3.8960114,3.8960114,3.4055803,2.7230926,2.6064866,3.2958336,4.4721823,3.683377,2.4658735,1.6084765,1.3478279,1.3443983,1.2106444,0.84367853,0.5178677,0.31895164,0.16119061,0.07888051,0.0274367,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.058302987,0.10288762,0.12689474,0.13032432,0.12689474,0.12689474,0.16119061,0.15433143,0.14747226,0.1371835,0.12346515,0.1097468,0.17490897,0.21263443,0.23664154,0.25721905,0.29151493,0.33609957,0.36696586,0.39783216,0.45613512,0.5658819,0.69963586,0.7956643,0.89855194,1.0528834,1.3169615,1.4438564,1.7559488,2.0131679,2.07833,1.9274281,1.646202,1.3684053,1.3272504,1.4095604,1.1729189,1.0288762,1.1214751,1.4507155,1.9480057,2.4795918,2.4898806,2.2498093,1.8588364,1.4335675,1.0940384,0.97057325,0.9259886,0.84024894,0.72707254,0.72364295,0.8025235,0.86082643,0.85739684,0.84367853,0.96714365,0.90541106,0.69963586,0.5212973,0.44927597,0.48700142,0.66533995,0.9842916,1.2415106,1.3203912,1.1866373,0.881404,0.6379033,0.4938606,0.47328308,0.59331864,0.7373613,0.8711152,1.0631721,1.3203912,1.5844694,1.8348293,2.2120838,2.5310357,2.8054025,3.2306714,3.2306714,3.093488,3.3472774,3.6936657,3.018037,3.3884325,4.2423997,5.0312047,5.6176643,6.293293,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.030866288,0.058302987,0.08916927,0.106317215,0.12346515,0.15090185,0.16804978,0.16804978,0.15090185,0.18519773,0.20577525,0.20234565,0.17833854,0.1371835,0.082310095,0.07545093,0.08916927,0.106317215,0.106317215,0.13375391,0.15776102,0.16119061,0.14747226,0.14404267,0.16119061,0.15433143,0.13032432,0.10288762,0.07545093,0.07888051,0.082310095,0.072021335,0.0548734,0.06859175,0.1371835,0.20234565,0.23664154,0.22635277,0.18862732,0.16119061,0.15090185,0.14061308,0.12346515,0.10288762,0.12003556,0.15090185,0.16462019,0.15090185,0.13032432,0.15090185,0.17147937,0.15090185,0.09259886,0.05144381,0.072021335,0.09945804,0.13032432,0.16119061,0.19548649,0.22292319,0.22978236,0.23664154,0.2469303,0.2469303,0.2194936,0.21263443,0.19548649,0.16804978,0.16119061,0.1097468,0.07545093,0.058302987,0.05144381,0.041155048,0.030866288,0.041155048,0.082310095,0.15433143,0.26407823,0.37382504,0.4664239,0.4629943,0.3806842,0.32924038,0.35324752,0.32238123,0.2503599,0.17833854,0.17147937,0.106317215,0.10288762,0.10288762,0.08573969,0.07888051,0.05144381,0.044584636,0.061732575,0.07888051,0.058302987,0.037725464,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.024007112,0.030866288,0.024007112,0.020577524,0.061732575,0.13032432,0.14747226,0.12003556,0.061732575,0.017147938,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.058302987,0.0548734,0.0034295875,0.0,0.0,0.006859175,0.0274367,0.0548734,0.072021335,0.024007112,0.010288762,0.01371835,0.037725464,0.1097468,0.274367,0.33952916,0.31552204,0.24007112,0.15776102,0.07888051,0.024007112,0.044584636,0.08916927,0.0,0.0,0.0,0.010288762,0.024007112,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.006859175,0.020577524,0.030866288,0.034295876,0.024007112,0.030866288,0.0548734,0.061732575,0.048014224,0.024007112,0.006859175,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.020577524,0.006859175,0.0,0.0,0.0,0.030866288,0.116605975,0.33266997,0.5727411,0.5624523,0.36010668,0.64476246,0.91227025,1.0734608,1.4644338,2.020027,2.0749004,1.5158776,0.8711152,1.3101025,1.1900668,1.1043272,0.9911508,0.84024894,0.7099246,0.7956643,0.5178677,0.31552204,0.29837412,0.2503599,0.16119061,0.14404267,0.18176813,0.21263443,0.14061308,0.09602845,0.16462019,0.32581082,0.5624523,0.8779744,1.2037852,1.7525192,2.0886188,2.2258022,2.627064,3.3266997,3.9474552,4.4859004,4.7088237,4.170378,4.7534084,4.98662,4.938606,4.8117113,4.9660425,5.6142344,6.392751,7.160979,7.7885933,8.141841,8.364764,8.110974,7.7542973,7.5245147,7.500508,8.378482,9.619993,10.693454,11.183885,10.803201,11.770344,12.994707,13.639469,13.392539,12.46312,11.537132,10.772334,10.240748,9.921797,9.719451,9.6988735,9.534253,9.112414,8.498518,7.9292064,6.914048,5.813151,4.870014,4.262977,4.0949273,3.707384,2.6236343,2.0097382,2.2635276,3.0214665,2.8980014,2.603057,2.5173173,2.627064,2.527606,1.9102802,1.3512574,0.88826317,0.5418748,0.31895164,0.18862732,0.07888051,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.017147938,0.044584636,0.07888051,0.12346515,0.12346515,0.13032432,0.14061308,0.18862732,0.31552204,0.34981793,0.37382504,0.33952916,0.2469303,0.15090185,0.14404267,0.18862732,0.2503599,0.30523327,0.34981793,0.44584638,0.58645946,0.6962063,0.7510797,0.77165717,0.90198153,1.039165,1.1660597,1.2792361,1.3992717,1.7216529,2.4761622,3.1826572,3.5118976,3.2615378,2.74367,2.1880767,1.8416885,1.7182233,1.5810398,1.4644338,1.4129901,1.5741806,1.978872,2.5173173,2.6956558,2.7093742,2.4898806,2.0920484,1.6873571,1.3375391,1.0768905,0.89855194,0.78537554,0.7442205,0.8162418,0.90884066,0.96714365,1.0220171,1.1934965,1.2415106,1.1180456,0.91227025,0.7407909,0.7305021,0.8676856,0.91227025,1.0597426,1.3032433,1.4095604,1.0288762,0.6756287,0.44927597,0.3806842,0.42526886,0.4629943,0.52472687,0.6344737,0.77508676,0.89169276,1.0288762,1.196926,1.3855534,1.6084765,1.8999915,1.8519772,1.7422304,1.646202,1.7559488,2.3801336,2.8225505,2.6133456,2.6887965,3.5564823,5.302142,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.034295876,0.082310095,0.16804978,0.20577525,0.22292319,0.20920484,0.18862732,0.21263443,0.274367,0.35324752,0.37382504,0.31895164,0.26064864,0.18519773,0.15090185,0.15090185,0.17833854,0.22978236,0.216064,0.18519773,0.17833854,0.216064,0.29151493,0.2777966,0.25721905,0.2194936,0.17490897,0.1371835,0.15090185,0.17147937,0.16462019,0.12689474,0.09259886,0.10288762,0.19891608,0.30866286,0.3841138,0.39783216,0.29837412,0.26407823,0.24007112,0.20234565,0.15090185,0.14061308,0.16462019,0.20234565,0.22978236,0.22978236,0.22978236,0.22978236,0.22292319,0.20920484,0.19891608,0.19891608,0.23664154,0.26407823,0.26750782,0.24350071,0.23321195,0.23664154,0.2503599,0.26064864,0.26064864,0.26064864,0.26750782,0.26407823,0.22292319,0.1371835,0.06516216,0.0548734,0.06859175,0.07888051,0.09259886,0.07888051,0.07545093,0.106317215,0.17833854,0.274367,0.39783216,0.45613512,0.38754338,0.24350071,0.18176813,0.20920484,0.20577525,0.18519773,0.15776102,0.12346515,0.048014224,0.020577524,0.01371835,0.017147938,0.030866288,0.041155048,0.044584636,0.044584636,0.044584636,0.044584636,0.034295876,0.01371835,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0034295875,0.01371835,0.0274367,0.030866288,0.017147938,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.017147938,0.06859175,0.082310095,0.037725464,0.0,0.048014224,0.14404267,0.216064,0.21263443,0.09259886,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.16462019,0.15776102,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.06859175,0.1097468,0.12346515,0.1097468,0.041155048,0.12689474,0.35324752,0.48700142,0.34295875,0.12346515,0.0,0.0,0.0,0.0,0.0,0.048014224,0.11317638,0.07545093,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.01371835,0.030866288,0.030866288,0.041155048,0.037725464,0.048014224,0.072021335,0.061732575,0.037725464,0.01371835,0.0,0.0,0.0,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.044584636,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.0034295875,0.017147938,0.07888051,0.23664154,0.5658819,1.5158776,1.2586586,0.8162418,0.6276145,0.5796003,0.32238123,0.22292319,0.24007112,0.28808534,0.21263443,0.14061308,0.11317638,0.13032432,0.2194936,0.42869842,0.58645946,0.72707254,0.91569984,1.2003556,1.6016173,2.2120838,2.8877127,3.2032347,3.2272418,3.508468,4.180667,4.7602673,5.144381,5.3432975,5.4770513,5.453044,5.9983487,6.6431108,7.130112,7.3839016,7.9086285,7.0443726,6.660259,7.281014,8.086967,9.1981535,10.419086,10.950673,10.669447,10.131001,10.912948,12.133881,13.337666,13.855534,12.816368,12.281353,11.506266,10.772334,10.329918,10.39165,10.782623,10.916377,10.813489,10.443094,9.736599,8.330468,6.7357097,5.24041,4.2183924,4.1189346,3.9371665,3.2032347,2.4795918,2.0577524,1.9823016,2.1915064,2.867135,3.1209247,2.9665933,3.2958336,2.8088322,2.0097382,1.2758065,0.8093826,0.6241849,0.3566771,0.16119061,0.058302987,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.020577524,0.048014224,0.12346515,0.13375391,0.15433143,0.19891608,0.2777966,0.4115505,0.59674823,0.7133542,0.6344737,0.39783216,0.21263443,0.16462019,0.17147937,0.20920484,0.29151493,0.47328308,0.8025235,1.1694894,1.2860953,1.1146159,0.8711152,0.83338976,0.9877212,1.2517995,1.5090185,1.6324836,2.0234566,2.6236343,3.3815732,3.9337368,3.6147852,2.9803114,2.4007113,2.1640697,2.3389788,2.7779658,2.8877127,2.8225505,2.8534167,3.0043187,3.0660512,2.6407824,2.3767042,1.9857311,1.4918705,1.2346514,1.0906088,0.9328478,0.8128122,0.7579388,0.7922347,0.805953,0.75450927,0.75450927,0.84024894,0.9602845,1.255229,1.6016173,1.529596,1.1797781,1.3272504,1.6324836,1.5261664,1.2517995,1.08032,1.313532,1.0666018,0.77851635,0.5521636,0.4355576,0.4115505,0.45956472,0.47328308,0.45613512,0.42869842,0.42869842,0.5727411,0.6276145,0.59674823,0.53501564,0.53501564,0.58302987,0.65162164,0.7305021,0.84367853,1.039165,1.5398848,1.8279701,1.8656956,1.8828435,2.3972816,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.010288762,0.037725464,0.09602845,0.15090185,0.24007112,0.28465575,0.2777966,0.26407823,0.25378948,0.24350071,0.2194936,0.2194936,0.34638834,0.3806842,0.3018037,0.216064,0.17833854,0.216064,0.274367,0.28808534,0.26750782,0.22292319,0.16804978,0.14747226,0.15776102,0.19548649,0.24007112,0.2709374,0.28465575,0.28465575,0.2709374,0.2469303,0.18862732,0.11317638,0.15776102,0.20920484,0.23664154,0.28808534,0.31552204,0.30866286,0.3018037,0.3018037,0.26407823,0.2194936,0.20234565,0.18519773,0.17147937,0.1920569,0.1920569,0.22978236,0.23321195,0.1920569,0.16119061,0.18176813,0.18519773,0.18862732,0.18862732,0.18176813,0.19891608,0.2194936,0.25721905,0.3018037,0.31895164,0.3018037,0.30523327,0.29837412,0.26750782,0.22292319,0.18862732,0.16119061,0.14404267,0.14404267,0.16462019,0.2194936,0.29494452,0.34295875,0.33952916,0.26407823,0.2469303,0.24350071,0.22978236,0.20920484,0.20920484,0.21263443,0.20577525,0.2194936,0.24007112,0.19548649,0.072021335,0.0274367,0.01371835,0.017147938,0.030866288,0.034295876,0.034295876,0.0274367,0.020577524,0.020577524,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0034295875,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.006859175,0.024007112,0.041155048,0.0548734,0.024007112,0.020577524,0.020577524,0.017147938,0.0,0.020577524,0.061732575,0.106317215,0.116605975,0.041155048,0.034295876,0.0274367,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.030866288,0.006859175,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.020577524,0.1097468,0.16462019,0.13032432,0.037725464,0.024007112,0.017147938,0.23664154,0.66876954,1.039165,0.7922347,0.29151493,0.0,0.0,0.0,0.0,0.037725464,0.07888051,0.09945804,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.024007112,0.024007112,0.024007112,0.030866288,0.034295876,0.0274367,0.06516216,0.05144381,0.044584636,0.058302987,0.06859175,0.08916927,0.11317638,0.1371835,0.14061308,0.09602845,0.10288762,0.15090185,0.15433143,0.09602845,0.048014224,0.030866288,0.020577524,0.01371835,0.010288762,0.0,0.010288762,0.01371835,0.006859175,0.006859175,0.020577524,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.010288762,0.041155048,0.09259886,0.15090185,0.37039545,0.35324752,0.274367,0.2194936,0.18862732,0.28465575,0.41840968,0.45956472,0.3806842,0.2503599,0.18519773,0.116605975,0.106317215,0.18176813,0.32924038,0.48700142,0.5624523,0.58988905,0.6859175,1.0288762,2.07833,3.117495,3.8137012,3.998899,3.7039545,3.2546785,3.8308492,4.386442,4.602506,4.8905916,5.0826488,5.2335505,5.4153185,5.672538,6.0052075,6.2967224,7.0923867,7.6925645,7.6685576,6.842027,7.298162,8.275595,9.259886,9.921797,10.106995,10.175586,10.436234,11.417097,12.63803,12.596875,12.120162,11.519984,11.06042,10.943813,11.30735,11.862943,12.0309925,11.753197,11.135871,10.467101,9.767465,8.515666,7.0786686,5.844017,5.219832,4.5853586,3.7691166,2.9563043,2.4384367,2.6167753,2.8054025,3.1106358,3.3061223,3.292404,3.07634,2.4795918,1.9754424,1.5227368,1.0837497,0.6379033,0.34981793,0.20234565,0.10288762,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.0274367,0.037725464,0.072021335,0.09602845,0.13375391,0.18519773,0.2709374,0.42526886,0.6379033,0.7613684,0.6824879,0.42526886,0.16462019,0.12689474,0.16462019,0.2777966,0.51100856,0.94999576,1.0837497,1.0357354,0.89169276,0.7476501,0.69963586,0.8196714,1.1214751,1.5810398,2.1743584,2.901431,3.340418,3.5461934,3.7348208,3.875434,3.666229,3.391862,3.1140654,3.0386145,3.2718265,3.8377085,4.338428,4.0057583,3.2718265,2.4795918,1.9068506,1.529596,1.2792361,1.097468,0.9842916,0.9911508,0.980862,0.90541106,0.8128122,0.7510797,0.7579388,0.7579388,0.72707254,0.7407909,0.805953,0.84024894,0.91569984,1.138623,1.1729189,0.9911508,0.864256,0.90541106,1.0048691,1.1592005,1.3478279,1.5330256,1.1214751,0.7990939,0.58302987,0.47328308,0.44927597,0.4972902,0.45956472,0.37725464,0.30523327,0.30523327,0.42183927,0.47671264,0.4424168,0.36010668,0.34981793,0.4081209,0.4355576,0.4698535,0.5624523,0.7579388,0.90541106,1.0117283,1.0631721,1.1043272,1.2346514,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.041155048,0.08573969,0.16119061,0.22978236,0.28122616,0.33952916,0.28465575,0.34295875,0.36353627,0.32238123,0.31209245,0.31209245,0.28122616,0.24007112,0.21263443,0.20577525,0.21263443,0.22292319,0.23664154,0.23321195,0.1920569,0.19548649,0.22635277,0.29494452,0.3841138,0.432128,0.30523327,0.29151493,0.33609957,0.37039545,0.32238123,0.21263443,0.16119061,0.1371835,0.13032432,0.17833854,0.216064,0.2503599,0.28465575,0.28808534,0.20920484,0.17490897,0.16462019,0.15776102,0.16462019,0.2194936,0.3018037,0.32238123,0.3841138,0.45270553,0.37382504,0.28808534,0.24007112,0.2469303,0.2709374,0.20577525,0.24350071,0.2709374,0.29837412,0.32924038,0.34638834,0.31209245,0.30866286,0.2709374,0.19891608,0.17147937,0.18176813,0.21263443,0.2503599,0.32581082,0.51100856,0.5041494,0.490431,0.4629943,0.39783216,0.23321195,0.17490897,0.17490897,0.18862732,0.19548649,0.18519773,0.17147937,0.1371835,0.13032432,0.14747226,0.12346515,0.061732575,0.0274367,0.01371835,0.017147938,0.020577524,0.0274367,0.030866288,0.024007112,0.01371835,0.01371835,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.030866288,0.041155048,0.058302987,0.15090185,0.15090185,0.048014224,0.0,0.0034295875,0.024007112,0.05144381,0.06859175,0.020577524,0.01371835,0.01371835,0.006859175,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.020577524,0.024007112,0.006859175,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.06859175,0.09259886,0.072021335,0.01371835,0.0034295875,0.0034295875,0.106317215,0.3018037,0.48014224,0.36353627,0.13375391,0.0,0.0,0.0,0.006859175,0.274367,0.5212973,0.5144381,0.06516216,0.020577524,0.010288762,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.020577524,0.0548734,0.08573969,0.13032432,0.10288762,0.09602845,0.116605975,0.07545093,0.08916927,0.14061308,0.16119061,0.13032432,0.08573969,0.07888051,0.08916927,0.09945804,0.09945804,0.08916927,0.116605975,0.16462019,0.16804978,0.11317638,0.061732575,0.044584636,0.030866288,0.030866288,0.058302987,0.12689474,0.06859175,0.05144381,0.048014224,0.037725464,0.006859175,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.017147938,0.041155048,0.072021335,0.09602845,0.12346515,0.20920484,0.6344737,0.7956643,0.70306545,0.44927597,0.18519773,0.12346515,0.08573969,0.072021335,0.09602845,0.15776102,0.22978236,0.28122616,0.32924038,0.42183927,0.65505123,1.2963841,1.8931323,2.3801336,2.750529,3.059192,3.0351849,3.3609958,3.5461934,3.6147852,4.1155047,5.206114,6.077229,6.1766872,5.7377,5.761707,5.8988905,6.3824625,6.6225333,6.3310184,5.5250654,5.686256,6.5196457,7.682276,8.838047,9.644,9.688584,9.650859,10.377932,11.598865,11.938394,11.72233,11.616013,11.543991,11.633161,12.212761,12.812939,13.049581,12.919256,12.542002,12.161317,11.159878,10.336777,9.499957,8.570539,7.579388,6.3447366,5.31929,4.180667,3.2409601,3.4535947,3.2992632,3.0146074,3.0420442,3.5770597,4.5853586,3.4227283,2.3629858,1.5673214,1.0837497,0.83338976,0.51100856,0.30523327,0.15776102,0.048014224,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.037725464,0.05144381,0.061732575,0.06859175,0.08573969,0.12689474,0.1920569,0.28122616,0.41840968,0.6379033,0.7888051,0.6962063,0.39783216,0.12346515,0.08916927,0.32238123,0.6756287,0.9774324,1.0323058,1.0494537,1.0185875,1.0048691,1.0700313,1.2586586,1.6976458,2.3835633,3.0626216,3.6627994,4.3007026,4.698535,4.839148,4.7945633,4.540774,3.9714622,3.6044965,3.3129816,3.1620796,3.1826572,3.3644254,3.457024,3.0557625,2.4624438,1.8999915,1.5261664,1.2998136,1.0768905,0.91912943,0.8711152,0.9568549,0.9534253,0.88826317,0.8128122,0.7682276,0.78537554,0.7922347,0.764798,0.77165717,0.8265306,0.89169276,0.980862,1.0940384,1.097468,0.97057325,0.8128122,0.7579388,0.83338976,1.0460242,1.3272504,1.5398848,1.155771,0.8265306,0.58645946,0.432128,0.3566771,0.33952916,0.26750782,0.19891608,0.16804978,0.18176813,0.24007112,0.26064864,0.23664154,0.19548649,0.21263443,0.26064864,0.29494452,0.33952916,0.42526886,0.5761707,0.64476246,0.6790583,0.70649505,0.7305021,0.75450927,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.020577524,0.05144381,0.10288762,0.17147937,0.25721905,0.36353627,0.33952916,0.41840968,0.4664239,0.42183927,0.31209245,0.26064864,0.2469303,0.24350071,0.24350071,0.2469303,0.22635277,0.20920484,0.216064,0.22978236,0.22292319,0.23664154,0.26407823,0.31895164,0.3806842,0.3841138,0.2469303,0.2709374,0.36010668,0.41840968,0.34295875,0.24350071,0.17147937,0.12689474,0.11317638,0.14061308,0.16804978,0.25378948,0.32924038,0.34638834,0.26407823,0.19891608,0.19891608,0.2194936,0.24350071,0.29151493,0.37725464,0.38754338,0.4389872,0.5178677,0.4698535,0.39440256,0.32924038,0.30523327,0.30866286,0.26407823,0.31552204,0.31895164,0.29837412,0.2709374,0.26064864,0.2469303,0.2709374,0.25378948,0.216064,0.274367,0.30523327,0.36696586,0.45956472,0.607037,0.86082643,0.7407909,0.6207553,0.5178677,0.41498008,0.2503599,0.16804978,0.15433143,0.15433143,0.14747226,0.1371835,0.1371835,0.1097468,0.09602845,0.106317215,0.1097468,0.07888051,0.044584636,0.024007112,0.01371835,0.01371835,0.024007112,0.0274367,0.024007112,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.010288762,0.01371835,0.058302987,0.09602845,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.017147938,0.048014224,0.14747226,0.14747226,0.044584636,0.0,0.0,0.006859175,0.024007112,0.041155048,0.0274367,0.01371835,0.017147938,0.020577524,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.0274367,0.0274367,0.006859175,0.006859175,0.010288762,0.01371835,0.010288762,0.010288762,0.010288762,0.01371835,0.020577524,0.024007112,0.01371835,0.006859175,0.006859175,0.0034295875,0.0034295875,0.010288762,0.0034295875,0.0034295875,0.006859175,0.010288762,0.024007112,0.048014224,0.29151493,0.5144381,0.4972902,0.06516216,0.030866288,0.020577524,0.020577524,0.01371835,0.006859175,0.0,0.0034295875,0.010288762,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.020577524,0.010288762,0.0,0.0,0.0,0.017147938,0.017147938,0.048014224,0.10288762,0.10288762,0.12346515,0.10288762,0.09602845,0.1097468,0.09945804,0.10288762,0.20234565,0.25721905,0.22292319,0.12689474,0.12346515,0.11317638,0.09945804,0.082310095,0.07545093,0.10288762,0.12003556,0.12689474,0.13375391,0.15776102,0.1920569,0.19891608,0.18519773,0.16462019,0.18176813,0.09602845,0.06859175,0.061732575,0.0548734,0.048014224,0.06859175,0.0548734,0.034295876,0.01371835,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.01371835,0.024007112,0.041155048,0.08573969,0.1920569,0.5693115,0.66533995,0.5590228,0.3566771,0.17833854,0.09945804,0.09602845,0.12003556,0.1371835,0.14061308,0.09945804,0.11317638,0.15776102,0.23664154,0.3806842,0.64476246,0.89512235,1.1900668,1.862266,3.5016088,4.5270553,4.5819287,4.012617,3.3884325,3.5153272,4.57164,5.9640527,6.5882373,6.416758,6.495639,6.697984,6.5230756,6.3207297,6.1149545,5.6073756,5.7068334,6.3310184,7.1232533,7.98408,9.057541,8.759167,8.597976,9.208443,10.439664,11.334786,10.988399,11.207891,11.502836,11.818358,12.542002,13.2690735,13.756075,14.1299,14.359683,14.260224,13.186764,12.329367,11.454823,10.401938,9.095266,7.7577267,6.591667,5.353586,4.2835546,4.1326528,3.6936657,3.1826572,3.059192,3.57363,4.73969,3.8685746,2.9460156,1.9308578,1.138623,1.2346514,0.99801,0.66191036,0.33266997,0.09602845,0.037725464,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.0274367,0.0548734,0.09259886,0.12003556,0.12003556,0.12003556,0.14747226,0.22292319,0.32924038,0.41840968,0.5555932,0.6859175,0.6344737,0.4046913,0.15433143,0.14404267,0.53501564,1.0185875,1.2826657,1.0254467,1.0871792,1.2517995,1.4541451,1.6804979,1.9514352,2.486451,3.2683969,4.0091877,4.523626,4.7499785,4.8597255,4.8494368,4.664239,4.266407,3.6456516,3.2512488,2.9665933,2.7813954,2.6613598,2.568761,2.3595562,2.0131679,1.6667795,1.4027013,1.2449403,1.1043272,0.9328478,0.7990939,0.7476501,0.805953,0.7990939,0.7579388,0.72021335,0.7133542,0.7407909,0.7407909,0.7099246,0.69963586,0.72707254,0.7990939,0.89855194,0.9568549,0.9842916,0.9842916,0.9568549,0.9294182,0.9568549,1.097468,1.3203912,1.5090185,1.2620882,1.0357354,0.83681935,0.6756287,0.5693115,0.48357183,0.31209245,0.18862732,0.16119061,0.18862732,0.22978236,0.22292319,0.20234565,0.1920569,0.20920484,0.20920484,0.2194936,0.2469303,0.29837412,0.3566771,0.42183927,0.4629943,0.48357183,0.4938606,0.490431,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.041155048,0.06859175,0.11317638,0.16804978,0.23664154,0.33266997,0.40126175,0.42526886,0.44927597,0.47328308,0.44927597,0.37382504,0.31209245,0.274367,0.2709374,0.31895164,0.31895164,0.2777966,0.24350071,0.23321195,0.23321195,0.22635277,0.23664154,0.2469303,0.24007112,0.1920569,0.17833854,0.2503599,0.33952916,0.3806842,0.29494452,0.2777966,0.22635277,0.17833854,0.15090185,0.15433143,0.1920569,0.31552204,0.41498008,0.4424168,0.39783216,0.29151493,0.29151493,0.33266997,0.36353627,0.3566771,0.36353627,0.3841138,0.38754338,0.3841138,0.42526886,0.4424168,0.39440256,0.32238123,0.2777966,0.32924038,0.3841138,0.35324752,0.28122616,0.20234565,0.16462019,0.18862732,0.2503599,0.28465575,0.31895164,0.48014224,0.5144381,0.58645946,0.70306545,0.8505377,0.9774324,0.82996017,0.6893471,0.5624523,0.4389872,0.30866286,0.18862732,0.1371835,0.11317638,0.09259886,0.09945804,0.13375391,0.14404267,0.14747226,0.15090185,0.16804978,0.12003556,0.072021335,0.037725464,0.017147938,0.01371835,0.01371835,0.024007112,0.024007112,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.020577524,0.020577524,0.01371835,0.0034295875,0.0,0.0034295875,0.010288762,0.017147938,0.024007112,0.01371835,0.0274367,0.11317638,0.1920569,0.037725464,0.006859175,0.0034295875,0.0034295875,0.006859175,0.010288762,0.020577524,0.030866288,0.044584636,0.058302987,0.06516216,0.072021335,0.08916927,0.06516216,0.01371835,0.0,0.0,0.0,0.0034295875,0.017147938,0.037725464,0.0274367,0.030866288,0.041155048,0.041155048,0.01371835,0.0034295875,0.006859175,0.01371835,0.017147938,0.01371835,0.006859175,0.017147938,0.020577524,0.01371835,0.01371835,0.024007112,0.041155048,0.05144381,0.044584636,0.01371835,0.01371835,0.010288762,0.01371835,0.017147938,0.01371835,0.01371835,0.017147938,0.01371835,0.006859175,0.0034295875,0.006859175,0.017147938,0.024007112,0.030866288,0.058302987,0.08573969,0.07888051,0.06516216,0.06516216,0.08573969,0.06516216,0.05144381,0.037725464,0.0274367,0.024007112,0.024007112,0.05144381,0.06516216,0.048014224,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.041155048,0.024007112,0.006859175,0.010288762,0.01371835,0.0274367,0.030866288,0.06516216,0.10288762,0.061732575,0.01371835,0.037725464,0.037725464,0.024007112,0.08916927,0.106317215,0.19548649,0.28465575,0.30866286,0.19548649,0.20920484,0.18519773,0.14404267,0.10288762,0.06859175,0.07545093,0.06516216,0.07888051,0.15433143,0.29494452,0.4115505,0.45270553,0.4046913,0.28122616,0.14404267,0.10288762,0.082310095,0.06516216,0.06516216,0.12346515,0.15090185,0.13375391,0.08916927,0.037725464,0.0,0.0034295875,0.0034295875,0.006859175,0.010288762,0.0,0.0,0.0034295875,0.010288762,0.0274367,0.044584636,0.0274367,0.030866288,0.034295876,0.0274367,0.006859175,0.006859175,0.010288762,0.017147938,0.017147938,0.017147938,0.024007112,0.01371835,0.010288762,0.024007112,0.0548734,0.12003556,0.16119061,0.21263443,0.29494452,0.41840968,0.32924038,0.31209245,0.31895164,0.31552204,0.26407823,0.14747226,0.12346515,0.1097468,0.106317215,0.18176813,0.38754338,0.6241849,0.90884066,1.7525192,4.15323,5.8508763,5.970912,5.086078,3.9303071,3.391862,3.6010668,4.839148,6.125243,7.0272245,7.6616983,8.008087,7.5279446,7.1952744,7.164408,6.783724,6.9346256,7.250148,7.3564653,7.407909,8.107545,7.3084507,7.133542,7.7542973,9.057541,10.652299,9.9698105,10.127572,10.556271,11.084427,11.965831,12.946692,13.872682,14.88441,15.731518,15.7966795,15.175924,14.177915,12.912396,11.434244,9.736599,8.611694,7.438775,6.416758,5.6176643,4.9523244,4.4584637,4.0091877,3.649081,3.4192986,3.340418,3.426158,3.316411,2.4761622,1.4061309,1.6496316,1.6084765,1.2620882,0.8265306,0.4629943,0.28465575,0.16804978,0.072021335,0.017147938,0.0034295875,0.0,0.0,0.0,0.020577524,0.041155048,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0274367,0.07888051,0.15433143,0.22292319,0.22635277,0.20234565,0.21263443,0.28122616,0.3806842,0.4115505,0.41840968,0.47328308,0.4938606,0.42183927,0.23664154,0.29837412,0.764798,1.2175035,1.371835,1.0940384,1.2860953,1.6256244,1.9582944,2.2120838,2.386993,2.6956558,3.1415021,3.6799474,4.108646,4.091498,3.875434,3.6147852,3.316411,3.0146074,2.767677,2.5447538,2.3629858,2.2326615,2.136633,2.0646117,1.937717,1.7113642,1.4472859,1.1934965,1.0048691,0.8471081,0.71678376,0.6276145,0.58302987,0.5693115,0.5693115,0.5555932,0.548734,0.5624523,0.58645946,0.5727411,0.5453044,0.5178677,0.50757897,0.53158605,0.5658819,0.61389613,0.7339317,0.91227025,1.0528834,1.0940384,1.1214751,1.1934965,1.3066728,1.3992717,1.3032433,1.2277923,1.1283343,1.0117283,0.939707,0.84367853,0.58988905,0.36353627,0.26750782,0.28465575,0.33266997,0.32238123,0.3018037,0.29151493,0.28122616,0.23321195,0.18176813,0.16119061,0.15776102,0.12346515,0.16804978,0.22978236,0.2709374,0.274367,0.26064864,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.041155048,0.09259886,0.12689474,0.18176813,0.20920484,0.22292319,0.31895164,0.4664239,0.4938606,0.5178677,0.607037,0.77851635,0.6927767,0.5418748,0.40126175,0.31895164,0.31895164,0.30866286,0.26064864,0.26064864,0.30523327,0.30523327,0.28122616,0.25721905,0.23321195,0.216064,0.22978236,0.216064,0.21263443,0.24350071,0.31895164,0.4424168,0.58988905,0.432128,0.23664154,0.13032432,0.106317215,0.14404267,0.28122616,0.34638834,0.31209245,0.274367,0.23664154,0.2469303,0.32581082,0.4046913,0.31895164,0.29494452,0.36353627,0.45613512,0.5212973,0.53501564,0.4355576,0.40126175,0.37725464,0.35324752,0.36696586,0.4389872,0.42183927,0.37382504,0.33609957,0.33609957,0.36010668,0.39440256,0.37039545,0.31895164,0.3806842,0.45613512,0.64819205,0.7990939,0.8162418,0.67219913,0.7682276,0.7579388,0.65162164,0.490431,0.31895164,0.16119061,0.13032432,0.14404267,0.15090185,0.1371835,0.16119061,0.17833854,0.15776102,0.12003556,0.106317215,0.12003556,0.08573969,0.048014224,0.0274367,0.01371835,0.01371835,0.024007112,0.017147938,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.0548734,0.09602845,0.10288762,0.06516216,0.01371835,0.0034295875,0.017147938,0.024007112,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.034295876,0.044584636,0.09602845,0.15090185,0.2194936,0.28465575,0.31895164,0.3566771,0.4389872,0.32238123,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.041155048,0.072021335,0.08916927,0.07545093,0.041155048,0.048014224,0.037725464,0.0,0.0,0.061732575,0.11317638,0.1371835,0.12346515,0.07545093,0.06516216,0.05144381,0.041155048,0.0274367,0.01371835,0.01371835,0.024007112,0.030866288,0.0274367,0.01371835,0.0274367,0.048014224,0.061732575,0.058302987,0.044584636,0.044584636,0.044584636,0.06859175,0.13375391,0.24350071,0.18176813,0.13032432,0.09602845,0.072021335,0.061732575,0.1097468,0.22292319,0.216064,0.08916927,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.0274367,0.048014224,0.061732575,0.037725464,0.030866288,0.024007112,0.01371835,0.0,0.0,0.037725464,0.048014224,0.041155048,0.07545093,0.06516216,0.116605975,0.2503599,0.36696586,0.24350071,0.20920484,0.14404267,0.08916927,0.058302987,0.044584636,0.020577524,0.024007112,0.037725464,0.08916927,0.26064864,0.4424168,0.48700142,0.4389872,0.32581082,0.16804978,0.16804978,0.17833854,0.15776102,0.12346515,0.12346515,0.2194936,0.19891608,0.12003556,0.037725464,0.0,0.024007112,0.020577524,0.010288762,0.0,0.0,0.0,0.010288762,0.058302987,0.14404267,0.22978236,0.14404267,0.07545093,0.044584636,0.041155048,0.030866288,0.030866288,0.020577524,0.020577524,0.030866288,0.030866288,0.0548734,0.041155048,0.024007112,0.030866288,0.09259886,0.17833854,0.24350071,0.44584638,0.78537554,1.1146159,1.1146159,0.94999576,0.71678376,0.48357183,0.29151493,0.1920569,0.22292319,0.22978236,0.17147937,0.12346515,0.26750782,0.37725464,0.5624523,0.8711152,1.2963841,2.2600982,3.2546785,3.9851806,4.2595477,3.9680326,4.417309,5.15467,6.0703697,7.1266828,8.347616,8.457363,7.81603,7.1987042,6.941485,6.941485,7.160979,7.181556,7.016936,6.6431108,5.9983487,5.8508763,6.169828,6.708273,7.5519514,9.139851,8.89635,8.615124,8.64599,9.208443,10.39165,11.622872,13.039291,14.359683,15.258235,15.3817,15.110763,15.110763,14.863832,13.862392,11.581717,9.956093,8.820899,8.069819,7.517656,6.883182,6.5024977,5.693115,4.6402316,3.6353626,3.0969174,3.0729103,2.8568463,2.393852,1.8588364,1.6633499,1.7971039,1.903421,1.9171394,1.7010754,1.0528834,0.6241849,0.24350071,0.048014224,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.12346515,0.26407823,0.3841138,0.39783216,0.33609957,0.34638834,0.35324752,0.33952916,0.34981793,0.32581082,0.31209245,0.31209245,0.31209245,0.274367,0.48357183,1.0288762,1.4541451,1.5330256,1.2517995,1.4335675,1.8005334,2.1297739,2.3252604,2.411,2.3389788,2.2360911,2.287535,2.5653315,3.0660512,3.1037767,2.8945718,2.5996273,2.3767042,2.3664153,2.2669573,2.1057668,1.9514352,1.8554068,1.8313997,1.8313997,1.786815,1.6804979,1.529596,1.3581166,1.1626302,0.9774324,0.823101,0.7133542,0.64133286,0.5555932,0.48700142,0.432128,0.39097297,0.36696586,0.39097297,0.39783216,0.3841138,0.36010668,0.33609957,0.31209245,0.34981793,0.47328308,0.65162164,0.8093826,0.8711152,0.89512235,0.91227025,0.9362774,0.9602845,0.91227025,0.864256,0.78537554,0.70649505,0.7339317,0.7442205,0.64819205,0.48357183,0.31895164,0.26064864,0.26064864,0.26064864,0.26064864,0.25721905,0.24350071,0.19548649,0.14747226,0.116605975,0.09945804,0.07545093,0.08916927,0.09945804,0.106317215,0.11317638,0.1371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.0548734,0.10288762,0.16462019,0.22292319,0.28465575,0.3806842,0.4115505,0.432128,0.48357183,0.58645946,0.71678376,0.7888051,0.6173257,0.44584638,0.39097297,0.48014224,0.44584638,0.32924038,0.2503599,0.26064864,0.32924038,0.33609957,0.274367,0.18519773,0.1097468,0.082310095,0.09945804,0.10288762,0.14404267,0.22292319,0.29494452,0.29494452,0.20577525,0.1097468,0.06516216,0.12003556,0.116605975,0.12003556,0.17833854,0.2709374,0.32238123,0.4046913,0.39097297,0.35324752,0.33266997,0.34638834,0.37039545,0.42526886,0.48014224,0.5041494,0.4972902,0.42869842,0.432128,0.3841138,0.29837412,0.32924038,0.42183927,0.4664239,0.4629943,0.42869842,0.4081209,0.3566771,0.36353627,0.40126175,0.45613512,0.52815646,0.65848076,0.823101,0.90198153,0.8676856,0.78194594,0.7407909,0.65848076,0.53501564,0.4115505,0.3566771,0.29494452,0.2469303,0.18519773,0.12346515,0.11317638,0.18519773,0.1920569,0.17833854,0.17833854,0.216064,0.18862732,0.13032432,0.072021335,0.0274367,0.01371835,0.01371835,0.017147938,0.010288762,0.0034295875,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.020577524,0.020577524,0.01371835,0.0034295875,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.006859175,0.010288762,0.020577524,0.030866288,0.06516216,0.106317215,0.11317638,0.1097468,0.14061308,0.1097468,0.034295876,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0034295875,0.044584636,0.072021335,0.06859175,0.07545093,0.06859175,0.072021335,0.06859175,0.061732575,0.061732575,0.12346515,0.14404267,0.106317215,0.041155048,0.041155048,0.16462019,0.20920484,0.18176813,0.106317215,0.01371835,0.006859175,0.01371835,0.0274367,0.044584636,0.05144381,0.07545093,0.08916927,0.09259886,0.082310095,0.06859175,0.1097468,0.13375391,0.14747226,0.18862732,0.31895164,0.432128,0.38754338,0.28808534,0.19548649,0.13375391,0.11317638,0.1371835,0.12003556,0.058302987,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.010288762,0.017147938,0.020577524,0.024007112,0.030866288,0.030866288,0.024007112,0.01371835,0.0,0.0,0.006859175,0.010288762,0.006859175,0.01371835,0.041155048,0.10288762,0.15433143,0.15776102,0.072021335,0.0548734,0.07888051,0.1097468,0.12346515,0.082310095,0.037725464,0.020577524,0.020577524,0.0274367,0.05144381,0.116605975,0.20920484,0.23321195,0.18176813,0.12003556,0.09945804,0.082310095,0.0548734,0.024007112,0.024007112,0.044584636,0.048014224,0.0548734,0.08916927,0.15776102,0.11317638,0.08573969,0.09945804,0.13032432,0.12346515,0.024007112,0.0034295875,0.010288762,0.0274367,0.044584636,0.0274367,0.01371835,0.010288762,0.010288762,0.017147938,0.037725464,0.061732575,0.09602845,0.14061308,0.18862732,0.12689474,0.1371835,0.274367,0.48700142,0.6173257,0.45613512,0.28808534,0.24007112,0.32581082,0.42869842,0.6241849,0.8093826,0.84024894,0.72364295,0.607037,0.5796003,0.64133286,0.75450927,0.91569984,1.1592005,1.1214751,0.7956643,0.52472687,0.490431,0.72364295,1.2860953,2.0165975,2.2635276,2.0097382,1.8931323,2.3732746,2.9631636,3.4810312,4.170378,5.672538,6.495639,6.9037595,7.181556,7.48336,7.8331776,7.449064,6.948344,6.4579134,6.042933,5.7274113,5.6485305,5.4976287,5.809721,6.7357097,8.028665,8.323608,8.052671,7.582818,7.500508,8.597976,10.055551,11.46854,12.758065,13.876111,14.805529,15.806969,16.678083,16.702091,15.621771,13.63261,11.794352,10.779194,10.179015,9.568549,8.505377,7.431916,6.4819202,5.6210938,4.6608095,3.2546785,2.3732746,2.3801336,2.5961976,2.4967396,1.7353712,2.0646117,2.0749004,1.8519772,1.471293,0.980862,0.65162164,0.5796003,0.5212973,0.37725464,0.19548649,0.048014224,0.01371835,0.01371835,0.010288762,0.0,0.058302987,0.08916927,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.0274367,0.041155048,0.072021335,0.14747226,0.25378948,0.33952916,0.31209245,0.41498008,0.4115505,0.35324752,0.29151493,0.26407823,0.24007112,0.33609957,0.490431,0.66876954,0.83681935,1.2003556,2.1160555,2.7470996,2.6750782,1.8862731,1.8348293,2.136633,2.5241764,2.8945718,3.3026927,3.3541365,3.0317552,2.7711067,2.8705647,3.457024,3.5804894,3.0557625,2.4555845,2.095478,2.0234566,2.054323,2.0749004,2.085189,2.0817597,2.0749004,2.0646117,2.0749004,2.1091962,2.1400626,2.1160555,1.7833855,1.3855534,1.0151579,0.72364295,0.5418748,0.4389872,0.36010668,0.28808534,0.22978236,0.19548649,0.17147937,0.18519773,0.19548649,0.18176813,0.17833854,0.17147937,0.20234565,0.274367,0.3841138,0.5041494,0.5727411,0.6379033,0.7099246,0.7922347,0.8745448,0.8265306,0.72021335,0.58302987,0.44584638,0.35324752,0.31895164,0.28122616,0.25378948,0.23321195,0.20920484,0.1920569,0.16462019,0.14404267,0.13375391,0.12346515,0.11317638,0.10288762,0.09259886,0.07888051,0.06516216,0.058302987,0.041155048,0.034295876,0.037725464,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.037725464,0.07545093,0.12689474,0.1920569,0.26750782,0.32581082,0.4046913,0.44927597,0.48700142,0.6001778,0.65848076,0.5658819,0.4629943,0.4664239,0.66533995,0.5041494,0.36696586,0.31209245,0.34981793,0.4629943,0.4972902,0.44927597,0.34295875,0.21263443,0.12003556,0.106317215,0.12003556,0.13032432,0.13032432,0.13032432,0.18176813,0.2194936,0.22635277,0.18862732,0.09602845,0.06859175,0.06516216,0.13032432,0.24350071,0.34638834,0.44584638,0.3841138,0.3018037,0.274367,0.29494452,0.28808534,0.28808534,0.32581082,0.4046913,0.5144381,0.59331864,0.66191036,0.64819205,0.53501564,0.37382504,0.36353627,0.36353627,0.36696586,0.37039545,0.3806842,0.37382504,0.39097297,0.45270553,0.5453044,0.61046654,0.69963586,0.89855194,0.9431366,0.78537554,0.6241849,0.61046654,0.6893471,0.7682276,0.7407909,0.51100856,0.36696586,0.26064864,0.18862732,0.15090185,0.15090185,0.20234565,0.2777966,0.31209245,0.29151493,0.25378948,0.25378948,0.30866286,0.24007112,0.06859175,0.006859175,0.006859175,0.006859175,0.006859175,0.010288762,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.024007112,0.020577524,0.024007112,0.024007112,0.010288762,0.006859175,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.006859175,0.010288762,0.01371835,0.0,0.0,0.030866288,0.048014224,0.058302987,0.11317638,0.12689474,0.09945804,0.06859175,0.06516216,0.08573969,0.10288762,0.09602845,0.058302987,0.017147938,0.030866288,0.19548649,0.21263443,0.16462019,0.10288762,0.041155048,0.024007112,0.0274367,0.05144381,0.09259886,0.12346515,0.16462019,0.17147937,0.15433143,0.17147937,0.34295875,0.4115505,0.4698535,0.58302987,0.78194594,1.0768905,0.83338976,0.607037,0.42869842,0.30523327,0.22635277,0.16119061,0.1097468,0.06516216,0.0274367,0.006859175,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.0274367,0.06859175,0.13032432,0.17490897,0.16119061,0.18862732,0.20234565,0.19891608,0.18519773,0.16462019,0.12003556,0.06516216,0.030866288,0.017147938,0.017147938,0.07545093,0.20234565,0.2469303,0.18519773,0.10288762,0.12003556,0.1920569,0.274367,0.31552204,0.26407823,0.17833854,0.116605975,0.08916927,0.09259886,0.1097468,0.06516216,0.09602845,0.12346515,0.13032432,0.15090185,0.16462019,0.1097468,0.13032432,0.19891608,0.1097468,0.044584636,0.058302987,0.13375391,0.22292319,0.25378948,0.15433143,0.106317215,0.09602845,0.09602845,0.061732575,0.01371835,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.048014224,0.06859175,0.09259886,0.058302987,0.06516216,0.13375391,0.24007112,0.29837412,0.21263443,0.12003556,0.07888051,0.09945804,0.14061308,0.28122616,0.44584638,0.4972902,0.4972902,0.72364295,0.70306545,0.5624523,0.5178677,0.6001778,0.66876954,0.61389613,0.42183927,0.42183927,0.7305021,1.2655178,1.0185875,1.3752645,1.4678634,1.1283343,0.8779744,1.1043272,1.4027013,1.7182233,2.153781,2.9803114,3.7176728,4.57164,5.7308407,7.058091,8.083538,8.220721,7.805741,7.1061053,6.4098988,6.0086374,5.802862,5.579939,5.5833683,5.9400454,6.6636887,7.654839,8.351046,7.936065,6.948344,7.2604365,8.416207,9.705732,11.015835,12.257345,13.354814,15.594335,17.051908,17.233677,16.19794,14.565458,13.749216,13.1421795,12.380811,11.266195,9.770895,8.556821,7.8091707,7.14726,6.2212715,4.715683,3.316411,2.6956558,2.8396983,3.0557625,1.9925903,2.1880767,2.2086544,1.9720128,1.5227368,1.0357354,0.9259886,1.0597426,1.0768905,0.86082643,0.5453044,0.39097297,0.21263443,0.08573969,0.06859175,0.16462019,0.22978236,0.17833854,0.082310095,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.030866288,0.06859175,0.1097468,0.16804978,0.22635277,0.30523327,0.41840968,0.5658819,0.4698535,0.432128,0.41498008,0.39097297,0.36353627,0.34638834,0.65505123,1.0563129,1.3752645,1.4987297,1.5501735,1.9857311,2.603057,2.9906003,2.5207467,2.294394,2.4212887,2.8945718,3.7348208,5.007198,4.938606,4.8254294,4.722542,4.650521,4.616225,4.184097,3.3712845,2.6922262,2.3595562,2.2566686,2.1880767,2.136633,2.1880767,2.3149714,2.3664153,2.352697,2.318401,2.270387,2.2086544,2.1126258,1.7250825,1.2963841,0.90198153,0.59331864,0.40126175,0.30523327,0.24350071,0.18862732,0.1371835,0.106317215,0.09945804,0.11317638,0.12003556,0.11317638,0.12003556,0.12689474,0.14061308,0.16804978,0.2194936,0.29837412,0.33609957,0.3841138,0.45270553,0.5453044,0.64476246,0.66191036,0.61046654,0.53158605,0.4389872,0.32238123,0.22978236,0.18862732,0.18176813,0.20234565,0.23664154,0.19548649,0.14061308,0.09945804,0.07888051,0.072021335,0.06516216,0.05144381,0.044584636,0.041155048,0.041155048,0.037725464,0.030866288,0.0274367,0.034295876,0.030866288,0.041155048,0.037725464,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.05144381,0.106317215,0.15090185,0.2503599,0.3566771,0.39783216,0.40126175,0.45956472,0.48357183,0.4355576,0.39783216,0.45270553,0.67219913,0.5590228,0.548734,0.5418748,0.5007198,0.4698535,0.45613512,0.47671264,0.51100856,0.47671264,0.20920484,0.13375391,0.13032432,0.11317638,0.06859175,0.034295876,0.09945804,0.17147937,0.21263443,0.18862732,0.06516216,0.041155048,0.05144381,0.09259886,0.15433143,0.22292319,0.29494452,0.274367,0.25721905,0.26750782,0.2709374,0.31209245,0.32581082,0.30866286,0.31209245,0.42526886,0.5521636,0.6207553,0.6276145,0.5624523,0.4046913,0.41840968,0.38754338,0.36010668,0.35324752,0.37382504,0.42183927,0.42183927,0.432128,0.4698535,0.51100856,0.5796003,0.75450927,0.77508676,0.6207553,0.5212973,0.53158605,0.66191036,0.7990939,0.8265306,0.58645946,0.4389872,0.29837412,0.19548649,0.15090185,0.15776102,0.18176813,0.2777966,0.4081209,0.5144381,0.52815646,0.53158605,0.5521636,0.37382504,0.07545093,0.006859175,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.024007112,0.010288762,0.0034295875,0.0,0.0034295875,0.017147938,0.0274367,0.030866288,0.024007112,0.017147938,0.030866288,0.034295876,0.030866288,0.020577524,0.010288762,0.006859175,0.0,0.006859175,0.010288762,0.017147938,0.017147938,0.037725464,0.05144381,0.0548734,0.06859175,0.12346515,0.13375391,0.09602845,0.08573969,0.12689474,0.17833854,0.116605975,0.058302987,0.024007112,0.017147938,0.030866288,0.17147937,0.16462019,0.106317215,0.06516216,0.048014224,0.044584636,0.06859175,0.116605975,0.16804978,0.20920484,0.24007112,0.22292319,0.1920569,0.39440256,1.2826657,1.3958421,1.2586586,1.2175035,1.3992717,1.7319417,1.1489118,0.77165717,0.5521636,0.432128,0.33609957,0.24007112,0.15090185,0.10288762,0.10288762,0.12689474,0.16804978,0.18862732,0.18176813,0.16119061,0.15090185,0.17490897,0.22292319,0.26407823,0.28122616,0.2709374,0.4115505,0.6927767,1.0014396,1.2175035,1.2277923,1.1180456,0.8128122,0.53158605,0.36696586,0.29837412,0.29494452,0.31895164,0.34981793,0.3566771,0.30523327,0.32581082,0.42183927,0.53844523,0.61046654,0.58302987,0.48700142,0.42526886,0.4046913,0.4046913,0.37382504,0.2709374,0.22292319,0.2194936,0.23664154,0.26750782,0.23664154,0.17147937,0.20234565,0.274367,0.15776102,0.072021335,0.082310095,0.15090185,0.216064,0.19891608,0.15433143,0.12689474,0.08573969,0.030866288,0.0,0.0034295875,0.010288762,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.024007112,0.024007112,0.030866288,0.048014224,0.08916927,0.14404267,0.16119061,0.20234565,0.4664239,0.44584638,0.2777966,0.17490897,0.17147937,0.106317215,0.08573969,0.06516216,0.2194936,0.58302987,1.039165,0.64133286,0.7579388,0.8265306,0.66533995,0.4698535,0.53844523,0.6241849,0.83681935,1.1694894,1.4987297,1.7902447,2.4590142,3.6627994,5.212973,6.5950966,7.514226,7.8263187,7.682276,7.3221693,7.0752387,6.8728933,6.680836,6.416758,6.138962,6.0326443,7.1061053,8.543102,8.759167,7.7714453,7.174697,7.81603,8.621983,9.561689,10.607714,11.760056,14.613472,17.137648,18.166525,17.62122,16.513464,16.191082,15.645778,14.634049,13.097594,11.1393,9.9801,9.174147,8.429926,7.5519514,6.4304767,4.822,3.7451096,3.4021509,3.3266997,2.3904223,2.311542,2.3081124,2.07833,1.6221949,1.2346514,1.1180456,1.1729189,1.196926,1.0768905,0.77851635,0.72364295,0.6310441,0.5418748,0.45270553,0.30523327,0.58645946,0.50757897,0.29151493,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.034295876,0.07545093,0.116605975,0.22292319,0.28122616,0.33952916,0.4629943,0.71678376,0.6379033,0.5796003,0.53158605,0.4938606,0.48357183,0.5178677,0.8471081,1.2998136,1.670209,1.7113642,1.529596,1.6084765,2.1503513,2.8637056,2.959734,3.2203827,3.5118976,3.9337368,4.636802,5.796003,6.101236,6.495639,6.7494283,6.7048435,6.245279,5.3158607,4.2595477,3.6079261,3.474172,3.5393343,3.3472774,2.9734523,2.633923,2.469303,2.5481834,2.6133456,2.5893385,2.4624438,2.2223728,1.879414,1.5364552,1.1866373,0.864256,0.6001778,0.4046913,0.3018037,0.2194936,0.15433143,0.11317638,0.09602845,0.09602845,0.10288762,0.11317638,0.12689474,0.15090185,0.15090185,0.15776102,0.16804978,0.19548649,0.23321195,0.23321195,0.25378948,0.29837412,0.36353627,0.4355576,0.48700142,0.4938606,0.47671264,0.4424168,0.37382504,0.29494452,0.26750782,0.2709374,0.2777966,0.2709374,0.20234565,0.1371835,0.09259886,0.06516216,0.061732575,0.048014224,0.034295876,0.024007112,0.020577524,0.024007112,0.024007112,0.0274367,0.034295876,0.037725464,0.030866288,0.08916927,0.07888051,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.06859175,0.09602845,0.19548649,0.26407823,0.31209245,0.33952916,0.33609957,0.34981793,0.3018037,0.30866286,0.4081209,0.5555932,0.61046654,0.7407909,0.7579388,0.607037,0.34638834,0.274367,0.3566771,0.548734,0.64133286,0.25378948,0.14404267,0.12003556,0.116605975,0.09945804,0.06516216,0.048014224,0.05144381,0.0548734,0.05144381,0.048014224,0.05144381,0.05144381,0.048014224,0.044584636,0.034295876,0.072021335,0.15090185,0.22292319,0.26064864,0.2469303,0.39097297,0.490431,0.4389872,0.28808534,0.24007112,0.28465575,0.31552204,0.32924038,0.34295875,0.39097297,0.5453044,0.58988905,0.5693115,0.53158605,0.5144381,0.5727411,0.5521636,0.47328308,0.39440256,0.36696586,0.44584638,0.52815646,0.53844523,0.5144381,0.59674823,0.6036074,0.607037,0.607037,0.59331864,0.53844523,0.48700142,0.35324752,0.22292319,0.14747226,0.15090185,0.20234565,0.29494452,0.48700142,0.7510797,0.9568549,0.939707,0.7613684,0.4046913,0.037725464,0.01371835,0.0034295875,0.0034295875,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0034295875,0.0,0.0,0.006859175,0.020577524,0.037725464,0.048014224,0.020577524,0.0034295875,0.0,0.006859175,0.037725464,0.058302987,0.06516216,0.048014224,0.030866288,0.061732575,0.0548734,0.041155048,0.030866288,0.024007112,0.01371835,0.006859175,0.0034295875,0.010288762,0.024007112,0.0548734,0.1097468,0.12003556,0.116605975,0.12346515,0.1371835,0.12003556,0.09259886,0.13032432,0.22292319,0.29151493,0.16462019,0.058302987,0.017147938,0.030866288,0.037725464,0.13032432,0.12346515,0.072021335,0.0274367,0.030866288,0.05144381,0.1097468,0.18862732,0.26064864,0.3018037,0.29151493,0.2469303,0.216064,0.6756287,2.5378947,2.767677,2.301253,1.8485477,1.7113642,1.8176813,1.2380811,0.8848336,0.70306545,0.6241849,0.5624523,0.45270553,0.32924038,0.26750782,0.28122616,0.34981793,0.45270553,0.5212973,0.5144381,0.45270553,0.41498008,0.4389872,0.45270553,0.4046913,0.32924038,0.31895164,0.5555932,1.138623,1.845118,2.4452958,2.702515,2.5756202,2.0097382,1.4575747,1.1283343,0.9911508,0.84024894,0.6344737,0.5727411,0.64133286,0.58988905,0.5555932,0.6276145,0.7407909,0.83338976,0.84367853,0.8025235,0.7922347,0.78194594,0.7407909,0.6173257,0.5453044,0.48014224,0.4424168,0.42869842,0.40126175,0.274367,0.2194936,0.21263443,0.20234565,0.1371835,0.082310095,0.072021335,0.07888051,0.07888051,0.061732575,0.12003556,0.1371835,0.08573969,0.006859175,0.006859175,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.0274367,0.044584636,0.048014224,0.044584636,0.034295876,0.024007112,0.01371835,0.020577524,0.030866288,0.037725464,0.037725464,0.0274367,0.024007112,0.024007112,0.024007112,0.01371835,0.024007112,0.048014224,0.09945804,0.14404267,0.09602845,0.12346515,0.16462019,0.22635277,0.31209245,0.42526886,0.51100856,0.5007198,0.59674823,0.8505377,1.1454822,1.1454822,1.3101025,1.7971039,2.6716487,3.8925817,5.2575574,6.5162163,7.486789,8.110974,8.460793,8.56368,8.498518,8.22758,7.654839,6.636252,7.1026754,8.556821,9.637141,9.589127,8.268735,8.419638,8.525954,8.745448,9.290752,10.415657,13.080446,16.726099,19.003344,19.294859,18.69811,17.936743,17.305698,16.403717,14.959861,12.809509,11.581717,10.340206,9.253027,8.447074,8.018375,6.6465406,5.6210938,4.7328305,3.8891523,3.1209247,2.6785078,2.4624438,2.1434922,1.7319417,1.5638919,1.2689474,1.0494537,1.0220171,1.0768905,0.8848336,0.89169276,1.039165,1.1146159,0.9294182,0.34638834,0.7956643,0.75450927,0.48357183,0.18176813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.01371835,0.041155048,0.06859175,0.07888051,0.20577525,0.274367,0.32581082,0.41840968,0.6241849,0.77851635,0.72364295,0.6001778,0.5144381,0.548734,0.67219913,0.8779744,1.1729189,1.4575747,1.5124481,1.3752645,1.4781522,1.8965619,2.5207467,3.0420442,4.383013,5.394741,5.892031,5.9914894,6.0978065,6.8043017,7.363324,7.8263187,8.107545,7.9737906,6.9860697,5.6793966,4.9008803,4.8597255,5.130663,4.928317,4.307562,3.5050385,2.8739944,2.884283,3.0523329,3.0351849,2.7642474,2.2669573,1.6770682,1.430138,1.1934965,0.9842916,0.7956643,0.607037,0.4424168,0.29494452,0.20234565,0.16804978,0.17833854,0.20577525,0.24007112,0.3018037,0.3841138,0.44927597,0.39097297,0.34295875,0.32924038,0.33609957,0.30866286,0.28808534,0.28465575,0.29494452,0.31552204,0.33952916,0.36696586,0.39097297,0.4046913,0.41498008,0.41840968,0.42526886,0.4664239,0.5041494,0.48700142,0.37725464,0.274367,0.19548649,0.14061308,0.09945804,0.07545093,0.058302987,0.05144381,0.05144381,0.044584636,0.034295876,0.0274367,0.034295876,0.034295876,0.030866288,0.0274367,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.16804978,0.15090185,0.16462019,0.23664154,0.274367,0.2503599,0.2709374,0.37382504,0.53158605,0.64133286,0.5796003,0.51100856,0.5041494,0.50757897,0.33609957,0.4081209,0.41840968,0.3566771,0.25378948,0.16804978,0.15433143,0.20920484,0.26407823,0.28465575,0.26064864,0.17490897,0.12346515,0.09602845,0.072021335,0.061732575,0.072021335,0.06859175,0.0548734,0.044584636,0.044584636,0.09602845,0.12346515,0.12003556,0.08916927,0.07545093,0.16119061,0.31895164,0.4046913,0.34981793,0.16804978,0.14404267,0.22978236,0.3018037,0.32924038,0.36696586,0.5007198,0.78194594,0.9774324,1.0048691,0.9294182,0.980862,1.0185875,0.9328478,0.7339317,0.548734,0.5624523,0.61046654,0.66533995,0.71678376,0.77851635,0.8745448,0.78194594,0.65848076,0.5727411,0.48700142,0.37725464,0.29494452,0.25378948,0.2503599,0.274367,0.432128,0.6824879,0.7682276,0.7613684,1.0528834,1.0768905,0.7888051,0.37039545,0.024007112,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.037725464,0.044584636,0.041155048,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.010288762,0.0,0.0,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.030866288,0.041155048,0.09259886,0.17833854,0.20920484,0.2194936,0.23664154,0.26064864,0.22292319,0.17833854,0.16462019,0.1920569,0.22978236,0.13032432,0.06859175,0.058302987,0.072021335,0.061732575,0.14747226,0.12346515,0.061732575,0.017147938,0.030866288,0.041155048,0.09259886,0.20920484,0.34981793,0.4115505,0.36353627,0.32238123,0.28808534,0.805953,2.9906003,3.4913201,2.9940298,2.2052248,1.5638919,1.2209331,1.0494537,0.9534253,0.9294182,0.9774324,1.097468,0.9877212,0.7510797,0.548734,0.45956472,0.47328308,0.58302987,0.72021335,0.7888051,0.7682276,0.7339317,0.70649505,0.6927767,0.6310441,0.52815646,0.4424168,0.45613512,0.65162164,1.1008976,1.8485477,2.8980014,2.8877127,2.5721905,2.2806756,2.1503513,2.1503513,1.8828435,1.5947582,1.3203912,1.0666018,0.8093826,0.6379033,0.59674823,0.6001778,0.6241849,0.6859175,0.77165717,0.78537554,0.6927767,0.5418748,0.45613512,0.5418748,0.58302987,0.5693115,0.51100856,0.42869842,0.31895164,0.26407823,0.24350071,0.23664154,0.19891608,0.11317638,0.082310095,0.06859175,0.061732575,0.061732575,0.061732575,0.06859175,0.058302987,0.030866288,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.05144381,0.216064,0.45613512,0.61046654,0.42869842,0.2194936,0.15090185,0.20920484,0.40126175,0.71678376,0.764798,0.65162164,0.47328308,0.37382504,0.53501564,0.97400284,0.9568549,0.980862,1.3409687,2.1194851,3.292404,4.804852,6.40304,7.864044,8.988949,9.6817255,10.179015,10.456812,10.14129,8.467651,8.2481575,9.208443,10.686595,11.427385,9.595985,9.427936,9.146709,8.858624,8.803751,9.352485,11.30735,14.486577,17.014183,17.977898,17.439453,16.269962,16.441442,16.657507,16.153357,14.723219,12.977559,11.362224,10.000677,9.263316,9.750318,9.39707,8.567109,7.4353456,6.111525,4.623084,3.6353626,2.8465576,2.3046827,2.0165975,1.9685832,1.7971039,1.471293,1.3306799,1.3478279,1.1283343,0.922559,0.9431366,0.9431366,0.7613684,0.31895164,0.1371835,0.0548734,0.037725464,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0274367,0.08916927,0.15090185,0.15090185,0.15090185,0.18862732,0.2503599,0.33266997,0.4424168,0.4664239,0.4629943,0.432128,0.42869842,0.548734,0.78194594,1.1146159,1.2723769,1.2929544,1.5261664,1.5638919,1.5981878,1.7216529,2.0303159,2.6407824,4.897451,7.191845,8.56025,8.80718,8.515666,7.939495,7.2295704,7.2775846,8.207003,9.352485,8.803751,7.1095347,5.6656785,5.055212,5.0826488,5.055212,4.90431,4.623084,4.2869844,4.0434837,4.15323,3.8514268,3.0523329,2.0406046,1.4815818,1.2860953,1.1249046,1.0460242,1.0117283,0.89855194,0.607037,0.41498008,0.31895164,0.31209245,0.39783216,0.59331864,0.77851635,0.9842916,1.2037852,1.3889829,1.155771,0.88826317,0.71678376,0.6379033,0.5041494,0.45613512,0.41498008,0.39097297,0.37382504,0.34981793,0.34981793,0.38754338,0.4424168,0.5041494,0.5658819,0.65162164,0.7613684,0.84367853,0.84367853,0.7339317,0.59674823,0.45613512,0.31895164,0.20920484,0.1371835,0.09945804,0.082310095,0.09602845,0.12003556,0.106317215,0.06859175,0.06859175,0.058302987,0.0274367,0.01371835,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.034295876,0.037725464,0.10288762,0.22635277,0.31209245,0.33609957,0.33266997,0.37382504,0.42526886,0.34638834,0.28808534,0.29151493,0.34295875,0.4046913,0.4081209,0.33609957,0.42526886,0.5212973,0.5521636,0.53501564,0.4355576,0.32581082,0.2469303,0.2194936,0.22292319,0.19548649,0.16804978,0.15433143,0.14404267,0.12346515,0.11317638,0.1097468,0.10288762,0.09259886,0.082310095,0.12003556,0.14061308,0.1371835,0.106317215,0.06516216,0.082310095,0.28122616,0.40126175,0.34981793,0.20577525,0.20920484,0.34638834,0.45270553,0.4698535,0.4389872,0.4972902,0.5521636,0.53158605,0.44584638,0.39440256,0.4424168,0.48357183,0.5144381,0.5418748,0.5727411,0.4389872,0.42869842,0.4698535,0.5453044,0.6927767,0.9842916,0.84367853,0.7339317,0.7990939,0.89169276,0.77165717,0.47328308,0.2709374,0.26064864,0.37382504,0.5418748,0.7579388,0.9945804,1.138623,0.9911508,0.6756287,0.39097297,0.16462019,0.0274367,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.030866288,0.09602845,0.16804978,0.14747226,0.07888051,0.010288762,0.0,0.006859175,0.037725464,0.05144381,0.037725464,0.01371835,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0034295875,0.010288762,0.020577524,0.024007112,0.024007112,0.017147938,0.006859175,0.0,0.0034295875,0.01371835,0.034295876,0.08573969,0.14404267,0.1920569,0.20234565,0.17833854,0.18176813,0.216064,0.2503599,0.2469303,0.24007112,0.26064864,0.31552204,0.33952916,0.18176813,0.082310095,0.09602845,0.17490897,0.26407823,0.28122616,0.12346515,0.05144381,0.037725464,0.058302987,0.07888051,0.061732575,0.12689474,0.23321195,0.33266997,0.36353627,0.35324752,0.36010668,0.3566771,0.48700142,1.0494537,1.1317638,1.1797781,1.5638919,1.9548649,1.3306799,1.1214751,1.0494537,1.1077567,1.2998136,1.6359133,1.6221949,1.4404267,1.2415106,1.1454822,1.2037852,1.5776103,2.1126258,2.4075704,2.3595562,2.1469216,1.879414,1.6359133,1.4164196,1.3615463,1.7250825,1.9891608,2.1332035,2.2463799,2.2738166,1.99602,2.1880767,2.3801336,2.5173173,2.5653315,2.5173173,2.3664153,2.1880767,1.9480057,1.6736387,1.4541451,1.430138,1.3889829,1.2003556,0.939707,0.89512235,0.97057325,0.980862,0.8505377,0.64819205,0.59331864,0.5521636,0.5007198,0.47328308,0.5212973,0.72021335,0.85396725,0.86082643,0.8093826,0.7305021,0.6241849,0.30523327,0.17147937,0.20920484,0.31209245,0.29151493,0.17490897,0.13375391,0.10288762,0.058302987,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0034295875,0.030866288,0.21263443,0.33609957,0.31552204,0.2194936,0.2469303,0.29494452,0.48014224,0.7133542,0.6790583,0.7476501,0.8505377,0.9842916,1.1694894,1.4267083,1.5124481,1.3786942,1.1866373,1.0940384,1.2312219,1.9445761,3.2272418,4.729401,6.193835,7.4627824,8.381912,9.626852,10.377932,10.278474,9.458802,9.160428,10.350495,11.914387,12.651748,11.269625,10.062409,9.098696,8.584257,8.673427,9.47595,10.6488695,13.059869,15.7795315,17.761833,17.881868,16.952452,16.163645,15.573756,15.158776,14.784951,14.376831,13.87954,13.046151,12.055,11.509696,11.194174,10.950673,10.419086,9.263316,7.1884155,5.161529,3.6696587,2.843128,2.7059445,3.1655092,2.3972816,1.6153357,1.1043272,0.9602845,1.0940384,1.0014396,1.0220171,0.9568549,0.71678376,0.3566771,0.29151493,0.274367,0.24007112,0.1920569,0.18176813,0.20234565,0.15776102,0.07888051,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.041155048,0.041155048,0.020577524,0.0,0.0,0.0,0.01371835,0.07545093,0.16119061,0.20234565,0.15090185,0.14747226,0.20234565,0.34638834,0.6001778,1.1043272,1.1180456,0.8196714,0.48700142,0.51100856,0.64819205,0.82996017,0.9602845,1.0220171,1.097468,1.4095604,1.4404267,1.4747226,1.7353712,2.3972816,4.420738,7.0375133,9.342196,10.686595,10.686595,8.56025,7.9017696,8.453933,9.506817,9.901219,8.707723,7.881192,7.56224,7.5519514,7.301592,7.64798,8.117833,8.498518,8.498518,7.716572,7.1129646,5.669108,3.841138,2.16064,1.2003556,1.1008976,1.0700313,1.0837497,1.1626302,1.3752645,1.611906,1.6599203,1.5638919,1.4129901,1.3615463,1.3306799,1.196926,1.0631721,1.0014396,1.0597426,0.9945804,0.7888051,0.58645946,0.47328308,0.45613512,0.4629943,0.4698535,0.4629943,0.44927597,0.42526886,0.42526886,0.432128,0.45613512,0.4938606,0.5144381,0.5418748,0.5693115,0.5796003,0.5624523,0.5007198,0.4629943,0.4046913,0.31895164,0.2194936,0.1371835,0.12003556,0.13032432,0.14747226,0.15433143,0.14404267,0.12689474,0.1097468,0.08573969,0.06516216,0.06516216,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.034295876,0.08916927,0.12689474,0.14404267,0.16119061,0.216064,0.28808534,0.31895164,0.37039545,0.42526886,0.44927597,0.4355576,0.3806842,0.28465575,0.30523327,0.36010668,0.4046913,0.4424168,0.40126175,0.32581082,0.2503599,0.1920569,0.15776102,0.16119061,0.15433143,0.15433143,0.15090185,0.12689474,0.116605975,0.106317215,0.09602845,0.082310095,0.0548734,0.06859175,0.10288762,0.12003556,0.106317215,0.07888051,0.058302987,0.13032432,0.18176813,0.16804978,0.11317638,0.13375391,0.2469303,0.4115505,0.5658819,0.6036074,0.6344737,0.6036074,0.4972902,0.34295875,0.21263443,0.21263443,0.2709374,0.34295875,0.41498008,0.5144381,0.58645946,0.51100856,0.42869842,0.44927597,0.67219913,0.9602845,0.94999576,0.805953,0.6859175,0.71678376,0.6173257,0.41840968,0.2777966,0.28122616,0.45956472,0.5727411,0.7510797,0.94656616,1.0494537,0.85739684,0.37382504,0.14061308,0.044584636,0.010288762,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.006859175,0.006859175,0.006859175,0.006859175,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.020577524,0.106317215,0.33266997,0.20577525,0.11317638,0.044584636,0.0034295875,0.0,0.020577524,0.06516216,0.072021335,0.037725464,0.006859175,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.006859175,0.01371835,0.020577524,0.010288762,0.010288762,0.024007112,0.048014224,0.06516216,0.058302987,0.030866288,0.01371835,0.006859175,0.006859175,0.034295876,0.072021335,0.16462019,0.26750782,0.33952916,0.34638834,0.30523327,0.30523327,0.30523327,0.29151493,0.2709374,0.29494452,0.36353627,0.45956472,0.4664239,0.18519773,0.08916927,0.15776102,0.3018037,0.37725464,0.18862732,0.072021335,0.0274367,0.0274367,0.048014224,0.06516216,0.0548734,0.12346515,0.23664154,0.36010668,0.48014224,0.58988905,0.6173257,0.53844523,0.42526886,0.44584638,0.48700142,0.72364295,1.2620882,1.7250825,1.2483698,1.1249046,1.3786942,1.8554068,2.2841053,2.311542,2.5721905,2.194936,1.7319417,1.529596,1.728512,2.253239,3.0454736,3.474172,3.3541365,2.9494452,2.4761622,2.0577524,1.8382589,1.8382589,1.9720128,2.0165975,1.9685832,1.8656956,1.7250825,1.5398848,1.5810398,1.7319417,1.9342873,2.1400626,2.3081124,2.294394,2.294394,2.0749004,1.6221949,1.1146159,1.0528834,1.0151579,0.8848336,0.69963586,0.6241849,0.66876954,0.7442205,0.7442205,0.6893471,0.70649505,0.7373613,0.77851635,0.8128122,0.9945804,1.6359133,2.0714707,2.1640697,1.9685832,1.5398848,0.9328478,0.4664239,0.26407823,0.22635277,0.24350071,0.20577525,0.15433143,0.16462019,0.18862732,0.18519773,0.14061308,0.07545093,0.030866288,0.01371835,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.017147938,0.01371835,0.017147938,0.024007112,0.010288762,0.010288762,0.01371835,0.01371835,0.017147938,0.0274367,0.13375391,0.26064864,0.35324752,0.42869842,0.5521636,0.6173257,0.52815646,0.51100856,0.61046654,0.67219913,0.8848336,1.1180456,1.9548649,3.2615378,4.201245,4.4275975,4.1600895,2.983741,1.5158776,1.4198492,1.5055889,1.9685832,2.8225505,4.029765,5.504488,7.332458,8.862054,9.770895,9.990388,9.73317,9.105555,10.244178,11.262765,11.194174,10.014396,8.995808,8.532814,8.4264965,8.735159,9.764035,10.666017,11.941824,14.006435,16.235666,16.96617,16.143068,14.908417,13.834956,13.310229,13.529722,14.188204,14.369971,13.920695,12.908967,11.626302,10.779194,10.861504,10.940384,10.398509,8.954653,6.9037595,5.271276,4.1772375,3.7279615,4.012617,3.4055803,2.4247184,1.6599203,1.313532,1.2037852,1.0837497,1.1180456,1.1489118,1.0117283,0.53158605,0.764798,0.7510797,0.64819205,0.5796003,0.6310441,0.5453044,0.36696586,0.2469303,0.2194936,0.20234565,0.041155048,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.030866288,0.024007112,0.006859175,0.0,0.0,0.01371835,0.11317638,0.2469303,0.26064864,0.16804978,0.13032432,0.17147937,0.28465575,0.42869842,2.318401,3.4398763,3.4021509,2.3732746,1.0700313,0.7476501,0.70649505,0.7956643,0.90884066,0.97400284,1.1454822,1.3032433,1.6599203,2.2463799,2.901431,4.1429415,5.90232,8.162418,10.124143,10.196163,8.378482,7.8263187,8.594546,9.877212,10.014396,9.184435,9.630281,10.950673,12.445972,13.13189,13.37882,13.313659,13.111313,12.836946,12.425395,11.485688,9.73317,7.4936485,5.219832,3.5016088,2.7470996,2.4007113,2.201795,2.1469216,2.4761622,2.8122618,2.9906003,2.9048605,2.5241764,1.8965619,1.4953002,1.0768905,0.7613684,0.61046654,0.6276145,0.5761707,0.48700142,0.4081209,0.36696586,0.38754338,0.4355576,0.4938606,0.53844523,0.5555932,0.5624523,0.58302987,0.6173257,0.6379033,0.64819205,0.65848076,0.6276145,0.6036074,0.6036074,0.6310441,0.66191036,0.66533995,0.58302987,0.45613512,0.32238123,0.22978236,0.20920484,0.22292319,0.22635277,0.20577525,0.17147937,0.15090185,0.14061308,0.13032432,0.12003556,0.10288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.06516216,0.13375391,0.22292319,0.3841138,0.5693115,0.70649505,0.77851635,0.8093826,0.6241849,0.45270553,0.33609957,0.29494452,0.3018037,0.29494452,0.25721905,0.20920484,0.16462019,0.12346515,0.1097468,0.10288762,0.10288762,0.106317215,0.08573969,0.072021335,0.06859175,0.06516216,0.05144381,0.024007112,0.024007112,0.05144381,0.07545093,0.07888051,0.072021335,0.061732575,0.0548734,0.058302987,0.058302987,0.041155048,0.058302987,0.11317638,0.24007112,0.39783216,0.4698535,0.52815646,0.5590228,0.5212973,0.4115505,0.26407823,0.17833854,0.23321195,0.28122616,0.28465575,0.3566771,0.5212973,0.45270553,0.32924038,0.34981793,0.7373613,0.97057325,0.9842916,0.7888051,0.5453044,0.5693115,0.51100856,0.42526886,0.35324752,0.33952916,0.44927597,0.45956472,0.53844523,0.6310441,0.65848076,0.5521636,0.18519773,0.044584636,0.010288762,0.0034295875,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.006859175,0.006859175,0.020577524,0.058302987,0.05144381,0.0034295875,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.017147938,0.09602845,0.29151493,0.13032432,0.041155048,0.006859175,0.0,0.006859175,0.024007112,0.048014224,0.048014224,0.020577524,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.006859175,0.01371835,0.0274367,0.041155048,0.041155048,0.05144381,0.06859175,0.07888051,0.058302987,0.0274367,0.020577524,0.024007112,0.030866288,0.058302987,0.082310095,0.14061308,0.20920484,0.26064864,0.26407823,0.2469303,0.26750782,0.274367,0.25378948,0.22292319,0.28465575,0.4081209,0.5178677,0.50757897,0.23664154,0.15776102,0.18519773,0.25378948,0.25378948,0.0548734,0.024007112,0.01371835,0.01371835,0.030866288,0.05144381,0.09602845,0.19548649,0.42869842,0.764798,1.0460242,1.138623,1.138623,0.89169276,0.5007198,0.36010668,0.548734,0.90884066,1.255229,1.3889829,1.1077567,1.0940384,1.4918705,2.1091962,2.5996273,2.4795918,2.6990852,2.294394,1.8279701,1.6427724,1.879414,2.3767042,3.2066643,3.7348208,3.74168,3.3952916,2.8705647,2.417859,2.1263442,1.9823016,1.8862731,1.8176813,1.7147937,1.5227368,1.3101025,1.2963841,1.2586586,1.2860953,1.3649758,1.5124481,1.7765263,2.0268862,2.0989075,1.9068506,1.5090185,1.1214751,0.9945804,0.96714365,0.9431366,0.9294182,1.0151579,1.2346514,1.1008976,0.9568549,0.9602845,1.0734608,1.5090185,2.0440342,1.9994495,1.6496316,2.253239,2.7573884,2.901431,2.651071,2.020027,1.0734608,0.5727411,0.32238123,0.20577525,0.14404267,0.09945804,0.09945804,0.13375391,0.17147937,0.17833854,0.14061308,0.07545093,0.034295876,0.017147938,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.010288762,0.017147938,0.017147938,0.010288762,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.017147938,0.01371835,0.017147938,0.024007112,0.010288762,0.01371835,0.020577524,0.017147938,0.01371835,0.034295876,0.13032432,0.18519773,0.26064864,0.39097297,0.5693115,0.85739684,0.9842916,1.0425946,1.0768905,1.0734608,1.3684053,1.5673214,2.2258022,3.2581081,3.9337368,4.331569,4.547633,3.6936657,2.2429502,2.0165975,1.6599203,1.313532,1.4438564,2.270387,3.765687,5.8543057,7.5382333,8.958082,9.952662,10.055551,9.362774,9.774324,10.010965,9.6988735,9.349055,9.06097,8.790032,8.652849,8.89635,9.884071,10.827208,11.231899,12.487128,14.5243025,15.817257,15.429714,13.989287,12.79922,12.5145645,13.118172,13.876111,14.006435,13.732068,12.950122,11.2421875,10.127572,10.155008,10.539123,10.765475,10.590566,9.146709,7.346176,5.6656785,4.5099077,4.214963,4.064061,3.0866287,2.1846473,1.7079345,1.4541451,1.3443983,1.1934965,1.255229,1.3546871,0.8711152,1.0048691,0.9842916,0.88826317,0.8711152,1.1249046,0.980862,0.66533995,0.3806842,0.23321195,0.21263443,0.041155048,0.07888051,0.14061308,0.116605975,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.006859175,0.0,0.0,0.017147938,0.12346515,0.28122616,0.34981793,0.24007112,0.16119061,0.15776102,0.216064,0.24007112,2.0474637,4.0537724,4.9488945,4.1772375,1.9239986,1.1454822,0.823101,0.78537554,0.8848336,0.99801,1.1043272,1.371835,2.0749004,3.0248961,3.5976372,4.081209,4.8905916,6.447624,8.210432,8.656279,8.090397,7.98065,8.584257,9.386781,9.122703,9.3936405,11.255906,13.934414,16.489456,17.823566,18.214539,18.142517,17.765263,17.2131,16.588915,14.839825,12.401388,9.942374,7.7920227,5.936616,4.7808447,4.201245,3.7519686,3.3609958,3.3232703,3.4535947,3.7142432,3.9371665,3.8685746,3.1895163,2.6990852,2.0474637,1.2963841,0.66533995,0.5007198,0.45270553,0.432128,0.42526886,0.42526886,0.42526886,0.432128,0.47671264,0.52472687,0.5624523,0.59331864,0.66876954,0.7956643,0.91912943,1.0082988,1.0494537,0.9602845,0.85396725,0.7990939,0.823101,0.91912943,0.939707,0.84367853,0.67219913,0.48357183,0.3566771,0.32238123,0.31895164,0.29837412,0.25378948,0.20234565,0.17147937,0.19548649,0.2194936,0.2194936,0.20234565,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.041155048,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.19891608,0.490431,0.7956643,1.0597426,1.2998136,1.0494537,0.75450927,0.52815646,0.4115505,0.35324752,0.30866286,0.2469303,0.19891608,0.17147937,0.1371835,0.07545093,0.05144381,0.044584636,0.041155048,0.034295876,0.020577524,0.020577524,0.024007112,0.020577524,0.01371835,0.01371835,0.01371835,0.020577524,0.037725464,0.037725464,0.061732575,0.07545093,0.082310095,0.072021335,0.0274367,0.041155048,0.061732575,0.07545093,0.08573969,0.106317215,0.1920569,0.31209245,0.39097297,0.39440256,0.32581082,0.19891608,0.22292319,0.22292319,0.17147937,0.19548649,0.24007112,0.22292319,0.17147937,0.24350071,0.7339317,0.90541106,0.82996017,0.6344737,0.4938606,0.64476246,0.61046654,0.52472687,0.4424168,0.39097297,0.37382504,0.33952916,0.33266997,0.33952916,0.33266997,0.26407823,0.14747226,0.06859175,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.010288762,0.010288762,0.0,0.0034295875,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.024007112,0.020577524,0.010288762,0.0,0.0,0.01371835,0.017147938,0.01371835,0.006859175,0.01371835,0.048014224,0.09945804,0.08573969,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.010288762,0.006859175,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0034295875,0.0,0.0034295875,0.010288762,0.034295876,0.082310095,0.07545093,0.06859175,0.06516216,0.058302987,0.034295876,0.017147938,0.034295876,0.0548734,0.06516216,0.06516216,0.0548734,0.037725464,0.030866288,0.030866288,0.0274367,0.041155048,0.09259886,0.14747226,0.17147937,0.14747226,0.22292319,0.36010668,0.44927597,0.42869842,0.29494452,0.2503599,0.17833854,0.08573969,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.0274367,0.058302987,0.17147937,0.32924038,0.69963586,1.2037852,1.5090185,1.3992717,1.3443983,1.0082988,0.52472687,0.4698535,0.88826317,1.3409687,1.4335675,1.1729189,0.96714365,1.039165,1.3341095,1.7593783,2.1297739,2.1743584,2.085189,1.920569,1.7833855,1.7456601,1.862266,2.1091962,2.6785078,3.1723683,3.3815732,3.2992632,2.9117198,2.5310357,2.1160555,1.762808,1.6907866,1.7353712,1.6839274,1.5021594,1.2655178,1.155771,1.1454822,1.1111864,1.1008976,1.1797781,1.4129901,1.8245405,1.8142518,1.6256244,1.4610043,1.4747226,1.4610043,1.5330256,1.670209,1.8965619,2.3081124,2.7333813,2.2600982,1.7696671,1.6530612,1.786815,2.527606,3.4055803,3.1723683,2.1674993,2.3424082,2.6304936,2.7162333,2.5996273,2.1469216,1.1077567,0.607037,0.32238123,0.18519773,0.13032432,0.09945804,0.07545093,0.072021335,0.06516216,0.048014224,0.0274367,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.020577524,0.030866288,0.030866288,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.020577524,0.017147938,0.0034295875,0.01371835,0.01371835,0.020577524,0.058302987,0.12689474,0.19548649,0.7510797,1.2998136,1.728512,1.920569,1.7833855,1.9171394,1.9068506,1.7182233,1.3992717,1.0666018,1.5090185,2.3664153,2.8328393,2.719663,2.4795918,1.8862731,1.1694894,0.8779744,1.3032433,2.469303,3.9886103,5.761707,7.881192,9.832627,10.484249,10.333347,9.928656,9.571979,9.5205345,10.014396,10.285333,9.736599,9.136421,9.016385,9.668007,10.604284,10.731179,11.495977,13.186764,14.949572,15.46401,14.116182,13.032433,13.035862,13.673765,13.924125,13.680624,13.4645605,13.011855,11.279913,10.120712,9.609704,9.846346,10.666017,11.64345,11.245617,9.602845,7.4181976,5.3913116,4.2218223,4.180667,3.3678548,2.5790498,2.1160555,1.7730967,1.6942163,1.2655178,1.214074,1.488441,1.2620882,1.0185875,0.9328478,0.8848336,0.9362774,1.3306799,1.1900668,0.91569984,0.59331864,0.32238123,0.22635277,0.13032432,0.2777966,0.36010668,0.26407823,0.07888051,0.10288762,0.08916927,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.08573969,0.21263443,0.3841138,0.34295875,0.24350071,0.18176813,0.16804978,0.15090185,0.64819205,2.5653315,4.2526884,4.4996185,2.5413244,1.488441,1.0563129,0.94656616,0.9774324,1.097468,1.2655178,1.5604624,2.4041407,3.57363,4.2115335,4.232111,4.355576,4.9214582,5.9160385,6.9792104,7.699424,8.237869,8.567109,8.546532,7.9292064,9.108984,11.64345,14.534592,16.986746,18.410025,20.251715,22.052248,23.19087,23.19773,21.753874,18.492336,14.7197895,11.784062,9.89093,8.107545,6.728851,5.9469047,5.40503,4.887162,4.32471,4.098357,4.2286816,4.712253,5.209543,5.0346346,4.5922174,3.8034124,2.5756202,1.3169615,0.94656616,0.939707,0.8505377,0.7407909,0.65162164,0.58645946,0.5041494,0.47328308,0.47328308,0.48700142,0.51100856,0.61389613,0.8196714,1.1043272,1.3786942,1.4987297,1.3786942,1.1797781,1.0117283,0.97057325,1.1214751,1.2209331,1.1866373,1.0185875,0.77165717,0.5521636,0.4629943,0.39783216,0.34295875,0.29151493,0.2469303,0.22978236,0.3018037,0.37039545,0.40126175,0.40126175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.12003556,0.12003556,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.0,0.0,0.06516216,0.18519773,0.34638834,0.5178677,0.59331864,0.61046654,0.6344737,0.67219913,0.67219913,0.58645946,0.5007198,0.41498008,0.31895164,0.19891608,0.08916927,0.05144381,0.041155048,0.034295876,0.044584636,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.041155048,0.044584636,0.041155048,0.01371835,0.041155048,0.12003556,0.14404267,0.09602845,0.044584636,0.034295876,0.041155048,0.044584636,0.058302987,0.106317215,0.106317215,0.08916927,0.106317215,0.17147937,0.24350071,0.23321195,0.1920569,0.16804978,0.19891608,0.31895164,0.39440256,0.36696586,0.36010668,0.45956472,0.71678376,0.65505123,0.5041494,0.37382504,0.33952916,0.4115505,0.58302987,0.66191036,0.66876954,0.607037,0.47328308,0.31552204,0.15433143,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.0034295875,0.01371835,0.0034295875,0.010288762,0.01371835,0.017147938,0.030866288,0.06859175,0.048014224,0.017147938,0.0,0.0,0.024007112,0.06859175,0.06859175,0.0274367,0.01371835,0.0274367,0.041155048,0.044584636,0.048014224,0.061732575,0.024007112,0.006859175,0.0,0.010288762,0.044584636,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.041155048,0.0274367,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.010288762,0.034295876,0.06859175,0.106317215,0.06859175,0.041155048,0.024007112,0.020577524,0.044584636,0.058302987,0.09602845,0.1097468,0.07545093,0.01371835,0.01371835,0.024007112,0.037725464,0.05144381,0.07545093,0.09945804,0.12346515,0.16804978,0.2194936,0.24350071,0.24350071,0.24350071,0.23664154,0.2469303,0.31895164,0.28465575,0.20234565,0.09602845,0.01371835,0.0,0.0,0.010288762,0.020577524,0.034295876,0.044584636,0.16804978,0.4081209,0.6036074,0.64133286,0.45613512,0.116605975,0.030866288,0.041155048,0.23664154,0.94656616,1.6667795,1.937717,1.6187652,1.0048691,0.8093826,0.9294182,1.2449403,1.6530612,2.0028791,2.0749004,2.0268862,2.1434922,2.2841053,2.3389788,2.2292318,2.0097382,1.961724,1.9823016,2.0063086,2.0303159,1.9068506,1.5844694,1.2723769,1.1043272,1.1283343,1.1523414,0.9294182,0.8265306,0.94999576,1.1454822,0.90198153,0.66533995,0.8848336,1.4987297,1.937717,1.8519772,1.6667795,1.4095604,1.1214751,0.84024894,1.3512574,1.8005334,2.3801336,3.1140654,3.8445675,3.9303071,3.6044965,3.1895163,2.8877127,2.7779658,2.7162333,2.435007,2.2086544,2.1812177,2.3664153,2.3424082,2.1983654,2.393852,2.5001693,1.2037852,0.5590228,0.26064864,0.15433143,0.1371835,0.1371835,0.09945804,0.072021335,0.048014224,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.024007112,0.12346515,0.31895164,0.6241849,1.1420527,1.7696671,2.1983654,1.7456601,1.4507155,1.4438564,1.5810398,1.4335675,1.9342873,2.061182,2.1091962,2.2258022,2.3972816,1.4815818,1.0768905,0.9431366,1.0151579,1.4198492,2.469303,4.0949273,6.1046658,8.275595,10.374502,11.561139,11.828648,11.454823,10.734609,9.962952,9.853205,9.753747,9.369633,8.9100685,9.095266,9.4862385,9.921797,10.782623,12.240198,14.267084,15.951012,15.412566,14.277372,13.478279,13.258785,13.821238,14.016724,14.003006,13.63604,12.449403,10.5597,8.951223,8.597976,9.469091,10.542552,11.64345,11.780633,10.295622,7.613684,5.2335505,4.098357,3.6147852,3.4604537,3.1517909,2.0303159,1.786815,1.4027013,1.1660597,1.1900668,1.4335675,1.3855534,1.0254467,0.83681935,0.8779744,0.7922347,0.58645946,0.83681935,1.2380811,1.4335675,1.0082988,0.6276145,0.58988905,0.4046913,0.14061308,0.39783216,0.50757897,0.4424168,0.22978236,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.07545093,0.07545093,0.048014224,0.041155048,0.07888051,0.15090185,0.3841138,0.37039545,0.2469303,0.12689474,0.09259886,0.90884066,1.5913286,2.1640697,2.469303,2.1503513,1.0288762,1.039165,1.2723769,1.3169615,1.2826657,1.2826657,1.4918705,2.218943,3.4295874,4.7602673,4.5784993,3.9097297,3.6113555,4.098357,5.3570156,6.5162163,7.390761,7.98408,8.30646,8.3922,8.735159,9.688584,10.683165,11.784062,13.687484,19.716698,26.277498,31.531628,34.01122,32.608517,27.467566,22.429502,18.272842,14.970149,11.674315,9.071259,7.490219,7.140401,7.473071,7.157549,6.6053853,6.012067,5.754848,5.830299,5.830299,4.839148,4.0880685,3.1689389,2.253239,2.1057668,2.1194851,1.7559488,1.3169615,0.9774324,0.7922347,0.6824879,0.6001778,0.5453044,0.51100856,0.47328308,0.45956472,0.548734,0.8676856,1.3169615,1.5707511,1.5090185,1.3032433,1.0597426,0.9602845,1.2655178,1.6324836,1.786815,1.6770682,1.3443983,0.9294182,0.6756287,0.47328308,0.34638834,0.29494452,0.31895164,0.3806842,0.48014224,0.58988905,0.6824879,0.7339317,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.037725464,0.044584636,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.010288762,0.030866288,0.06516216,0.1097468,0.16462019,0.2194936,0.25378948,0.29837412,0.35324752,0.39097297,0.40126175,0.4081209,0.4115505,0.3841138,0.2709374,0.14061308,0.072021335,0.034295876,0.024007112,0.044584636,0.041155048,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.006859175,0.0034295875,0.017147938,0.0274367,0.034295876,0.0274367,0.010288762,0.017147938,0.01371835,0.010288762,0.020577524,0.058302987,0.08573969,0.13375391,0.1920569,0.2503599,0.29151493,0.24007112,0.20577525,0.19548649,0.21263443,0.2469303,0.23321195,0.21263443,0.2709374,0.4081209,0.5590228,0.45956472,0.36353627,0.28808534,0.25721905,0.3018037,0.37382504,0.39440256,0.3806842,0.34295875,0.2777966,0.216064,0.15433143,0.08916927,0.030866288,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.0034295875,0.020577524,0.020577524,0.024007112,0.041155048,0.0548734,0.072021335,0.0548734,0.030866288,0.010288762,0.0,0.024007112,0.06859175,0.09602845,0.1097468,0.1371835,0.2194936,0.28465575,0.29494452,0.24007112,0.14747226,0.15776102,0.16119061,0.15433143,0.12346515,0.034295876,0.020577524,0.006859175,0.0,0.0034295875,0.01371835,0.030866288,0.020577524,0.006859175,0.0034295875,0.0034295875,0.006859175,0.006859175,0.0034295875,0.0034295875,0.0034295875,0.05144381,0.14404267,0.29494452,0.4355576,0.4046913,0.3841138,0.432128,0.5041494,0.51100856,0.3018037,0.20577525,0.15090185,0.116605975,0.10288762,0.106317215,0.07888051,0.058302987,0.041155048,0.034295876,0.05144381,0.12003556,0.16804978,0.18519773,0.18862732,0.22292319,0.23664154,0.20234565,0.17147937,0.17833854,0.23321195,0.2503599,0.25721905,0.2503599,0.25378948,0.30866286,0.29151493,0.25721905,0.20234565,0.13032432,0.061732575,0.05144381,0.034295876,0.024007112,0.020577524,0.020577524,0.0548734,0.09259886,0.12003556,0.12689474,0.09259886,0.05144381,0.15090185,0.82996017,1.7353712,1.7525192,1.1626302,0.7407909,0.48700142,0.42869842,0.61389613,0.939707,1.2312219,1.3924125,1.529596,1.9514352,2.0508933,2.277246,2.486451,2.503599,2.1297739,1.704505,1.4164196,1.2277923,1.1008976,1.0151579,0.7956643,0.77165717,0.8162418,0.864256,0.89855194,0.7956643,0.58302987,0.5693115,0.7339317,0.75450927,0.64476246,0.7305021,1.155771,1.9239986,2.901431,2.503599,1.8897027,1.4644338,1.4472859,1.8416885,2.1674993,2.8328393,3.5873485,4.1189346,4.040054,3.5873485,3.4227283,3.3438478,3.2375305,3.069481,3.0489032,2.7985435,2.7642474,2.8739944,2.5481834,1.8588364,1.5810398,1.6187652,1.670209,1.2175035,0.7956643,0.4355576,0.22292319,0.16804978,0.19891608,0.20920484,0.18176813,0.116605975,0.048014224,0.0274367,0.044584636,0.06516216,0.07888051,0.08573969,0.08573969,0.06516216,0.030866288,0.006859175,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0274367,0.024007112,0.030866288,0.020577524,0.0,0.0,0.010288762,0.01371835,0.006859175,0.0,0.0,0.01371835,0.01371835,0.0274367,0.05144381,0.048014224,0.020577524,0.0034295875,0.0,0.010288762,0.048014224,0.23321195,0.8745448,2.428148,4.3761535,5.212973,4.4104495,3.525616,3.0626216,2.9563043,2.6064866,1.9239986,1.4267083,1.2346514,1.3786942,1.7730967,1.4541451,1.2449403,1.1283343,1.0871792,1.0906088,1.728512,2.651071,3.9337368,5.579939,7.5450926,9.860064,11.578287,12.367092,12.281353,11.746337,11.283342,11.375941,11.077567,10.182446,9.205012,8.951223,9.263316,9.897789,10.882081,12.507706,13.872682,14.30481,14.174485,13.656617,12.723769,12.747777,12.850664,13.073587,13.29994,13.2690735,11.492548,10.683165,10.607714,10.926665,11.190743,11.273054,10.39508,9.355915,8.399059,7.1987042,6.15268,5.07236,3.998899,2.976882,2.07833,1.7662375,1.4781522,1.155771,0.9328478,1.1283343,1.1763484,1.0700313,0.96714365,0.8505377,0.5007198,0.4389872,0.5007198,0.61389613,0.67219913,0.5178677,0.23664154,0.17147937,0.29151493,0.5796003,1.0323058,1.2209331,0.88826317,0.6276145,0.5521636,0.31895164,0.072021335,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.037725464,0.041155048,0.044584636,0.061732575,0.116605975,0.2503599,0.37039545,0.32238123,0.1371835,0.030866288,0.32238123,1.0082988,1.8073926,2.3149714,2.0165975,1.4610043,1.5981878,1.7147937,1.5638919,1.3786942,1.5741806,1.9720128,2.5721905,3.5153272,5.0895076,6.3035817,6.495639,6.427047,6.625963,7.394191,7.881192,7.949784,8.011517,8.255017,8.673427,9.22902,10.48082,12.490558,15.505165,19.949911,25.032558,29.106909,31.706535,32.471333,31.154373,29.35727,28.235794,27.121178,25.121729,21.133118,16.060759,12.161317,9.839486,8.97866,8.913498,9.115844,8.488229,7.857185,7.596536,7.6342616,6.8626046,6.2898636,5.597087,4.8014226,4.2526884,4.040054,3.4021509,2.6613598,2.0268862,1.5981878,1.155771,0.9774324,0.89855194,0.84024894,0.8025235,0.8196714,0.8196714,0.980862,1.2689474,1.4369972,1.3066728,1.1420527,0.89169276,0.65505123,0.65505123,1.0220171,1.4129901,1.605047,1.5158776,1.1866373,0.84367853,0.5761707,0.4115505,0.35324752,0.37039545,0.5658819,0.77851635,0.9568549,1.08032,1.1489118,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.017147938,0.01371835,0.01371835,0.0274367,0.0274367,0.0274367,0.017147938,0.0,0.0,0.0,0.0,0.01371835,0.041155048,0.0548734,0.0548734,0.034295876,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.030866288,0.041155048,0.058302987,0.07888051,0.106317215,0.14061308,0.17490897,0.20234565,0.23321195,0.25378948,0.2469303,0.18176813,0.10288762,0.06859175,0.05144381,0.044584636,0.044584636,0.037725464,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.0274367,0.058302987,0.1097468,0.15776102,0.18862732,0.19548649,0.14061308,0.12689474,0.13375391,0.15090185,0.15433143,0.14061308,0.15090185,0.19891608,0.26407823,0.29837412,0.24007112,0.20920484,0.18176813,0.15433143,0.14747226,0.17490897,0.18862732,0.19548649,0.20577525,0.22978236,0.22292319,0.20920484,0.17833854,0.13375391,0.08916927,0.037725464,0.010288762,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.024007112,0.017147938,0.020577524,0.01371835,0.01371835,0.030866288,0.05144381,0.058302987,0.044584636,0.030866288,0.024007112,0.017147938,0.020577524,0.037725464,0.05144381,0.061732575,0.07545093,0.22635277,0.2777966,0.22635277,0.116605975,0.06859175,0.07545093,0.07888051,0.07545093,0.061732575,0.01371835,0.006859175,0.020577524,0.030866288,0.041155048,0.05144381,0.061732575,0.058302987,0.044584636,0.034295876,0.017147938,0.017147938,0.01371835,0.01371835,0.037725464,0.12003556,0.30523327,0.5007198,0.64133286,0.6927767,0.65162164,0.59674823,0.5418748,0.47671264,0.3806842,0.22292319,0.17833854,0.15433143,0.14747226,0.15776102,0.18519773,0.1920569,0.15090185,0.12346515,0.15090185,0.25378948,0.39783216,0.432128,0.4115505,0.3806842,0.34981793,0.32581082,0.32581082,0.34981793,0.4046913,0.4938606,0.490431,0.432128,0.36696586,0.32924038,0.33266997,0.31895164,0.35324752,0.39097297,0.39440256,0.33266997,0.2194936,0.12003556,0.0548734,0.0274367,0.034295876,0.044584636,0.048014224,0.048014224,0.0548734,0.0548734,0.06859175,0.18862732,0.52815646,0.90198153,0.8093826,0.44927597,0.21263443,0.1371835,0.26064864,0.6276145,1.0014396,1.2586586,1.2998136,1.3306799,1.8588364,2.1915064,2.4590142,2.5893385,2.4967396,2.0886188,1.5604624,1.0460242,0.72021335,0.6001778,0.5418748,0.51100856,0.5418748,0.61389613,0.70649505,0.7922347,0.78537554,0.59674823,0.5144381,0.5693115,0.5453044,0.5521636,0.7888051,1.4267083,2.2258022,2.5310357,2.4041407,2.3252604,2.2292318,2.3389788,3.1346428,3.707384,4.2698364,4.6848164,4.8322887,4.602506,4.016047,3.765687,3.5118976,3.07634,2.4384367,2.6819375,2.3629858,2.0920484,2.054323,1.9891608,1.9342873,1.9411465,1.8382589,1.5844694,1.2758065,1.0700313,0.97057325,0.78194594,0.5144381,0.4046913,0.42183927,0.42869842,0.36696586,0.2469303,0.15090185,0.13032432,0.16119061,0.20920484,0.24007112,0.216064,0.14747226,0.082310095,0.037725464,0.017147938,0.010288762,0.020577524,0.01371835,0.010288762,0.006859175,0.0,0.0,0.01371835,0.024007112,0.024007112,0.020577524,0.0274367,0.041155048,0.0274367,0.006859175,0.0274367,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.037725464,0.05144381,0.030866288,0.01371835,0.010288762,0.010288762,0.020577524,0.09602845,0.6927767,2.1091962,4.040054,5.5833683,6.3378778,5.9571934,5.3501563,4.787704,3.9165888,2.901431,2.5241764,2.2635276,2.0234566,2.1023371,2.218943,2.4247184,2.4795918,2.311542,2.0234566,1.8725548,1.9411465,2.4761622,3.566771,5.1512403,8.001227,10.268185,11.8115,12.644889,12.915827,12.891819,12.943263,12.555719,11.55771,10.120712,9.126132,9.112414,9.287323,9.534253,10.422516,11.513125,12.247057,12.418536,12.171606,12.010415,12.003556,11.869802,12.133881,12.895248,13.848674,13.509145,13.173045,12.703192,12.411677,13.063298,14.188204,13.238208,11.430815,9.671436,8.532814,7.2432885,6.0703697,5.0106273,4.0709205,3.2718265,2.6853669,2.2395205,1.7936742,1.3855534,1.2449403,1.1660597,1.0871792,1.0700313,1.0220171,0.70306545,0.5590228,0.48700142,0.48700142,0.47671264,0.29494452,0.6036074,0.72707254,0.6344737,0.58645946,1.1077567,1.196926,0.9534253,0.7339317,0.6276145,0.45956472,0.13375391,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.010288762,0.0274367,0.044584636,0.061732575,0.08916927,0.1920569,0.28465575,0.25378948,0.11317638,0.006859175,0.08573969,0.490431,1.1489118,1.7388009,1.6804979,1.529596,1.6804979,1.8348293,1.8073926,1.5124481,1.9857311,2.7059445,3.6353626,4.8597255,6.5813785,8.56368,9.366203,9.335337,8.923786,8.700864,8.790032,8.766026,8.903209,9.201583,9.403929,9.770895,11.149589,13.934414,18.008764,22.741594,26.130028,27.584171,27.357819,25.886526,23.78076,23.328054,23.76704,24.230036,23.996824,22.491234,19.147387,15.786391,12.730629,10.398509,9.3079,10.4533825,10.63858,10.628291,10.597425,10.110424,8.443645,7.4765005,6.7631464,6.029215,5.1855364,4.4413157,3.5804894,2.7813954,2.1091962,1.5261664,1.2655178,1.0494537,0.9259886,0.90884066,0.96714365,1.0666018,1.155771,1.313532,1.5055889,1.587899,1.3443983,1.1146159,0.8745448,0.64476246,0.5212973,0.7339317,1.0734608,1.3169615,1.3649758,1.2517995,1.0597426,0.8162418,0.5761707,0.4115505,0.41840968,0.71678376,1.0220171,1.1866373,1.1832076,1.1317638,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.017147938,0.020577524,0.0274367,0.05144381,0.030866288,0.0274367,0.017147938,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.037725464,0.05144381,0.037725464,0.030866288,0.034295876,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.020577524,0.034295876,0.044584636,0.058302987,0.061732575,0.08573969,0.10288762,0.10288762,0.07545093,0.048014224,0.037725464,0.037725464,0.034295876,0.0274367,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0274367,0.06859175,0.09945804,0.106317215,0.10288762,0.07545093,0.06859175,0.07545093,0.082310095,0.07545093,0.082310095,0.106317215,0.12689474,0.13032432,0.12346515,0.10288762,0.09945804,0.09602845,0.08573969,0.072021335,0.14061308,0.20234565,0.25378948,0.29494452,0.33266997,0.3018037,0.2777966,0.24350071,0.18519773,0.09945804,0.034295876,0.006859175,0.0034295875,0.006859175,0.006859175,0.0,0.010288762,0.034295876,0.061732575,0.06859175,0.05144381,0.034295876,0.024007112,0.030866288,0.041155048,0.034295876,0.030866288,0.030866288,0.030866288,0.030866288,0.024007112,0.017147938,0.01371835,0.017147938,0.020577524,0.12003556,0.14061308,0.082310095,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.020577524,0.034295876,0.037725464,0.041155048,0.05144381,0.072021335,0.1097468,0.15090185,0.17833854,0.15776102,0.20234565,0.2777966,0.31552204,0.32238123,0.39440256,0.53844523,0.764798,0.9774324,1.0151579,0.6379033,0.48700142,0.36696586,0.26407823,0.18176813,0.15433143,0.17833854,0.2469303,0.32581082,0.39097297,0.42869842,0.41840968,0.32581082,0.26750782,0.28122616,0.34981793,0.4424168,0.5144381,0.5178677,0.4629943,0.40126175,0.41840968,0.5693115,0.7990939,0.980862,0.90884066,0.77851635,0.6344737,0.5007198,0.39097297,0.30866286,0.33609957,0.432128,0.53501564,0.5624523,0.42869842,0.2777966,0.16462019,0.10288762,0.09945804,0.15090185,0.19548649,0.25721905,0.31552204,0.34981793,0.33609957,0.25721905,0.25721905,0.20920484,0.106317215,0.05144381,0.0548734,0.048014224,0.061732575,0.17833854,0.53844523,0.8745448,1.097468,1.138623,1.214074,1.8279701,2.3801336,2.6922262,2.7230926,2.4624438,1.9342873,1.4815818,0.864256,0.44927597,0.32581082,0.31895164,0.39440256,0.41840968,0.45270553,0.52815646,0.64133286,0.77165717,0.8196714,0.8676856,0.90198153,0.8162418,0.6756287,0.7888051,1.2998136,1.978872,2.2292318,2.6476414,3.069481,3.292404,3.5187566,4.341858,5.2335505,5.686256,5.528495,4.98662,4.6745276,4.187526,3.940596,3.6627994,3.1826572,2.4384367,2.1812177,1.704505,1.3478279,1.2655178,1.4232788,1.6290541,1.728512,1.6359133,1.430138,1.3306799,1.4678634,1.7490896,1.8073926,1.5604624,1.2106444,0.90541106,0.77165717,0.7099246,0.64476246,0.5521636,0.5658819,0.61046654,0.5453044,0.4046913,0.37039545,0.28465575,0.20920484,0.14404267,0.08916927,0.05144381,0.041155048,0.0274367,0.020577524,0.01371835,0.0,0.0,0.010288762,0.024007112,0.030866288,0.0274367,0.034295876,0.034295876,0.030866288,0.0274367,0.044584636,0.0274367,0.0274367,0.020577524,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.041155048,0.0274367,0.0274367,0.041155048,0.06859175,0.11317638,0.082310095,0.38754338,1.0837497,2.095478,3.2032347,4.3452873,4.4516044,4.184097,3.940596,3.8857226,5.4633327,5.504488,4.9077396,4.3349986,4.2389703,4.5784993,4.448175,4.0674906,3.7005248,3.642222,3.3952916,2.8465576,2.6373527,3.000889,3.765687,5.888602,7.966932,10.007536,11.838936,13.111313,13.54687,13.6086035,13.275933,12.476839,11.094715,10.14129,9.633711,9.1981535,8.89635,9.239308,9.6988735,10.175586,10.4533825,10.696883,11.4754,12.171606,11.948683,12.113303,13.111313,14.531162,15.165636,14.668345,13.612033,12.956982,14.057879,16.108772,16.331696,15.097044,13.090735,11.327928,9.4862385,7.798882,6.166398,4.7191124,3.8137012,3.3712845,3.0283258,2.651071,2.201795,1.728512,1.4815818,1.3752645,1.3855534,1.3924125,1.196926,0.91227025,0.9431366,1.0494537,1.0185875,0.6927767,0.8745448,1.2037852,1.0940384,0.70306545,0.9362774,0.881404,0.7305021,0.6207553,0.548734,0.3806842,0.1371835,0.058302987,0.034295876,0.010288762,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.037725464,0.044584636,0.17833854,0.28465575,0.2469303,0.09259886,0.006859175,0.017147938,0.15433143,0.5144381,0.9945804,1.2963841,1.2860953,1.3238207,1.4232788,1.5021594,1.4095604,2.2292318,3.450165,4.938606,6.5882373,8.323608,10.168727,10.875222,10.535692,9.56512,8.694004,8.868914,9.414218,10.199594,10.799771,10.501397,10.189304,11.008976,13.275933,16.722668,20.488356,22.10712,21.719578,19.929333,17.504614,15.3817,15.182784,15.584045,16.064188,16.338554,16.338554,15.343974,13.687484,11.609154,9.633711,8.549961,9.938945,10.786053,11.286773,11.345076,10.573419,8.903209,8.06296,7.822889,7.7783046,7.3701835,6.1766872,4.6573796,3.3884325,2.750529,2.952875,3.210094,2.8808534,2.3149714,1.8245405,1.7182233,1.937717,2.3629858,2.8259802,3.0523329,2.6476414,2.1297739,1.670209,1.2517995,0.8745448,0.5418748,0.6207553,0.8093826,0.9774324,1.0666018,1.0940384,1.0528834,0.8711152,0.6344737,0.44584638,0.4424168,0.70649505,1.0048691,1.1043272,0.99801,0.88826317,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.030866288,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.08916927,0.09945804,0.037725464,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.0274367,0.024007112,0.024007112,0.0034295875,0.010288762,0.024007112,0.037725464,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.041155048,0.0548734,0.05144381,0.061732575,0.061732575,0.0548734,0.044584636,0.034295876,0.024007112,0.034295876,0.05144381,0.058302987,0.0548734,0.06859175,0.058302987,0.048014224,0.05144381,0.06859175,0.09602845,0.22292319,0.36696586,0.490431,0.5658819,0.5727411,0.4698535,0.39440256,0.31552204,0.2194936,0.09945804,0.044584636,0.020577524,0.020577524,0.030866288,0.0274367,0.01371835,0.017147938,0.048014224,0.09259886,0.09945804,0.082310095,0.061732575,0.048014224,0.041155048,0.0274367,0.017147938,0.020577524,0.024007112,0.024007112,0.0274367,0.0274367,0.020577524,0.01371835,0.017147938,0.0274367,0.006859175,0.0034295875,0.006859175,0.01371835,0.020577524,0.010288762,0.006859175,0.010288762,0.020577524,0.037725464,0.06516216,0.06516216,0.048014224,0.034295876,0.048014224,0.09602845,0.17833854,0.26407823,0.32238123,0.29494452,0.3806842,0.53844523,0.61389613,0.58302987,0.5693115,0.5418748,0.6859175,0.9774324,1.097468,0.42183927,0.22292319,0.17147937,0.19548649,0.26064864,0.33952916,0.36696586,0.490431,0.6241849,0.71678376,0.7339317,0.66191036,0.52815646,0.42183927,0.36696586,0.29494452,0.2503599,0.40126175,0.48700142,0.4424168,0.42869842,0.5590228,0.84024894,1.2175035,1.4747226,1.2037852,0.97400284,0.8025235,0.64476246,0.4938606,0.37382504,0.4081209,0.48014224,0.53158605,0.4972902,0.28465575,0.20234565,0.16462019,0.18176813,0.25378948,0.37382504,0.48357183,0.64133286,0.7922347,0.8848336,0.85739684,0.65848076,0.490431,0.33952916,0.19891608,0.10288762,0.06859175,0.044584636,0.030866288,0.082310095,0.29837412,0.5521636,0.72707254,0.83338976,1.0597426,1.7696671,2.5584722,2.9220085,2.860276,2.4212887,1.7113642,1.3512574,0.77851635,0.34981793,0.18519773,0.17490897,0.20920484,0.24350071,0.2777966,0.32924038,0.4046913,0.5727411,0.881404,1.1694894,1.313532,1.1934965,0.84024894,0.8196714,1.039165,1.5261664,2.4247184,3.2649672,3.7725463,4.108646,4.48933,5.171818,6.1458206,6.5162163,5.9400454,4.856296,4.4996185,4.197815,4.012617,3.8377085,3.5839188,3.1689389,1.9548649,1.3101025,1.0563129,1.0254467,1.0528834,0.9911508,0.9877212,1.2175035,1.7182233,2.411,2.5584722,3.3061223,3.8891523,3.865145,3.1140654,1.9685832,1.3855534,1.2517995,1.3684053,1.4472859,1.4953002,1.3066728,0.90884066,0.4972902,0.45956472,0.4355576,0.4081209,0.3566771,0.28122616,0.18862732,0.12346515,0.082310095,0.044584636,0.01371835,0.0034295875,0.0034295875,0.006859175,0.020577524,0.037725464,0.041155048,0.05144381,0.030866288,0.030866288,0.048014224,0.041155048,0.030866288,0.048014224,0.044584636,0.010288762,0.0034295875,0.0,0.010288762,0.017147938,0.020577524,0.034295876,0.030866288,0.048014224,0.08573969,0.14404267,0.22978236,0.17833854,0.18862732,0.18862732,0.14404267,0.034295876,0.14061308,0.34638834,0.607037,1.1660597,2.534465,6.9654922,7.291303,6.4098988,5.892031,5.9640527,6.1046658,5.3501563,4.4687524,4.0091877,4.314421,4.4584637,3.8342788,3.2512488,3.0111778,2.8980014,3.5839188,5.0826488,7.291303,9.788043,11.849225,12.686044,13.090735,13.138749,12.754636,11.736049,11.338216,10.446524,9.56512,9.108984,9.424506,8.999237,8.848335,9.098696,9.798331,10.923236,12.442543,12.576297,12.902108,13.992717,15.429714,16.146498,15.364552,14.044161,13.166186,13.7526455,15.367981,17.000465,17.55263,16.606062,14.445422,12.336226,10.271614,7.7440085,5.130663,3.690236,3.3712845,3.199805,3.0077481,2.6819375,2.1503513,1.8725548,1.7730967,1.7147937,1.6256244,1.4815818,1.1900668,1.4267083,1.6770682,1.6359133,1.2209331,0.77165717,1.1249046,1.2483698,0.9431366,0.8265306,0.64476246,0.5041494,0.48357183,0.47328308,0.18176813,0.106317215,0.15776102,0.15090185,0.0548734,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.18862732,0.37039545,0.32581082,0.09945804,0.01371835,0.006859175,0.024007112,0.106317215,0.33609957,0.83681935,0.823101,0.764798,0.7305021,0.805953,1.0940384,2.2978237,3.882293,5.6793966,7.514226,9.218731,10.868362,11.629731,11.513125,10.844356,10.254466,10.6488695,11.38623,12.21619,12.586586,11.619442,10.545981,10.425946,11.201033,12.71691,14.726648,14.87755,13.773223,12.05843,10.340206,9.1981535,8.851766,8.570539,8.200144,7.7131424,7.1849856,7.274155,7.116394,6.8557453,6.6465406,6.6636887,7.740579,8.676856,9.1981535,9.191295,8.724871,8.158989,7.936065,8.529384,9.685155,10.401938,9.225591,6.9860697,5.099797,4.5510626,5.892031,6.7048435,6.385892,5.3673043,4.2046742,3.5839188,3.7451096,4.386442,5.0826488,5.254128,4.170378,3.175798,2.3389788,1.6153357,0.9877212,0.48357183,0.53501564,0.607037,0.6859175,0.7510797,0.8025235,0.8265306,0.72707254,0.58988905,0.48700142,0.48357183,0.6207553,0.823101,0.881404,0.8025235,0.7922347,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.17490897,0.3806842,0.16119061,0.061732575,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.030866288,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.020577524,0.044584636,0.034295876,0.041155048,0.058302987,0.082310095,0.106317215,0.16804978,0.37382504,0.6241849,0.82996017,0.91569984,0.78194594,0.64819205,0.53158605,0.42869842,0.31895164,0.18519773,0.106317215,0.082310095,0.08916927,0.07545093,0.06516216,0.041155048,0.024007112,0.01371835,0.01371835,0.01371835,0.01371835,0.020577524,0.0274367,0.01371835,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.010288762,0.034295876,0.06859175,0.106317215,0.044584636,0.030866288,0.030866288,0.037725464,0.061732575,0.1097468,0.15776102,0.17147937,0.15776102,0.18176813,0.23321195,0.25378948,0.22978236,0.16119061,0.07545093,0.05144381,0.044584636,0.05144381,0.06859175,0.106317215,0.106317215,0.09602845,0.09602845,0.12689474,0.21263443,0.29837412,0.44927597,0.6310441,0.8162418,0.9602845,0.864256,0.7922347,0.7579388,0.7476501,0.7476501,0.72364295,0.6790583,0.5761707,0.41840968,0.26064864,0.22292319,0.37725464,0.47671264,0.490431,0.6241849,0.78537554,0.88826317,0.9294182,0.9328478,0.94656616,0.9842916,0.96371406,0.8848336,0.8128122,0.8848336,0.72707254,0.5212973,0.31895164,0.17490897,0.1371835,0.17490897,0.23664154,0.34638834,0.4938606,0.64133286,0.7990939,1.0494537,1.2998136,1.4678634,1.4815818,1.2586586,1.0323058,0.77508676,0.50757897,0.274367,0.15090185,0.11317638,0.09602845,0.09259886,0.15090185,0.23664154,0.31552204,0.48357183,0.84367853,1.4644338,2.6716487,3.0386145,2.819121,2.2738166,1.6633499,1.0288762,0.58645946,0.31895164,0.17490897,0.07545093,0.15090185,0.18519773,0.19891608,0.19891608,0.19891608,0.16119061,0.18862732,0.32238123,0.5212973,0.65505123,0.64476246,1.0906088,1.5604624,1.961724,2.5481834,3.2306714,3.642222,4.0057583,4.537344,5.4153185,5.977771,6.0737996,5.7068334,5.2472687,5.4153185,5.271276,4.822,4.166949,3.532475,3.2649672,2.277246,1.5638919,1.1043272,0.8196714,0.5658819,1.039165,1.371835,2.3835633,4.2766957,6.6225333,5.4153185,6.831738,8.207003,8.165848,6.6533995,4.0537724,2.651071,2.3046827,2.644212,3.083199,2.8877127,1.7319417,0.75450927,0.38754338,0.34981793,0.47328308,0.61389613,0.69963586,0.6790583,0.5178677,0.3841138,0.26064864,0.13032432,0.0274367,0.01371835,0.01371835,0.041155048,0.061732575,0.0548734,0.030866288,0.06859175,0.048014224,0.017147938,0.0034295875,0.01371835,0.06516216,0.041155048,0.010288762,0.0034295875,0.01371835,0.0034295875,0.010288762,0.020577524,0.034295876,0.044584636,0.082310095,0.1097468,0.12346515,0.12003556,0.106317215,0.15433143,0.23321195,0.18862732,0.06859175,0.106317215,0.34981793,0.6036074,0.84367853,1.08032,1.371835,1.5193073,1.5570327,1.5741806,1.6804979,1.9823016,1.1283343,1.3649758,1.7319417,1.7388009,1.371835,0.8745448,0.94999576,1.0906088,1.08032,1.0082988,1.313532,2.386993,4.139512,6.3207297,8.529384,10.31277,11.674315,12.466551,12.590015,11.993267,11.2593355,10.6488695,10.017825,9.740028,10.679735,9.729739,8.831187,8.546532,8.944365,9.626852,10.628291,11.859513,13.337666,14.942713,16.417435,17.261114,17.408587,16.681513,15.206791,13.413116,12.936404,13.87954,14.63062,14.459141,13.519434,12.579727,12.325937,10.628291,7.4113383,4.65395,2.9563043,2.1469216,1.8313997,1.7353712,1.7250825,1.7010754,1.6496316,1.4164196,1.0425946,0.7613684,0.8128122,0.90541106,0.9294182,0.8162418,0.548734,0.59674823,0.59331864,0.6344737,0.7888051,1.0837497,0.8162418,0.7373613,0.6276145,0.40126175,0.12346515,0.12346515,0.37039545,0.4046913,0.17147937,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.216064,0.34981793,0.31895164,0.15090185,0.01371835,0.01371835,0.006859175,0.006859175,0.030866288,0.09259886,0.274367,0.4115505,0.48357183,0.5796003,0.8848336,2.4590142,3.6044965,4.7259717,6.1321025,8.011517,11.317638,14.479718,17.055338,18.811287,19.713268,19.593233,18.097933,16.05733,14.003006,12.147599,11.108434,10.840926,10.834066,10.686595,10.100135,9.187865,8.23444,7.5690994,7.1952744,6.8043017,6.3893213,5.9297566,5.312431,4.4859004,3.450165,3.1689389,3.2546785,3.4124396,3.4878905,3.4638834,4.8425775,5.4633327,5.888602,6.3310184,6.636252,6.7357097,6.4579134,7.239859,9.170717,11.002116,10.683165,8.8929205,7.4456344,7.1849856,7.98065,8.958082,9.31133,9.030104,8.176137,6.8797526,6.368744,6.3035817,6.245279,5.7925735,4.6093655,3.0077481,1.7662375,0.8745448,0.34638834,0.21263443,0.32238123,0.4046913,0.47328308,0.53501564,0.59674823,0.66876954,0.66876954,0.6379033,0.6173257,0.64133286,0.7510797,0.8779744,1.0082988,1.1592005,1.4027013,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.020577524,0.01371835,0.01371835,0.061732575,0.14061308,0.18862732,0.19891608,0.2194936,0.24007112,0.13375391,0.0548734,0.06516216,0.12346515,0.16804978,0.14747226,0.09259886,0.030866288,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.010288762,0.006859175,0.024007112,0.041155048,0.058302987,0.082310095,0.14404267,0.25721905,0.36353627,0.44927597,0.52472687,0.53844523,0.5418748,0.5041494,0.42183927,0.33266997,0.2194936,0.11317638,0.06516216,0.07545093,0.09945804,0.1371835,0.14404267,0.106317215,0.048014224,0.0274367,0.017147938,0.01371835,0.017147938,0.01371835,0.0034295875,0.01371835,0.006859175,0.0,0.0,0.0034295875,0.0034295875,0.010288762,0.01371835,0.01371835,0.0034295875,0.010288762,0.020577524,0.044584636,0.10288762,0.216064,0.33266997,0.16804978,0.041155048,0.06516216,0.14747226,0.20577525,0.18176813,0.14061308,0.14061308,0.24350071,0.3018037,0.29837412,0.2194936,0.1097468,0.05144381,0.06516216,0.11317638,0.1920569,0.26407823,0.24007112,0.1920569,0.16462019,0.15433143,0.16804978,0.21263443,0.29837412,0.4115505,0.4972902,0.52815646,0.51100856,0.45956472,0.44584638,0.44927597,0.45270553,0.4424168,0.39783216,0.34981793,0.31209245,0.31209245,0.4046913,0.61389613,0.8676856,0.91569984,0.7613684,0.65162164,0.65162164,0.70306545,0.72021335,0.7339317,0.8711152,0.939707,0.94999576,0.90884066,0.8471081,0.8128122,0.65162164,0.47671264,0.32924038,0.22635277,0.16119061,0.22635277,0.38754338,0.5796003,0.75450927,0.8711152,0.91569984,1.1283343,1.4232788,1.6907866,1.8108221,1.5810398,1.3032433,0.9842916,0.66191036,0.42183927,0.28808534,0.22635277,0.18862732,0.15776102,0.14061308,0.16804978,0.19891608,0.29151493,0.5178677,0.96371406,1.471293,2.1434922,2.4075704,2.1846473,1.8965619,1.5536032,1.214074,0.9259886,0.7373613,0.69963586,0.607037,0.53501564,0.4972902,0.5144381,0.61389613,0.9294182,1.2723769,1.6736387,2.095478,2.4247184,2.3561265,2.4795918,2.6990852,2.9734523,3.3061223,3.6456516,4.0880685,5.3227196,7.2432885,8.930646,9.513676,9.239308,8.834618,8.532814,8.090397,7.514226,6.773435,6.0052075,5.096367,3.7039545,2.959734,2.3595562,1.6324836,0.9294182,0.8196714,2.0989075,2.6407824,2.6579304,2.4590142,2.4487255,3.9131594,5.768566,7.4044795,8.450503,8.766026,7.610255,5.9400454,4.9180284,4.787704,4.863155,3.683377,2.287535,1.2037852,0.6344737,0.45956472,0.5521636,0.5693115,0.5555932,0.53158605,0.4698535,0.37382504,0.26064864,0.15433143,0.08573969,0.06516216,0.06516216,0.034295876,0.01371835,0.010288762,0.006859175,0.041155048,0.061732575,0.06516216,0.061732575,0.06516216,0.044584636,0.017147938,0.0034295875,0.0,0.0034295875,0.0,0.0034295875,0.020577524,0.048014224,0.06859175,0.09602845,0.26750782,0.37725464,0.36010668,0.29151493,0.24007112,0.17490897,0.11317638,0.07888051,0.09602845,0.21263443,0.36696586,0.47328308,0.6824879,1.3855534,2.3801336,3.2958336,3.789694,4.122364,5.1683884,5.1066556,4.9008803,4.6573796,4.9831905,6.989499,4.2423997,2.503599,1.5844694,1.155771,0.7510797,1.1454822,1.8588364,2.726522,3.6525106,4.6127954,6.5024977,8.40249,9.997248,11.159878,11.955542,12.377381,11.677745,10.923236,10.590566,10.583707,10.449953,10.690024,10.871792,10.72775,10.14129,9.551401,9.379922,9.836057,10.827208,11.962401,13.341095,14.342535,15.021593,15.319967,15.059319,14.095605,14.095605,14.184773,13.735497,12.397959,13.018714,13.413116,12.686044,10.63858,7.740579,6.2487082,5.0243454,3.9543142,3.0111778,2.2360911,1.762808,1.6942163,1.5947582,1.3032433,0.9328478,0.5418748,0.45613512,0.44584638,0.4355576,0.48700142,0.4972902,0.36353627,0.48700142,0.8265306,0.9259886,0.8505377,0.65505123,0.4424168,0.29837412,0.28122616,0.4972902,0.5624523,0.44584638,0.2709374,0.30523327,0.13032432,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.20577525,0.33266997,0.31552204,0.16804978,0.01371835,0.034295876,0.044584636,0.044584636,0.041155048,0.041155048,0.12003556,0.19891608,0.26750782,0.34638834,0.4938606,1.1626302,1.9823016,2.726522,3.4638834,4.5819287,6.5127864,8.48137,10.690024,13.090735,15.3817,16.108772,15.666355,13.896688,11.290202,8.995808,7.589677,6.948344,6.7871537,6.697984,6.169828,5.312431,4.6676683,4.2252517,3.9440255,3.7794054,3.8137012,4.0263357,4.197815,4.064061,3.3369887,3.1552205,2.9220085,2.9048605,3.07634,3.1106358,3.3472774,3.9371665,4.5167665,5.096367,6.077229,6.7219915,6.9620624,7.06838,7.2535777,7.6685576,8.268735,8.251588,7.7440085,6.948344,6.1492505,5.826869,5.6965446,5.5559316,5.3501563,5.161529,5.038064,5.363875,5.658819,5.3227196,3.6182148,2.6956558,2.2738166,1.8931323,1.3992717,0.922559,1.0597426,1.1660597,1.2175035,1.2517995,1.3512574,1.3272504,1.3032433,1.2483698,1.1694894,1.1180456,1.1592005,1.2175035,1.3409687,1.5638919,1.9171394,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.006859175,0.006859175,0.044584636,0.09259886,0.13032432,0.15776102,0.20920484,0.22635277,0.12346515,0.034295876,0.017147938,0.041155048,0.09259886,0.08916927,0.06859175,0.0548734,0.061732575,0.041155048,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.024007112,0.041155048,0.08573969,0.14404267,0.18862732,0.23321195,0.33609957,0.4081209,0.45270553,0.51100856,0.5590228,0.51100856,0.33952916,0.19548649,0.116605975,0.1097468,0.12346515,0.16804978,0.17833854,0.14404267,0.08573969,0.030866288,0.017147938,0.01371835,0.01371835,0.01371835,0.010288762,0.01371835,0.006859175,0.0,0.0034295875,0.010288762,0.0034295875,0.0034295875,0.006859175,0.0034295875,0.0,0.01371835,0.020577524,0.030866288,0.06516216,0.12346515,0.18862732,0.09945804,0.048014224,0.14061308,0.37039545,0.4389872,0.31209245,0.15090185,0.06859175,0.13032432,0.22292319,0.25378948,0.20920484,0.12003556,0.09259886,0.1097468,0.13032432,0.15433143,0.16804978,0.14747226,0.17490897,0.15776102,0.13032432,0.12003556,0.15090185,0.20577525,0.28465575,0.33952916,0.35324752,0.34295875,0.37039545,0.37039545,0.36353627,0.36353627,0.3566771,0.32924038,0.2709374,0.2503599,0.29837412,0.4046913,0.53501564,0.607037,0.5761707,0.48014224,0.45613512,0.53501564,0.67219913,0.8265306,0.96714365,1.0666018,0.99801,0.8711152,0.7373613,0.6241849,0.5555932,0.4389872,0.31209245,0.20234565,0.13375391,0.10288762,0.1920569,0.34981793,0.58302987,0.8848336,1.2517995,1.7182233,1.7216529,1.5810398,1.4541451,1.3443983,1.1763484,1.1797781,1.1249046,0.94656616,0.7682276,0.6344737,0.4698535,0.36010668,0.31209245,0.28465575,0.28122616,0.30523327,0.36353627,0.47671264,0.6756287,0.8779744,1.3032433,1.6804979,1.9582944,2.2909644,2.4418662,2.510458,2.5550427,2.5824795,2.5653315,2.411,2.3218307,2.3389788,2.486451,2.7779658,3.1792276,3.3541365,3.4913201,3.7108135,4.0674906,4.40702,4.7808447,5.1169443,5.377593,5.579939,5.802862,6.2418494,7.2432885,8.604835,9.571979,9.770895,9.962952,10.323058,10.751757,10.864933,10.14472,8.597976,7.1678376,6.169828,5.2781353,4.6676683,3.865145,2.6545007,1.5398848,1.7353712,2.3561265,2.5927682,2.469303,2.1126258,1.7422304,3.3952916,6.094377,8.748878,10.14472,8.944365,8.152129,7.6788464,7.438775,7.1198235,6.169828,4.3452873,2.7916842,1.6221949,0.8711152,0.48700142,0.35324752,0.4938606,0.6824879,0.85739684,1.1077567,1.2346514,0.7682276,0.35324752,0.20920484,0.14061308,0.10288762,0.044584636,0.010288762,0.017147938,0.0548734,0.09945804,0.14061308,0.11317638,0.048014224,0.048014224,0.06516216,0.058302987,0.034295876,0.0,0.0,0.0,0.0,0.01371835,0.048014224,0.09602845,0.14061308,0.2777966,0.35324752,0.30866286,0.17147937,0.12003556,0.07888051,0.0548734,0.05144381,0.06516216,0.11317638,0.2777966,0.41840968,0.69963586,1.6084765,2.7951138,3.4364467,3.549623,3.5976372,4.5030484,4.979761,5.137522,5.0277753,5.271276,7.0272245,5.874883,4.664239,3.6936657,2.867135,1.7216529,1.2586586,1.1249046,1.3169615,1.8519772,2.7711067,4.166949,5.9400454,7.9017696,9.692014,10.792912,11.581717,11.499407,11.201033,10.960961,10.659158,10.607714,10.666017,10.686595,10.587136,10.343636,9.750318,9.088407,8.944365,9.455373,10.347065,11.756626,12.6586075,13.275933,13.831526,14.54831,14.575747,14.260224,13.954991,13.474849,12.116733,12.418536,12.823228,12.919256,12.240198,10.261326,9.489669,8.776315,7.9257765,6.800872,5.329579,3.8137012,2.8156912,2.1160555,1.5707511,1.1214751,0.6962063,0.50757897,0.42183927,0.3841138,0.44584638,0.7682276,0.5693115,0.4389872,0.52472687,0.53844523,0.48357183,0.45956472,0.37382504,0.25721905,0.2469303,0.45613512,0.6241849,0.53844523,0.29494452,0.26407823,0.14404267,0.12346515,0.15776102,0.17147937,0.0548734,0.041155048,0.048014224,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.16462019,0.29837412,0.31209245,0.19548649,0.041155048,0.037725464,0.05144381,0.0548734,0.041155048,0.030866288,0.058302987,0.09602845,0.1371835,0.18519773,0.26064864,0.4629943,0.78537554,1.0700313,1.3169615,1.6804979,2.3081124,3.0626216,4.108646,5.429037,6.8283086,7.7440085,8.604835,9.177576,9.235879,8.573969,7.366754,6.077229,4.955754,4.105216,3.4776018,3.2203827,3.3026927,3.4227283,3.4295874,3.340418,3.4227283,3.532475,3.5461934,3.3747141,2.9631636,2.8911421,2.884283,2.6853669,2.3218307,2.1160555,2.2120838,2.651071,3.1620796,3.7176728,4.5339146,5.212973,5.579939,5.5833683,5.381023,5.3261495,5.6793966,5.8234396,5.5730796,5.0414934,4.619654,4.4859004,4.636802,4.9180284,5.188966,5.3261495,5.381023,5.638242,5.7891436,5.4084597,3.957744,3.3026927,3.3472774,3.2546785,2.6922262,1.8313997,1.670209,1.6804979,1.6530612,1.5673214,1.605047,1.6359133,1.5398848,1.3478279,1.1420527,1.0151579,1.039165,1.1008976,1.2277923,1.4438564,1.7422304,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.037725464,0.06516216,0.11317638,0.116605975,0.06859175,0.030866288,0.020577524,0.030866288,0.041155048,0.041155048,0.048014224,0.07545093,0.10288762,0.10288762,0.07545093,0.048014224,0.0274367,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0274367,0.06859175,0.10288762,0.12003556,0.17490897,0.37725464,0.4698535,0.5658819,0.7305021,0.86082643,0.7099246,0.45613512,0.2709374,0.18176813,0.16804978,0.16804978,0.22292319,0.23664154,0.20234565,0.12689474,0.030866288,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.010288762,0.006859175,0.006859175,0.006859175,0.01371835,0.006859175,0.006859175,0.0034295875,0.0,0.006859175,0.024007112,0.034295876,0.037725464,0.037725464,0.044584636,0.041155048,0.030866288,0.07545093,0.21263443,0.490431,0.5007198,0.31895164,0.1371835,0.048014224,0.06516216,0.20234565,0.26407823,0.22978236,0.14404267,0.12689474,0.12003556,0.106317215,0.08573969,0.06859175,0.061732575,0.116605975,0.106317215,0.082310095,0.082310095,0.1371835,0.24350071,0.2709374,0.26407823,0.25378948,0.274367,0.37382504,0.42183927,0.42869842,0.4115505,0.4115505,0.41840968,0.36353627,0.34295875,0.37039545,0.37382504,0.3566771,0.29151493,0.26750782,0.3566771,0.6001778,0.8676856,1.1317638,1.4164196,1.5604624,1.2243627,0.9774324,0.75450927,0.5521636,0.39097297,0.32238123,0.24350071,0.15776102,0.08916927,0.048014224,0.037725464,0.09602845,0.1920569,0.3566771,0.607037,0.9568549,1.4815818,1.4781522,1.2415106,0.96371406,0.72707254,0.61046654,0.7476501,0.90198153,0.97400284,0.9945804,0.9911508,1.0871792,1.039165,0.83338976,0.6927767,0.65505123,0.65162164,0.7888051,0.9877212,0.9842916,0.94999576,0.9911508,1.1900668,1.5570327,2.054323,2.4315774,2.7985435,3.1826572,3.57363,3.8960114,4.0229063,4.2115335,4.5339146,5.0449233,5.778855,6.2555676,6.2727156,6.0737996,5.874883,5.857735,6.2692857,6.7357097,7.1095347,7.332458,7.407909,7.459353,7.750868,8.2481575,8.772884,9.023245,9.006097,9.489669,10.179015,10.868362,11.4205265,10.998687,9.119273,7.1781263,5.9812007,5.7377,5.552502,4.856296,3.542764,2.294394,2.5653315,3.0317552,3.5153272,3.724532,3.82399,4.4413157,4.880303,6.355026,8.289313,9.760606,9.482809,8.477941,8.412778,8.577398,8.158989,6.2692857,4.8288593,3.3232703,1.961724,0.939707,0.4389872,0.23664154,0.3566771,0.6036074,0.9328478,1.4541451,2.1091962,1.6667795,1.0940384,0.77851635,0.52472687,0.28808534,0.12689474,0.044584636,0.030866288,0.072021335,0.12689474,0.32238123,0.31552204,0.106317215,0.041155048,0.058302987,0.058302987,0.034295876,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.082310095,0.12003556,0.17490897,0.21263443,0.19891608,0.1097468,0.06859175,0.048014224,0.044584636,0.05144381,0.06859175,0.08573969,0.24007112,0.4115505,0.70306545,1.4267083,2.3492675,2.860276,2.942586,2.8877127,3.3232703,3.99204,4.6676683,5.206114,5.7411294,6.697984,6.550512,6.0635104,5.3501563,4.506478,3.6182148,2.843128,1.5364552,0.8848336,1.214074,1.99602,2.7711067,4.0057583,5.9297566,8.114404,9.47595,10.4705305,10.988399,11.218181,11.214751,10.916377,10.840926,10.539123,10.189304,9.952662,9.983529,9.80862,9.355915,9.191295,9.534253,10.264755,11.30049,11.835506,12.164746,12.6586075,13.773223,15.011304,15.289101,15.107333,14.483148,12.956982,12.000127,11.852654,12.686044,13.852104,13.88297,13.560589,12.542002,11.002116,9.235879,7.6445503,6.1321025,4.7019644,3.316411,2.1263442,1.4472859,0.99801,0.7373613,0.59674823,0.52815646,0.51100856,0.83338976,0.6927767,0.4664239,0.33952916,0.29151493,0.2503599,0.33266997,0.34981793,0.274367,0.26064864,0.36696586,0.5144381,0.5007198,0.3566771,0.32238123,0.16804978,0.19548649,0.2709374,0.29494452,0.18862732,0.09602845,0.09945804,0.09259886,0.048014224,0.017147938,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.10288762,0.26064864,0.3566771,0.32924038,0.18176813,0.072021335,0.048014224,0.0548734,0.061732575,0.0548734,0.05144381,0.058302987,0.072021335,0.08916927,0.12003556,0.14404267,0.16119061,0.18862732,0.216064,0.22292319,0.216064,0.31209245,0.5212973,0.8162418,1.1249046,1.6633499,2.6167753,4.040054,5.593657,6.543653,6.7357097,6.001778,4.804852,3.525616,2.4555845,2.294394,2.609916,2.877424,2.8568463,2.5790498,2.4452958,2.3835633,2.311542,2.2086544,2.1400626,2.1915064,2.3492675,2.153781,1.646202,1.3752645,1.5090185,1.7902447,2.1846473,2.6407824,3.0900583,3.4878905,3.758828,3.8548563,3.758828,3.4878905,3.275256,3.0626216,2.7985435,2.5790498,2.644212,2.884283,3.2649672,3.765687,4.314421,4.770556,5.192395,5.662249,5.926327,5.7308407,4.835718,4.2835546,4.3178506,4.256118,3.7691166,2.8877127,2.3732746,2.2395205,2.1263442,1.9582944,1.9239986,2.0474637,2.061182,1.8382589,1.4610043,1.2003556,1.1900668,1.255229,1.3752645,1.5570327,1.8348293,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.010288762,0.0034295875,0.0034295875,0.010288762,0.020577524,0.01371835,0.010288762,0.017147938,0.0274367,0.01371835,0.0274367,0.07888051,0.1371835,0.14061308,0.09602845,0.06516216,0.058302987,0.072021335,0.09945804,0.14061308,0.14404267,0.116605975,0.072021335,0.037725464,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.05144381,0.12003556,0.15433143,0.15776102,0.20920484,0.47671264,0.66533995,0.82996017,1.0048691,1.0666018,0.7579388,0.5041494,0.32581082,0.23321195,0.216064,0.23664154,0.40126175,0.4389872,0.36696586,0.22292319,0.061732575,0.034295876,0.030866288,0.0274367,0.01371835,0.0034295875,0.0034295875,0.010288762,0.01371835,0.017147938,0.020577524,0.020577524,0.020577524,0.017147938,0.017147938,0.030866288,0.048014224,0.06859175,0.06859175,0.0548734,0.061732575,0.05144381,0.0548734,0.1097468,0.22978236,0.4115505,0.36353627,0.22292319,0.12346515,0.09602845,0.09259886,0.28808534,0.36696586,0.32581082,0.22292319,0.16462019,0.15090185,0.20577525,0.26407823,0.28465575,0.23664154,0.12003556,0.06516216,0.058302987,0.10288762,0.22292319,0.4698535,0.48700142,0.40126175,0.31209245,0.28465575,0.39440256,0.53501564,0.58302987,0.53501564,0.5178677,0.5521636,0.5453044,0.548734,0.53844523,0.42869842,0.30523327,0.20920484,0.24007112,0.45613512,0.8745448,1.2243627,1.5090185,1.7765263,1.7971039,1.0597426,0.75450927,0.5761707,0.41498008,0.26750782,0.22978236,0.15433143,0.08916927,0.048014224,0.0274367,0.010288762,0.010288762,0.0274367,0.058302987,0.106317215,0.17147937,0.29494452,0.432128,0.48357183,0.42183927,0.29151493,0.21263443,0.30866286,0.58302987,0.9568549,1.2380811,1.3306799,1.9754424,2.153781,1.7662375,1.6221949,1.7113642,1.4164196,1.3992717,1.6667795,1.5638919,1.3478279,1.1900668,1.1351935,1.2003556,1.3684053,1.6393428,2.0337453,2.5824795,3.2889743,4.1360826,4.7774153,5.48734,6.3618846,7.449064,8.721441,9.362774,9.458802,9.160428,8.656279,8.169277,8.134981,8.200144,8.22758,8.128122,7.8606143,7.630832,7.73372,8.056101,8.495089,8.947794,9.294182,9.3593445,9.294182,9.246168,9.373062,9.259886,7.6685576,5.8200097,4.6745276,4.914599,5.6142344,5.2026844,4.149801,3.223812,3.5016088,4.5819287,5.5662203,6.001778,6.307011,7.7748747,7.058091,6.2555676,6.478491,8.069819,10.604284,9.256456,8.368194,8.069819,7.5862474,5.24041,4.7191124,3.5633414,2.2086544,1.0528834,0.48357183,0.490431,0.4698535,0.53844523,0.8025235,1.3581166,2.5413244,2.6133456,2.270387,1.862266,1.3992717,0.922559,0.48014224,0.17490897,0.037725464,0.044584636,0.08573969,0.42183927,0.47671264,0.20234565,0.07545093,0.030866288,0.006859175,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.010288762,0.044584636,0.05144381,0.058302987,0.08916927,0.1371835,0.16804978,0.13032432,0.09602845,0.09259886,0.11317638,0.12346515,0.12346515,0.2194936,0.3841138,0.65848076,1.1626302,1.8519772,2.6579304,3.1655092,3.3369887,3.525616,3.8102717,4.40359,5.2506986,6.1629686,6.807731,6.48535,6.1492505,5.6348124,5.2026844,5.5490727,5.5730796,3.2546785,1.5570327,1.3924125,1.6221949,1.9068506,2.5138876,3.9303071,5.9126086,7.4799304,8.738589,9.743458,10.590566,11.170166,11.166737,11.166737,10.813489,10.240748,9.650859,9.3079,9.211872,9.153569,9.369633,9.863494,10.408798,10.88894,11.173596,11.492548,12.103014,13.296511,15.419425,17.034761,17.751545,17.247395,15.271953,12.943263,11.938394,12.950122,15.395418,17.391438,17.765263,16.064188,13.21763,10.281903,8.450503,7.39762,6.2864337,4.8425775,3.309552,2.452155,1.8005334,1.5638919,1.3992717,1.155771,0.86082643,0.70649505,0.7305021,0.7099246,0.58645946,0.4664239,0.39783216,0.37725464,0.36353627,0.35324752,0.37725464,0.3841138,0.33609957,0.34981793,0.4389872,0.5178677,0.26750782,0.2709374,0.32924038,0.34638834,0.32581082,0.15090185,0.13032432,0.1371835,0.13375391,0.16804978,0.08573969,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.1920569,0.3806842,0.48700142,0.3841138,0.16119061,0.061732575,0.048014224,0.07888051,0.09259886,0.06859175,0.058302987,0.058302987,0.061732575,0.05144381,0.034295876,0.020577524,0.017147938,0.030866288,0.061732575,0.06516216,0.08916927,0.11317638,0.11317638,0.041155048,0.030866288,0.07545093,0.4355576,1.2655178,2.6064866,4.1943855,4.7019644,4.389872,3.4844608,2.2155135,1.7662375,1.7593783,1.7353712,1.4781522,1.0254467,0.7339317,0.72021335,0.82996017,0.980862,1.1523414,1.3066728,1.4232788,1.4095604,1.2758065,1.1420527,1.1249046,1.2483698,1.4953002,1.7799559,1.9480057,2.0406046,2.1915064,2.386993,2.452155,2.0474637,1.5433143,1.1249046,0.83338976,0.6927767,0.72364295,1.0048691,1.3341095,1.7971039,2.4590142,3.3369887,4.180667,5.055212,5.6656785,5.8371577,5.48734,5.051782,4.852866,4.73969,4.547633,4.0949273,3.4844608,3.2615378,3.1243541,2.983741,2.9494452,3.1277838,3.3266997,3.175798,2.6819375,2.2292318,2.0817597,2.1057668,2.2086544,2.3767042,2.6476414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.06859175,0.048014224,0.017147938,0.010288762,0.044584636,0.106317215,0.07545093,0.034295876,0.01371835,0.01371835,0.0034295875,0.010288762,0.20577525,0.50757897,0.5796003,0.31209245,0.14404267,0.05144381,0.01371835,0.01371835,0.06516216,0.15776102,0.16462019,0.08573969,0.061732575,0.048014224,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.041155048,0.07545093,0.22292319,0.2777966,0.26407823,0.23321195,0.24350071,0.805953,0.94656616,0.82996017,0.61046654,0.42869842,0.47671264,0.38754338,0.2709374,0.22635277,0.33609957,0.8128122,0.91227025,0.7476501,0.45270553,0.18176813,0.14747226,0.12003556,0.07545093,0.0274367,0.01371835,0.01371835,0.01371835,0.01371835,0.020577524,0.044584636,0.044584636,0.037725464,0.041155048,0.06859175,0.09259886,0.07888051,0.08573969,0.09259886,0.09602845,0.12346515,0.12346515,0.12346515,0.12689474,0.14404267,0.16804978,0.26407823,0.28122616,0.21263443,0.116605975,0.09259886,0.34638834,0.51100856,0.5555932,0.4698535,0.274367,0.36010668,0.7305021,1.0700313,1.1763484,0.9294182,0.30866286,0.08916927,0.07545093,0.17490897,0.3806842,0.78537554,0.9568549,0.89855194,0.6859175,0.5041494,0.52815646,0.72707254,0.7888051,0.66533995,0.5796003,0.6036074,0.72021335,0.823101,0.83338976,0.6859175,0.45613512,0.2503599,0.15776102,0.18862732,0.274367,0.32238123,0.33609957,0.32924038,0.31552204,0.29151493,0.2777966,0.274367,0.25721905,0.24007112,0.29151493,0.20577525,0.1097468,0.048014224,0.034295876,0.044584636,0.044584636,0.0274367,0.01371835,0.024007112,0.061732575,0.048014224,0.0274367,0.01371835,0.020577524,0.044584636,0.09602845,0.39097297,0.9945804,1.7147937,2.1057668,1.7765263,2.6819375,3.1209247,2.9288676,3.4776018,4.2115335,2.9220085,1.7662375,1.4815818,1.3581166,1.3443983,1.371835,1.3649758,1.3443983,1.4027013,1.5501735,1.8245405,2.3149714,3.0351849,3.9508848,4.866585,6.0497923,7.5759587,9.270175,10.710602,11.5645685,11.934964,11.917816,11.684605,11.489118,10.926665,10.175586,9.259886,8.213862,7.0786686,6.5539417,6.7528577,7.6376915,9.105555,10.984968,12.524854,11.406808,9.441654,7.6514096,6.2727156,5.4667625,4.07435,3.1415021,3.2889743,4.729401,6.7185616,5.8988905,4.804852,4.722542,5.675967,6.725421,6.7494283,6.5367937,6.420188,6.2864337,6.262427,6.660259,8.158989,10.103564,10.484249,9.016385,7.425057,6.6876955,6.2418494,3.981751,3.2272418,2.7882545,2.3801336,1.8039631,0.9602845,1.3272504,1.4541451,1.3889829,1.2963841,1.4815818,2.4555845,3.059192,3.3026927,3.216953,2.8396983,2.4590142,1.4507155,0.52815646,0.058302987,0.044584636,0.010288762,0.010288762,0.058302987,0.12346515,0.1371835,0.05144381,0.01371835,0.0,0.0034295875,0.01371835,0.0274367,0.01371835,0.0,0.010288762,0.044584636,0.06859175,0.07545093,0.082310095,0.09602845,0.106317215,0.12003556,0.14061308,0.19548649,0.24350071,0.18176813,0.19548649,0.2709374,0.44927597,0.9294182,2.0920484,3.3369887,4.1120753,4.523626,4.8425775,5.5387836,4.5270553,3.5393343,2.9254382,2.9391565,3.7691166,5.3330083,5.209543,4.7808447,4.9248877,6.012067,7.599966,5.2301207,2.6064866,1.4129901,1.3272504,1.2895249,1.5741806,1.8485477,2.1332035,2.7916842,4.197815,6.0669403,8.210432,10.127572,11.032983,10.984968,10.714031,10.367643,9.89436,9.0644,8.344186,8.052671,8.522525,9.3593445,9.445084,9.554831,9.774324,10.14129,10.868362,12.343085,15.189643,18.296848,20.954779,21.921923,19.469769,16.37971,14.658057,14.280802,15.073037,16.70895,19.795578,19.689262,17.364002,13.735497,9.657719,6.691125,5.7754254,5.65539,5.5422134,5.127233,4.064061,4.15666,3.9474552,2.9734523,1.7388009,0.97057325,1.1626302,1.4507155,1.4438564,1.2346514,0.89512235,0.607037,0.48357183,0.5007198,0.48700142,0.4629943,0.31895164,0.29494452,0.4081209,0.45613512,0.4698535,0.47328308,0.4972902,0.48357183,0.29151493,0.1920569,0.13032432,0.09602845,0.1920569,0.65505123,0.34981793,0.1097468,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.17490897,0.3841138,0.45613512,0.32238123,0.13375391,0.024007112,0.030866288,0.09259886,0.07888051,0.07545093,0.09945804,0.12346515,0.07545093,0.041155048,0.01371835,0.0,0.0,0.0,0.01371835,0.024007112,0.037725464,0.041155048,0.01371835,0.01371835,0.034295876,0.13032432,0.31209245,0.5178677,0.44584638,0.37382504,0.36010668,0.42183927,0.5178677,0.7133542,0.6344737,0.5624523,0.59674823,0.67219913,0.7682276,0.8745448,0.84367853,0.72707254,0.7613684,0.9328478,1.1214751,1.2517995,1.2380811,1.0082988,0.77508676,0.6344737,0.548734,0.4938606,0.45956472,0.5796003,0.8128122,1.1283343,1.3752645,1.2655178,1.0837497,0.864256,0.65162164,0.52815646,0.6241849,0.85739684,1.2175035,1.7422304,2.4487255,3.3266997,3.974892,4.5201964,4.9214582,5.144381,5.1580997,4.98662,4.972902,5.1100855,5.3398676,5.5250654,5.4016004,5.305572,5.2644167,5.2918534,5.4016004,5.5730796,5.579939,5.3844523,4.976331,4.3795834,3.8788633,3.7622573,3.8960114,4.1017866,4.149801,0.037725464,0.06516216,0.06516216,0.041155048,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.0274367,0.01371835,0.0034295875,0.010288762,0.058302987,0.07888051,0.048014224,0.020577524,0.020577524,0.041155048,0.048014224,0.020577524,0.044584636,0.13375391,0.22635277,0.21263443,0.15776102,0.082310095,0.017147938,0.0274367,0.048014224,0.09602845,0.15090185,0.19891608,0.23321195,0.16119061,0.1097468,0.072021335,0.041155048,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.041155048,0.07888051,0.106317215,0.13032432,0.16462019,0.25721905,0.6241849,0.6859175,0.59674823,0.4664239,0.34295875,0.274367,0.22978236,0.20577525,0.21263443,0.26407823,0.45613512,0.6173257,0.6962063,0.66191036,0.5007198,0.33609957,0.2469303,0.17147937,0.08916927,0.0274367,0.006859175,0.010288762,0.01371835,0.020577524,0.034295876,0.044584636,0.058302987,0.08573969,0.13375391,0.22635277,0.17490897,0.11317638,0.09259886,0.116605975,0.12346515,0.12346515,0.18176813,0.28122616,0.4046913,0.5453044,0.52815646,0.40126175,0.28122616,0.2777966,0.50757897,0.82996017,0.8676856,0.7339317,0.5418748,0.39783216,0.71678376,1.1729189,1.4095604,1.2655178,0.7956643,0.22292319,0.058302987,0.09602845,0.22635277,0.45613512,0.77851635,0.7373613,0.6344737,0.607037,0.6001778,0.65505123,0.77851635,0.88826317,0.9568549,1.0185875,1.0940384,1.1763484,1.2277923,1.1934965,1.0288762,0.7476501,0.47328308,0.32581082,0.32238123,0.36010668,0.4389872,0.47328308,0.432128,0.33266997,0.24007112,0.20920484,0.18519773,0.17490897,0.16462019,0.15433143,0.18862732,0.18176813,0.16804978,0.18862732,0.2777966,0.13032432,0.0548734,0.024007112,0.017147938,0.024007112,0.01371835,0.006859175,0.0034295875,0.0034295875,0.010288762,0.037725464,0.16119061,0.52472687,1.0494537,1.4232788,1.2209331,1.2483698,1.8485477,2.9288676,3.9680326,4.5922174,5.055212,4.9591837,4.355576,3.724532,3.1963756,2.7402403,2.4212887,2.1812177,1.8313997,1.6942163,1.8108221,1.9857311,2.201795,2.609916,3.457024,4.671098,6.183546,7.8537555,9.489669,10.062409,10.302481,10.463672,10.6488695,10.792912,10.943813,10.978109,10.844356,10.508256,9.949233,8.944365,8.14527,7.764586,7.9943686,8.995808,10.858074,10.611144,9.369633,7.874333,6.5162163,5.5833683,5.1340923,5.1855364,5.6793966,6.475061,7.1266828,7.0478024,7.459353,8.690575,10.179015,11.005547,10.329918,9.592556,9.266746,8.848335,7.9189177,6.118384,6.728851,9.678296,11.533703,11.153018,9.242738,7.5279446,6.4716315,5.288424,4.962613,4.65395,3.8342788,2.4898806,1.1214751,1.0871792,1.4369972,1.8759843,2.2223728,2.3972816,3.0111778,3.4638834,3.6010668,3.3438478,2.6922262,3.0660512,2.726522,1.5021594,0.09602845,0.082310095,0.034295876,0.18862732,0.37382504,0.5144381,0.6241849,0.36353627,0.17147937,0.0548734,0.01371835,0.01371835,0.017147938,0.030866288,0.037725464,0.048014224,0.09602845,0.19548649,0.31209245,0.39097297,0.41840968,0.40126175,0.32238123,0.2709374,0.274367,0.3018037,0.26750782,0.2503599,0.31209245,0.4664239,0.7510797,1.2483698,1.7799559,2.1229146,2.1229146,1.9308578,2.0097382,1.8588364,2.1126258,3.3815732,5.528495,7.6857057,8.086967,7.56567,6.831738,6.138962,5.2918534,5.686256,5.1100855,4.2081037,3.2306714,2.0234566,2.085189,2.194936,2.1812177,2.0440342,1.961724,2.9254382,3.8891523,5.3432975,7.425057,9.908078,10.796341,11.084427,10.840926,10.192734,9.331907,9.091836,8.423067,7.98408,7.9086285,7.798882,7.5931067,8.073249,9.026674,10.1481495,11.050131,12.428825,15.004445,17.806417,20.313446,22.450079,22.906214,21.472647,19.682402,18.1288,16.46545,16.496315,16.87014,17.641798,17.926455,15.920145,12.88496,10.590566,9.335337,8.841476,8.237869,7.706283,7.5245147,7.2432885,6.4579134,4.8151407,3.998899,3.6593697,3.5153272,3.391862,3.2135234,2.9494452,2.3389788,1.7079345,1.2586586,1.0494537,0.66533995,0.3806842,0.22292319,0.16119061,0.09259886,0.2709374,0.2777966,0.274367,0.33952916,0.4972902,0.8505377,0.7305021,0.5693115,0.607037,0.9259886,1.155771,0.69963586,0.2469303,0.06859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.044584636,0.12003556,0.20234565,0.16462019,0.116605975,0.1097468,0.1371835,0.12689474,0.1371835,0.09945804,0.06516216,0.048014224,0.041155048,0.041155048,0.030866288,0.01371835,0.0,0.0,0.01371835,0.017147938,0.020577524,0.017147938,0.0034295875,0.0034295875,0.006859175,0.030866288,0.08573969,0.16462019,0.18862732,0.20577525,0.20234565,0.18862732,0.18862732,0.2469303,0.274367,0.28465575,0.28808534,0.29151493,0.31209245,0.37039545,0.48014224,0.64133286,0.823101,0.96714365,1.138623,1.3409687,1.488441,1.4232788,1.2380811,1.0597426,0.8711152,0.66191036,0.4081209,0.30523327,0.29151493,0.33609957,0.38754338,0.37382504,0.34981793,0.31552204,0.28465575,0.3018037,0.41840968,0.6001778,0.8471081,1.2106444,1.7319417,2.435007,3.0729103,3.7348208,4.091498,4.1463714,4.2183924,5.305572,5.892031,6.252138,6.5813785,6.989499,7.394191,7.922347,8.196714,8.179566,8.172707,8.666568,8.899779,8.601405,7.864044,7.15069,6.883182,6.495639,6.3378778,6.451054,6.5779486,0.072021335,0.08916927,0.07545093,0.05144381,0.024007112,0.0274367,0.034295876,0.048014224,0.044584636,0.024007112,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0034295875,0.017147938,0.05144381,0.09259886,0.106317215,0.1097468,0.1097468,0.082310095,0.07888051,0.058302987,0.048014224,0.06859175,0.12689474,0.22978236,0.22292319,0.15090185,0.07545093,0.06859175,0.10288762,0.17833854,0.24007112,0.2503599,0.20920484,0.13375391,0.11317638,0.09602845,0.061732575,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.034295876,0.044584636,0.082310095,0.15090185,0.23321195,0.38754338,0.45270553,0.42183927,0.33266997,0.23664154,0.15433143,0.12003556,0.12346515,0.15433143,0.19891608,0.31895164,0.5453044,0.85739684,1.0906088,0.9568549,0.69963586,0.5007198,0.37039545,0.29494452,0.21263443,0.15090185,0.10288762,0.058302987,0.024007112,0.020577524,0.034295876,0.0548734,0.082310095,0.116605975,0.16804978,0.12003556,0.07888051,0.072021335,0.08916927,0.06859175,0.10288762,0.22292319,0.432128,0.7133542,1.0425946,0.59331864,0.32581082,0.25721905,0.40126175,0.77508676,1.2346514,1.2895249,1.0734608,0.7407909,0.4355576,0.5796003,0.9911508,1.2483698,1.1763484,0.83681935,0.34638834,0.23321195,0.32581082,0.5144381,0.7373613,0.91912943,0.78537554,0.72021335,0.84367853,1.0185875,1.2415106,1.4747226,1.4610043,1.2380811,1.1763484,1.5673214,2.1160555,1.9480057,1.1660597,0.85739684,0.6756287,0.5178677,0.432128,0.41840968,0.4355576,0.5007198,0.51100856,0.42869842,0.28808534,0.1920569,0.14747226,0.11317638,0.08916927,0.07545093,0.058302987,0.10288762,0.16119061,0.21263443,0.2469303,0.26407823,0.3806842,0.29151493,0.13375391,0.020577524,0.034295876,0.01371835,0.01371835,0.020577524,0.030866288,0.037725464,0.037725464,0.07545093,0.24007112,0.51100856,0.7305021,0.64476246,0.58988905,0.9774324,1.8005334,2.6167753,3.316411,4.280125,4.513337,3.9543142,3.4673128,3.093488,2.4452958,2.201795,2.369845,2.2841053,2.0337453,1.7490896,1.5810398,1.5947582,1.7422304,2.294394,3.1723683,4.3349986,5.6313825,6.831738,7.3564653,7.6616983,7.915488,8.282454,8.916927,9.671436,10.412228,11.118723,11.756626,12.284782,11.228469,10.199594,9.431366,8.985519,8.766026,9.3936405,9.043822,8.186425,7.208993,6.4133286,6.0326443,6.0223556,6.2041235,6.447624,6.6636887,6.910619,7.15069,8.049242,9.671436,11.509696,12.0138445,12.435684,13.306799,14.188204,13.684054,10.933525,8.200144,7.548522,8.944365,10.230459,10.443094,9.547972,8.501947,7.6959944,6.941485,6.307011,5.3501563,4.383013,3.3644254,1.8999915,1.6496316,2.3286898,2.5138876,2.095478,2.2566686,3.0557625,3.998899,4.6402316,4.681387,3.981751,3.357566,2.5207467,1.2895249,0.106317215,0.06516216,0.082310095,0.35324752,0.6756287,1.0494537,1.6907866,1.9068506,1.6667795,1.1523414,0.7099246,0.85739684,0.85739684,0.7922347,0.64819205,0.42526886,0.15090185,0.4355576,0.69963586,0.8779744,0.9328478,0.85739684,0.61389613,0.5624523,0.61389613,0.70306545,0.77508676,0.86082643,0.83681935,0.9877212,1.3992717,1.9720128,2.6613598,3.216953,3.426158,3.3541365,3.3644254,3.5770597,4.15323,5.1580997,6.6533995,8.711152,9.818909,10.017825,9.740028,9.136421,8.069819,7.2124224,6.461343,6.200694,5.967482,4.4413157,3.6010668,2.8739944,2.369845,1.9857311,1.3786942,1.7353712,2.2635276,3.2581081,5.051782,8.025234,9.938945,11.393089,12.277924,12.38767,11.441104,11.063849,10.521975,10.14129,9.877212,9.318189,8.522525,8.176137,8.303031,8.735159,9.098696,9.530824,11.108434,13.296511,15.902997,19.082224,21.647556,22.899355,23.170294,22.559826,20.934202,18.495766,16.911295,16.516893,16.650646,15.638919,13.214201,11.375941,10.535692,10.422516,10.052121,9.438225,8.7317295,8.090397,7.517656,6.848886,6.7219915,6.550512,6.2144127,5.703404,5.1100855,4.3658648,3.3747141,2.3664153,1.6016173,1.3443983,1.0837497,0.8093826,0.51100856,0.24007112,0.12003556,0.19891608,0.23321195,0.30866286,0.5007198,0.8711152,0.8711152,0.6756287,0.48014224,0.38754338,0.39783216,0.6893471,0.52815646,0.24007112,0.034295876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.06516216,0.08916927,0.09259886,0.10288762,0.12003556,0.12003556,0.12346515,0.08916927,0.044584636,0.01371835,0.01371835,0.024007112,0.024007112,0.01371835,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0034295875,0.010288762,0.030866288,0.05144381,0.072021335,0.07545093,0.06516216,0.061732575,0.08573969,0.13032432,0.16462019,0.17147937,0.15090185,0.15090185,0.20234565,0.32581082,0.5144381,0.7476501,0.85396725,0.94999576,1.0837497,1.214074,1.2415106,1.138623,0.99801,0.82996017,0.6379033,0.4046913,0.23321195,0.13032432,0.07888051,0.06516216,0.06859175,0.07545093,0.07888051,0.08573969,0.116605975,0.20920484,0.36010668,0.5555932,0.8196714,1.1900668,1.7079345,2.3801336,3.1277838,3.5050385,3.4776018,3.4227283,4.6882463,5.813151,6.584808,7.0752387,7.6205435,7.9086285,8.347616,8.652849,8.64599,8.289313,8.570539,8.769455,8.666568,8.272165,7.8434668,7.7748747,7.8537555,8.176137,8.738589,9.448513,0.072021335,0.06859175,0.05144381,0.034295876,0.020577524,0.0274367,0.041155048,0.0548734,0.05144381,0.037725464,0.048014224,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.041155048,0.1097468,0.15090185,0.17833854,0.18519773,0.15090185,0.1371835,0.09602845,0.06859175,0.07888051,0.116605975,0.20577525,0.2194936,0.17147937,0.10288762,0.072021335,0.12346515,0.22978236,0.29494452,0.2777966,0.17490897,0.09602845,0.08573969,0.07888051,0.0548734,0.037725464,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.017147938,0.048014224,0.10288762,0.15776102,0.19891608,0.24350071,0.2469303,0.19891608,0.13375391,0.07545093,0.05144381,0.05144381,0.072021335,0.106317215,0.20920484,0.39783216,0.6893471,0.9945804,1.1146159,0.8711152,0.6001778,0.44584638,0.42869842,0.4698535,0.3806842,0.28122616,0.19548649,0.13032432,0.09602845,0.09259886,0.07888051,0.072021335,0.07545093,0.082310095,0.06859175,0.072021335,0.08573969,0.09259886,0.0548734,0.116605975,0.33609957,0.59331864,0.8196714,0.97057325,0.44927597,0.2709374,0.31209245,0.4972902,0.7922347,1.1592005,1.2758065,1.1660597,0.9259886,0.7099246,0.88826317,1.3478279,1.5604624,1.3581166,0.939707,0.45270553,0.32924038,0.44584638,0.6927767,1.0014396,1.3684053,1.6770682,1.8039631,1.762808,1.7147937,1.6770682,1.6907866,1.5947582,1.430138,1.4541451,1.7696671,2.1263442,1.7799559,0.91569984,0.66876954,0.58645946,0.52815646,0.490431,0.4664239,0.42869842,0.42526886,0.39097297,0.30866286,0.20920484,0.16119061,0.12346515,0.082310095,0.048014224,0.024007112,0.01371835,0.061732575,0.1371835,0.20234565,0.22978236,0.17833854,0.33952916,0.2709374,0.12346515,0.01371835,0.0274367,0.017147938,0.017147938,0.024007112,0.037725464,0.061732575,0.07888051,0.1097468,0.15776102,0.21263443,0.2469303,0.22635277,0.37039545,0.805953,1.4404267,1.9445761,1.9754424,2.3492675,2.3972816,2.0508933,1.8176813,1.7079345,1.4164196,1.4507155,1.821111,2.0234566,1.9239986,1.5604624,1.2689474,1.1797781,1.2346514,1.529596,2.0097382,2.6956558,3.4947495,4.197815,4.65395,5.038064,5.4839106,6.121814,7.051232,8.131552,9.239308,10.31277,11.355364,12.452832,11.766914,10.950673,10.251037,9.619993,8.738589,8.772884,8.591117,8.186425,7.654839,7.174697,7.377043,7.514226,7.5382333,7.473071,7.421627,7.5725293,7.888051,8.683716,10.007536,11.653738,11.96926,12.912396,14.376831,15.683503,15.570327,13.138749,11.677745,10.854645,10.288762,9.551401,8.783174,8.81404,8.652849,7.953213,7.010077,6.1732574,5.254128,4.537344,3.8102717,2.3664153,1.6530612,2.277246,2.435007,1.9480057,2.2635276,3.7108135,6.0703697,7.274155,6.7700057,5.5387836,3.8479972,2.0337453,0.70306545,0.08573969,0.041155048,0.08573969,0.44927597,1.0460242,1.8073926,2.6613598,2.8019729,2.301253,1.6016173,1.1351935,1.2963841,1.2586586,1.1454822,0.96371406,0.6893471,0.2503599,0.66533995,1.0940384,1.3958421,1.4644338,1.2243627,1.2346514,1.2895249,1.255229,1.08032,0.7922347,0.9774324,1.1317638,1.6187652,2.6064866,4.046913,3.7691166,4.125794,4.705394,5.2506986,5.6348124,6.2247014,7.051232,7.682276,8.255017,9.462232,11.0981455,12.325937,12.97413,12.9707,12.370522,11.074138,9.379922,8.237869,7.531374,6.0806584,5.079219,3.9200184,3.0660512,2.5173173,1.7936742,1.6873571,1.8588364,2.3218307,3.426158,5.871454,8.337327,10.7586155,13.015285,14.534592,14.291091,13.845244,13.502286,13.433694,13.320518,12.343085,11.207891,10.155008,9.297611,8.597976,7.8777623,7.881192,8.64599,9.839486,11.489118,13.954991,16.722668,19.658396,22.316326,24.161444,24.572994,21.86362,19.274282,17.144508,15.395418,13.543441,11.434244,10.196163,9.702303,9.623423,9.424506,9.692014,9.5205345,9.187865,8.916927,8.862054,8.848335,8.690575,8.203573,7.3873315,6.420188,5.2918534,4.400161,3.5770597,2.8225505,2.3286898,1.821111,1.5570327,1.2929544,0.980862,0.75450927,0.5212973,0.52472687,0.5418748,0.53501564,0.6756287,0.5212973,0.48700142,0.47328308,0.41840968,0.29151493,0.48700142,0.50757897,0.30523327,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.044584636,0.058302987,0.07888051,0.10288762,0.106317215,0.07888051,0.05144381,0.0274367,0.01371835,0.024007112,0.030866288,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.017147938,0.034295876,0.06859175,0.11317638,0.14747226,0.14747226,0.15776102,0.1920569,0.2503599,0.34638834,0.5041494,0.5693115,0.58645946,0.61046654,0.64476246,0.66876954,0.6276145,0.5624523,0.48014224,0.3806842,0.2709374,0.14747226,0.072021335,0.030866288,0.01371835,0.010288762,0.010288762,0.010288762,0.01371835,0.034295876,0.08916927,0.2194936,0.5590228,0.9294182,1.2175035,1.3615463,1.7113642,2.386993,2.867135,2.976882,2.8739944,3.4844608,4.3487167,5.3913116,6.420188,7.15069,7.414768,7.720001,8.045813,8.134981,7.48336,7.274155,7.466212,7.9086285,8.354475,8.453933,8.618553,9.153569,9.983529,11.012405,12.109874,0.044584636,0.041155048,0.024007112,0.010288762,0.0,0.0,0.010288762,0.01371835,0.01371835,0.024007112,0.06516216,0.0274367,0.006859175,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.010288762,0.037725464,0.106317215,0.13375391,0.15776102,0.18519773,0.20234565,0.18519773,0.106317215,0.06516216,0.09259886,0.15090185,0.16804978,0.17833854,0.16462019,0.12346515,0.072021335,0.12346515,0.23321195,0.31552204,0.32238123,0.23664154,0.1371835,0.08573969,0.061732575,0.0548734,0.048014224,0.044584636,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.061732575,0.082310095,0.082310095,0.082310095,0.08573969,0.058302987,0.024007112,0.01371835,0.006859175,0.0034295875,0.01371835,0.07545093,0.15090185,0.24007112,0.42526886,0.84024894,0.70306545,0.4972902,0.39097297,0.4355576,0.58988905,0.5144381,0.42183927,0.35324752,0.31552204,0.29494452,0.24007112,0.16804978,0.11317638,0.09259886,0.09945804,0.12346515,0.1371835,0.1371835,0.12346515,0.09259886,0.1371835,0.41840968,0.65162164,0.6893471,0.48700142,0.3566771,0.48357183,0.64819205,0.7476501,0.8128122,0.89855194,1.0288762,1.0940384,1.1146159,1.2277923,1.646202,2.0646117,2.0989075,1.6976458,1.1077567,0.6310441,0.5007198,0.64476246,1.0014396,1.5330256,2.4624438,3.649081,3.8788633,3.1106358,2.486451,1.9411465,1.5261664,1.4267083,1.7147937,2.3458378,2.1229146,1.4404267,0.864256,0.6276145,0.64476246,0.6344737,0.58302987,0.5212973,0.45270553,0.37725464,0.29151493,0.21263443,0.16119061,0.14061308,0.14747226,0.12346515,0.08916927,0.05144381,0.024007112,0.020577524,0.07888051,0.13375391,0.17147937,0.16804978,0.09945804,0.041155048,0.010288762,0.0,0.0034295875,0.0,0.010288762,0.0034295875,0.006859175,0.024007112,0.061732575,0.12346515,0.18519773,0.20234565,0.15433143,0.07888051,0.082310095,0.4115505,1.1043272,1.8759843,2.1332035,1.1111864,0.607037,0.37725464,0.25721905,0.16119061,0.16804978,0.42869842,0.6824879,0.85739684,1.0837497,1.2312219,1.138623,0.96714365,0.8471081,0.90884066,1.1008976,1.3341095,1.6530612,2.0474637,2.4795918,2.867135,3.3266997,4.029765,4.955754,5.874883,6.958633,8.035523,8.916927,9.637141,10.446524,10.357354,10.100135,9.945804,9.962952,10.0041065,10.734609,11.2421875,11.406808,11.238758,10.868362,11.077567,10.80663,10.175586,9.510246,9.349055,9.373062,9.56512,9.928656,10.456812,11.135871,11.187314,11.598865,12.308789,13.121602,13.708061,13.612033,14.568888,14.911846,14.003006,12.22305,9.122703,8.704293,8.378482,7.130112,5.518206,4.763697,4.4584637,4.07435,3.3061223,2.07833,1.1523414,1.3821237,1.7730967,2.1332035,3.0797696,6.200694,9.417647,10.1481495,8.347616,6.509357,4.9934793,2.2155135,0.40126175,0.06859175,0.041155048,0.05144381,0.39440256,1.2998136,2.486451,3.1449318,2.7916842,2.294394,1.9925903,1.9274281,1.8588364,1.6736387,1.5433143,1.2998136,0.9911508,0.8711152,1.5638919,2.277246,2.486451,2.136633,1.6324836,2.3767042,2.8911421,2.7299516,1.8999915,0.8676856,0.89855194,1.2449403,2.0474637,3.532475,6.025785,4.40702,4.15323,4.8185706,5.8817425,6.7665763,7.6651278,8.635701,9.253027,9.510246,9.832627,11.14273,13.049581,14.668345,15.563468,15.731518,14.970149,12.840376,10.398509,8.296172,6.783724,6.258997,5.381023,4.6093655,4.057202,3.4878905,2.8808534,2.503599,2.3149714,2.5721905,3.8342788,6.0978065,9.071259,12.445972,15.374841,16.503176,16.187653,15.947581,16.081335,16.249386,15.481158,14.723219,13.519434,12.065289,10.408798,8.460793,8.049242,8.2481575,8.587687,9.119273,10.425946,12.061859,14.671775,18.159666,21.78474,24.154585,23.235455,21.805317,19.582945,16.530611,12.850664,10.323058,8.999237,8.162418,7.534804,7.2775846,8.700864,9.657719,10.316199,10.714031,10.748327,10.39508,10.048691,9.47595,8.625413,7.6376915,6.3310184,5.7308407,5.40503,4.979761,4.1635194,2.9734523,2.4727325,2.2463799,2.1057668,2.07833,1.430138,1.488441,1.587899,1.2929544,0.40126175,0.2469303,0.40126175,0.61046654,0.70649505,0.61046654,0.9602845,0.8676856,0.47671264,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.06516216,0.10288762,0.09602845,0.037725464,0.010288762,0.010288762,0.034295876,0.058302987,0.061732575,0.041155048,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.07545093,0.14061308,0.20234565,0.2469303,0.2503599,0.22978236,0.20234565,0.20577525,0.22978236,0.20577525,0.16462019,0.12003556,0.09259886,0.08573969,0.082310095,0.07888051,0.06859175,0.06516216,0.0274367,0.017147938,0.017147938,0.01371835,0.0,0.0,0.0034295875,0.01371835,0.034295876,0.06859175,0.19891608,0.6756287,1.1694894,1.4198492,1.214074,1.0666018,1.5021594,2.0406046,2.3835633,2.4384367,2.3492675,2.4418662,3.275256,4.5990767,5.3741636,5.895461,6.3618846,6.8626046,7.140401,6.5779486,6.0875177,6.3653145,7.3358874,8.621983,9.544542,10.31277,11.153018,12.140739,13.251926,14.363112,0.044584636,0.06859175,0.041155048,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.01371835,0.0,0.0,0.0,0.01371835,0.034295876,0.034295876,0.024007112,0.061732575,0.061732575,0.041155048,0.041155048,0.07888051,0.15090185,0.116605975,0.061732575,0.07888051,0.18519773,0.31895164,0.30866286,0.2777966,0.2777966,0.28122616,0.18176813,0.24350071,0.33266997,0.4046913,0.4424168,0.4424168,0.29494452,0.19548649,0.15090185,0.13375391,0.061732575,0.037725464,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.020577524,0.034295876,0.044584636,0.020577524,0.006859175,0.0,0.0,0.0,0.024007112,0.06859175,0.13375391,0.216064,0.29151493,0.29151493,0.35324752,0.42183927,0.41840968,0.26064864,0.2709374,0.274367,0.31895164,0.42869842,0.6241849,0.4424168,0.32238123,0.26750782,0.2709374,0.31895164,0.34638834,0.26750782,0.17147937,0.10288762,0.09259886,0.07888051,0.20577525,0.3566771,0.48700142,0.61046654,0.82996017,1.2517995,1.5090185,1.5090185,1.4335675,1.4335675,1.4541451,1.4404267,1.4575747,1.6770682,1.9239986,1.5981878,1.4164196,1.5090185,1.4507155,1.3169615,1.3375391,1.6359133,2.253239,3.1415021,4.7191124,6.584808,6.245279,4.0023284,2.976882,2.585909,2.311542,2.136633,2.5173173,4.4104495,3.7382503,1.9308578,0.70649505,0.53501564,0.65505123,0.75450927,0.72364295,0.5521636,0.36696586,0.42869842,0.32924038,0.24007112,0.17833854,0.14747226,0.12346515,0.1097468,0.09602845,0.07888051,0.058302987,0.044584636,0.09602845,0.12346515,0.13032432,0.09945804,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.0,0.0,0.0,0.006859175,0.024007112,0.061732575,0.12346515,0.16462019,0.18862732,0.20234565,0.21263443,0.274367,0.6927767,1.1008976,1.255229,1.0220171,0.216064,0.01371835,0.010288762,0.0034295875,0.01371835,0.041155048,0.1097468,0.18176813,0.24007112,0.29151493,0.33952916,0.34295875,0.34638834,0.39783216,0.5178677,0.7373613,0.9945804,1.2895249,1.6256244,2.0303159,2.5893385,3.2992632,4.0606318,4.8254294,5.56965,6.39961,7.2021337,7.7028537,7.870903,7.9189177,8.261876,9.033533,10.371073,12.603734,16.266533,18.12194,19.095943,19.634388,20.02193,20.399187,19.497204,17.514904,14.747226,12.1921835,11.519984,11.30049,11.118723,10.813489,10.182446,8.988949,8.073249,8.337327,9.3936405,10.731179,11.718901,12.706621,14.116182,16.009314,18.28999,20.70442,15.45715,12.048141,9.424506,6.958633,4.4550343,3.5633414,2.7642474,2.037175,1.4438564,1.1146159,1.6153357,1.6942163,1.670209,2.311542,4.835718,11.856084,12.089295,9.685155,7.3530354,6.3618846,7.181556,3.7794054,0.8779744,0.12346515,0.07545093,0.041155048,0.07545093,0.97400284,2.4247184,3.0214665,3.216953,4.3007026,5.171818,5.3261495,4.835718,4.3109913,4.081209,3.1586502,2.0920484,2.9460156,4.616225,5.967482,5.3844523,3.3781435,2.609916,4.184097,5.960623,6.077229,4.4927597,2.9906003,2.270387,1.9891608,2.0131679,2.767677,5.2335505,5.381023,5.195825,5.195825,5.65539,6.6053853,7.0958166,7.181556,7.016936,6.842027,6.989499,7.829748,9.517105,11.633161,13.704632,15.182784,15.426285,14.682064,13.169616,11.105004,8.711152,7.407909,7.0443726,7.0203657,6.869464,6.2727156,4.4516044,3.199805,2.4247184,2.0886188,2.1983654,3.5050385,7.016936,11.012405,14.342535,16.417435,16.016174,15.868701,16.071047,16.654078,17.593784,18.348293,17.192522,15.385129,13.536582,11.595435,9.791472,9.163857,9.414218,10.096705,10.621432,11.427385,13.035862,15.172495,17.329706,18.78385,19.809298,20.724997,20.817596,19.28457,15.244516,11.691463,9.613133,8.134981,7.010077,6.608815,6.4990683,6.90033,8.31675,10.261326,11.2593355,11.688034,11.72233,11.369082,10.7757635,10.237319,8.529384,7.298162,6.883182,6.8969,6.2247014,4.6265135,3.3198407,2.5824795,2.7128036,4.0434837,3.0420442,3.6147852,4.770556,4.8940215,1.7696671,0.6962063,0.36353627,0.36353627,0.36696586,0.12346515,1.3786942,1.1626302,0.48357183,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.037725464,0.061732575,0.061732575,0.024007112,0.006859175,0.020577524,0.044584636,0.058302987,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.041155048,0.116605975,0.274367,0.39783216,0.40126175,0.31552204,0.1920569,0.106317215,0.09602845,0.082310095,0.082310095,0.09259886,0.09259886,0.116605975,0.11317638,0.106317215,0.09945804,0.07545093,0.041155048,0.030866288,0.024007112,0.01371835,0.0,0.0,0.010288762,0.01371835,0.034295876,0.106317215,0.26407823,0.32238123,0.432128,0.6036074,0.70306545,0.64133286,0.7990939,1.0425946,1.3409687,1.7559488,2.2292318,2.3492675,2.1846473,1.9823016,2.1503513,2.860276,3.7862647,4.629943,5.212973,5.4941993,5.627953,5.936616,6.608815,7.922347,10.254466,12.572867,14.05102,14.819247,15.350834,16.448301,0.020577524,0.037725464,0.024007112,0.020577524,0.020577524,0.01371835,0.030866288,0.030866288,0.020577524,0.010288762,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0274367,0.06859175,0.09602845,0.08573969,0.0548734,0.044584636,0.05144381,0.06859175,0.10288762,0.048014224,0.037725464,0.06859175,0.11317638,0.15090185,0.16804978,0.24007112,0.29151493,0.274367,0.15776102,0.10288762,0.13375391,0.18176813,0.20920484,0.19891608,0.15776102,0.13032432,0.1371835,0.16462019,0.17147937,0.12689474,0.07888051,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.048014224,0.09602845,0.15433143,0.22978236,0.18176813,0.17490897,0.1920569,0.20920484,0.19891608,0.15090185,0.13375391,0.17490897,0.28808534,0.45613512,0.47671264,0.5555932,0.607037,0.6001778,0.53844523,0.3806842,0.23321195,0.1371835,0.08916927,0.06859175,0.09259886,0.3018037,0.6344737,0.9842916,1.1832076,1.1489118,1.0768905,0.97400284,0.8676856,0.77508676,0.77508676,0.9328478,1.2483698,1.605047,1.7765263,1.7662375,1.6221949,1.4472859,1.3478279,1.4267083,1.5536032,1.6873571,1.8725548,2.095478,2.2635276,2.4830213,2.6853669,2.2978237,1.5090185,1.255229,1.2449403,1.3752645,1.6873571,2.0886188,2.3595562,1.845118,1.1180456,0.66533995,0.58645946,0.58302987,0.6036074,0.5521636,0.42526886,0.3018037,0.34295875,0.29151493,0.2469303,0.20577525,0.16804978,0.13375391,0.11317638,0.08916927,0.072021335,0.06859175,0.09602845,0.17147937,0.23321195,0.25721905,0.2194936,0.06516216,0.07545093,0.058302987,0.041155048,0.0274367,0.024007112,0.044584636,0.08573969,0.22978236,0.4938606,0.84367853,0.77508676,0.50757897,0.2469303,0.20920484,0.64133286,2.7813954,2.4452958,1.4232788,0.66191036,0.26407823,0.09602845,0.05144381,0.06859175,0.106317215,0.1371835,0.10288762,0.13032432,0.18176813,0.26064864,0.38754338,0.52472687,0.4698535,0.4664239,0.5693115,0.65162164,0.764798,1.1934965,1.5913286,1.8108221,1.8828435,1.9857311,2.3664153,3.018037,3.7725463,4.3109913,4.8288593,5.4804807,6.0154963,6.3138704,6.392751,6.6293926,7.239859,8.652849,11.036412,14.335675,17.21653,19.418324,20.227707,19.79901,19.13024,17.87501,16.407146,15.138199,14.339106,14.095605,13.749216,13.29994,12.761495,12.250486,11.989838,11.036412,10.580277,10.875222,11.928105,13.512574,13.38911,13.413116,13.783512,14.232788,14.040731,13.313659,12.024134,9.9698105,7.431916,5.164959,4.633373,3.940596,3.100347,2.1915064,1.3443983,1.3958421,1.3649758,1.5193073,2.253239,4.0674906,8.772884,9.56512,8.628842,7.3255987,6.1904054,4.149801,2.719663,2.1057668,2.0714707,1.9445761,0.71678376,1.0048691,1.9102802,2.719663,2.8980014,2.253239,2.1400626,1.99602,1.6324836,1.2106444,1.1454822,1.2929544,1.546744,2.1263442,3.5564823,5.871454,7.7440085,8.011517,7.1266828,7.1369715,8.23444,8.718011,7.2192817,4.8322887,5.127233,7.2192817,7.3564653,7.239859,7.490219,7.6514096,7.377043,7.4765005,7.431916,6.9517736,5.960623,5.802862,5.6176643,5.5559316,5.6313825,5.720552,6.142391,6.9963584,8.303031,10.000677,11.934964,12.737488,12.8197975,12.356804,11.341646,9.602845,8.659708,8.056101,7.514226,6.7700057,5.576509,5.055212,5.0140567,5.086078,4.73969,3.309552,3.5221863,4.9523244,7.1232533,9.887501,13.426835,14.596324,15.076467,15.261664,15.45715,15.909856,16.859852,16.20137,14.836395,13.519434,12.830087,11.080997,10.683165,11.05356,11.664027,12.010415,12.79922,13.605173,14.308239,14.774663,14.891269,14.918706,15.71094,16.698662,17.189093,16.341984,12.271064,10.957532,10.984968,11.441104,11.917816,11.406808,10.875222,10.436234,10.093276,9.746887,9.938945,10.069269,10.168727,10.251037,10.299051,9.839486,9.119273,8.8929205,8.98209,8.251588,6.701414,6.169828,5.353586,4.166949,3.7519686,3.4638834,3.4981792,4.647091,5.7136927,3.5153272,1.4747226,1.1043272,0.89169276,0.3566771,0.072021335,0.48014224,0.7476501,0.5590228,0.08916927,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.037725464,0.0548734,0.048014224,0.0274367,0.020577524,0.034295876,0.044584636,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.037725464,0.07888051,0.12346515,0.14404267,0.1371835,0.10288762,0.058302987,0.0548734,0.05144381,0.048014224,0.044584636,0.0548734,0.07888051,0.09259886,0.09945804,0.09945804,0.07545093,0.041155048,0.030866288,0.024007112,0.01371835,0.01371835,0.0034295875,0.0034295875,0.006859175,0.024007112,0.058302987,0.1371835,0.21263443,0.29494452,0.38754338,0.4938606,0.70649505,1.1900668,1.6256244,1.9068506,2.1572106,2.428148,2.311542,2.5584722,3.3266997,4.190956,4.8117113,4.633373,4.7499785,5.470192,6.2864337,6.790583,6.835168,7.2947326,8.56025,10.511685,13.306799,15.944152,17.254255,17.415445,17.936743,0.01371835,0.020577524,0.034295876,0.041155048,0.034295876,0.006859175,0.037725464,0.048014224,0.037725464,0.020577524,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.010288762,0.030866288,0.05144381,0.06516216,0.09259886,0.16119061,0.18862732,0.16119061,0.12689474,0.06859175,0.030866288,0.037725464,0.06516216,0.061732575,0.06516216,0.11317638,0.22292319,0.32924038,0.2709374,0.14061308,0.06859175,0.06516216,0.09602845,0.09259886,0.07888051,0.09602845,0.14747226,0.20920484,0.23664154,0.15090185,0.08916927,0.058302987,0.044584636,0.017147938,0.017147938,0.030866288,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.0548734,0.10288762,0.16804978,0.14404267,0.11317638,0.09945804,0.1097468,0.12689474,0.10288762,0.08916927,0.10288762,0.14747226,0.20920484,0.2469303,0.33266997,0.42526886,0.4938606,0.5418748,0.5007198,0.4046913,0.31552204,0.26750782,0.23664154,0.2777966,0.4424168,0.7442205,1.0906088,1.2723769,1.196926,0.9774324,0.805953,0.7476501,0.7373613,0.77508676,0.8711152,1.0220171,1.214074,1.4267083,1.4404267,1.2723769,1.1454822,1.1523414,1.255229,1.3169615,1.3341095,1.3409687,1.4027013,1.587899,1.5536032,1.371835,1.1111864,0.89169276,0.89855194,0.805953,0.7476501,0.8265306,1.0288762,1.2346514,1.0871792,0.90198153,0.805953,0.77165717,0.64819205,0.5212973,0.4081209,0.31552204,0.2503599,0.22978236,0.20577525,0.1920569,0.17833854,0.17490897,0.17490897,0.15090185,0.12003556,0.09602845,0.082310095,0.05144381,0.09259886,0.14404267,0.18176813,0.18176813,0.12346515,0.14061308,0.13375391,0.12003556,0.12003556,0.14061308,0.30523327,0.58988905,0.91912943,1.2175035,1.4027013,1.0631721,0.72021335,0.44927597,0.34295875,0.5007198,1.471293,1.214074,0.64476246,0.2469303,0.08573969,0.10288762,0.07888051,0.058302987,0.058302987,0.06859175,0.048014224,0.058302987,0.082310095,0.116605975,0.18176813,0.2469303,0.21263443,0.22978236,0.32581082,0.42183927,0.5658819,0.864256,1.097468,1.1832076,1.1763484,1.2106444,1.5158776,2.0268862,2.6304936,3.1552205,3.7039545,4.2698364,4.729401,5.0243454,5.161529,5.4324665,6.0669403,7.051232,8.522525,10.789482,13.457702,15.923574,17.226818,17.339994,17.165085,16.62321,15.951012,15.453721,15.343974,15.738377,15.782962,15.46401,14.839825,14.201921,14.068168,13.776653,13.708061,13.927555,14.647768,16.204802,16.37285,16.112202,15.570327,14.544881,12.504276,12.085866,11.526843,10.477389,9.033533,7.747438,6.9071894,5.693115,4.149801,2.5619018,1.4404267,1.4438564,1.6187652,2.0063086,2.719663,3.9680326,5.3913116,6.025785,6.3824625,6.385892,5.353586,3.3987212,2.7299516,2.784825,2.9906003,2.7402403,1.903421,1.9548649,2.301253,2.5310357,2.393852,2.2841053,2.170929,1.937717,1.5604624,1.1283343,0.7956643,1.1420527,2.1023371,3.5770597,5.4016004,4.8254294,4.90431,4.8117113,4.4447455,4.4241676,4.962613,5.5319247,5.24041,4.431027,4.65395,5.7582774,5.967482,6.169828,6.5882373,6.7802944,6.783724,6.883182,6.5950966,5.7754254,4.636802,4.602506,4.537344,4.506478,4.540774,4.605936,4.7671266,4.9214582,5.597087,6.8969,8.488229,9.705732,10.981539,12.445972,13.581166,13.224489,11.753197,10.113853,8.453933,7.116394,6.6465406,7.0306544,7.9875093,8.615124,8.279024,6.6053853,5.4016004,4.8254294,5.3227196,7.181556,10.501397,13.001566,15.138199,16.153357,16.307688,16.88043,17.881868,17.775553,15.9578705,13.330807,12.322508,11.489118,11.46854,11.8115,12.05157,11.691463,11.739478,11.921246,12.367092,12.912396,13.111313,12.943263,13.2862215,13.858963,14.472859,15.0250225,12.30536,10.847785,10.257896,10.281903,10.799771,11.201033,11.324498,11.245617,10.882081,10.010965,9.163857,8.724871,8.697433,9.071259,9.829198,9.56512,8.923786,8.467651,8.258447,7.888051,7.630832,7.582818,7.133542,6.2144127,5.2781353,4.0503426,3.2512488,3.4844608,4.232111,3.8788633,2.627064,1.8588364,1.3546871,1.0151579,0.8848336,0.64819205,0.85739684,0.8505377,0.4698535,0.037725464,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.030866288,0.030866288,0.024007112,0.017147938,0.020577524,0.041155048,0.034295876,0.01371835,0.006859175,0.0274367,0.06516216,0.058302987,0.0274367,0.0034295875,0.010288762,0.0034295875,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.020577524,0.030866288,0.048014224,0.06859175,0.10288762,0.14747226,0.18176813,0.19891608,0.1920569,0.17490897,0.16462019,0.16804978,0.16462019,0.15776102,0.13032432,0.08573969,0.048014224,0.034295876,0.024007112,0.01371835,0.006859175,0.0,0.0,0.006859175,0.020577524,0.037725464,0.09602845,0.19891608,0.31209245,0.4046913,0.432128,0.53158605,0.82996017,1.1592005,1.4061309,1.5158776,1.6770682,1.7422304,2.2155135,3.2032347,4.4241676,5.2506986,5.6485305,5.9571934,6.385892,7.016936,8.05953,8.652849,9.256456,10.264755,12.010415,15.193072,17.823566,18.897026,18.502625,17.826996,0.010288762,0.020577524,0.044584636,0.05144381,0.0274367,0.0,0.020577524,0.034295876,0.030866288,0.017147938,0.010288762,0.010288762,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.041155048,0.082310095,0.14747226,0.17490897,0.15090185,0.12346515,0.09945804,0.072021335,0.0548734,0.048014224,0.030866288,0.024007112,0.0274367,0.1097468,0.22635277,0.22978236,0.13032432,0.041155048,0.01371835,0.037725464,0.041155048,0.044584636,0.08573969,0.16804978,0.24007112,0.20577525,0.11317638,0.06516216,0.05144381,0.05144381,0.017147938,0.034295876,0.06859175,0.08573969,0.06859175,0.037725464,0.030866288,0.034295876,0.030866288,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.044584636,0.082310095,0.08573969,0.06516216,0.05144381,0.0548734,0.061732575,0.061732575,0.061732575,0.06516216,0.072021335,0.07545093,0.082310095,0.12689474,0.1920569,0.2709374,0.3566771,0.42183927,0.42183927,0.42183927,0.4355576,0.4355576,0.4938606,0.6173257,0.78194594,0.9328478,0.9842916,0.9328478,0.83338976,0.922559,1.155771,1.1832076,1.097468,1.0014396,0.89512235,0.82996017,0.88826317,0.90884066,0.78194594,0.7305021,0.8025235,0.881404,0.881404,0.83338976,0.75450927,0.7305021,0.90884066,0.91569984,0.8093826,0.6962063,0.65505123,0.7613684,0.6241849,0.4424168,0.34638834,0.4389872,0.823101,0.9602845,0.9602845,0.8711152,0.7373613,0.59331864,0.42869842,0.31209245,0.2469303,0.21263443,0.16119061,0.15433143,0.15090185,0.15776102,0.17147937,0.1920569,0.17147937,0.14404267,0.116605975,0.08573969,0.0274367,0.034295876,0.07888051,0.14404267,0.216064,0.28122616,0.274367,0.26750782,0.30523327,0.42526886,0.67219913,1.6942163,2.4898806,2.8877127,2.7745364,2.1126258,1.4164196,0.97400284,0.6962063,0.5144381,0.37725464,0.19891608,0.1097468,0.06516216,0.05144381,0.061732575,0.09259886,0.08573969,0.08916927,0.12346515,0.16462019,0.072021335,0.030866288,0.020577524,0.017147938,0.024007112,0.030866288,0.020577524,0.041155048,0.106317215,0.20234565,0.39097297,0.5693115,0.70649505,0.7990939,0.8779744,0.9877212,1.1420527,1.4369972,1.8828435,2.3972816,2.9288676,3.5290456,3.9337368,4.091498,4.1600895,4.383013,4.8768735,5.4941993,6.416758,8.1384115,10.587136,13.039291,14.7197895,15.4914465,15.834405,15.700651,15.309678,14.87755,14.695783,15.134769,15.512024,15.62863,15.350834,14.904987,14.891269,15.230798,15.71094,16.0539,16.420864,17.412016,18.012194,18.180243,17.662374,16.29397,14.023583,13.101024,12.634601,11.866373,10.744898,9.901219,8.704293,7.1198235,5.295283,3.5770597,2.5070283,2.4212887,2.5481834,2.7711067,3.0969174,3.6319332,3.3747141,3.5187566,3.865145,4.029765,3.4535947,2.5378947,2.1674993,2.3046827,2.6476414,2.6476414,2.5447538,2.5653315,2.6133456,2.620205,2.5378947,3.0660512,3.3061223,3.2821152,2.935727,2.136633,1.5021594,1.7388009,2.7368107,3.9783216,4.554492,3.6593697,3.1346428,2.6647894,2.16064,1.7696671,2.7470996,3.7519686,4.413879,4.4927597,3.8788633,3.6353626,3.6216443,3.8685746,4.3178506,4.835718,5.192395,5.394741,5.302142,4.996909,4.763697,5.4839106,5.627953,5.4804807,5.3090014,5.360445,5.7102633,5.645101,5.8474464,6.5539417,7.5588107,9.304471,11.595435,14.054449,16.112202,17.007324,16.434584,14.538021,12.0309925,9.692014,8.330468,8.944365,11.262765,12.672326,12.243628,10.707172,8.985519,7.4627824,6.773435,7.222711,8.786603,10.840926,13.810948,16.12935,17.257685,17.689812,17.562918,17.21996,15.6526375,13.275933,11.924676,10.995257,11.163307,11.859513,12.46312,12.30193,11.80464,11.153018,11.286773,12.229909,13.114742,13.313659,12.740917,12.421966,12.823228,13.838386,12.994707,11.492548,9.877212,8.718011,8.597976,9.534253,10.38479,11.159878,11.588576,11.146159,10.103564,9.211872,8.573969,8.440215,9.211872,8.97866,8.433355,7.8606143,7.425057,7.181556,7.4627824,7.4765005,7.490219,7.346176,6.444195,4.705394,3.532475,3.1895163,3.4398763,3.532475,3.1415021,2.6853669,2.318401,2.0303159,1.6599203,1.2003556,1.2209331,1.3375391,1.2415106,0.7339317,0.48700142,0.17490897,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.010288762,0.01371835,0.01371835,0.0548734,0.061732575,0.041155048,0.024007112,0.06516216,0.15433143,0.12346515,0.061732575,0.017147938,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.030866288,0.06516216,0.1371835,0.24350071,0.33952916,0.41498008,0.44927597,0.4389872,0.4081209,0.36353627,0.30866286,0.2469303,0.17147937,0.09259886,0.05144381,0.030866288,0.020577524,0.01371835,0.0,0.0,0.0,0.0034295875,0.010288762,0.017147938,0.06859175,0.15090185,0.24350071,0.31552204,0.31209245,0.3566771,0.53158605,0.7613684,0.9534253,0.99801,1.1008976,1.2998136,1.6976458,2.335549,3.1723683,3.8377085,4.6093655,5.271276,5.895461,6.8557453,8.772884,10.813489,12.373952,13.516005,14.96672,17.473747,19.521212,20.436913,20.073376,18.807858,0.0,0.037725464,0.061732575,0.048014224,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.01371835,0.0034295875,0.0,0.0,0.0,0.0034295875,0.024007112,0.0274367,0.01371835,0.01371835,0.034295876,0.061732575,0.106317215,0.12346515,0.09945804,0.0548734,0.041155048,0.048014224,0.034295876,0.020577524,0.020577524,0.044584636,0.0548734,0.030866288,0.006859175,0.0034295875,0.01371835,0.037725464,0.07888051,0.15433143,0.20920484,0.12346515,0.082310095,0.061732575,0.05144381,0.037725464,0.01371835,0.041155048,0.09945804,0.14404267,0.14061308,0.08573969,0.106317215,0.11317638,0.09602845,0.058302987,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0274367,0.041155048,0.05144381,0.061732575,0.06516216,0.07888051,0.09602845,0.10288762,0.11317638,0.15433143,0.22978236,0.33266997,0.4355576,0.5007198,0.5727411,0.6790583,0.72021335,0.66533995,0.5624523,0.5212973,0.6036074,0.9842916,1.4678634,1.4575747,1.2106444,0.9842916,0.8093826,0.65848076,0.4424168,0.39783216,0.4046913,0.4081209,0.4046913,0.42869842,0.48700142,0.5007198,0.4389872,0.33952916,0.31895164,0.33266997,0.33266997,0.30523327,0.30523327,0.45613512,0.432128,0.37725464,0.3806842,0.4972902,0.7613684,0.94999576,0.96371406,0.7888051,0.5453044,0.4629943,0.35324752,0.274367,0.22292319,0.18176813,0.14404267,0.14404267,0.14404267,0.15090185,0.16119061,0.16462019,0.16119061,0.14747226,0.12003556,0.08916927,0.048014224,0.048014224,0.12003556,0.2503599,0.432128,0.66533995,0.59331864,0.5555932,0.66876954,1.0597426,1.8416885,3.99204,5.188966,5.4016004,4.6676683,3.0729103,1.9891608,1.3272504,0.91569984,0.64133286,0.432128,0.24350071,0.12689474,0.061732575,0.030866288,0.017147938,0.041155048,0.06859175,0.14061308,0.26064864,0.37382504,0.15776102,0.058302987,0.024007112,0.017147938,0.01371835,0.030866288,0.020577524,0.020577524,0.05144381,0.116605975,0.28122616,0.4355576,0.607037,0.7956643,0.97400284,1.1214751,1.0734608,1.1694894,1.5055889,1.937717,2.335549,2.9631636,3.3884325,3.5016088,3.4981792,3.4398763,3.6147852,4.105216,5.0757895,6.7940125,9.22902,11.537132,13.272504,14.291091,14.740367,14.565458,14.04759,13.406258,12.915827,12.88496,13.330807,13.876111,14.150477,14.205351,14.507155,15.158776,16.064188,16.647217,16.822126,17.014183,17.370861,17.895588,17.977898,17.401728,16.341984,15.6697855,15.21022,14.167625,12.596875,11.406808,9.932085,8.364764,6.848886,5.5593615,4.695105,4.3041325,4.0057583,3.6010668,3.1380725,2.901431,2.7402403,2.3149714,1.7319417,1.2415106,1.2620882,1.1489118,1.0014396,1.1351935,1.6427724,2.3972816,2.6647894,2.8705647,2.935727,2.9185789,3.0146074,3.5290456,3.858286,3.981751,3.7313912,2.7711067,2.417859,2.8054025,4.122364,5.3844523,4.431027,5.4016004,5.288424,4.6573796,3.858286,3.0214665,4.5853586,5.6313825,6.166398,5.9640527,4.5922174,3.9028704,3.542764,3.5221863,3.7211025,3.8960114,4.256118,4.5442033,4.8117113,5.212973,6.0052075,7.3187394,7.5759587,7.3393173,7.1061053,7.298162,8.080108,8.347616,8.553391,9.026674,10.007536,11.934964,14.483148,16.599203,18.073925,19.521212,20.96164,20.220848,18.145947,15.1862135,11.38966,11.516555,14.606613,16.86671,16.839275,15.402277,14.13333,12.319078,10.377932,8.937505,8.827758,9.4862385,11.732618,14.4145565,16.362562,16.37285,14.942713,14.167625,13.828096,13.437123,12.236768,10.175586,10.062409,11.043272,12.30536,13.070158,13.176475,12.089295,11.574858,12.181894,13.245067,13.834956,12.689473,12.006986,12.542002,13.601744,14.369971,13.63604,11.924676,9.942374,8.580828,8.951223,9.740028,10.751757,11.64345,11.921246,11.526843,10.762046,9.73317,8.844906,8.820899,8.419638,8.008087,7.582818,7.160979,6.776865,6.6568294,6.591667,6.8969,7.205563,6.468202,5.06893,4.081209,3.7862647,3.7965534,3.083199,2.942586,3.3198407,3.3850029,2.8534167,1.9994495,1.6084765,1.5158776,1.762808,2.0714707,1.8691251,1.2483698,0.5212973,0.08573969,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.06516216,0.082310095,0.06516216,0.041155048,0.07888051,0.18519773,0.14747226,0.09259886,0.058302987,0.0274367,0.006859175,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.034295876,0.072021335,0.14404267,0.2503599,0.37382504,0.5007198,0.5761707,0.58988905,0.5693115,0.4938606,0.39783216,0.29494452,0.18862732,0.08916927,0.041155048,0.017147938,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.05144381,0.072021335,0.09602845,0.12346515,0.25378948,0.490431,0.7476501,0.94999576,1.0220171,1.0700313,1.1797781,1.2929544,1.371835,1.4198492,1.5638919,1.9480057,2.6167753,3.642222,5.120374,7.4696417,10.607714,13.3033695,15.241087,17.021042,18.938183,20.910194,22.319756,22.686722,21.664703,0.0,0.09602845,0.11317638,0.06859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.01371835,0.01371835,0.0,0.08573969,0.08916927,0.06516216,0.05144381,0.07545093,0.11317638,0.08573969,0.041155048,0.020577524,0.044584636,0.14404267,0.10288762,0.037725464,0.0,0.0,0.037725464,0.037725464,0.041155048,0.072021335,0.12346515,0.17147937,0.16462019,0.12689474,0.08916927,0.07545093,0.05144381,0.09945804,0.12346515,0.09602845,0.061732575,0.20920484,0.216064,0.16119061,0.09259886,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.024007112,0.024007112,0.01371835,0.01371835,0.0274367,0.06859175,0.1097468,0.15776102,0.24350071,0.31895164,0.37382504,0.42183927,0.4389872,0.36696586,0.31895164,0.31552204,0.37382504,0.44584638,0.39783216,0.3841138,0.42869842,0.53158605,0.58988905,0.3806842,0.4046913,0.42183927,0.37382504,0.26750782,0.18176813,0.32924038,0.40126175,0.33609957,0.19548649,0.18176813,0.35324752,0.45270553,0.432128,0.34638834,0.33609957,0.34638834,0.37039545,0.4046913,0.45613512,0.5178677,0.53158605,0.5796003,0.64133286,0.67219913,0.61046654,0.4389872,0.30523327,0.21263443,0.15433143,0.106317215,0.106317215,0.116605975,0.12346515,0.116605975,0.09259886,0.116605975,0.13032432,0.13032432,0.1097468,0.061732575,0.061732575,0.18862732,0.45270553,0.86082643,1.4335675,1.2758065,1.1249046,1.3101025,2.1126258,3.782835,5.8337283,6.495639,6.200694,5.31929,4.1360826,2.6716487,1.7010754,1.0666018,0.65162164,0.39783216,0.274367,0.16119061,0.082310095,0.041155048,0.030866288,0.041155048,0.044584636,0.07545093,0.14404267,0.22978236,0.06859175,0.020577524,0.020577524,0.0274367,0.01371835,0.041155048,0.017147938,0.0,0.006859175,0.030866288,0.07888051,0.14747226,0.24350071,0.36353627,0.47328308,0.47328308,0.5658819,0.7305021,0.9602845,1.2655178,1.6942163,2.020027,2.5207467,3.1312134,3.450165,2.8259802,2.8088322,3.1723683,3.875434,5.0346346,6.866034,8.532814,9.911508,10.967821,11.749766,12.140739,12.13731,11.873232,11.5645685,11.506266,11.931535,12.343085,12.665466,12.946692,13.337666,14.143619,15.724659,16.993607,17.439453,17.134218,16.245956,15.848124,16.060759,16.647217,17.014183,17.075916,16.907866,16.496315,15.680074,14.1299,12.079007,10.621432,9.345626,8.134981,7.1712675,6.3893213,5.6348124,4.396731,2.9494452,2.3664153,1.8519772,0.90198153,0.38754338,0.490431,0.6859175,0.8093826,0.82996017,0.8676856,1.3992717,3.2649672,3.3747141,3.292404,2.9803114,2.527606,2.136633,1.7833855,1.546744,1.6564908,2.0886188,2.5619018,3.625074,5.6485305,9.702303,14.38026,15.806969,13.9138365,11.382801,10.089847,9.880642,8.573969,8.100685,8.327039,9.084977,9.513676,8.073249,6.924337,6.355026,6.4133286,6.619104,5.936616,5.6793966,5.442755,5.020916,4.7602673,5.5559316,5.871454,6.060081,6.200694,6.5059276,7.3255987,8.093826,9.026674,10.364213,12.264205,14.815818,15.426285,16.859852,18.320856,19.473198,20.460918,22.096832,23.623,24.380938,23.218307,18.492336,17.61436,18.410025,20.755863,22.933651,21.650986,20.735287,17.487467,12.80608,9.156999,10.573419,12.05157,12.394529,12.092726,11.698323,11.794352,11.917816,12.607163,13.399398,13.666906,12.603734,10.209882,9.081548,8.862054,9.211872,9.81205,12.679185,13.149038,12.332796,11.180455,10.497967,10.669447,11.087856,11.729189,12.528283,13.38225,15.261664,16.564907,16.657507,15.162207,11.962401,10.88894,10.621432,10.772334,10.957532,10.772334,10.2236,10.30591,10.401938,10.065839,9.002667,7.2947326,6.6636887,6.3961806,6.142391,5.936616,6.118384,6.495639,6.7185616,6.5779486,5.967482,4.48933,3.724532,3.391862,3.2409601,3.083199,2.9220085,3.1860867,3.1860867,2.7059445,1.9994495,1.5090185,1.3443983,1.6427724,2.1846473,2.3801336,1.5261664,0.90884066,0.3841138,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.01371835,0.01371835,0.030866288,0.030866288,0.017147938,0.06859175,0.12346515,0.1371835,0.07545093,0.0274367,0.006859175,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.01371835,0.006859175,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.0274367,0.0548734,0.09259886,0.116605975,0.13032432,0.15090185,0.17833854,0.21263443,0.23664154,0.22635277,0.18862732,0.1371835,0.07545093,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.037725464,0.061732575,0.13375391,0.29151493,0.6310441,1.0597426,1.2655178,1.2037852,1.097468,1.0014396,0.91912943,0.8093826,0.7476501,0.7510797,0.823101,0.9842916,1.2517995,1.9102802,3.2203827,5.4667625,8.803751,13.258785,17.923023,21.891056,24.717037,25.972265,25.252052,0.0,0.020577524,0.024007112,0.01371835,0.0034295875,0.0,0.010288762,0.01371835,0.006859175,0.0,0.0,0.0,0.0034295875,0.017147938,0.041155048,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.030866288,0.07545093,0.072021335,0.041155048,0.024007112,0.017147938,0.041155048,0.11317638,0.18862732,0.12003556,0.08573969,0.13032432,0.15433143,0.1371835,0.07545093,0.0274367,0.01371835,0.01371835,0.030866288,0.017147938,0.01371835,0.030866288,0.061732575,0.09945804,0.14404267,0.1371835,0.09602845,0.11317638,0.09945804,0.06859175,0.044584636,0.037725464,0.048014224,0.16462019,0.29837412,0.2777966,0.12689474,0.06859175,0.044584636,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.08916927,0.106317215,0.07545093,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.01371835,0.037725464,0.05144381,0.048014224,0.041155048,0.048014224,0.072021335,0.08573969,0.10288762,0.12346515,0.15776102,0.22635277,0.31209245,0.40126175,0.44927597,0.36010668,0.38754338,0.41840968,0.45613512,0.52815646,0.66191036,0.5796003,0.45613512,0.33609957,0.2503599,0.24350071,0.39097297,0.4698535,0.44927597,0.36353627,0.34295875,0.39440256,0.44927597,0.4938606,0.5178677,0.4938606,0.4389872,0.39097297,0.36353627,0.36353627,0.3841138,0.39783216,0.41498008,0.4424168,0.48357183,0.548734,0.52472687,0.41840968,0.28465575,0.17490897,0.15433143,0.1371835,0.14061308,0.19548649,0.31209245,0.4938606,0.75450927,1.0254467,1.1660597,1.0048691,0.34295875,0.19548649,0.23664154,0.4355576,0.75450927,1.1420527,1.646202,2.2566686,2.9288676,3.6216443,4.297273,5.1855364,4.931747,4.122364,3.2649672,2.8054025,2.3149714,1.7799559,1.2586586,0.7956643,0.42183927,0.28808534,0.17490897,0.1097468,0.106317215,0.15090185,0.1371835,0.15433143,0.16462019,0.14747226,0.106317215,0.13375391,0.16119061,0.15433143,0.106317215,0.01371835,0.020577524,0.017147938,0.01371835,0.010288762,0.006859175,0.017147938,0.044584636,0.116605975,0.2469303,0.4355576,0.61046654,0.607037,0.6276145,0.78194594,1.1077567,1.6530612,1.9925903,2.218943,2.352697,2.3389788,2.1640697,2.2292318,2.469303,2.8980014,3.6079261,4.9694724,6.036074,6.90033,7.6445503,8.30646,8.913498,9.1981535,9.544542,10.117283,10.844356,11.410237,11.897239,12.298501,12.6586075,13.080446,13.797231,15.316538,16.918156,18.091074,18.54035,17.463459,16.448301,15.9921665,16.160215,16.575195,16.88043,17.679523,18.389448,18.45461,17.353712,14.29452,12.133881,10.257896,8.453933,6.9037595,5.8371577,4.911169,3.6627994,2.1880767,1.1454822,0.8848336,0.8745448,0.89855194,0.8505377,0.72364295,0.65848076,1.0460242,1.9754424,3.1860867,4.057202,3.5530527,3.6456516,3.8034124,3.7485392,3.4535947,3.0111778,3.1209247,3.216953,3.4673128,4.773986,6.694555,5.6142344,5.003768,6.0737996,7.7748747,9.575408,9.870353,9.585697,9.321619,9.345626,9.571979,8.40249,7.795452,8.152129,8.303031,8.152129,7.3187394,6.3721733,5.6519604,5.2506986,5.2506986,4.9591837,4.616225,4.465323,4.7602673,4.9523244,4.822,4.8185706,5.096367,5.5422134,6.0978065,6.8283086,8.220721,10.220171,12.264205,13.687484,15.059319,16.444872,17.748116,18.728977,19.174824,19.572655,19.757853,19.654966,19.288,19.795578,21.78817,23.924803,26.03057,29.08633,29.782537,26.099161,18.718689,10.731179,7.6445503,7.658269,6.9963584,6.783724,7.363324,8.292743,9.702303,11.63659,13.9309845,15.892709,16.314548,15.162207,13.529722,11.8115,10.669447,11.043272,12.075578,12.445972,12.411677,11.924676,10.655728,9.908078,9.5205345,8.999237,8.772884,10.182446,11.674315,12.689473,13.293081,13.495427,13.245067,12.6586075,12.147599,12.483699,13.505715,14.092175,13.876111,13.155897,11.96926,10.566559,9.403929,8.759167,8.368194,7.6033955,6.3790326,5.164959,4.870014,5.0312047,5.3878818,5.593657,5.195825,4.3658648,3.7348208,3.4227283,3.4398763,3.6799474,3.100347,2.8328393,3.223812,3.758828,3.059192,2.6887965,2.3767042,2.020027,1.6873571,1.5981878,1.4953002,1.3375391,0.9945804,0.53501564,0.23321195,0.09602845,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.010288762,0.030866288,0.048014224,0.048014224,0.044584636,0.037725464,0.01371835,0.006859175,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.010288762,0.01371835,0.010288762,0.0,0.0034295875,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.0274367,0.041155048,0.06859175,0.10288762,0.1371835,0.13375391,0.13375391,0.15433143,0.20234565,0.2469303,0.2469303,0.21263443,0.15776102,0.07545093,0.037725464,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.08573969,0.18862732,0.33609957,0.5555932,0.823101,1.0700313,1.3238207,1.5810398,1.8142518,1.9102802,1.6633499,1.5433143,1.605047,1.7456601,1.8828435,1.9480057,2.0886188,2.3972816,2.983741,3.9646032,5.4599032,7.407909,11.797781,15.110763,17.04848,20.515793,0.010288762,0.0034295875,0.020577524,0.08573969,0.1371835,0.0548734,0.024007112,0.01371835,0.010288762,0.0,0.0,0.006859175,0.010288762,0.020577524,0.037725464,0.037725464,0.030866288,0.0274367,0.034295876,0.048014224,0.0548734,0.034295876,0.017147938,0.030866288,0.06516216,0.06516216,0.024007112,0.024007112,0.044584636,0.06859175,0.06859175,0.09259886,0.061732575,0.0548734,0.09945804,0.14747226,0.12003556,0.07545093,0.030866288,0.006859175,0.006859175,0.010288762,0.0034295875,0.0034295875,0.01371835,0.037725464,0.06516216,0.10288762,0.1097468,0.08916927,0.08573969,0.072021335,0.041155048,0.020577524,0.017147938,0.017147938,0.06859175,0.15776102,0.17490897,0.12003556,0.10288762,0.14404267,0.14747226,0.106317215,0.048014224,0.017147938,0.010288762,0.010288762,0.006859175,0.006859175,0.0274367,0.0274367,0.017147938,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.0034295875,0.0034295875,0.01371835,0.034295876,0.05144381,0.061732575,0.044584636,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.044584636,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0,0.010288762,0.01371835,0.006859175,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.034295876,0.030866288,0.0274367,0.024007112,0.017147938,0.030866288,0.034295876,0.041155048,0.048014224,0.05144381,0.09945804,0.15433143,0.22635277,0.29837412,0.33266997,0.28808534,0.2469303,0.2194936,0.23321195,0.32924038,0.32924038,0.28465575,0.22635277,0.19548649,0.21263443,0.3806842,0.48700142,0.51100856,0.48700142,0.5007198,0.59674823,0.61046654,0.5624523,0.48014224,0.39783216,0.36010668,0.32238123,0.30523327,0.31895164,0.36010668,0.3806842,0.39783216,0.42183927,0.45270553,0.4972902,0.51100856,0.53844523,0.53158605,0.4389872,0.22292319,0.18519773,0.28808534,0.4664239,0.65848076,0.7888051,0.89855194,1.1351935,1.3032433,1.1866373,0.5212973,0.3018037,0.26750782,0.53844523,1.2380811,2.486451,3.4878905,4.4687524,5.2987127,5.857735,6.036074,5.127233,3.9474552,2.8122618,2.0028791,1.7662375,1.5536032,1.3684053,1.2106444,1.0837497,0.9945804,1.1694894,1.0151579,0.70306545,0.3806842,0.16462019,0.13375391,0.15090185,0.17490897,0.15433143,0.06859175,0.08916927,0.09945804,0.08916927,0.061732575,0.034295876,0.020577524,0.010288762,0.017147938,0.041155048,0.06516216,0.0274367,0.020577524,0.07545093,0.216064,0.44584638,0.5761707,0.58302987,0.58302987,0.64819205,0.8025235,1.2209331,1.7216529,2.1297739,2.3321195,2.2806756,2.277246,2.2292318,2.2155135,2.3321195,2.6819375,3.5016088,4.0880685,4.623084,5.2335505,5.970912,6.5642304,7.366754,8.255017,9.105555,9.791472,10.676306,11.341646,11.780633,12.017275,12.099585,12.435684,13.502286,14.918706,16.39,17.689812,18.173384,17.62465,16.911295,16.482597,16.39,16.0539,16.756964,17.79613,18.567787,18.550638,15.9921665,13.937843,11.97269,9.938945,7.936065,6.1972647,4.5784993,3.093488,1.8519772,1.0494537,0.86082643,1.2655178,1.546744,1.3752645,0.7888051,0.7442205,1.1111864,1.8554068,2.7333813,3.2581081,2.651071,2.8637056,3.4295874,4.170378,5.1752477,7.874333,8.927217,9.22216,9.547972,10.607714,12.178465,10.4533825,8.762596,8.700864,10.096705,11.729189,12.079007,11.533703,10.590566,9.839486,9.054111,7.239859,5.9400454,5.7274113,6.1732574,7.0478024,6.8043017,6.0497923,5.2472687,4.695105,4.6916757,4.396731,4.149801,4.105216,4.2252517,4.184097,3.9268777,3.7725463,3.8685746,4.197815,5.2335505,6.101236,7.1266828,8.303031,9.283894,9.729739,10.532263,11.818358,13.540011,15.484588,16.599203,16.925014,16.976458,17.168514,17.826996,19.174824,21.517231,23.400076,24.675882,26.52443,27.556736,26.675331,22.8582,17.29541,13.419975,13.903547,11.324498,9.253027,8.64942,7.874333,7.394191,8.923786,11.667457,14.644339,16.684942,16.345413,15.011304,13.4474125,12.367092,12.449403,13.516005,14.071597,14.195063,13.852104,12.88496,12.120162,11.14273,9.818909,8.621983,8.632272,9.184435,9.592556,10.106995,10.768905,11.4033785,11.211322,10.991828,11.043272,11.290202,11.290202,10.978109,11.074138,10.744898,9.918367,9.266746,9.160428,8.543102,7.8091707,7.1129646,6.3653145,5.2266912,4.5510626,4.4241676,4.6127954,4.602506,4.1635194,3.707384,3.7176728,4.2389703,4.8837323,4.5784993,3.858286,3.6696587,4.0537724,4.149801,4.48933,4.715683,4.1600895,2.9322972,1.9171394,1.5536032,1.4507155,1.3924125,1.2586586,1.0048691,0.548734,0.22978236,0.0548734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07888051,0.041155048,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.034295876,0.13032432,0.19891608,0.09945804,0.0274367,0.030866288,0.017147938,0.010288762,0.01371835,0.020577524,0.024007112,0.01371835,0.0034295875,0.0034295875,0.006859175,0.0034295875,0.0,0.006859175,0.010288762,0.020577524,0.034295876,0.034295876,0.037725464,0.041155048,0.044584636,0.058302987,0.07888051,0.1097468,0.11317638,0.13032432,0.16804978,0.216064,0.26407823,0.26750782,0.22292319,0.14404267,0.06859175,0.037725464,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.030866288,0.037725464,0.0548734,0.12003556,0.22292319,0.3806842,0.58302987,0.8128122,1.0906088,1.3855534,1.6221949,1.728512,1.6393428,1.5844694,1.670209,1.8554068,2.0508933,2.1194851,2.1023371,2.0886188,2.170929,2.4212887,2.877424,3.673088,5.871454,7.7268605,9.355915,12.723769,0.01371835,0.006859175,0.048014224,0.13375391,0.19548649,0.09259886,0.044584636,0.0274367,0.01371835,0.006859175,0.006859175,0.01371835,0.024007112,0.030866288,0.034295876,0.024007112,0.030866288,0.048014224,0.07888051,0.1097468,0.12689474,0.08573969,0.061732575,0.058302987,0.061732575,0.058302987,0.06859175,0.058302987,0.061732575,0.06516216,0.024007112,0.01371835,0.01371835,0.024007112,0.041155048,0.07888051,0.1097468,0.09259886,0.044584636,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.037725464,0.061732575,0.07888051,0.08916927,0.08573969,0.058302987,0.041155048,0.030866288,0.024007112,0.01371835,0.030866288,0.06516216,0.116605975,0.16462019,0.19548649,0.23321195,0.23321195,0.18176813,0.09259886,0.024007112,0.01371835,0.020577524,0.0274367,0.0274367,0.044584636,0.044584636,0.048014224,0.05144381,0.044584636,0.01371835,0.0274367,0.0274367,0.017147938,0.0034295875,0.0,0.01371835,0.010288762,0.010288762,0.017147938,0.020577524,0.030866288,0.030866288,0.0274367,0.020577524,0.010288762,0.010288762,0.010288762,0.006859175,0.0,0.006859175,0.020577524,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.034295876,0.082310095,0.034295876,0.0274367,0.030866288,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.044584636,0.034295876,0.0274367,0.024007112,0.017147938,0.030866288,0.034295876,0.041155048,0.041155048,0.01371835,0.017147938,0.034295876,0.072021335,0.13375391,0.22292319,0.15776102,0.09602845,0.0548734,0.037725464,0.048014224,0.10288762,0.14061308,0.16804978,0.1920569,0.23321195,0.33609957,0.47328308,0.5727411,0.607037,0.5796003,0.64476246,0.6036074,0.5007198,0.3841138,0.31895164,0.29494452,0.2709374,0.26750782,0.29494452,0.34295875,0.36696586,0.40126175,0.48700142,0.66876954,0.99801,0.83338976,0.7922347,0.77508676,0.6893471,0.4355576,0.36353627,0.48357183,0.72021335,0.9945804,1.2209331,1.2655178,1.4918705,1.6564908,1.488441,0.71678376,0.4664239,0.4115505,0.67219913,1.3821237,2.6819375,4.166949,5.3261495,6.1149545,6.492209,6.427047,4.5442033,3.069481,2.0063086,1.3512574,1.0940384,0.96714365,0.922559,0.9431366,1.0254467,1.2037852,1.4781522,1.430138,1.2037852,0.91569984,0.66533995,0.490431,0.36696586,0.28122616,0.22635277,0.18176813,0.24007112,0.216064,0.14061308,0.061732575,0.034295876,0.024007112,0.030866288,0.05144381,0.07545093,0.07545093,0.044584636,0.030866288,0.06859175,0.17490897,0.35324752,0.41840968,0.45613512,0.50757897,0.6001778,0.75450927,1.0220171,1.4404267,1.8142518,2.0165975,1.9857311,1.862266,1.7147937,1.6221949,1.6427724,1.821111,2.4041407,2.8225505,3.2032347,3.6319332,4.1600895,5.0414934,6.217842,7.3839016,8.333898,8.97523,10.161868,11.012405,11.543991,11.794352,11.838936,11.914387,12.487128,13.457702,14.778092,16.441442,17.682953,17.717249,17.189093,16.561478,16.12935,15.659496,16.016174,16.842705,17.826996,18.680964,17.573206,16.184223,14.352823,12.092726,9.595985,7.740579,5.9914894,4.506478,3.350707,2.503599,2.0165975,2.0063086,2.0406046,2.0337453,2.2223728,2.8945718,3.2409601,3.1895163,2.8705647,2.6133456,2.644212,3.1106358,3.8857226,5.195825,7.5931067,12.408247,14.243076,14.359683,13.845244,13.612033,14.582606,13.526293,12.202472,11.859513,13.224489,13.985858,13.588025,12.401388,11.043272,10.39508,9.235879,7.6274023,6.3001523,5.6039457,5.5387836,6.3310184,6.3173003,5.8543057,5.219832,4.623084,4.4927597,4.190956,3.9337368,3.82399,3.8445675,3.6970954,3.4810312,3.3301294,3.3815732,3.7794054,4.863155,5.6656785,6.2830043,6.715132,6.8591747,6.358455,6.4098988,7.023795,8.213862,10.0041065,11.338216,11.808069,11.756626,11.89038,13.2690735,15.244516,17.78927,20.004784,21.397196,21.884197,22.498095,23.1943,22.408924,20.560377,20.056227,22.083115,20.217419,17.645227,15.505165,12.878101,9.925226,9.815479,10.81006,12.315649,14.87755,15.930434,15.693792,14.730078,13.759505,13.653188,14.308239,14.860402,15.354263,15.673215,15.532601,15.114192,14.020154,12.421966,10.731179,9.585697,8.927217,8.4264965,8.320179,8.591117,8.98209,9.081548,9.362774,9.578837,9.4862385,8.827758,8.244728,8.64599,9.078118,9.105555,8.796892,8.635701,7.9772205,7.500508,7.31531,6.9654922,5.7754254,4.7945633,4.2286816,4.1326528,4.3933015,4.190956,3.8857226,3.865145,4.2423997,4.839148,5.5422134,5.40503,5.099797,4.9831905,5.096367,5.6999745,6.2144127,5.977771,4.8322887,3.1243541,2.3321195,1.9720128,1.9274281,1.9651536,1.7113642,1.313532,0.8676856,0.48700142,0.23664154,0.12689474,0.06516216,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07888051,0.041155048,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.037725464,0.15090185,0.22292319,0.106317215,0.024007112,0.030866288,0.024007112,0.01371835,0.010288762,0.01371835,0.017147938,0.010288762,0.006859175,0.0034295875,0.0034295875,0.006859175,0.01371835,0.010288762,0.010288762,0.020577524,0.034295876,0.041155048,0.034295876,0.037725464,0.037725464,0.037725464,0.048014224,0.06516216,0.06859175,0.08573969,0.12003556,0.15433143,0.19548649,0.19891608,0.16462019,0.10288762,0.0548734,0.030866288,0.01371835,0.006859175,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.030866288,0.030866288,0.024007112,0.05144381,0.09259886,0.17490897,0.3018037,0.4389872,0.61389613,0.8025235,0.939707,1.0151579,1.039165,1.0254467,1.0871792,1.2483698,1.4644338,1.6393428,1.7490896,1.8485477,1.9891608,2.177788,2.3972816,2.7093742,3.1380725,3.5873485,4.32128,5.9469047,0.020577524,0.020577524,0.058302987,0.11317638,0.14747226,0.106317215,0.08573969,0.058302987,0.037725464,0.034295876,0.041155048,0.037725464,0.048014224,0.0548734,0.048014224,0.037725464,0.05144381,0.082310095,0.13032432,0.17833854,0.19891608,0.14061308,0.11317638,0.09259886,0.07888051,0.06859175,0.11317638,0.082310095,0.048014224,0.030866288,0.020577524,0.006859175,0.010288762,0.01371835,0.01371835,0.01371835,0.09259886,0.08916927,0.048014224,0.0034295875,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0274367,0.058302987,0.09602845,0.11317638,0.06516216,0.058302987,0.058302987,0.044584636,0.034295876,0.044584636,0.072021335,0.13032432,0.21263443,0.26407823,0.2194936,0.1920569,0.16462019,0.116605975,0.041155048,0.01371835,0.0274367,0.048014224,0.058302987,0.0548734,0.06516216,0.08573969,0.106317215,0.106317215,0.06859175,0.07545093,0.06516216,0.041155048,0.020577524,0.01371835,0.041155048,0.0274367,0.01371835,0.017147938,0.0274367,0.048014224,0.06516216,0.058302987,0.034295876,0.01371835,0.01371835,0.017147938,0.017147938,0.020577524,0.024007112,0.048014224,0.05144381,0.037725464,0.017147938,0.006859175,0.0,0.01371835,0.024007112,0.0274367,0.020577524,0.020577524,0.01371835,0.017147938,0.037725464,0.07888051,0.037725464,0.05144381,0.06516216,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.034295876,0.0548734,0.05144381,0.034295876,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.058302987,0.058302987,0.041155048,0.024007112,0.01371835,0.017147938,0.017147938,0.020577524,0.024007112,0.017147938,0.01371835,0.017147938,0.0274367,0.041155048,0.06859175,0.06516216,0.048014224,0.030866288,0.024007112,0.030866288,0.058302987,0.10288762,0.15776102,0.216064,0.26750782,0.29837412,0.42869842,0.5658819,0.6310441,0.5624523,0.4938606,0.4046913,0.33609957,0.31209245,0.33609957,0.30866286,0.30523327,0.31552204,0.33609957,0.35324752,0.5041494,0.548734,0.64133286,0.939707,1.5947582,1.4507155,1.3341095,1.2003556,1.0048691,0.7305021,0.64819205,0.7442205,0.9774324,1.2963841,1.6496316,1.9274281,2.2292318,2.3801336,2.201795,1.5261664,1.1763484,1.039165,1.0906088,1.3032433,1.6427724,3.0489032,3.99204,4.5201964,4.6916757,4.5682106,3.199805,2.2978237,1.6976458,1.2346514,0.7133542,0.72021335,0.6962063,0.6824879,0.7305021,0.88826317,0.9568549,1.0631721,1.1866373,1.2929544,1.3341095,1.0323058,0.72707254,0.47328308,0.32581082,0.34638834,0.5521636,0.5727411,0.45270553,0.26407823,0.07545093,0.061732575,0.07545093,0.09259886,0.08916927,0.041155048,0.05144381,0.061732575,0.08573969,0.12346515,0.16804978,0.21263443,0.28122616,0.39783216,0.58645946,0.8471081,1.0185875,1.1317638,1.1866373,1.2037852,1.2380811,0.90884066,0.7476501,0.7510797,0.881404,1.08032,1.6873571,2.1297739,2.4041407,2.5550427,2.6476414,3.9303071,5.2575574,6.574519,7.7268605,8.453933,9.897789,11.012405,11.766914,12.199042,12.394529,12.517994,12.836946,13.419975,14.421415,16.108772,16.777542,16.877,16.513464,16.016174,15.940722,16.12935,16.335125,16.678083,17.350283,18.605513,19.085653,18.62266,17.117071,14.726648,11.852654,10.278474,8.923786,7.699424,6.4819202,5.1169443,4.105216,3.549623,3.7176728,4.40359,4.897451,5.874883,6.077229,5.394741,4.1155047,2.9322972,3.8479972,4.588788,5.206114,6.615674,10.587136,15.038741,16.86671,16.407146,14.671775,13.365103,13.72178,13.337666,12.493987,12.0309925,13.361672,13.87954,13.227919,11.852654,10.628291,10.844356,10.22703,9.297611,8.333898,7.4799304,6.7391396,6.468202,6.046363,5.597087,5.178677,4.791134,4.540774,4.2286816,3.8720043,3.57363,3.4844608,3.3952916,3.316411,3.3061223,3.4604537,3.9200184,4.4756117,4.9591837,5.3501563,5.56965,5.4736214,4.846007,4.331569,3.9131594,3.7553983,4.197815,4.8494368,5.3707337,5.2301207,5.1340923,7.016936,9.095266,11.616013,14.404267,16.80498,17.682953,18.04649,18.53692,18.584934,19.188541,22.923363,25.958548,26.908543,25.85566,23.293758,20.155685,16.269962,14.517444,12.874671,11.657167,13.516005,15.927004,17.178804,16.852993,15.608052,15.155347,14.616901,14.79524,15.450292,16.252815,16.767254,16.79469,16.180794,14.987297,13.481709,12.133881,10.477389,9.139851,8.272165,7.846896,7.6376915,7.7920227,8.22758,8.882631,9.331907,8.800322,8.141841,7.7748747,8.038953,8.56368,8.268735,7.699424,7.181556,6.910619,6.7974424,6.4544835,6.0669403,5.5250654,4.846007,4.3109913,4.4721823,4.3933015,4.280125,3.9886103,3.6456516,3.6696587,5.099797,6.4064693,6.9346256,6.684266,6.327589,6.6396813,6.8145905,7.058091,6.9723516,5.5559316,4.5853586,3.4913201,2.8465576,2.6064866,2.1126258,2.020027,1.6599203,1.1660597,0.6962063,0.4081209,0.23664154,0.07888051,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.06516216,0.09259886,0.048014224,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.010288762,0.0034295875,0.0034295875,0.01371835,0.024007112,0.0034295875,0.0,0.0034295875,0.01371835,0.024007112,0.01371835,0.020577524,0.024007112,0.020577524,0.034295876,0.030866288,0.020577524,0.020577524,0.030866288,0.041155048,0.058302987,0.06516216,0.058302987,0.048014224,0.037725464,0.017147938,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0274367,0.020577524,0.024007112,0.044584636,0.07545093,0.1371835,0.19891608,0.25721905,0.3018037,0.30866286,0.2777966,0.3018037,0.39097297,0.5555932,0.7922347,1.097468,1.4095604,1.6907866,1.9102802,2.0646117,2.2326615,2.352697,2.3218307,2.2395205,2.428148,0.044584636,0.034295876,0.048014224,0.07888051,0.12003556,0.16804978,0.16804978,0.11317638,0.08916927,0.11317638,0.1371835,0.12346515,0.11317638,0.09602845,0.08573969,0.12346515,0.19548649,0.20577525,0.22292319,0.26064864,0.26064864,0.17490897,0.106317215,0.06516216,0.041155048,0.030866288,0.017147938,0.024007112,0.037725464,0.044584636,0.044584636,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.08916927,0.07545093,0.0274367,0.05144381,0.06859175,0.058302987,0.044584636,0.010288762,0.0,0.037725464,0.09259886,0.09259886,0.017147938,0.0,0.048014224,0.12689474,0.15090185,0.0548734,0.020577524,0.034295876,0.06859175,0.09259886,0.14061308,0.09602845,0.09602845,0.16462019,0.21263443,0.10288762,0.048014224,0.037725464,0.05144381,0.07545093,0.05144381,0.0274367,0.01371835,0.01371835,0.01371835,0.0274367,0.048014224,0.06859175,0.07545093,0.07545093,0.07545093,0.08573969,0.09259886,0.08573969,0.061732575,0.024007112,0.08916927,0.12003556,0.07888051,0.030866288,0.006859175,0.072021335,0.12689474,0.13032432,0.106317215,0.106317215,0.06859175,0.034295876,0.017147938,0.030866288,0.017147938,0.024007112,0.024007112,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.16462019,0.274367,0.21263443,0.15090185,0.09602845,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.06516216,0.07545093,0.072021335,0.061732575,0.037725464,0.030866288,0.024007112,0.017147938,0.030866288,0.0548734,0.05144381,0.044584636,0.044584636,0.044584636,0.06859175,0.06859175,0.0548734,0.041155048,0.030866288,0.07888051,0.09259886,0.09259886,0.09602845,0.12346515,0.31895164,0.31895164,0.29494452,0.34295875,0.48700142,0.39097297,0.3018037,0.25378948,0.26407823,0.33609957,0.34638834,0.4424168,0.5212973,0.548734,0.548734,1.196926,1.2106444,0.97400284,0.77508676,0.823101,1.8245405,2.3321195,2.3321195,1.8279701,0.84024894,0.8745448,1.1763484,1.5090185,1.6770682,1.5398848,2.335549,2.568761,2.6853669,3.0626216,4.029765,3.309552,2.7711067,2.393852,2.1434922,1.9823016,1.5090185,1.2243627,1.1077567,1.1249046,1.2346514,1.7113642,2.1057668,2.1743584,1.6770682,0.39783216,0.53158605,0.72021335,0.8711152,0.88826317,0.65505123,0.51100856,0.44584638,0.47671264,0.6241849,0.9294182,0.9431366,0.78194594,0.53158605,0.31209245,0.274367,0.66533995,0.9259886,1.0014396,0.8196714,0.31895164,0.19891608,0.10288762,0.041155048,0.0274367,0.07545093,0.08916927,0.12689474,0.17147937,0.16804978,0.044584636,0.06859175,0.17833854,0.33609957,0.4698535,0.45613512,0.53158605,0.5418748,0.51100856,0.5555932,0.8848336,0.70306545,0.5555932,0.5418748,0.70306545,1.0082988,1.4472859,1.6564908,1.6496316,1.5501735,1.587899,2.4795918,3.9200184,5.7479887,7.366754,7.720001,9.513676,11.207891,12.404818,12.871242,12.542002,12.956982,13.481709,14.116182,15.217079,17.487467,17.70696,17.065628,15.88242,15.138199,16.479168,17.271402,17.600643,17.490896,17.580065,19.11995,20.19341,20.591244,19.857311,17.96761,15.319967,13.1593275,11.547421,10.429376,9.403929,7.706283,6.4098988,6.866034,9.544542,11.670886,7.2158523,5.360445,4.695105,4.65395,4.65395,4.105216,4.9214582,5.528495,5.4187484,6.608815,13.625751,16.592344,17.106783,16.194511,15.148488,15.501736,14.733508,13.543441,12.761495,12.566009,12.4802685,12.88496,13.059869,12.754636,11.88352,10.528833,9.575408,8.906639,8.200144,7.373613,6.591667,5.675967,4.852866,4.479041,4.4859004,4.3624353,4.1429415,3.8514268,3.474172,3.1072063,2.959734,2.9494452,3.000889,3.0729103,3.1860867,3.4192986,3.7108135,4.040054,4.461893,4.8905916,5.096367,4.9248877,4.4516044,3.642222,2.8054025,2.609916,3.0969174,3.7862647,3.9165888,3.3781435,2.7299516,3.415869,4.8322887,7.1026754,9.613133,11.015835,12.641459,14.493437,16.609491,18.79757,20.62897,21.729866,23.046827,23.533829,22.793037,21.071384,19.459478,18.087645,16.688372,15.786391,16.678083,18.190533,20.52951,21.249723,19.963629,18.341434,17.463459,17.003895,15.96816,14.63062,14.5585985,15.13134,15.621771,15.638919,14.977009,13.612033,11.828648,10.449953,9.434795,8.711152,8.162418,7.857185,7.31531,7.3873315,8.155559,8.9100685,8.886061,7.682276,7.4113383,8.172707,8.025234,7.2192817,6.385892,6.0395036,6.1972647,6.392751,6.601956,6.560801,5.950334,4.9831905,4.4104495,4.3624353,4.695105,4.73969,4.256118,3.4638834,3.2821152,5.56965,7.425057,8.073249,8.865483,9.170717,8.549961,8.64256,9.595985,10.086417,9.1810055,6.4579134,4.2835546,3.2821152,2.318401,1.9651536,1.786815,1.5158776,1.1180456,0.7613684,0.5418748,0.19548649,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.034295876,0.044584636,0.034295876,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.020577524,0.010288762,0.0034295875,0.01371835,0.0274367,0.041155048,0.044584636,0.041155048,0.01371835,0.01371835,0.05144381,0.11317638,0.19548649,0.30523327,0.5144381,0.6824879,0.82996017,0.96714365,1.1146159,1.6496316,2.0063086,2.1880767,2.3081124,2.5619018,0.3018037,0.22292319,0.16119061,0.14747226,0.216064,0.4115505,0.4115505,0.34295875,0.24350071,0.16804978,0.17490897,0.26064864,0.28465575,0.24350071,0.17147937,0.15776102,0.2503599,0.274367,0.20920484,0.116605975,0.1371835,0.13032432,0.10288762,0.06516216,0.034295876,0.041155048,0.09945804,0.14404267,0.13032432,0.07888051,0.06859175,0.0548734,0.044584636,0.044584636,0.048014224,0.041155048,0.0274367,0.0274367,0.0274367,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.024007112,0.041155048,0.0274367,0.006859175,0.024007112,0.0274367,0.01371835,0.020577524,0.044584636,0.07888051,0.12003556,0.14747226,0.12689474,0.08573969,0.05144381,0.037725464,0.034295876,0.030866288,0.030866288,0.044584636,0.05144381,0.08916927,0.2503599,0.28122616,0.13032432,0.030866288,0.05144381,0.09259886,0.15776102,0.3018037,0.31895164,0.20920484,0.17490897,0.13032432,0.072021335,0.044584636,0.05144381,0.05144381,0.06516216,0.072021335,0.06516216,0.058302987,0.07545093,0.09602845,0.08916927,0.06516216,0.048014224,0.061732575,0.17147937,0.4046913,0.50757897,0.4355576,0.34638834,0.274367,0.16119061,0.09259886,0.08573969,0.082310095,0.082310095,0.07545093,0.05144381,0.0274367,0.030866288,0.037725464,0.048014224,0.044584636,0.024007112,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.024007112,0.07545093,0.116605975,0.12346515,0.16804978,0.15776102,0.07888051,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.024007112,0.037725464,0.037725464,0.030866288,0.030866288,0.030866288,0.0274367,0.030866288,0.024007112,0.024007112,0.020577524,0.024007112,0.034295876,0.0274367,0.034295876,0.034295876,0.030866288,0.017147938,0.048014224,0.14404267,0.29837412,0.47671264,0.59674823,0.4424168,0.37039545,0.33609957,0.31552204,0.30523327,0.36353627,0.3806842,0.41840968,0.5178677,0.6790583,0.7476501,0.7099246,0.6241849,0.53501564,0.47671264,0.72364295,0.84367853,0.85396725,0.78537554,0.6790583,0.7510797,0.7922347,0.9568549,1.3169615,1.8416885,1.2998136,1.2689474,1.3786942,1.3615463,1.0528834,1.2312219,1.1934965,1.1317638,1.2003556,1.5398848,1.7250825,1.5981878,1.3238207,1.0460242,0.89855194,0.6962063,0.6036074,0.5796003,0.58645946,0.58988905,0.8779744,1.4678634,1.9548649,1.8554068,0.59331864,0.41498008,0.34981793,0.34981793,0.37382504,0.37382504,0.36696586,0.5041494,0.7305021,0.9259886,0.91912943,0.91227025,0.7442205,0.5041494,0.34638834,0.50757897,0.72021335,0.764798,0.66533995,0.5555932,0.65162164,0.6241849,0.4972902,0.28465575,0.106317215,0.17490897,0.24350071,0.32238123,0.3841138,0.3841138,0.24007112,0.216064,0.22978236,0.2709374,0.32238123,0.34638834,0.3806842,0.4046913,0.41840968,0.45956472,0.6036074,0.91912943,1.1523414,1.1763484,0.96714365,0.6173257,0.6344737,0.72707254,0.8093826,0.86082643,0.9294182,1.3786942,2.2120838,3.5290456,5.1169443,6.427047,8.261876,10.14129,11.869802,12.929544,12.4802685,12.253916,12.418536,13.317088,14.887839,16.681513,17.075916,16.698662,15.96816,15.580616,16.503176,17.521763,18.228258,18.091074,17.851004,19.486916,21.983656,24.319204,24.970827,23.451519,20.323736,17.734396,16.023033,14.661487,13.426835,12.394529,10.971251,9.115844,7.8846216,7.6274023,7.9875093,8.405919,7.5759587,6.601956,5.8337283,4.8734436,5.4667625,7.870903,11.756626,15.477728,16.091625,14.390549,13.845244,13.155897,12.267634,12.377381,12.555719,12.394529,12.360233,12.449403,12.188754,11.869802,11.941824,11.533703,10.542552,9.637141,8.762596,7.442205,6.509357,6.1458206,5.871454,5.4153185,4.479041,3.758828,3.474172,3.3644254,3.3987212,3.3232703,3.093488,2.7779658,2.5447538,2.4555845,2.4590142,2.6304936,2.9185789,3.1620796,3.2786856,3.5942078,3.8891523,4.016047,3.9131594,3.508468,3.333559,3.1346428,2.8568463,2.6819375,2.6716487,2.877424,3.216953,3.5942078,3.9028704,4.1189346,4.65395,5.223262,5.6828265,6.060081,6.8557453,7.795452,9.451943,11.7086115,13.7938,14.171056,16.832415,19.137098,20.36832,21.743584,21.764162,21.002794,21.294308,22.220297,21.109112,18.091074,19.44919,20.718138,19.912186,17.549198,15.429714,14.771234,14.572317,14.441993,14.592895,15.059319,15.011304,15.011304,15.237658,15.501736,13.749216,12.349944,11.207891,10.261326,9.458802,8.879202,7.6651278,6.725421,6.543653,7.2021337,7.548522,7.599966,7.64798,7.6171136,7.051232,6.7802944,6.200694,5.6313825,5.288424,5.271276,6.0532217,6.077229,5.579939,4.863155,4.2869844,4.3452873,5.23698,6.1972647,6.550512,5.6965446,4.5167665,4.523626,5.0449233,5.861165,7.191845,9.695444,10.607714,10.816919,11.365653,13.454271,15.090185,13.344524,9.623423,5.874883,4.5784993,3.1586502,2.201795,1.5810398,1.1249046,0.6036074,0.77508676,0.7510797,0.5555932,0.26407823,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.010288762,0.01371835,0.020577524,0.034295876,0.044584636,0.034295876,0.020577524,0.010288762,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.017147938,0.0274367,0.044584636,0.0548734,0.041155048,0.048014224,0.06516216,0.09259886,0.12346515,0.14747226,0.17833854,0.20234565,0.22635277,0.26407823,0.33266997,0.58645946,0.89169276,1.2689474,1.7113642,2.1743584,0.3018037,0.3566771,0.29151493,0.23321195,0.25721905,0.37382504,0.39440256,0.28808534,0.216064,0.23321195,0.28465575,0.26064864,0.28122616,0.31209245,0.33609957,0.33266997,0.24007112,0.19548649,0.1371835,0.08573969,0.116605975,0.18519773,0.16462019,0.106317215,0.058302987,0.0548734,0.07545093,0.09259886,0.07888051,0.0548734,0.058302987,0.09602845,0.1097468,0.11317638,0.116605975,0.12003556,0.12003556,0.12689474,0.116605975,0.07888051,0.010288762,0.030866288,0.030866288,0.034295876,0.058302987,0.09945804,0.041155048,0.024007112,0.034295876,0.041155048,0.006859175,0.0,0.006859175,0.006859175,0.0034295875,0.01371835,0.10288762,0.13375391,0.13032432,0.10288762,0.06516216,0.048014224,0.034295876,0.020577524,0.0034295875,0.0,0.010288762,0.024007112,0.0274367,0.041155048,0.12346515,0.28122616,0.274367,0.18862732,0.1097468,0.116605975,0.18176813,0.29151493,0.33609957,0.2777966,0.17147937,0.1371835,0.11317638,0.08916927,0.07545093,0.08916927,0.09259886,0.082310095,0.06516216,0.044584636,0.041155048,0.09259886,0.13375391,0.12003556,0.06859175,0.041155048,0.10288762,0.2777966,0.34638834,0.28122616,0.22635277,0.24350071,0.2469303,0.20920484,0.15433143,0.17833854,0.21263443,0.22292319,0.16804978,0.082310095,0.06859175,0.06516216,0.072021335,0.058302987,0.024007112,0.006859175,0.006859175,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.010288762,0.030866288,0.07888051,0.14061308,0.16462019,0.14747226,0.10288762,0.05144381,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.034295876,0.048014224,0.06516216,0.061732575,0.058302987,0.058302987,0.06859175,0.06859175,0.07545093,0.072021335,0.072021335,0.11317638,0.19548649,0.216064,0.18176813,0.12003556,0.07888051,0.14747226,0.22978236,0.30866286,0.37039545,0.41498008,0.37725464,0.31209245,0.274367,0.2777966,0.28808534,0.26750782,0.31209245,0.39783216,0.50757897,0.65162164,0.8196714,0.65848076,0.4389872,0.3018037,0.26407823,0.32581082,0.38754338,0.42869842,0.432128,0.40126175,0.37725464,0.37039545,0.5453044,0.97400284,1.6496316,1.6564908,1.6564908,1.5707511,1.3341095,0.922559,1.0425946,0.96714365,0.7990939,0.6310441,0.5590228,0.8265306,0.864256,0.7990939,0.7339317,0.7613684,0.7373613,0.7339317,0.84024894,1.1729189,1.8725548,1.7216529,1.5844694,1.3924125,1.0563129,0.45613512,0.5178677,0.53158605,0.50757897,0.4664239,0.45956472,0.4355576,0.4664239,0.5212973,0.5521636,0.4938606,0.5041494,0.4972902,0.5007198,0.5590228,0.7305021,0.7305021,0.64476246,0.5212973,0.4698535,0.6310441,0.7133542,0.71678376,0.65162164,0.5418748,0.4081209,0.3566771,0.39440256,0.5521636,0.7613684,0.85739684,0.6379033,0.36696586,0.21263443,0.20234565,0.2469303,0.2709374,0.30866286,0.34638834,0.42183927,0.607037,0.8265306,0.9602845,0.9877212,0.88826317,0.61046654,0.4664239,0.39097297,0.4115505,0.52472687,0.70649505,1.1008976,1.7456601,2.7779658,4.0880685,5.3158607,6.9620624,8.98209,11.211322,13.13189,13.848674,14.675205,16.03675,16.904436,17.051908,17.082775,16.753534,16.410576,16.431154,16.897577,17.600643,18.293419,19.023922,19.737276,20.577524,21.894485,23.372639,24.998262,25.745913,25.351511,24.284908,23.256033,21.53095,19.682402,18.28656,17.940172,17.826996,14.935853,11.694893,9.489669,8.628842,8.186425,8.608265,8.793462,8.597976,8.848335,11.201033,12.05843,13.687484,15.909856,16.077906,14.613472,13.6086035,12.346515,10.868362,9.959522,10.343636,10.611144,10.655728,10.364213,9.626852,8.838047,8.800322,8.872343,8.81404,8.772884,7.9909387,6.8043017,5.8543057,5.3398676,5.0312047,4.9694724,4.5613513,4.1635194,3.9028704,3.6970954,3.4878905,3.1380725,2.6819375,2.1846473,1.7456601,1.605047,1.6324836,1.8005334,2.020027,2.1469216,2.2978237,2.620205,2.959734,3.2032347,3.2683969,2.959734,2.7162333,2.4384367,2.0989075,1.7662375,1.5947582,1.6736387,2.0165975,2.5619018,3.1620796,3.9200184,4.32471,4.3590055,4.32128,4.8322887,4.3624353,4.372724,5.171818,6.7048435,8.549961,9.054111,10.847785,12.857523,14.894698,17.662374,17.278261,17.021042,18.224829,20.70785,22.793037,21.829325,22.710728,24.741043,25.917393,22.933651,18.598652,15.422854,13.745787,13.540011,14.38369,15.553179,16.444872,17.240536,17.669235,17.000465,15.227368,13.718349,12.641459,11.746337,10.367643,9.410788,8.31332,7.1232533,6.341307,6.893471,7.414768,7.7680154,7.8846216,7.6788464,7.0443726,6.615674,6.025785,5.4187484,5.0414934,5.209543,5.830299,6.029215,5.7651367,5.1752477,4.5956473,4.5339146,5.1409516,6.355026,7.6342616,7.966932,7.7131424,7.5039372,6.783724,6.0154963,6.6739774,9.719451,12.977559,14.88098,15.419425,16.12935,16.678083,16.719238,14.119612,9.637141,6.910619,5.055212,3.9474552,2.860276,1.6427724,0.7373613,0.7888051,0.9294182,0.881404,0.607037,0.29151493,0.13032432,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.0,0.0,0.01371835,0.020577524,0.0274367,0.030866288,0.037725464,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0034295875,0.010288762,0.010288762,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.006859175,0.01371835,0.030866288,0.05144381,0.06859175,0.06516216,0.07545093,0.082310095,0.09602845,0.11317638,0.106317215,0.09602845,0.09259886,0.09945804,0.106317215,0.1097468,0.17490897,0.30866286,0.5041494,0.7407909,0.96714365,0.2709374,0.40126175,0.39440256,0.39440256,0.4081209,0.32238123,0.29151493,0.17490897,0.15090185,0.23664154,0.28465575,0.20920484,0.20234565,0.2709374,0.35324752,0.34638834,0.18519773,0.1097468,0.08916927,0.09259886,0.116605975,0.17833854,0.15776102,0.116605975,0.07888051,0.072021335,0.06516216,0.048014224,0.030866288,0.030866288,0.058302987,0.12003556,0.1371835,0.1371835,0.14404267,0.16119061,0.18519773,0.19891608,0.18519773,0.13375391,0.044584636,0.048014224,0.05144381,0.07545093,0.116605975,0.15433143,0.082310095,0.05144381,0.072021335,0.116605975,0.116605975,0.1097468,0.058302987,0.01371835,0.0034295875,0.020577524,0.12346515,0.14747226,0.12003556,0.061732575,0.010288762,0.010288762,0.010288762,0.006859175,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.010288762,0.16462019,0.24350071,0.216064,0.13375391,0.12346515,0.20920484,0.23664154,0.2503599,0.2469303,0.18862732,0.18519773,0.1920569,0.16804978,0.116605975,0.08916927,0.08916927,0.07545093,0.05144381,0.0274367,0.010288762,0.05144381,0.09602845,0.10288762,0.06516216,0.024007112,0.034295876,0.12003556,0.15090185,0.116605975,0.12346515,0.18862732,0.26750782,0.26750782,0.20577525,0.18862732,0.22978236,0.2469303,0.20920484,0.13032432,0.09602845,0.07545093,0.072021335,0.0548734,0.0274367,0.01371835,0.01371835,0.01371835,0.017147938,0.024007112,0.0274367,0.024007112,0.017147938,0.030866288,0.06859175,0.12689474,0.14404267,0.09602845,0.0548734,0.044584636,0.044584636,0.06859175,0.10288762,0.12346515,0.12689474,0.116605975,0.08573969,0.048014224,0.0274367,0.034295876,0.048014224,0.072021335,0.07888051,0.07888051,0.09602845,0.15090185,0.20920484,0.216064,0.26407823,0.35324752,0.42526886,0.4424168,0.4424168,0.37382504,0.25721905,0.17147937,0.20920484,0.2503599,0.2709374,0.28122616,0.31209245,0.42869842,0.4938606,0.48357183,0.41840968,0.37725464,0.33609957,0.34981793,0.4629943,0.64133286,0.7682276,0.6824879,0.4698535,0.26750782,0.14404267,0.11317638,0.1371835,0.15776102,0.22978236,0.37725464,0.5658819,0.70306545,0.70306545,0.7682276,0.980862,1.3409687,1.4610043,1.4644338,1.4027013,1.3203912,1.2449403,1.5947582,1.471293,1.1077567,0.6893471,0.34981793,0.50757897,0.548734,0.5624523,0.607037,0.7339317,0.70649505,0.7099246,0.8676856,1.3238207,2.2635276,1.7799559,1.2517995,0.7613684,0.4115505,0.28808534,0.47671264,0.59674823,0.64476246,0.6379033,0.607037,0.5521636,0.45956472,0.34295875,0.2503599,0.25721905,0.34981793,0.4424168,0.5178677,0.5658819,0.5658819,0.48357183,0.4698535,0.5796003,0.8093826,1.0940384,1.1626302,1.1351935,1.1283343,1.1420527,1.08032,0.91912943,0.78194594,0.77851635,0.90541106,1.0597426,0.91227025,0.7579388,0.7990939,0.9534253,0.85739684,0.65162164,0.4698535,0.4046913,0.47328308,0.61389613,0.66191036,0.6756287,0.69963586,0.7339317,0.72021335,0.64819205,0.53501564,0.48700142,0.5590228,0.7613684,1.1111864,1.5981878,2.318401,3.223812,4.1155047,5.453044,7.332458,9.640571,12.017275,13.841815,15.704081,18.135658,19.514353,19.490345,18.999914,18.420315,19.03764,20.313446,21.654415,22.415783,22.463799,22.223726,22.518671,23.386356,24.089422,24.466677,25.097721,25.632736,25.955118,26.1849,25.76649,24.384367,22.683292,21.256582,20.656404,20.893047,18.687822,15.9613,13.625751,11.588576,10.127572,10.542552,11.0981455,11.38623,12.308789,13.725209,12.795791,12.315649,13.3033695,14.990726,14.13333,12.788932,11.063849,9.1981535,7.5416627,7.706283,8.052671,8.172707,7.8503256,7.0752387,6.2864337,6.1149545,6.341307,6.800872,7.363324,7.023795,6.3721733,5.641671,4.98662,4.513337,4.5682106,4.5682106,4.4996185,4.3795834,4.273266,3.8857226,3.4295874,2.976882,2.5138876,1.9514352,1.6770682,1.5741806,1.5570327,1.5398848,1.4369972,1.488441,1.6942163,2.0680413,2.4898806,2.7059445,2.6407824,2.4590142,2.1091962,1.6496316,1.2586586,1.0666018,1.0734608,1.2620882,1.6153357,2.1126258,3.1072063,3.707384,3.9303071,3.9851806,4.2698364,3.2786856,2.7985435,2.8739944,3.5564823,4.931747,5.6828265,6.5710897,7.73029,9.325048,11.523414,11.38623,12.240198,14.016724,16.599203,19.833303,20.920483,22.44322,25.893385,29.693369,29.206367,25.444109,21.832754,19.723558,18.934752,17.744686,18.722118,18.526632,18.269413,18.060207,17.014183,15.937293,14.421415,13.502286,13.118172,12.106443,10.950673,10.213311,9.14328,7.9017696,7.5519514,7.2467184,7.3427467,7.5210853,7.56224,7.3427467,6.8454566,6.2898636,5.768566,5.435896,5.4770513,5.4633327,5.6245236,5.658819,5.4907694,5.2918534,5.641671,5.686256,6.2864337,7.64798,9.328478,10.792912,11.324498,10.686595,9.379922,8.639131,10.796341,13.872682,15.659496,15.3817,13.704632,13.841815,14.832966,13.828096,10.864933,8.879202,7.6376915,6.5882373,5.188966,3.457024,1.9651536,1.4232788,1.1420527,0.9431366,0.7613684,0.6241849,0.37725464,0.18519773,0.058302987,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.006859175,0.01371835,0.017147938,0.017147938,0.017147938,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.006859175,0.01371835,0.010288762,0.006859175,0.0034295875,0.01371835,0.024007112,0.034295876,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.017147938,0.017147938,0.024007112,0.020577524,0.0034295875,0.0,0.006859175,0.030866288,0.061732575,0.082310095,0.08916927,0.09259886,0.07888051,0.07888051,0.08916927,0.082310095,0.07545093,0.07888051,0.082310095,0.082310095,0.06859175,0.0548734,0.06859175,0.09259886,0.116605975,0.1371835,0.274367,0.31895164,0.38754338,0.50757897,0.58302987,0.38754338,0.24007112,0.14061308,0.1371835,0.1920569,0.19548649,0.17147937,0.14747226,0.17490897,0.22635277,0.19891608,0.12346515,0.082310095,0.08573969,0.1097468,0.116605975,0.10288762,0.09602845,0.09945804,0.10288762,0.10288762,0.09945804,0.06859175,0.034295876,0.024007112,0.06516216,0.1097468,0.11317638,0.116605975,0.13375391,0.15090185,0.17833854,0.1920569,0.1920569,0.16804978,0.10288762,0.061732575,0.07545093,0.116605975,0.15433143,0.14404267,0.12003556,0.09945804,0.14404267,0.24350071,0.31895164,0.29151493,0.15090185,0.037725464,0.01371835,0.037725464,0.09945804,0.11317638,0.09259886,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.048014224,0.06516216,0.072021335,0.072021335,0.22978236,0.24350071,0.21263443,0.19891608,0.24350071,0.23664154,0.25378948,0.24007112,0.17147937,0.06859175,0.058302987,0.048014224,0.030866288,0.01371835,0.0,0.0,0.0,0.01371835,0.0274367,0.020577524,0.044584636,0.082310095,0.09945804,0.09945804,0.13375391,0.19548649,0.22978236,0.23664154,0.20577525,0.13032432,0.13032432,0.14061308,0.15090185,0.14747226,0.106317215,0.07888051,0.06516216,0.05144381,0.037725464,0.037725464,0.037725464,0.030866288,0.030866288,0.041155048,0.05144381,0.044584636,0.034295876,0.0274367,0.037725464,0.072021335,0.072021335,0.06516216,0.061732575,0.06516216,0.08916927,0.20577525,0.34981793,0.41840968,0.39097297,0.33266997,0.28465575,0.20920484,0.12346515,0.061732575,0.0548734,0.06859175,0.07545093,0.08573969,0.13032432,0.25721905,0.37725464,0.39097297,0.490431,0.6824879,0.764798,0.64476246,0.6173257,0.5693115,0.4629943,0.35324752,0.2777966,0.2469303,0.2709374,0.35324752,0.5007198,0.6893471,0.8265306,0.7990939,0.64133286,0.5144381,0.548734,0.5453044,0.65848076,0.85739684,0.94656616,0.5693115,0.4115505,0.32238123,0.24350071,0.18519773,0.24350071,0.34981793,0.5624523,0.8745448,1.2243627,1.4198492,1.2517995,1.0734608,1.0460242,1.1420527,0.84367853,0.7682276,0.881404,1.1489118,1.5398848,2.0474637,1.862266,1.3615463,0.8196714,0.4115505,0.48700142,0.45613512,0.40126175,0.3806842,0.45613512,0.35324752,0.34295875,0.44927597,0.69963586,1.1317638,0.66876954,0.40126175,0.3018037,0.28808534,0.2503599,0.34981793,0.47671264,0.58988905,0.64819205,0.59674823,0.53844523,0.4355576,0.31209245,0.22978236,0.2777966,0.4424168,0.5144381,0.4664239,0.31895164,0.17147937,0.14747226,0.28465575,0.64133286,1.1420527,1.5981878,1.587899,1.4335675,1.3581166,1.4575747,1.7182233,1.6599203,1.4472859,1.1283343,0.8265306,0.7442205,0.8196714,1.039165,1.5021594,1.9342873,1.7182233,1.2483698,0.7407909,0.4938606,0.52472687,0.5418748,0.58302987,0.6173257,0.64476246,0.6962063,0.85396725,0.97057325,0.9602845,0.91912943,0.91912943,1.0185875,1.2106444,1.4164196,1.728512,2.1983654,2.819121,3.806842,5.377593,7.442205,9.784613,12.037852,14.054449,16.753534,19.157675,20.78673,21.674994,21.990515,24.11,26.455837,28.126047,28.904564,28.208357,26.36324,24.953678,24.572994,24.809635,25.210897,25.69104,26.26378,26.83995,27.203487,25.893385,24.806206,23.657295,22.395206,21.191422,20.406046,19.637817,18.79071,17.840714,16.822126,15.138199,13.9309845,13.214201,13.022143,13.409687,11.777204,10.484249,10.285333,11.38623,13.419975,11.993267,10.353925,8.64599,7.006647,5.5730796,5.3673043,5.501058,5.7274113,5.8337283,5.6348124,5.2575574,5.003768,4.9214582,5.099797,5.638242,5.7994323,5.6485305,5.2609873,4.7499785,4.266407,4.2081037,4.2252517,4.1943855,4.166949,4.3521466,4.15323,3.9680326,3.9200184,3.8479972,3.316411,2.8328393,2.5138876,2.2635276,1.9925903,1.6359133,1.3855534,1.3341095,1.5844694,2.0063086,2.2258022,2.4144297,2.4658735,2.2463799,1.8348293,1.5124481,1.2998136,1.2037852,1.2106444,1.3409687,1.6427724,2.3458378,3.2272418,3.8788633,4.0503426,3.6696587,3.000889,2.5001693,2.0920484,1.9994495,2.726522,3.4227283,4.098357,4.7088237,5.2781353,5.8988905,6.81802,9.009526,11.334786,13.289652,14.997586,15.87213,18.245405,22.683292,28.204927,32.299854,32.43704,30.739393,29.59391,28.59247,24.51469,24.329493,21.503513,18.735836,17.28169,16.952452,16.897577,15.412566,14.280802,14.068168,14.119612,13.251926,12.775213,11.921246,10.511685,8.985519,7.380472,6.975781,7.1849856,7.606825,8.014946,7.8434668,7.380472,6.790583,6.307011,6.210983,5.871454,5.9914894,6.042933,5.970912,6.2144127,7.2467184,7.0306544,6.715132,7.239859,9.349055,12.027563,13.529722,14.174485,13.841815,11.965831,12.325937,12.761495,12.764925,11.664027,8.625413,9.462232,10.127572,10.2921915,10.254466,10.933525,10.947243,10.1652975,8.793462,7.023795,5.0106273,3.549623,2.294394,1.4987297,1.1592005,1.0048691,0.7956643,0.59674823,0.39097297,0.21263443,0.13032432,0.048014224,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.006859175,0.0034295875,0.0,0.0,0.0,0.0034295875,0.017147938,0.041155048,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0034295875,0.01371835,0.034295876,0.041155048,0.037725464,0.0274367,0.01371835,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.010288762,0.020577524,0.030866288,0.037725464,0.048014224,0.0548734,0.0548734,0.041155048,0.020577524,0.006859175,0.0034295875,0.024007112,0.0548734,0.07888051,0.09602845,0.082310095,0.0548734,0.037725464,0.037725464,0.037725464,0.037725464,0.037725464,0.030866288,0.024007112,0.024007112,0.017147938,0.01371835,0.006859175,0.0,0.0,0.21263443,0.09259886,0.13375391,0.274367,0.4355576,0.53501564,0.33952916,0.22635277,0.17833854,0.18176813,0.24350071,0.2194936,0.20577525,0.19891608,0.19891608,0.19891608,0.12346515,0.09602845,0.10288762,0.12689474,0.15090185,0.12689474,0.12346515,0.12689474,0.14061308,0.15090185,0.12689474,0.08573969,0.037725464,0.0034295875,0.01371835,0.041155048,0.09259886,0.13375391,0.15090185,0.1371835,0.1371835,0.1371835,0.15433143,0.17833854,0.15090185,0.14061308,0.17490897,0.18519773,0.16804978,0.16804978,0.1920569,0.20920484,0.26407823,0.35324752,0.42869842,0.35324752,0.16119061,0.041155048,0.037725464,0.061732575,0.08573969,0.044584636,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.061732575,0.20920484,0.30866286,0.34638834,0.31895164,0.24350071,0.1097468,0.14061308,0.18176813,0.16804978,0.106317215,0.044584636,0.030866288,0.024007112,0.01371835,0.0,0.0,0.0,0.01371835,0.034295876,0.044584636,0.058302987,0.041155048,0.030866288,0.024007112,0.0,0.15776102,0.22635277,0.23321195,0.216064,0.22978236,0.16804978,0.13375391,0.12346515,0.12003556,0.106317215,0.12003556,0.11317638,0.09602845,0.072021335,0.061732575,0.061732575,0.061732575,0.061732575,0.06516216,0.07545093,0.08916927,0.082310095,0.07545093,0.09602845,0.18176813,0.18176813,0.14747226,0.09602845,0.06516216,0.07545093,0.37039545,0.71678376,0.84024894,0.69963586,0.5041494,0.5658819,0.6173257,0.4629943,0.18862732,0.15090185,0.12689474,0.09602845,0.09945804,0.17147937,0.30523327,0.41498008,0.4698535,0.4938606,0.5212973,0.59674823,0.66876954,0.70649505,0.77851635,0.85396725,0.7922347,0.61046654,0.42869842,0.32238123,0.37725464,0.67219913,1.039165,0.7613684,0.53158605,0.5658819,0.6241849,0.6379033,0.77851635,0.77165717,0.6036074,0.5178677,0.823101,0.84367853,0.75450927,0.66191036,0.6241849,0.66191036,1.0666018,1.4918705,1.7730967,1.9068506,1.920569,1.2998136,0.6962063,0.42183927,0.45613512,0.53158605,0.6241849,0.70306545,0.7476501,0.7476501,0.881404,0.86082643,0.7510797,0.607037,0.47328308,0.31552204,0.20920484,0.14404267,0.09945804,0.07545093,0.11317638,0.15776102,0.19548649,0.18176813,0.044584636,0.06859175,0.13032432,0.20920484,0.29837412,0.39783216,0.6036074,0.72021335,0.70649505,0.5590228,0.29151493,0.20577525,0.17490897,0.16804978,0.15433143,0.106317215,0.14404267,0.17147937,0.14061308,0.1097468,0.24350071,0.26750782,0.26407823,0.28465575,0.34295875,0.42869842,0.5144381,0.58988905,0.64476246,0.75450927,1.0837497,1.5227368,1.8897027,1.6633499,0.96371406,0.548734,0.34295875,0.34638834,0.6207553,1.0220171,1.2037852,1.0460242,0.59674823,0.32581082,0.37382504,0.5178677,0.66533995,0.72021335,0.77508676,0.89169276,1.097468,1.2826657,1.3992717,1.4610043,1.4815818,1.4953002,1.5193073,1.3992717,1.3375391,1.4404267,1.7079345,2.3424082,3.8857226,5.9914894,8.292743,10.39165,11.684605,14.188204,17.21653,20.320305,23.300617,25.6053,27.85854,29.494452,30.286688,30.334702,28.990303,26.26721,23.983105,23.11542,23.773901,25.385807,26.43869,27.481285,28.863409,30.732533,28.877127,26.956558,25.413242,24.548986,24.535269,22.961088,21.925352,21.407484,21.37319,21.78817,19.62753,17.130789,14.644339,12.737488,12.175035,11.249047,11.228469,11.808069,12.199042,11.122152,9.414218,7.8434668,6.4579134,5.5490727,5.645101,5.1580997,4.6779575,4.448175,4.6093655,5.219832,5.3398676,5.223262,5.0003386,4.773986,4.6402316,4.4550343,4.262977,4.0880685,3.923448,3.7553983,3.6559403,3.532475,3.309552,3.1792276,3.5702004,3.9371665,4.173808,4.664239,5.147811,4.746549,4.1360826,3.8720043,3.6593697,3.333559,2.867135,2.3424082,1.9823016,1.8485477,1.9548649,2.2738166,2.627064,2.7059445,2.5241764,2.1743584,1.8313997,1.5364552,1.3992717,1.4198492,1.5913286,1.9239986,2.6545007,3.8445675,4.6573796,4.8288593,4.6676683,4.2183924,3.7485392,2.8122618,1.7113642,1.4815818,1.6873571,2.16064,2.6545007,3.0317552,3.2512488,3.6525106,5.9331865,8.964942,12.212761,15.717799,16.191082,17.19938,19.572655,23.671013,29.35727,34.045513,32.7457,31.298416,31.387585,30.533617,29.799686,27.26522,23.996824,21.311457,20.735287,20.45406,18.746124,16.187653,14.009865,14.085316,14.328816,13.865822,13.176475,12.377381,11.231899,9.705732,8.793462,8.718011,9.283894,9.856634,10.2236,9.637141,8.330468,7.3221693,8.405919,9.345626,10.175586,9.328478,7.3839016,7.0786686,7.798882,8.217292,8.004657,7.579388,8.117833,10.034973,12.397959,14.033872,14.29795,13.077017,11.550851,10.381361,10.621432,11.444533,10.161868,9.417647,9.239308,10.55284,12.88839,14.387119,15.083325,15.21365,14.29795,12.4802685,10.528833,8.06296,5.778855,4.0949273,2.9322972,1.7250825,1.5055889,1.4850113,1.3752645,1.0700313,0.65505123,0.24007112,0.072021335,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.044584636,0.106317215,0.058302987,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.0548734,0.05144381,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.030866288,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.024007112,0.030866288,0.0274367,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.010288762,0.0274367,0.048014224,0.061732575,0.08573969,0.09259886,0.07888051,0.0548734,0.030866288,0.017147938,0.01371835,0.01371835,0.020577524,0.044584636,0.034295876,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.0,0.0,0.0,0.26407823,0.18862732,0.22978236,0.25721905,0.2469303,0.2777966,0.28808534,0.30523327,0.3018037,0.26407823,0.20920484,0.13375391,0.13032432,0.12689474,0.1097468,0.09945804,0.09602845,0.09945804,0.10288762,0.09259886,0.07888051,0.06516216,0.061732575,0.072021335,0.09259886,0.10288762,0.08916927,0.072021335,0.048014224,0.020577524,0.0034295875,0.006859175,0.024007112,0.044584636,0.0548734,0.05144381,0.082310095,0.08916927,0.106317215,0.14404267,0.18862732,0.18519773,0.20920484,0.2194936,0.19891608,0.13032432,0.116605975,0.12346515,0.14404267,0.16462019,0.15776102,0.11317638,0.0548734,0.034295876,0.07888051,0.18176813,0.15776102,0.08573969,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.10288762,0.26750782,0.3566771,0.274367,0.16804978,0.12003556,0.13375391,0.15776102,0.18176813,0.216064,0.22978236,0.16804978,0.058302987,0.017147938,0.0034295875,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.024007112,0.044584636,0.037725464,0.017147938,0.006859175,0.006859175,0.01371835,0.072021335,0.1097468,0.11317638,0.10288762,0.09602845,0.10288762,0.106317215,0.1097468,0.11317638,0.13032432,0.15433143,0.17147937,0.18176813,0.17490897,0.13375391,0.11317638,0.1097468,0.12346515,0.15776102,0.20920484,0.20234565,0.17147937,0.13375391,0.12346515,0.17147937,0.19891608,0.17147937,0.106317215,0.058302987,0.08916927,0.15776102,0.24350071,0.29837412,0.32238123,0.3806842,0.4424168,0.45613512,0.38754338,0.26750782,0.20234565,0.20577525,0.25378948,0.37725464,0.48357183,0.35324752,0.33609957,0.41840968,0.5555932,0.6824879,0.71678376,0.72364295,0.70649505,0.7442205,0.8128122,0.78194594,0.65505123,0.48014224,0.31895164,0.24007112,0.32924038,0.48014224,0.432128,0.41498008,0.48014224,0.5041494,0.45613512,0.53844523,0.50757897,0.37725464,0.4081209,0.70306545,0.96371406,1.2449403,1.4918705,1.5536032,1.2689474,1.5227368,1.7216529,1.6496316,1.4918705,1.5055889,1.0254467,0.5727411,0.3806842,0.39783216,0.36353627,0.36696586,0.42869842,0.53844523,0.6756287,0.7099246,0.6207553,0.48357183,0.34638834,0.24007112,0.13032432,0.09259886,0.082310095,0.082310095,0.07545093,0.044584636,0.044584636,0.0548734,0.06516216,0.058302987,0.32581082,0.44927597,0.45613512,0.4081209,0.39783216,0.37039545,0.31895164,0.24007112,0.15433143,0.082310095,0.06516216,0.07545093,0.09602845,0.11317638,0.082310095,0.061732575,0.058302987,0.05144381,0.058302987,0.13375391,0.16804978,0.2194936,0.32581082,0.4389872,0.42869842,0.51100856,0.69963586,0.9294182,1.1592005,1.3512574,1.7319417,2.3252604,2.6133456,2.301253,1.3306799,0.4115505,0.17490897,0.34295875,0.64819205,0.8505377,0.91569984,0.84367853,0.71678376,0.6001778,0.53158605,0.5212973,0.5212973,0.66533995,0.91912943,1.097468,1.0666018,1.0940384,1.3272504,1.7147937,2.020027,1.8382589,1.5433143,1.3238207,1.2723769,1.3546871,1.5810398,2.6887965,4.3658648,6.3447366,8.412778,9.911508,12.723769,16.12249,19.634388,23.03311,25.056566,25.859089,25.6053,24.487255,22.731306,22.734735,21.61326,20.37175,19.905325,21.013083,23.44466,25.27606,26.713057,28.078033,29.779108,30.42387,30.358707,29.655643,28.68507,28.136335,25.965406,23.749893,21.819035,20.845032,21.825895,19.637817,16.63007,13.742357,11.941824,12.250486,12.277924,12.329367,12.284782,11.928105,10.9541025,9.585697,8.172707,7.0375133,6.3790326,6.279575,5.9400454,5.377593,4.839148,4.506478,4.5099077,4.5442033,4.530485,4.4275975,4.249259,4.064061,3.841138,3.5461934,3.4776018,3.5976372,3.532475,3.2992632,3.059192,3.000889,3.175798,3.508468,3.7691166,3.8034124,4.0434837,4.4859004,4.695105,4.8082814,4.4550343,4.0263357,3.707384,3.4673128,3.3129816,3.2889743,3.391862,3.57363,3.7142432,3.6182148,3.5359046,3.3266997,2.942586,2.417859,1.8416885,1.529596,1.5193073,1.8073926,2.3629858,2.4487255,3.5016088,5.0449233,6.776865,8.56368,6.245279,4.945465,4.5819287,4.1360826,1.6393428,1.4953002,1.5227368,1.8965619,2.5241764,3.0043187,3.3301294,4.081209,5.2747054,7.5279446,12.065289,14.514014,16.184223,17.556059,19.411465,22.813616,25.920822,27.374968,27.289227,27.35096,30.801125,32.99949,33.054363,31.946608,30.749681,30.622786,29.806545,27.59789,23.70188,19.363451,17.353712,17.802988,19.425184,18.886738,16.0539,13.989287,12.188754,11.207891,10.6488695,10.185875,9.589127,8.930646,8.021805,7.0032177,6.200694,6.125243,6.56766,8.14527,9.369633,9.73317,9.692014,8.529384,8.080108,7.6171136,7.1061053,7.2021337,8.4264965,9.914937,10.861504,10.823778,9.719451,8.916927,8.110974,7.630832,7.4353456,7.1095347,9.22902,10.439664,11.938394,14.188204,16.938732,17.29541,17.12393,16.506605,15.649208,14.898128,13.944703,12.260776,10.405369,8.80718,7.7680154,5.5730796,4.4996185,4.3795834,4.605936,4.122364,2.9940298,1.5947582,0.50757897,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.058302987,0.048014224,0.0274367,0.12003556,0.13032432,0.082310095,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.041155048,0.11317638,0.18176813,0.20234565,0.12689474,0.15090185,0.16462019,0.15433143,0.11317638,0.024007112,0.0034295875,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.006859175,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.017147938,0.017147938,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.024007112,0.01371835,0.020577524,0.034295876,0.048014224,0.061732575,0.09602845,0.12003556,0.12003556,0.10288762,0.07888051,0.058302987,0.037725464,0.024007112,0.020577524,0.034295876,0.13032432,0.12003556,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.3018037,0.28465575,0.29151493,0.2709374,0.22635277,0.23321195,0.2777966,0.33266997,0.36353627,0.34981793,0.2709374,0.22292319,0.20577525,0.16462019,0.09259886,0.058302987,0.0548734,0.07545093,0.10288762,0.12003556,0.08916927,0.0548734,0.030866288,0.024007112,0.037725464,0.06516216,0.05144381,0.041155048,0.037725464,0.037725464,0.0274367,0.01371835,0.006859175,0.024007112,0.0548734,0.07545093,0.11317638,0.09945804,0.09602845,0.12689474,0.18176813,0.216064,0.22635277,0.2194936,0.18862732,0.13032432,0.09259886,0.07888051,0.08573969,0.08916927,0.072021335,0.037725464,0.030866288,0.041155048,0.061732575,0.09602845,0.15433143,0.1371835,0.09945804,0.058302987,0.017147938,0.010288762,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.048014224,0.07888051,0.116605975,0.17490897,0.30523327,0.32238123,0.25721905,0.17147937,0.17147937,0.19548649,0.20577525,0.19891608,0.17147937,0.1097468,0.048014224,0.01371835,0.0034295875,0.010288762,0.01371835,0.0034295875,0.0,0.0034295875,0.006859175,0.017147938,0.01371835,0.0034295875,0.006859175,0.024007112,0.041155048,0.072021335,0.08573969,0.09945804,0.12003556,0.15090185,0.18519773,0.20577525,0.19891608,0.17147937,0.17490897,0.22635277,0.22635277,0.216064,0.20577525,0.17147937,0.12346515,0.17490897,0.22978236,0.2469303,0.22635277,0.15433143,0.11317638,0.08573969,0.082310095,0.10288762,0.1097468,0.10288762,0.08916927,0.08573969,0.12689474,0.14061308,0.13375391,0.1371835,0.17147937,0.2503599,0.33952916,0.38754338,0.3841138,0.34981793,0.31552204,0.30523327,0.36696586,0.5178677,0.70306545,0.7888051,0.7442205,0.7442205,0.8093826,0.96371406,1.214074,1.2106444,1.097468,1.0254467,0.99801,0.8779744,0.7407909,0.6173257,0.53844523,0.52472687,0.6207553,0.6790583,0.6173257,0.5590228,0.52472687,0.42869842,0.31552204,0.31552204,0.83338976,1.728512,2.294394,2.2429502,1.4575747,1.1249046,1.430138,1.529596,1.1317638,1.2895249,1.4781522,1.4610043,1.2895249,1.0425946,0.7922347,0.61046654,0.53158605,0.52815646,0.5178677,0.6927767,0.86082643,0.9431366,0.96714365,1.0220171,0.97057325,0.8093826,0.548734,0.20920484,0.09259886,0.044584636,0.030866288,0.030866288,0.041155048,0.0274367,0.058302987,0.106317215,0.15433143,0.17147937,0.22292319,0.23664154,0.22292319,0.216064,0.26750782,0.21263443,0.14061308,0.072021335,0.0274367,0.041155048,0.030866288,0.030866288,0.041155048,0.048014224,0.041155048,0.024007112,0.0274367,0.044584636,0.06859175,0.06859175,0.07888051,0.11317638,0.18862732,0.2709374,0.26407823,0.28122616,0.35324752,0.47328308,0.61389613,0.70649505,0.8676856,1.1180456,1.2689474,1.1832076,0.77508676,0.39440256,0.2709374,0.3841138,0.64819205,0.89855194,1.1317638,1.3512574,1.4507155,1.430138,1.3958421,1.4267083,1.3032433,1.1900668,1.1489118,1.1351935,1.2758065,1.3238207,1.4438564,1.670209,1.8862731,1.9411465,1.8005334,1.6427724,1.5604624,1.5673214,1.471293,2.0268862,3.0557625,4.420738,6.0052075,7.9429245,10.199594,12.740917,15.772673,19.713268,21.990515,22.94737,22.847912,22.093403,21.232576,21.236006,20.546658,19.44919,18.509483,18.567787,20.53637,22.597551,24.401514,25.862518,27.134895,28.067743,28.530739,28.541027,28.27352,28.067743,26.85367,25.228045,23.310905,21.61326,21.03023,19.03078,16.496315,14.123041,12.4974165,12.120162,11.766914,11.173596,10.408798,9.599416,8.940934,8.443645,7.8434668,7.281014,6.848886,6.584808,6.310441,6.1492505,5.8474464,5.363875,4.8734436,4.372724,4.2183924,4.190956,4.170378,4.149801,4.0194764,3.8171308,3.7005248,3.673088,3.5702004,3.4844608,3.3438478,3.223812,3.1277838,2.9906003,3.3472774,3.357566,3.292404,3.2649672,3.2272418,3.9474552,4.0503426,3.8960114,3.7725463,3.9200184,4.297273,4.629943,4.9523244,5.4187484,6.307011,6.166398,5.809721,5.284994,4.5819287,3.642222,2.7333813,2.07833,1.7559488,1.8965619,2.6922262,3.000889,3.6765177,4.8151407,6.3618846,8.128122,6.800872,5.188966,4.413879,4.273266,3.2066643,3.1655092,1.9411465,1.4335675,2.1674993,3.309552,3.625074,4.1429415,4.636802,5.597087,8.23444,10.744898,12.809509,14.493437,16.62664,20.814167,22.967947,24.799347,25.228045,25.063425,27.01486,29.950588,30.434158,30.272968,30.615927,31.943178,34.09696,32.296425,28.486153,24.463247,21.87048,22.20315,23.256033,23.201159,21.85333,20.70099,19.603521,16.496315,12.843805,10.151579,9.9801,10.000677,9.22902,7.922347,6.4819202,5.470192,5.363875,6.3035817,7.579388,8.457363,8.176137,7.051232,6.4716315,6.2041235,6.2075534,6.6431108,7.4799304,8.532814,9.637141,10.247607,9.431366,8.529384,7.579388,6.9071894,6.81802,7.6205435,8.937505,9.170717,10.425946,12.830087,14.54831,15.175924,16.208231,16.846134,16.842705,16.496315,15.563468,13.831526,12.05157,10.604284,9.513676,7.846896,6.848886,6.433906,6.3001523,5.9331865,5.3227196,3.683377,2.0680413,0.9911508,0.4115505,0.082310095,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.030866288,0.020577524,0.010288762,0.048014224,0.058302987,0.037725464,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.08916927,0.14747226,0.18862732,0.14404267,0.14061308,0.15433143,0.16804978,0.14404267,0.10288762,0.08916927,0.07888051,0.0548734,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.037725464,0.037725464,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.006859175,0.006859175,0.0034295875,0.0034295875,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.037725464,0.05144381,0.06516216,0.06516216,0.061732575,0.061732575,0.058302987,0.07545093,0.09259886,0.10288762,0.09945804,0.09602845,0.106317215,0.12003556,0.13032432,0.12689474,0.1097468,0.072021335,0.041155048,0.020577524,0.010288762,0.020577524,0.06859175,0.061732575,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.31895164,0.34638834,0.29837412,0.2469303,0.23664154,0.274367,0.37382504,0.38754338,0.37039545,0.33952916,0.26407823,0.24007112,0.21263443,0.15433143,0.07888051,0.034295876,0.041155048,0.058302987,0.08573969,0.10288762,0.07545093,0.048014224,0.024007112,0.01371835,0.020577524,0.044584636,0.05144381,0.048014224,0.041155048,0.034295876,0.041155048,0.020577524,0.010288762,0.020577524,0.048014224,0.07545093,0.09945804,0.07888051,0.08573969,0.1371835,0.216064,0.26750782,0.25721905,0.21263443,0.16462019,0.14404267,0.12003556,0.12003556,0.11317638,0.09259886,0.061732575,0.024007112,0.037725464,0.05144381,0.061732575,0.106317215,0.26750782,0.30523327,0.2469303,0.14404267,0.041155048,0.020577524,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.0548734,0.09259886,0.12003556,0.12003556,0.20577525,0.28808534,0.29151493,0.2194936,0.15090185,0.18519773,0.19891608,0.17147937,0.1097468,0.048014224,0.030866288,0.020577524,0.0274367,0.034295876,0.01371835,0.006859175,0.006859175,0.0034295875,0.0,0.006859175,0.024007112,0.041155048,0.041155048,0.034295876,0.041155048,0.058302987,0.072021335,0.08916927,0.1097468,0.14061308,0.16119061,0.18862732,0.2194936,0.23664154,0.23664154,0.26064864,0.23321195,0.20577525,0.1920569,0.17833854,0.14404267,0.19548649,0.23321195,0.22292319,0.17147937,0.106317215,0.07888051,0.06516216,0.058302987,0.06859175,0.058302987,0.06859175,0.09945804,0.15776102,0.23321195,0.2194936,0.18519773,0.15776102,0.15090185,0.17833854,0.26407823,0.33609957,0.4081209,0.48700142,0.6001778,0.6344737,0.88826317,1.2277923,1.4644338,1.3375391,1.3101025,1.2517995,1.1866373,1.2037852,1.4472859,1.5433143,1.5330256,1.488441,1.3958421,1.1523414,1.0185875,0.99801,1.0871792,1.2003556,1.1626302,1.1077567,0.97400284,0.7510797,0.5007198,0.34638834,0.37382504,0.58988905,1.3958421,2.49331,2.867135,2.469303,1.5570327,1.155771,1.3889829,1.4747226,1.2209331,1.2689474,1.2963841,1.1797781,1.0014396,0.8093826,0.7990939,0.7956643,0.7510797,0.7613684,0.980862,1.1146159,1.1694894,1.1523414,1.0837497,1.0906088,0.99801,0.8128122,0.548734,0.22978236,0.1097468,0.05144381,0.034295876,0.048014224,0.09602845,0.17833854,0.20234565,0.18176813,0.15433143,0.15090185,0.072021335,0.0274367,0.017147938,0.044584636,0.116605975,0.08916927,0.058302987,0.034295876,0.0274367,0.041155048,0.0274367,0.020577524,0.01371835,0.017147938,0.0274367,0.030866288,0.037725464,0.05144381,0.058302987,0.041155048,0.048014224,0.07545093,0.116605975,0.15776102,0.17147937,0.16119061,0.14747226,0.14404267,0.17147937,0.25378948,0.36696586,0.4389872,0.48014224,0.51100856,0.5658819,0.6344737,0.66876954,0.8128122,1.0837497,1.3581166,1.5810398,1.8999915,2.1263442,2.2052248,2.201795,2.1434922,1.9925903,1.821111,1.6976458,1.6599203,1.6907866,1.7010754,1.7216529,1.7525192,1.7696671,1.9891608,2.0303159,2.0097382,2.0131679,2.0886188,1.9651536,2.1846473,2.6922262,3.433017,4.3624353,5.9914894,7.449064,9.050681,11.375941,15.265094,17.833855,19.476627,20.262003,20.587814,21.177702,21.342323,20.995934,20.059656,18.866161,18.176813,19.301718,21.085104,22.77932,23.986534,24.662163,25.01884,25.19032,25.26234,25.348082,25.59501,25.61559,25.084003,24.147726,23.063976,22.20658,21.187992,19.469769,17.556059,15.762384,14.21564,12.771784,11.321068,9.993818,8.937505,8.30646,7.949784,7.5450926,7.14726,6.8145905,6.608815,6.3378778,6.341307,6.2658563,5.9880595,5.593657,4.938606,4.671098,4.588788,4.557922,4.5339146,4.465323,4.273266,4.0057583,3.7108135,3.474172,3.3781435,3.2203827,2.983741,2.74367,2.6785078,3.192946,3.3884325,3.309552,3.1037767,3.0043187,3.7348208,4.081209,4.1189346,4.149801,4.705394,5.4496145,6.0223556,6.447624,7.016936,8.268735,8.707723,8.841476,8.443645,7.431916,5.871454,4.187526,3.1072063,2.5207467,2.4624438,3.093488,3.7108135,4.372724,5.223262,6.2864337,7.455923,7.0478024,5.7754254,4.9523244,4.996909,5.422178,5.8680243,3.8960114,2.2120838,1.9754424,2.7813954,3.2135234,3.7794054,4.180667,4.5784993,5.5902276,7.1678376,8.899779,10.669447,12.977559,16.94902,18.845583,20.580954,21.541239,22.158566,23.893936,26.047716,26.418112,26.521,27.460707,29.971165,33.630535,33.49335,31.709965,29.42929,26.795366,25.965406,25.084003,24.298628,23.914513,24.391226,24.398085,21.019941,16.163645,12.113303,11.509696,11.382801,10.703742,9.56512,8.210432,7.051232,6.276145,6.0497923,6.4887795,7.2124224,7.3701835,7.4970784,6.6876955,5.950334,5.8645945,6.5779486,7.7851634,8.793462,9.853205,10.569988,9.89436,8.488229,7.8949103,7.64798,7.6925645,8.364764,8.947794,8.522525,9.012956,10.511685,11.245617,11.873232,13.327377,14.7026415,15.656067,16.396858,15.580616,14.119612,12.548861,10.981539,9.105555,8.381912,7.8537555,7.3598948,6.866034,6.4579134,6.121814,4.8288593,3.3026927,1.9823016,1.0048691,0.39440256,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0274367,0.048014224,0.041155048,0.0274367,0.01371835,0.017147938,0.041155048,0.061732575,0.082310095,0.09602845,0.13375391,0.18519773,0.21263443,0.14061308,0.09602845,0.07545093,0.072021335,0.082310095,0.030866288,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.030866288,0.030866288,0.020577524,0.01371835,0.01371835,0.024007112,0.010288762,0.017147938,0.034295876,0.05144381,0.0548734,0.044584636,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.01371835,0.010288762,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.006859175,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.006859175,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.010288762,0.024007112,0.044584636,0.06859175,0.09945804,0.1097468,0.1097468,0.106317215,0.09945804,0.13375391,0.15433143,0.16119061,0.15090185,0.13375391,0.12346515,0.11317638,0.1097468,0.10288762,0.08573969,0.05144381,0.0274367,0.010288762,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0034295875,0.006859175,0.017147938,0.01371835,0.0034295875,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.26407823,0.3018037,0.22292319,0.16119061,0.18176813,0.26750782,0.432128,0.4046913,0.32581082,0.26750782,0.21263443,0.18519773,0.14747226,0.10288762,0.061732575,0.020577524,0.05144381,0.0548734,0.048014224,0.037725464,0.030866288,0.030866288,0.0274367,0.030866288,0.037725464,0.048014224,0.08916927,0.09602845,0.06516216,0.024007112,0.024007112,0.01371835,0.01371835,0.01371835,0.01371835,0.0274367,0.0274367,0.020577524,0.058302987,0.14747226,0.25378948,0.3018037,0.2777966,0.21263443,0.15433143,0.16462019,0.18176813,0.20577525,0.18519773,0.12003556,0.06859175,0.037725464,0.0548734,0.06859175,0.10288762,0.22978236,0.4081209,0.4355576,0.34981793,0.20577525,0.08573969,0.0548734,0.034295876,0.017147938,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.020577524,0.06516216,0.12003556,0.16804978,0.15433143,0.17490897,0.20234565,0.19891608,0.08916927,0.1371835,0.16119061,0.14747226,0.09602845,0.034295876,0.020577524,0.030866288,0.048014224,0.0548734,0.024007112,0.024007112,0.020577524,0.017147938,0.017147938,0.037725464,0.06859175,0.09259886,0.072021335,0.0274367,0.0274367,0.030866288,0.05144381,0.058302987,0.041155048,0.0274367,0.030866288,0.0548734,0.13032432,0.22635277,0.23664154,0.19548649,0.16462019,0.15433143,0.15776102,0.17147937,0.18519773,0.17147937,0.15090185,0.14061308,0.13375391,0.14747226,0.14061308,0.13032432,0.12346515,0.12346515,0.116605975,0.12346515,0.16462019,0.24007112,0.33266997,0.30523327,0.28465575,0.25378948,0.21263443,0.18862732,0.25721905,0.36353627,0.5041494,0.6893471,0.9294182,1.0460242,1.5398848,2.1194851,2.3972816,1.8862731,1.8725548,1.8245405,1.670209,1.4644338,1.371835,1.5776103,1.7833855,1.903421,1.8485477,1.5398848,1.4678634,1.5055889,1.6359133,1.728512,1.5193073,1.3615463,1.2277923,0.9431366,0.6173257,0.64133286,0.88826317,1.3306799,1.8176813,2.0749004,1.7079345,1.2175035,1.1694894,1.3032433,1.4369972,1.4815818,1.4678634,1.430138,1.2106444,0.8676856,0.66876954,0.8162418,1.0288762,1.1043272,1.0425946,1.0425946,1.4335675,1.3375391,1.1454822,1.0254467,0.9328478,0.7305021,0.5212973,0.3566771,0.26407823,0.25721905,0.17833854,0.16119061,0.17147937,0.19548649,0.21263443,0.34981793,0.31209245,0.17490897,0.034295876,0.017147938,0.017147938,0.006859175,0.0,0.006859175,0.017147938,0.0034295875,0.010288762,0.030866288,0.048014224,0.0274367,0.020577524,0.017147938,0.020577524,0.024007112,0.041155048,0.0548734,0.061732575,0.048014224,0.030866288,0.041155048,0.07888051,0.12346515,0.16119061,0.18176813,0.1920569,0.19891608,0.19891608,0.17490897,0.17833854,0.31552204,0.53844523,0.70649505,0.82996017,0.9259886,0.99801,1.0597426,1.1763484,1.371835,1.6153357,1.821111,1.8965619,2.136633,2.3321195,2.3767042,2.277246,2.0474637,1.9823016,2.0268862,2.1469216,2.3286898,2.095478,2.1023371,2.194936,2.2395205,2.1194851,2.2292318,2.3389788,2.486451,2.668219,2.8568463,2.8465576,2.901431,3.0454736,3.316411,3.765687,4.4996185,5.3432975,6.4064693,8.124693,11.269625,13.786942,15.7966795,17.243965,18.37573,19.737276,20.556948,20.872469,20.491785,19.661825,19.071936,19.44576,20.580954,21.760733,22.573545,22.909645,22.875349,22.724447,22.60098,22.679861,23.170294,23.725885,23.869928,24.065414,24.507832,25.114868,25.574434,24.710178,23.03654,20.875898,18.37916,15.913286,13.872682,12.260776,10.984968,9.873782,8.669997,7.7028537,7.06838,6.783724,6.776865,6.478491,6.23499,6.0703697,6.0223556,6.142391,5.830299,5.5902276,5.4153185,5.2918534,5.192395,5.1100855,4.822,4.355576,3.82399,3.4124396,3.1140654,2.8465576,2.5927682,2.527606,3.0214665,3.683377,4.2766957,4.547633,4.5613513,4.6882463,4.8768735,5.020916,5.0312047,5.127233,5.830299,6.5470824,7.1095347,7.4181976,7.7131424,8.570539,10.155008,11.47197,11.670886,10.494537,8.275595,5.8405876,4.523626,3.9097297,3.7622573,4.033195,4.6608095,5.4496145,6.2418494,6.989499,7.7268605,7.5245147,7.023795,6.660259,6.715132,7.298162,8.052671,6.358455,4.1600895,2.5619018,1.8416885,2.417859,2.877424,3.3266997,3.8548563,4.547633,5.096367,5.9228973,7.034084,8.56368,10.748327,12.6929035,14.527733,16.033321,17.79613,21.19828,21.980227,22.388348,22.796469,23.911083,26.77479,29.192648,30.465025,31.226395,31.370436,30.074053,28.976585,26.791937,24.61415,23.537258,24.665592,25.420103,23.465237,19.661825,15.4914465,13.039291,11.478829,10.63858,10.113853,9.654288,9.167287,8.107545,7.1884155,6.910619,7.39762,8.3922,9.860064,9.06097,7.7440085,7.0203657,7.3564653,8.89635,9.815479,10.398509,10.611144,10.103564,8.388771,8.255017,8.484799,8.4093485,7.9086285,8.543102,8.40249,8.097256,8.134981,8.923786,9.369633,10.028113,11.201033,12.9707,15.199932,15.275383,14.726648,13.594885,11.849225,9.362774,8.899779,8.501947,8.06296,7.5553813,7.0203657,6.385892,5.6176643,4.554492,3.2889743,2.170929,1.3066728,0.67219913,0.33952916,0.216064,0.06859175,0.06859175,0.0548734,0.061732575,0.07888051,0.06516216,0.058302987,0.034295876,0.01371835,0.0034295875,0.006859175,0.024007112,0.034295876,0.030866288,0.020577524,0.034295876,0.048014224,0.048014224,0.044584636,0.037725464,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.010288762,0.0,0.0,0.010288762,0.024007112,0.037725464,0.041155048,0.017147938,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.01371835,0.0548734,0.09602845,0.08916927,0.07545093,0.0548734,0.06516216,0.10288762,0.13032432,0.16804978,0.14747226,0.116605975,0.09259886,0.06516216,0.030866288,0.024007112,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0034295875,0.006859175,0.024007112,0.048014224,0.07888051,0.07888051,0.058302987,0.041155048,0.034295876,0.0548734,0.034295876,0.024007112,0.0274367,0.030866288,0.041155048,0.05144381,0.037725464,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.01371835,0.01371835,0.010288762,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.020577524,0.041155048,0.037725464,0.017147938,0.006859175,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0034295875,0.010288762,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.034295876,0.0548734,0.08916927,0.11317638,0.12346515,0.12346515,0.12346515,0.14404267,0.16119061,0.17147937,0.16804978,0.15090185,0.14404267,0.12346515,0.09602845,0.072021335,0.041155048,0.024007112,0.01371835,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.041155048,0.0274367,0.010288762,0.0,0.0034295875,0.0034295875,0.006859175,0.017147938,0.024007112,0.0274367,0.024007112,0.044584636,0.034295876,0.020577524,0.01371835,0.024007112,0.061732575,0.09602845,0.16119061,0.24007112,0.31209245,0.33609957,0.28808534,0.22978236,0.16119061,0.09602845,0.044584636,0.044584636,0.037725464,0.024007112,0.017147938,0.030866288,0.030866288,0.020577524,0.0274367,0.048014224,0.061732575,0.12346515,0.12003556,0.08916927,0.048014224,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.0274367,0.058302987,0.106317215,0.20577525,0.22978236,0.19891608,0.16462019,0.21263443,0.2503599,0.2503599,0.18862732,0.10288762,0.09259886,0.09259886,0.09945804,0.106317215,0.12003556,0.16804978,0.18176813,0.14747226,0.12689474,0.14747226,0.18176813,0.17147937,0.10288762,0.048014224,0.0274367,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.017147938,0.058302987,0.106317215,0.17833854,0.17147937,0.17833854,0.20920484,0.19891608,0.09945804,0.10288762,0.12346515,0.106317215,0.044584636,0.034295876,0.01371835,0.006859175,0.024007112,0.061732575,0.061732575,0.041155048,0.041155048,0.072021335,0.12346515,0.08573969,0.048014224,0.024007112,0.0274367,0.07545093,0.08916927,0.09259886,0.06859175,0.0274367,0.01371835,0.0274367,0.041155048,0.034295876,0.01371835,0.01371835,0.01371835,0.024007112,0.061732575,0.12346515,0.18176813,0.20920484,0.15776102,0.13375391,0.17147937,0.24350071,0.30523327,0.274367,0.26750782,0.30866286,0.31895164,0.28465575,0.274367,0.25721905,0.23664154,0.26064864,0.31895164,0.4081209,0.42183927,0.34638834,0.274367,0.42183927,0.64133286,0.83681935,0.939707,0.91569984,1.0117283,1.3203912,1.7319417,2.1434922,2.4727325,2.4590142,2.4007113,2.2669573,2.0063086,1.5570327,1.5913286,1.7593783,1.9651536,2.0646117,1.845118,1.8691251,1.7490896,1.4061309,1.0563129,1.1900668,1.1763484,1.1832076,1.2586586,1.5090185,2.1057668,2.2155135,1.9857311,1.6873571,1.4541451,1.2826657,1.1214751,0.864256,0.7476501,0.7956643,0.8093826,0.7956643,0.8025235,0.75450927,0.66876954,0.65505123,0.8162418,1.2586586,1.5330256,1.5090185,1.371835,1.2758065,1.2312219,1.1900668,1.0940384,0.8848336,0.31209245,0.10288762,0.10288762,0.20920484,0.36696586,0.36696586,0.48357183,0.5693115,0.50757897,0.21263443,0.116605975,0.0548734,0.024007112,0.017147938,0.030866288,0.017147938,0.006859175,0.006859175,0.017147938,0.030866288,0.006859175,0.010288762,0.020577524,0.0274367,0.01371835,0.0274367,0.030866288,0.037725464,0.041155048,0.030866288,0.041155048,0.06516216,0.07545093,0.07888051,0.09259886,0.12689474,0.17490897,0.18519773,0.16804978,0.16804978,0.15433143,0.13375391,0.17147937,0.2777966,0.4115505,0.5590228,0.59674823,0.65505123,0.7888051,0.9602845,1.1694894,1.3581166,1.4850113,1.529596,1.4815818,1.4678634,1.5844694,1.6256244,1.4953002,1.1900668,1.1180456,1.1249046,1.255229,1.5364552,1.9994495,2.2909644,2.6579304,3.0317552,3.2649672,3.1449318,2.959734,3.0797696,3.4707425,3.9200184,4.029765,3.7348208,3.3609958,3.0557625,3.0351849,3.5702004,4.15666,4.7979927,5.5422134,6.728851,8.988949,10.830637,12.253916,13.536582,14.781522,15.916716,17.03819,18.060207,18.499195,18.327715,17.974468,17.744686,18.087645,18.962189,20.11453,21.102251,21.61669,22.175713,22.923363,23.78076,24.428951,24.123718,23.965958,24.288338,25.176601,26.459267,27.728214,27.807095,26.77479,24.747904,21.880768,19.377169,17.490896,15.841265,14.119612,12.068718,9.774324,8.467651,7.956643,7.9120584,7.888051,7.5588107,7.0375133,6.4133286,5.970912,6.1801167,6.1321025,6.0086374,5.967482,6.0978065,6.4407654,6.3653145,6.0635104,5.446185,4.6676683,4.1189346,3.8034124,3.7039545,3.6799474,3.7794054,4.2423997,5.0586414,6.23499,7.010077,7.1541195,6.958633,6.5779486,6.385892,6.444195,6.6705475,6.8043017,6.975781,7.1849856,7.0203657,6.677407,6.958633,9.911508,12.089295,12.668896,11.451392,8.851766,6.9689217,6.0806584,5.720552,5.7308407,6.2555676,6.608815,6.625963,6.5470824,6.6396813,7.2021337,8.141841,8.285883,7.846896,7.346176,7.613684,7.431916,6.807731,6.1629686,5.164959,2.7470996,3.1723683,3.5564823,3.799983,4.0229063,4.547633,4.852866,5.0003386,5.223262,5.9160385,7.6616983,9.136421,10.707172,11.859513,12.651748,13.704632,13.7526455,14.064738,15.769243,18.660385,21.208569,22.065966,21.11597,21.568676,24.411804,28.42785,32.553646,32.467903,30.855999,29.192648,27.741934,27.909983,24.85079,20.584383,16.191082,11.794352,9.170717,7.9737906,7.449064,7.3255987,7.8126,7.936065,7.9086285,7.936065,8.1487,8.635701,10.014396,10.97468,11.180455,10.618003,9.568549,9.349055,9.294182,9.544542,10.007536,10.360784,9.297611,7.9429245,7.455923,7.5931067,6.715132,5.871454,5.5593615,5.4736214,5.8234396,7.3255987,8.484799,8.546532,9.211872,10.9541025,13.015285,14.517444,15.230798,15.073037,14.356253,13.7938,12.80608,11.46854,10.539123,10.172156,9.901219,9.208443,8.738589,7.891481,6.5162163,4.928317,3.391862,2.393852,1.6976458,1.0837497,0.34981793,0.33952916,0.28122616,0.31209245,0.39440256,0.31895164,0.28465575,0.17490897,0.06859175,0.017147938,0.030866288,0.12689474,0.17833854,0.15090185,0.09602845,0.16804978,0.24007112,0.23321195,0.22635277,0.19548649,0.0,0.0,0.0,0.01371835,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.07888051,0.048014224,0.0,0.0,0.044584636,0.12003556,0.18862732,0.21263443,0.07888051,0.0274367,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.09945804,0.14061308,0.14061308,0.106317215,0.044584636,0.082310095,0.12689474,0.116605975,0.05144381,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.041155048,0.030866288,0.017147938,0.041155048,0.06859175,0.07888051,0.09259886,0.09259886,0.09945804,0.07545093,0.030866288,0.030866288,0.06859175,0.06859175,0.048014224,0.0274367,0.01371835,0.0274367,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.020577524,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.11317638,0.12003556,0.07888051,0.030866288,0.006859175,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.017147938,0.030866288,0.0548734,0.06859175,0.07545093,0.07545093,0.07545093,0.07545093,0.10288762,0.12346515,0.12346515,0.1371835,0.16119061,0.17833854,0.17147937,0.1371835,0.07545093,0.05144381,0.037725464,0.024007112,0.01371835,0.0,0.0,0.010288762,0.010288762,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.01371835,0.041155048,0.044584636,0.058302987,0.072021335,0.061732575,0.034295876,0.020577524,0.044584636,0.07888051,0.08573969,0.024007112,0.030866288,0.05144381,0.08573969,0.12689474,0.15090185,0.2194936,0.22978236,0.17490897,0.10288762,0.082310095,0.09259886,0.09259886,0.072021335,0.037725464,0.030866288,0.030866288,0.0274367,0.058302987,0.106317215,0.09602845,0.12003556,0.11317638,0.07545093,0.020577524,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.0274367,0.020577524,0.017147938,0.0274367,0.044584636,0.08573969,0.17490897,0.22635277,0.2194936,0.20234565,0.26750782,0.30523327,0.30523327,0.3018037,0.34638834,0.30866286,0.29494452,0.28122616,0.2503599,0.1920569,0.1371835,0.07888051,0.0548734,0.06859175,0.08573969,0.10288762,0.09259886,0.06516216,0.0274367,0.01371835,0.006859175,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.017147938,0.0274367,0.044584636,0.061732575,0.072021335,0.08573969,0.09259886,0.09945804,0.1097468,0.12003556,0.09602845,0.05144381,0.020577524,0.010288762,0.010288762,0.01371835,0.017147938,0.024007112,0.044584636,0.037725464,0.024007112,0.01371835,0.024007112,0.06516216,0.07888051,0.082310095,0.09945804,0.1371835,0.082310095,0.05144381,0.037725464,0.030866288,0.0274367,0.020577524,0.0274367,0.020577524,0.006859175,0.01371835,0.024007112,0.037725464,0.048014224,0.0548734,0.048014224,0.0548734,0.06516216,0.13032432,0.22292319,0.25721905,0.3566771,0.45956472,0.48357183,0.4355576,0.41840968,0.39097297,0.33266997,0.30523327,0.31209245,0.29494452,0.29837412,0.3806842,0.48357183,0.5761707,0.64133286,0.6893471,0.65848076,0.6344737,0.66191036,0.7442205,0.94999576,1.1832076,1.3615463,1.4644338,1.5330256,1.7936742,1.9925903,2.0749004,1.9651536,1.5810398,1.6359133,2.1640697,2.8808534,3.4638834,3.5564823,2.8088322,2.294394,2.095478,2.0886188,1.9582944,1.7319417,1.7662375,2.2052248,2.6785078,2.287535,1.920569,1.5570327,1.2689474,1.1489118,1.3306799,1.786815,2.311542,1.9891608,1.0048691,0.6379033,0.6859175,0.7922347,0.7579388,0.59674823,0.53501564,0.6241849,0.9259886,1.0940384,1.0494537,0.9842916,1.0014396,0.9945804,0.96371406,0.88826317,0.7510797,0.45956472,0.3018037,0.22978236,0.20920484,0.2194936,0.19891608,0.29151493,0.36696586,0.33952916,0.15090185,0.09259886,0.072021335,0.06516216,0.05144381,0.006859175,0.0034295875,0.006859175,0.006859175,0.006859175,0.017147938,0.01371835,0.006859175,0.01371835,0.034295876,0.05144381,0.06516216,0.058302987,0.06516216,0.08573969,0.09259886,0.10288762,0.13375391,0.19891608,0.26407823,0.23664154,0.16804978,0.09945804,0.08573969,0.12003556,0.12003556,0.09602845,0.14061308,0.24007112,0.37382504,0.4972902,0.59674823,0.65505123,0.7990939,1.039165,1.2792361,1.3203912,1.4610043,1.6324836,1.7936742,1.920569,1.8485477,1.7010754,1.5158776,1.3203912,1.1420527,1.155771,1.1934965,1.2723769,1.4404267,1.7662375,1.9720128,2.3149714,2.8294096,3.3747141,3.642222,3.940596,4.3452873,4.7671266,5.137522,5.4324665,5.2472687,4.7945633,4.3521466,4.098357,4.108646,4.3041325,4.7431192,5.147811,5.5079174,6.108095,7.0032177,8.532814,10.038403,11.235329,12.202472,13.042721,14.112752,15.361122,16.561478,17.29198,16.79469,17.147938,18.070496,19.281141,20.505503,21.047379,21.496655,21.77788,21.85676,21.733295,22.559826,23.139427,23.506393,23.588703,23.211449,23.845922,24.521551,25.073713,25.056566,23.749893,21.743584,19.613811,17.326277,14.990726,12.850664,11.30735,10.329918,9.836057,9.599416,9.242738,8.64942,7.997798,7.442205,7.0135064,6.5950966,6.1732574,5.844017,5.7822843,5.9812007,6.2555676,6.4373355,6.5059276,6.3378778,6.012067,5.802862,5.703404,5.6793966,5.813151,6.1286726,6.6225333,7.1952744,7.298162,7.0546613,6.5985265,6.090947,5.8680243,6.1972647,6.5367937,6.5710897,6.2075534,6.094377,5.7994323,5.3844523,5.06893,5.212973,8.292743,9.952662,10.254466,9.56512,8.556821,9.030104,9.1981535,8.453933,7.1198235,6.4133286,6.5642304,7.1952744,7.8846216,8.4264965,8.81404,9.205012,9.352485,8.800322,7.9429245,8.004657,8.14527,8.224151,8.124693,7.6033955,6.310441,5.909179,5.2335505,4.647091,4.3452873,4.3521466,4.431027,4.5030484,4.647091,4.99005,5.7308407,6.7871537,8.800322,10.971251,12.950122,14.850114,14.829536,15.645778,17.490896,20.131678,22.919933,21.928782,19.229696,16.750105,16.287111,19.490345,25.814505,29.720804,31.50762,31.401302,29.545897,29.504742,29.106909,27.982004,25.416672,20.340883,15.536031,11.423956,8.766026,7.507367,6.773435,6.5059276,6.5299344,6.9346256,7.407909,7.233,7.284444,7.500508,9.407358,12.044711,11.97269,9.877212,8.995808,8.611694,8.244728,7.6514096,6.6465406,6.5367937,6.8557453,6.9963584,6.2144127,5.06893,3.8308492,3.2272418,3.5804894,4.8082814,6.0566516,6.48535,7.2707253,8.934075,11.317638,12.4802685,13.128461,13.039291,12.281353,11.231899,11.382801,10.9198065,10.151579,9.637141,10.158438,10.216741,9.9801,9.424506,8.56025,7.431916,6.848886,6.5813785,6.0532217,4.945465,3.2066643,1.9754424,1.3615463,0.90884066,0.47328308,0.22292319,0.1371835,0.09602845,0.12346515,0.25378948,0.53158605,0.64819205,0.4629943,0.4664239,0.6962063,0.7305021,0.2469303,0.12003556,0.12003556,0.09945804,0.01371835,0.0034295875,0.2709374,0.41840968,0.30866286,0.05144381,0.030866288,0.030866288,0.05144381,0.06859175,0.048014224,0.010288762,0.0,0.0,0.09602845,0.47671264,0.33952916,0.2194936,0.12003556,0.05144381,0.061732575,0.45270553,0.5727411,0.3841138,0.06859175,0.041155048,0.10288762,0.1371835,0.116605975,0.06516216,0.061732575,0.020577524,0.020577524,0.020577524,0.037725464,0.1371835,0.28122616,0.32238123,0.2709374,0.16804978,0.058302987,0.0274367,0.024007112,0.024007112,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.048014224,0.048014224,0.041155048,0.0548734,0.08573969,0.09259886,0.1097468,0.12003556,0.12689474,0.12003556,0.041155048,0.024007112,0.020577524,0.024007112,0.024007112,0.006859175,0.01371835,0.020577524,0.037725464,0.0548734,0.05144381,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.058302987,0.11317638,0.16462019,0.21263443,0.09259886,0.024007112,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.020577524,0.041155048,0.058302987,0.06859175,0.08916927,0.08916927,0.09259886,0.10288762,0.11317638,0.12346515,0.15090185,0.17147937,0.18519773,0.17490897,0.12346515,0.082310095,0.0548734,0.030866288,0.01371835,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0034295875,0.0,0.0,0.006859175,0.01371835,0.0034295875,0.017147938,0.0274367,0.041155048,0.05144381,0.048014224,0.020577524,0.017147938,0.024007112,0.037725464,0.041155048,0.006859175,0.01371835,0.030866288,0.048014224,0.06516216,0.08916927,0.1920569,0.20234565,0.16462019,0.12003556,0.09945804,0.11317638,0.106317215,0.07888051,0.05144381,0.030866288,0.024007112,0.0548734,0.1097468,0.14404267,0.08916927,0.116605975,0.11317638,0.06516216,0.0034295875,0.0,0.006859175,0.01371835,0.0274367,0.037725464,0.020577524,0.01371835,0.006859175,0.01371835,0.024007112,0.030866288,0.06859175,0.17490897,0.24007112,0.24007112,0.22635277,0.26407823,0.32238123,0.34638834,0.34295875,0.37382504,0.3841138,0.36353627,0.32581082,0.2777966,0.20920484,0.15776102,0.12003556,0.10288762,0.09945804,0.08916927,0.06859175,0.05144381,0.030866288,0.010288762,0.006859175,0.0,0.006859175,0.017147938,0.0274367,0.024007112,0.030866288,0.034295876,0.041155048,0.06859175,0.14061308,0.21263443,0.26064864,0.26407823,0.2469303,0.28808534,0.23664154,0.12003556,0.037725464,0.017147938,0.006859175,0.017147938,0.034295876,0.030866288,0.017147938,0.024007112,0.048014224,0.034295876,0.01371835,0.0,0.0,0.024007112,0.034295876,0.037725464,0.05144381,0.08916927,0.13375391,0.09259886,0.041155048,0.01371835,0.01371835,0.01371835,0.020577524,0.030866288,0.06859175,0.15090185,0.09259886,0.058302987,0.041155048,0.034295876,0.024007112,0.024007112,0.034295876,0.06859175,0.11317638,0.13032432,0.2469303,0.36010668,0.38754338,0.34638834,0.34981793,0.39097297,0.42526886,0.4389872,0.4355576,0.432128,0.48700142,0.6207553,0.70649505,0.7099246,0.70649505,0.67219913,0.5796003,0.53158605,0.5693115,0.65505123,0.8162418,1.0528834,1.255229,1.3786942,1.4541451,1.5913286,1.7388009,1.9102802,2.0817597,2.1915064,2.3321195,2.7642474,3.391862,4.122364,4.8322887,3.6970954,3.0043187,2.7059445,2.5927682,2.2806756,2.819121,3.1689389,3.2889743,3.2306714,3.1312134,2.6716487,2.07833,1.4507155,1.0288762,1.196926,1.4027013,1.5844694,1.2963841,0.6962063,0.5418748,0.64476246,0.77508676,0.72707254,0.5418748,0.47671264,0.53501564,0.70306545,0.7922347,0.77508676,0.78537554,0.922559,1.1008976,1.3306799,1.529596,1.5330256,0.864256,0.5521636,0.37382504,0.22292319,0.1097468,0.17490897,0.2469303,0.28122616,0.23664154,0.09945804,0.07545093,0.0548734,0.044584636,0.030866288,0.0,0.006859175,0.01371835,0.010288762,0.0034295875,0.01371835,0.01371835,0.017147938,0.024007112,0.034295876,0.05144381,0.058302987,0.048014224,0.058302987,0.09259886,0.12346515,0.1371835,0.12346515,0.13375391,0.15776102,0.12689474,0.09602845,0.082310095,0.08573969,0.10288762,0.12346515,0.15776102,0.2194936,0.31552204,0.432128,0.5555932,0.6927767,0.90541106,1.0734608,1.1283343,1.0563129,0.99801,1.0768905,1.2415106,1.4472859,1.6633499,1.5330256,1.4781522,1.5433143,1.762808,2.1743584,2.2395205,2.3286898,2.486451,2.5996273,2.4315774,2.5653315,2.867135,3.2889743,3.8137012,4.465323,4.887162,5.2575574,5.960623,6.800872,7.010077,6.660259,6.042933,5.48734,5.038064,4.461893,3.974892,3.99204,4.2423997,4.547633,4.8082814,5.15467,6.1629686,7.274155,8.217292,9.043822,9.753747,10.621432,11.876661,13.474849,15.107333,15.700651,16.407146,17.326277,18.550638,20.162544,20.419764,20.543228,20.502073,20.340883,20.169403,21.04395,21.712719,22.076254,21.956219,21.091963,21.602972,22.789608,24.552416,26.003132,25.471546,23.736176,21.44864,18.972477,16.592344,14.510585,12.97413,11.8115,11.091286,10.64201,10.041832,9.263316,8.505377,7.9909387,7.740579,7.531374,7.390761,6.9689217,6.584808,6.3310184,6.0806584,5.73427,5.720552,5.796003,5.895461,6.125243,6.632822,6.526505,6.3173003,6.3618846,6.869464,6.5539417,5.844017,4.9523244,4.108646,3.5221863,3.3987212,3.7485392,4.314421,4.955754,5.645101,5.456474,4.928317,4.413879,4.273266,4.8597255,6.7185616,7.7748747,7.7097125,7.0958166,7.394191,8.1487,7.932636,7.4627824,7.239859,7.5450926,8.299602,8.858624,9.074688,8.995808,8.868914,8.89635,9.328478,9.537683,9.451943,9.530824,9.177576,9.671436,10.415657,10.933525,10.871792,8.724871,7.349606,6.138962,4.955754,4.139512,3.9440255,3.9063,3.9954693,4.170378,4.3795834,4.804852,5.7377,7.2535777,10.463672,17.490896,17.78927,17.61436,18.36544,19.8676,20.361462,19.473198,17.916164,15.553179,13.88297,16.012743,20.745575,24.957108,28.369547,30.334702,29.823692,29.062325,29.624777,29.864847,28.661062,25.44068,21.19485,16.228807,12.281353,9.873782,8.337327,7.421627,7.349606,7.56224,7.658269,7.366754,8.742019,9.0644,9.9698105,11.543991,12.343085,10.477389,9.242738,8.292743,7.4627824,6.773435,6.684266,6.632822,6.1492505,5.504488,5.7136927,4.880303,3.806842,3.1586502,3.0146074,2.8637056,3.3266997,3.9954693,4.787704,5.909179,7.857185,9.414218,11.019264,11.72233,11.279913,10.158438,9.434795,9.078118,8.9100685,8.920357,9.242738,9.078118,9.462232,9.582268,9.095266,8.1487,7.3873315,7.689135,8.028665,7.7577267,6.5950966,3.7005248,2.07833,1.1763484,0.71678376,0.7099246,0.3566771,0.2194936,0.26750782,0.44927597,0.6756287,0.607037,0.4081209,0.34295875,0.5178677,0.88826317,0.59674823,0.36353627,0.18519773,0.07545093,0.041155048,0.030866288,0.17833854,0.31209245,0.31209245,0.13375391,0.06516216,0.058302987,0.08916927,0.13375391,0.16119061,0.12689474,0.106317215,0.061732575,0.048014224,0.23664154,0.16804978,0.15433143,0.13032432,0.09945804,0.13032432,0.39097297,0.48014224,0.36010668,0.13032432,0.0274367,0.072021335,0.08916927,0.07888051,0.0548734,0.041155048,0.034295876,0.037725464,0.041155048,0.072021335,0.19548649,0.24350071,0.22978236,0.16462019,0.07888051,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.006859175,0.0,0.006859175,0.01371835,0.017147938,0.030866288,0.08916927,0.15433143,0.18862732,0.1920569,0.16804978,0.15090185,0.16119061,0.116605975,0.07545093,0.05144381,0.020577524,0.020577524,0.017147938,0.0274367,0.037725464,0.0274367,0.034295876,0.034295876,0.037725464,0.037725464,0.024007112,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.017147938,0.044584636,0.07545093,0.10288762,0.044584636,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0274367,0.044584636,0.0548734,0.048014224,0.05144381,0.061732575,0.072021335,0.07545093,0.09259886,0.106317215,0.12003556,0.13032432,0.12003556,0.09259886,0.061732575,0.034295876,0.017147938,0.024007112,0.030866288,0.01371835,0.0034295875,0.010288762,0.010288762,0.017147938,0.030866288,0.041155048,0.05144381,0.044584636,0.0274367,0.017147938,0.01371835,0.020577524,0.0274367,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.0,0.01371835,0.0274367,0.034295876,0.037725464,0.05144381,0.116605975,0.12003556,0.10288762,0.08916927,0.08916927,0.106317215,0.09602845,0.072021335,0.041155048,0.017147938,0.017147938,0.082310095,0.1371835,0.13375391,0.05144381,0.07545093,0.07545093,0.044584636,0.006859175,0.01371835,0.024007112,0.058302987,0.09259886,0.09259886,0.0274367,0.01371835,0.0034295875,0.010288762,0.024007112,0.030866288,0.06516216,0.12689474,0.16462019,0.16804978,0.17833854,0.19891608,0.2469303,0.2709374,0.2709374,0.28465575,0.31895164,0.31209245,0.28122616,0.2469303,0.2194936,0.20234565,0.19891608,0.17833854,0.13375391,0.09945804,0.061732575,0.030866288,0.01371835,0.010288762,0.006859175,0.006859175,0.01371835,0.030866288,0.048014224,0.048014224,0.037725464,0.07545093,0.116605975,0.14404267,0.16462019,0.22978236,0.274367,0.2709374,0.2469303,0.274367,0.19891608,0.072021335,0.0,0.0034295875,0.01371835,0.048014224,0.06516216,0.048014224,0.010288762,0.017147938,0.037725464,0.024007112,0.006859175,0.006859175,0.030866288,0.034295876,0.017147938,0.0034295875,0.006859175,0.0274367,0.116605975,0.13375391,0.09602845,0.034295876,0.0,0.01371835,0.024007112,0.044584636,0.09259886,0.18862732,0.13375391,0.082310095,0.05144381,0.044584636,0.0548734,0.044584636,0.041155048,0.041155048,0.037725464,0.044584636,0.18176813,0.25721905,0.25378948,0.20577525,0.216064,0.25721905,0.31209245,0.32924038,0.31895164,0.32924038,0.41840968,0.5590228,0.6241849,0.6001778,0.61389613,0.6036074,0.5521636,0.52815646,0.5624523,0.66876954,0.8265306,1.1008976,1.313532,1.4335675,1.5570327,1.7113642,2.1503513,2.5173173,2.6887965,2.7642474,2.6579304,2.819121,3.1895163,3.7862647,4.6676683,4.6745276,4.5442033,4.2938433,3.8617156,3.1106358,3.8891523,4.3109913,4.245829,3.8891523,3.7519686,3.1963756,2.5413244,1.8862731,1.4164196,1.3992717,1.2826657,1.0871792,0.8025235,0.59674823,0.7888051,0.96714365,1.0220171,0.8676856,0.6001778,0.47671264,0.48700142,0.5624523,0.6344737,0.6927767,0.7613684,0.89512235,1.1763484,1.4507155,1.5981878,1.5261664,0.89512235,0.5658819,0.36696586,0.20920484,0.09602845,0.15776102,0.18519773,0.18176813,0.14404267,0.06859175,0.072021335,0.072021335,0.07545093,0.07545093,0.06859175,0.0548734,0.041155048,0.024007112,0.01371835,0.020577524,0.0274367,0.037725464,0.05144381,0.06516216,0.08916927,0.07545093,0.041155048,0.034295876,0.0548734,0.08916927,0.09602845,0.06859175,0.06859175,0.09602845,0.09259886,0.07888051,0.14061308,0.17147937,0.15776102,0.17490897,0.26064864,0.32924038,0.40126175,0.490431,0.59331864,0.7373613,0.96371406,1.097468,1.0666018,0.89169276,0.8711152,0.94999576,1.1008976,1.2929544,1.4987297,1.4610043,1.546744,1.762808,2.1297739,2.6990852,2.877424,3.07634,3.3198407,3.5118976,3.4467354,3.57363,3.6868064,3.7862647,3.9646032,4.417309,4.506478,4.3624353,4.7328305,5.4907694,5.641671,5.504488,5.4633327,5.3913116,5.137522,4.530485,3.724532,3.6456516,3.957744,4.386442,4.722542,4.715683,5.020916,5.4736214,5.9983487,6.6122446,7.377043,8.107545,9.0644,10.374502,12.055,13.402828,14.318527,15.110763,16.204802,18.142517,18.886738,19.349733,19.473198,19.418324,19.53493,20.083664,20.474638,20.467777,20.066517,19.517782,20.073376,21.28402,23.077694,24.734184,24.871368,24.085993,22.724447,20.875898,18.807858,16.945591,15.563468,14.356253,13.365103,12.504276,11.5645685,10.837497,9.914937,9.177576,8.786603,8.673427,8.844906,8.611694,8.186425,7.658269,6.9860697,5.9640527,5.453044,5.2644167,5.267846,5.40503,5.809721,5.5833683,5.1992545,5.0414934,5.3878818,4.8288593,4.098357,3.3026927,2.5790498,2.0989075,2.0131679,2.2498093,2.784825,3.6559403,4.9694724,5.284994,5.0483527,4.7534084,4.7945633,5.4976287,6.3001523,6.7802944,6.2830043,5.23698,5.15467,5.5662203,5.641671,5.8680243,6.341307,6.7494283,7.5416627,8.080108,8.30646,8.279024,8.165848,8.591117,9.146709,9.551401,9.856634,10.4533825,10.14472,10.899229,12.346515,13.852104,14.555169,12.764925,11.495977,9.400499,6.543653,4.413879,3.525616,3.1792276,3.350707,3.724532,3.724532,3.5839188,3.5599117,4.4275975,7.922347,16.715809,20.063087,18.79757,17.61436,17.754974,17.024471,16.520323,15.844694,14.507155,13.334236,14.445422,16.767254,19.723558,23.046827,26.00999,27.43327,27.282368,28.239223,28.911423,28.52731,26.908543,24.730755,20.762722,16.173935,12.188754,10.106995,8.841476,8.573969,8.707723,8.790032,8.519095,10.079557,10.6488695,10.467101,10.120712,10.532263,9.582268,8.659708,7.81603,7.1232533,6.667118,6.8728933,6.711703,5.9434752,5.0757895,5.360445,4.5990767,4.1429415,3.806842,3.340418,2.4247184,2.2635276,2.7985435,3.4055803,4.0057583,5.079219,6.6053853,8.940934,10.88894,11.921246,12.1921835,12.277924,12.212761,11.657167,10.940384,11.074138,11.934964,13.4645605,14.150477,13.38225,11.461681,9.472521,8.748878,9.088407,9.788043,9.650859,6.9654922,4.5647807,2.719663,1.5776103,1.1763484,0.7579388,1.3512574,1.5741806,1.0666018,0.48014224,0.3566771,0.25378948,0.28122616,0.5453044,1.155771,1.0631721,0.7442205,0.42526886,0.23321195,0.19548649,0.12003556,0.2194936,0.40126175,0.48014224,0.19548649,0.116605975,0.116605975,0.16804978,0.22978236,0.25378948,0.24350071,0.274367,0.31895164,0.28465575,0.0,0.0,0.048014224,0.16804978,0.29837412,0.32581082,0.36353627,0.37039545,0.34981793,0.29494452,0.18519773,0.07545093,0.041155048,0.041155048,0.044584636,0.01371835,0.024007112,0.0274367,0.030866288,0.0548734,0.12689474,0.12003556,0.08573969,0.041155048,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.037725464,0.082310095,0.12346515,0.14061308,0.14061308,0.15090185,0.24350071,0.30523327,0.26407823,0.15776102,0.116605975,0.12003556,0.07545093,0.030866288,0.01371835,0.01371835,0.024007112,0.034295876,0.041155048,0.037725464,0.0274367,0.034295876,0.030866288,0.024007112,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.010288762,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.020577524,0.041155048,0.030866288,0.024007112,0.0274367,0.034295876,0.041155048,0.041155048,0.048014224,0.05144381,0.06859175,0.09259886,0.09945804,0.08916927,0.06516216,0.041155048,0.024007112,0.030866288,0.037725464,0.020577524,0.006859175,0.010288762,0.010288762,0.017147938,0.030866288,0.041155048,0.048014224,0.05144381,0.034295876,0.017147938,0.0034295875,0.0034295875,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.01371835,0.017147938,0.017147938,0.01371835,0.01371835,0.020577524,0.0274367,0.024007112,0.020577524,0.05144381,0.072021335,0.072021335,0.0548734,0.0274367,0.010288762,0.030866288,0.106317215,0.13032432,0.07888051,0.01371835,0.01371835,0.01371835,0.01371835,0.017147938,0.0274367,0.041155048,0.09602845,0.14061308,0.13032432,0.041155048,0.030866288,0.01371835,0.010288762,0.017147938,0.0274367,0.041155048,0.041155048,0.041155048,0.048014224,0.06859175,0.10288762,0.12003556,0.13375391,0.15433143,0.16804978,0.18176813,0.20577525,0.20920484,0.20234565,0.2194936,0.22978236,0.24350071,0.20920484,0.13375391,0.09259886,0.06859175,0.034295876,0.020577524,0.020577524,0.01371835,0.01371835,0.020577524,0.030866288,0.041155048,0.061732575,0.020577524,0.09602845,0.16804978,0.16462019,0.072021335,0.0548734,0.06516216,0.072021335,0.058302987,0.041155048,0.017147938,0.006859175,0.010288762,0.024007112,0.048014224,0.09259886,0.09602845,0.05144381,0.0,0.0,0.010288762,0.006859175,0.0034295875,0.017147938,0.06516216,0.072021335,0.037725464,0.006859175,0.0034295875,0.01371835,0.041155048,0.12346515,0.1371835,0.06859175,0.0034295875,0.01371835,0.030866288,0.044584636,0.061732575,0.09602845,0.11317638,0.09602845,0.08916927,0.10288762,0.12689474,0.09259886,0.07545093,0.06859175,0.061732575,0.058302987,0.18176813,0.216064,0.17490897,0.106317215,0.09602845,0.07545093,0.061732575,0.0548734,0.061732575,0.09602845,0.16462019,0.25378948,0.31552204,0.36696586,0.48357183,0.5521636,0.5555932,0.5418748,0.6001778,0.8676856,1.08032,1.2312219,1.3649758,1.5398848,1.8348293,2.301253,3.2203827,3.7965534,3.7485392,3.309552,2.6407824,2.527606,2.74367,3.175798,3.8137012,5.3981705,6.125243,6.200694,5.7582774,4.852866,4.945465,4.9248877,4.7945633,4.513337,3.981751,3.3952916,2.9494452,2.651071,2.3801336,1.8965619,1.5501735,1.2689474,0.96714365,0.7888051,1.1214751,1.3066728,1.2517995,1.0151579,0.71678376,0.52472687,0.4629943,0.4629943,0.5658819,0.7373613,0.8848336,0.9774324,1.1797781,1.2209331,1.039165,0.7922347,0.7305021,0.490431,0.2709374,0.16462019,0.1371835,0.1097468,0.10288762,0.10288762,0.106317215,0.106317215,0.13032432,0.16462019,0.19891608,0.2194936,0.21263443,0.15776102,0.11317638,0.07545093,0.05144381,0.05144381,0.07545093,0.09602845,0.13032432,0.16804978,0.18176813,0.14404267,0.08573969,0.044584636,0.034295876,0.058302987,0.06859175,0.07545093,0.13375391,0.22635277,0.2709374,0.25378948,0.34295875,0.38754338,0.36353627,0.3566771,0.45270553,0.52815646,0.59674823,0.66876954,0.7476501,0.84367853,0.939707,1.0254467,1.0837497,1.097468,1.2860953,1.4369972,1.546744,1.6221949,1.6942163,1.7662375,1.8382589,1.9308578,2.0817597,2.3732746,2.6887965,2.9871707,3.2649672,3.5770597,4.057202,4.2115335,4.0880685,3.8514268,3.625074,3.4947495,3.1346428,2.4144297,2.0234566,2.1091962,2.2635276,2.620205,3.549623,4.2869844,4.523626,4.4104495,3.8685746,4.0194764,4.4241676,4.8082814,5.0826488,4.938606,4.8151407,4.8151407,4.996909,5.3878818,6.193835,6.866034,7.514226,8.258447,9.242738,10.436234,11.303921,11.96926,12.871242,14.778092,16.499744,17.864721,18.663815,19.058218,19.576086,19.881319,19.901896,19.384027,18.653526,18.62266,19.082224,19.819586,20.670124,21.503513,22.216867,22.8582,23.18744,22.597551,21.184563,19.733847,18.893597,17.899017,16.722668,15.433144,14.205351,13.577737,12.476839,11.369082,10.55284,10.1652975,10.388221,10.439664,10.247607,9.764035,8.961512,7.596536,6.5196457,5.7102633,5.1100855,4.647091,4.266407,3.923448,3.673088,3.5530527,3.6079261,3.4776018,3.2478194,2.9906003,2.7368107,2.4795918,2.4007113,2.5173173,2.7813954,3.2718265,4.197815,5.206114,5.456474,5.4839106,5.6176643,5.977771,6.3721733,6.5470824,5.9880595,4.715683,3.309552,3.4947495,4.431027,5.15467,5.1752477,4.4756117,4.537344,5.103226,5.994919,6.9552035,7.623973,8.762596,9.088407,8.937505,8.934075,9.962952,10.189304,10.882081,12.439114,14.4145565,15.529172,16.232237,16.12592,14.05102,10.439664,7.3118806,4.633373,3.1620796,3.1106358,3.858286,3.940596,3.4227283,3.0111778,3.5633414,6.108095,11.845795,19.517782,18.495766,15.693792,14.363112,14.088745,14.092175,13.481709,12.782072,12.38767,12.566009,13.13532,14.603184,16.760393,19.456049,22.60098,24.295198,25.492125,26.19176,26.222626,25.241764,24.881657,22.576975,18.269413,13.454271,11.173596,9.884071,9.441654,9.678296,10.065839,9.716022,9.695444,10.199594,9.908078,8.827758,8.268735,7.953213,7.623973,7.31531,7.0135064,6.6533995,6.392751,6.2555676,5.9880595,5.56965,5.1752477,4.3487167,4.3109913,4.2526884,3.8445675,3.2375305,3.1072063,3.40901,3.7691166,4.012617,4.1772375,5.0826488,7.281014,9.983529,12.699762,15.258235,17.854433,18.30028,16.914726,15.134769,15.498305,17.864721,19.997925,20.60839,19.233126,16.252815,13.2690735,10.796341,10.113853,10.964391,11.55428,11.005547,8.899779,6.3824625,4.098357,2.1983654,1.5776103,3.0214665,3.782835,3.1243541,2.318401,2.0337453,1.5536032,1.1592005,1.1351935,1.7593783,1.8588364,1.7730967,1.5981878,1.3855534,1.1523414,0.77165717,0.70649505,0.7888051,0.7613684,0.2709374,0.22978236,0.25378948,0.31552204,0.36696586,0.34638834,0.39783216,0.5212973,0.70649505,0.70649505,0.044584636,0.09259886,0.08573969,0.23321195,0.47328308,0.47671264,0.39783216,0.34295875,0.33609957,0.36010668,0.33609957,0.10288762,0.041155048,0.044584636,0.041155048,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.01371835,0.017147938,0.034295876,0.0548734,0.05144381,0.041155048,0.0274367,0.01371835,0.0,0.0,0.0034295875,0.0034295875,0.017147938,0.07545093,0.16119061,0.22978236,0.26750782,0.25378948,0.17490897,0.22978236,0.29494452,0.24350071,0.106317215,0.037725464,0.05144381,0.07545093,0.06859175,0.037725464,0.024007112,0.020577524,0.041155048,0.041155048,0.020577524,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.017147938,0.034295876,0.0548734,0.041155048,0.041155048,0.041155048,0.037725464,0.037725464,0.037725464,0.044584636,0.05144381,0.06859175,0.08573969,0.08573969,0.07888051,0.06859175,0.05144381,0.037725464,0.037725464,0.034295876,0.024007112,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.017147938,0.006859175,0.0034295875,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.030866288,0.024007112,0.01371835,0.01371835,0.041155048,0.037725464,0.017147938,0.0034295875,0.01371835,0.01371835,0.024007112,0.037725464,0.044584636,0.044584636,0.106317215,0.15090185,0.12003556,0.041155048,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0274367,0.041155048,0.041155048,0.0274367,0.01371835,0.01371835,0.024007112,0.024007112,0.01371835,0.01371835,0.0274367,0.020577524,0.020577524,0.034295876,0.044584636,0.058302987,0.06859175,0.07545093,0.082310095,0.106317215,0.13032432,0.15433143,0.18176813,0.19548649,0.18176813,0.18176813,0.16462019,0.13375391,0.10288762,0.09259886,0.06859175,0.034295876,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.030866288,0.024007112,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.0034295875,0.017147938,0.0548734,0.09602845,0.12346515,0.14747226,0.106317215,0.044584636,0.0,0.0,0.0,0.010288762,0.020577524,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.01371835,0.061732575,0.061732575,0.034295876,0.010288762,0.0034295875,0.01371835,0.01371835,0.01371835,0.020577524,0.034295876,0.044584636,0.034295876,0.08573969,0.17147937,0.2503599,0.274367,0.18862732,0.14061308,0.12346515,0.12003556,0.106317215,0.082310095,0.06859175,0.061732575,0.058302987,0.044584636,0.044584636,0.072021335,0.116605975,0.17833854,0.29151493,0.34981793,0.3841138,0.40126175,0.4115505,0.4115505,0.40126175,0.37725464,0.432128,0.70649505,1.4027013,1.5501735,1.1111864,1.1660597,1.9685832,2.9460156,3.82399,4.417309,4.7774153,4.846007,4.4550343,3.3678548,3.0317552,3.309552,3.9851806,4.791134,5.0346346,5.470192,6.0532217,6.708273,7.3530354,6.550512,5.5422134,4.633373,4.1292233,4.3487167,4.3487167,4.3487167,4.262977,3.724532,2.0920484,1.1489118,0.6310441,0.5590228,0.7305021,0.71678376,0.6790583,0.6344737,0.65162164,0.6962063,0.61046654,0.48700142,0.3566771,0.45613512,0.7888051,1.1283343,1.3992717,1.371835,1.2517995,1.1592005,1.1592005,1.3786942,0.89512235,0.37039545,0.11317638,0.07545093,0.08916927,0.15433143,0.23664154,0.29151493,0.29151493,0.3018037,0.34295875,0.39783216,0.432128,0.39783216,0.31209245,0.24350071,0.18176813,0.1371835,0.1371835,0.19891608,0.26750782,0.34295875,0.37725464,0.30523327,0.25721905,0.216064,0.17833854,0.16804978,0.22978236,0.29151493,0.31552204,0.3806842,0.5041494,0.6241849,0.7339317,0.78194594,0.8128122,0.84367853,0.8711152,0.90541106,0.9877212,1.0940384,1.2003556,1.2963841,1.3341095,1.4164196,1.5261664,1.6359133,1.7079345,2.2566686,2.5138876,2.4727325,2.2292318,1.9994495,1.7662375,1.5913286,1.5055889,1.6187652,2.1057668,2.411,2.633923,2.867135,3.117495,3.3266997,3.4124396,3.3129816,3.1552205,3.0043187,2.884283,2.7368107,2.369845,2.037175,1.862266,1.862266,2.177788,2.9460156,3.6765177,4.15323,4.4104495,4.496189,4.664239,4.791134,4.8151407,4.729401,4.8768735,5.1066556,5.4153185,5.778855,6.135532,6.5367937,6.958633,7.390761,7.8263187,8.255017,8.951223,9.729739,10.583707,11.540562,12.665466,14.201921,15.9613,17.63151,19.017063,20.004784,20.347742,20.155685,19.764713,19.414894,19.257133,19.219408,19.349733,19.500635,19.713268,20.2037,21.45893,22.607841,23.156574,22.94394,22.12427,21.795029,20.86218,19.658396,18.45461,17.439453,16.45173,15.333686,14.188204,13.193623,12.617453,12.655178,12.572867,12.274493,11.718901,10.926665,9.863494,8.783174,7.610255,6.4407654,5.5387836,4.856296,4.3624353,4.149801,4.1189346,3.998899,3.74168,3.4227283,3.2066643,3.1380725,3.1140654,3.07634,2.976882,2.9700227,3.1449318,3.525616,4.232111,4.245829,4.1360826,4.184097,4.3795834,4.48933,5.020916,5.6073756,5.7891436,5.020916,5.1066556,5.144381,5.127233,4.9660425,4.5030484,4.07435,3.9680326,4.773986,6.4407654,8.268735,8.988949,8.776315,8.423067,8.268735,8.193284,7.997798,7.8023114,8.433355,10.021255,12.024134,14.366542,16.554619,18.221397,18.6158,16.599203,10.045261,5.56965,4.0263357,4.6848164,5.2335505,4.4996185,3.532475,3.0900583,3.865145,6.4407654,14.459141,16.46545,14.30481,10.940384,10.4533825,12.418536,13.111313,12.195613,10.39508,9.489669,8.964942,9.201583,10.336777,12.7272,16.938732,19.634388,20.62897,21.129688,21.578964,21.650986,20.543228,18.413456,16.04018,13.88297,12.099585,10.6488695,10.220171,10.203023,10.096705,9.5205345,8.680285,8.632272,8.700864,8.742019,9.170717,8.669997,8.279024,7.840037,7.239859,6.4098988,6.138962,5.73427,5.164959,4.7362604,5.0655007,5.079219,4.5784993,4.0949273,3.8720043,3.8617156,4.372724,5.1238036,5.5079174,5.3878818,5.0826488,5.593657,6.773435,8.1487,10.045261,13.612033,16.722668,16.997036,16.894148,17.449741,18.279701,18.890167,18.804428,18.108221,17.024471,15.899568,14.640909,12.843805,11.38623,10.844356,11.506266,12.871242,13.104454,12.229909,9.935514,5.552502,3.4776018,3.4913201,5.3227196,8.213862,10.923236,9.544542,7.157549,4.2423997,2.0508933,2.6236343,3.625074,4.671098,5.2266912,5.0483527,4.180667,2.9494452,1.7799559,0.97400284,0.6001778,0.5041494,0.490431,0.5144381,0.52815646,0.53158605,0.5796003,0.77508676,0.9431366,0.9431366,0.70649505,0.22978236,0.45956472,0.42869842,0.28808534,0.15776102,0.12346515,0.024007112,0.0,0.0,0.017147938,0.09259886,0.041155048,0.020577524,0.010288762,0.0,0.0,0.0,0.0,0.0,0.010288762,0.044584636,0.06859175,0.048014224,0.07888051,0.17833854,0.274367,0.2503599,0.19891608,0.1371835,0.072021335,0.0,0.0,0.017147938,0.024007112,0.01371835,0.01371835,0.05144381,0.07888051,0.1097468,0.11317638,0.01371835,0.0034295875,0.09945804,0.22292319,0.26750782,0.12346515,0.14747226,0.216064,0.18519773,0.072021335,0.061732575,0.048014224,0.037725464,0.017147938,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.037725464,0.0548734,0.09259886,0.07888051,0.07545093,0.06859175,0.061732575,0.061732575,0.09602845,0.09602845,0.07888051,0.061732575,0.061732575,0.072021335,0.06859175,0.06859175,0.072021335,0.061732575,0.048014224,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.0034295875,0.0,0.0034295875,0.01371835,0.0274367,0.058302987,0.072021335,0.06516216,0.06516216,0.08916927,0.06516216,0.024007112,0.0034295875,0.01371835,0.024007112,0.044584636,0.06516216,0.08573969,0.09602845,0.106317215,0.09945804,0.06516216,0.024007112,0.041155048,0.030866288,0.0274367,0.024007112,0.017147938,0.0274367,0.030866288,0.041155048,0.048014224,0.048014224,0.0274367,0.0274367,0.037725464,0.037725464,0.0274367,0.0274367,0.041155048,0.034295876,0.034295876,0.044584636,0.058302987,0.061732575,0.0548734,0.058302987,0.06859175,0.09602845,0.09945804,0.10288762,0.1097468,0.1097468,0.09602845,0.08916927,0.082310095,0.07888051,0.07545093,0.0548734,0.041155048,0.024007112,0.01371835,0.010288762,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.010288762,0.01371835,0.006859175,0.01371835,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0,0.034295876,0.08916927,0.14747226,0.17147937,0.1371835,0.082310095,0.037725464,0.01371835,0.01371835,0.020577524,0.034295876,0.034295876,0.0274367,0.01371835,0.0034295875,0.006859175,0.01371835,0.024007112,0.072021335,0.082310095,0.06516216,0.030866288,0.0034295875,0.01371835,0.01371835,0.024007112,0.034295876,0.044584636,0.044584636,0.034295876,0.048014224,0.09945804,0.17833854,0.2503599,0.26407823,0.22292319,0.24350071,0.33266997,0.40126175,0.36696586,0.33952916,0.30866286,0.2709374,0.22978236,0.17147937,0.16119061,0.18519773,0.22978236,0.3018037,0.36353627,0.42526886,0.48357183,0.5178677,0.51100856,0.4972902,0.5624523,0.77508676,1.0666018,1.2449403,1.5570327,1.8862731,2.1194851,2.452155,3.3609958,4.3281393,4.98662,5.192395,5.003768,4.698535,4.3933015,4.7088237,5.144381,5.5113473,5.926327,6.444195,6.9860697,7.205563,6.989499,6.464772,5.5422134,4.9523244,4.5853586,4.3692946,4.2869844,3.758828,3.5702004,3.590778,3.5187566,2.860276,2.4658735,2.054323,1.5810398,1.138623,0.94999576,0.84367853,0.8265306,0.97400284,1.1729189,1.0871792,0.9945804,0.980862,1.2037852,1.6427724,2.0920484,2.4007113,2.2463799,1.9925903,1.7902447,1.5741806,1.3169615,0.97400284,0.6790583,0.48700142,0.3806842,0.23664154,0.17833854,0.17490897,0.20234565,0.24007112,0.36010668,0.4355576,0.490431,0.52815646,0.53158605,0.53501564,0.52472687,0.50757897,0.490431,0.490431,0.52472687,0.548734,0.5144381,0.4355576,0.39097297,0.37039545,0.36696586,0.40126175,0.47671264,0.59674823,0.7442205,0.8848336,1.0323058,1.1626302,1.2346514,1.2277923,1.1934965,1.155771,1.1283343,1.1146159,1.1592005,1.2895249,1.4953002,1.7765263,2.1263442,2.3492675,2.486451,2.5550427,2.5961976,2.6476414,2.7573884,2.7368107,2.5721905,2.3629858,2.3149714,2.2292318,2.1126258,1.9445761,1.8108221,1.8965619,1.9994495,2.061182,2.1812177,2.3732746,2.568761,2.8225505,3.1620796,3.210094,2.9391565,2.651071,2.5447538,2.5173173,2.585909,2.7162333,2.8122618,2.4384367,2.633923,3.0454736,3.4604537,3.82399,3.8788633,4.149801,4.557922,5.0620713,5.669108,5.7582774,5.9640527,6.3447366,6.7700057,6.9380555,7.2364297,7.5553813,7.822889,7.98408,8.011517,8.285883,8.755736,9.438225,10.268185,11.077567,12.079007,13.440554,14.959861,16.414005,17.549198,17.981327,17.902447,17.974468,18.4649,19.233126,19.555508,19.44576,19.181683,18.962189,18.883308,20.052797,21.383478,22.686722,23.760181,24.394655,23.44123,22.343761,21.308027,20.172834,18.416885,17.4566,16.588915,15.604623,14.63062,14.143619,13.996146,13.941273,13.718349,13.245067,12.596875,11.8869505,10.9369545,9.551401,7.966932,6.869464,6.324159,5.967482,5.535354,4.938606,4.290414,3.7519686,3.4913201,3.3609958,3.275256,3.223812,3.4021509,3.3747141,3.3026927,3.3232703,3.5873485,3.5702004,3.724532,4.190956,4.856296,5.3570156,5.446185,5.56965,6.012067,6.475061,6.0566516,5.4599032,4.911169,5.003768,5.5490727,5.562791,5.144381,4.8288593,5.3673043,6.708273,8.001227,8.927217,9.702303,10.446524,11.146159,11.646879,11.667457,10.984968,10.319629,9.997248,9.949233,11.149589,12.775213,14.30481,15.440002,16.101913,13.814379,11.80121,8.320179,4.5682106,4.695105,4.5613513,4.331569,4.07435,4.15323,5.254128,9.6817255,13.87954,14.081886,11.197603,10.80663,12.010415,13.214201,14.071597,14.284232,13.615462,11.372512,9.990388,9.949233,11.327928,13.810948,17.065628,18.084215,18.1288,17.984756,17.940172,17.768692,17.346853,16.585485,15.477728,14.126471,13.05301,12.274493,11.447963,10.645439,10.364213,10.000677,9.626852,9.14328,9.074688,10.587136,10.8958,10.131001,9.119273,8.364764,8.032094,7.0032177,6.375603,6.3001523,6.451054,6.018926,5.2575574,4.8425775,4.5819287,4.3452873,4.081209,3.7039545,4.262977,5.1169443,5.8371577,6.217842,6.7974424,7.8126,9.122703,10.666017,12.46312,13.732068,14.335675,14.781522,14.96329,14.143619,13.502286,12.788932,11.873232,10.847785,10.017825,8.954653,7.6171136,6.142391,5.0586414,5.267846,6.6053853,8.412778,9.9801,10.72775,10.192734,8.625413,7.1026754,6.8728933,8.169277,10.206452,12.339656,10.487679,7.0306544,3.8960114,2.5756202,4.5030484,6.9826403,9.067829,10.076128,9.599416,6.7940125,4.149801,2.1880767,1.1008976,0.7476501,0.6379033,0.44584638,0.274367,0.16804978,0.12689474,0.216064,0.29837412,0.33609957,0.28808534,0.09602845,0.10288762,0.09259886,0.07545093,0.0548734,0.048014224,0.010288762,0.0,0.0034295875,0.017147938,0.030866288,0.041155048,0.0548734,0.072021335,0.072021335,0.01371835,0.061732575,0.07888051,0.05144381,0.0034295875,0.010288762,0.034295876,0.048014224,0.05144381,0.044584636,0.0548734,0.07888051,0.11317638,0.15433143,0.16462019,0.072021335,0.06516216,0.0274367,0.010288762,0.01371835,0.01371835,0.024007112,0.0274367,0.030866288,0.024007112,0.01371835,0.041155048,0.06859175,0.17147937,0.30523327,0.30523327,0.1920569,0.11317638,0.061732575,0.037725464,0.037725464,0.01371835,0.01371835,0.024007112,0.048014224,0.08916927,0.07888051,0.058302987,0.037725464,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.006859175,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0034295875,0.0274367,0.058302987,0.06859175,0.0548734,0.05144381,0.0548734,0.06516216,0.08573969,0.12346515,0.12346515,0.09945804,0.072021335,0.072021335,0.06516216,0.06859175,0.07545093,0.07888051,0.09602845,0.07545093,0.082310095,0.09602845,0.09259886,0.024007112,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.006859175,0.0274367,0.0548734,0.072021335,0.01371835,0.006859175,0.0034295875,0.0,0.0034295875,0.01371835,0.020577524,0.048014224,0.09259886,0.12003556,0.07545093,0.07888051,0.06516216,0.0548734,0.0548734,0.05144381,0.041155048,0.037725464,0.058302987,0.09602845,0.106317215,0.09259886,0.06516216,0.037725464,0.030866288,0.0548734,0.06516216,0.044584636,0.024007112,0.017147938,0.030866288,0.037725464,0.044584636,0.044584636,0.041155048,0.041155048,0.030866288,0.034295876,0.030866288,0.0274367,0.048014224,0.037725464,0.020577524,0.017147938,0.030866288,0.05144381,0.06516216,0.072021335,0.082310095,0.10288762,0.12003556,0.10288762,0.09602845,0.09602845,0.09945804,0.09602845,0.082310095,0.061732575,0.048014224,0.037725464,0.0274367,0.024007112,0.017147938,0.01371835,0.01371835,0.0,0.006859175,0.006859175,0.006859175,0.006859175,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.024007112,0.020577524,0.01371835,0.006859175,0.0,0.0,0.006859175,0.030866288,0.0548734,0.072021335,0.082310095,0.06859175,0.048014224,0.037725464,0.044584636,0.05144381,0.048014224,0.05144381,0.048014224,0.037725464,0.024007112,0.01371835,0.01371835,0.01371835,0.020577524,0.048014224,0.0548734,0.048014224,0.041155048,0.041155048,0.05144381,0.07545093,0.09259886,0.09602845,0.07888051,0.072021335,0.061732575,0.06859175,0.1097468,0.17833854,0.23664154,0.25721905,0.24350071,0.34638834,0.5418748,0.6276145,0.5761707,0.5418748,0.5144381,0.5007198,0.5041494,0.5178677,0.58302987,0.66876954,0.764798,0.85396725,0.8711152,0.9294182,1.0048691,1.0666018,1.0837497,1.0288762,1.0563129,1.1934965,1.3958421,1.5536032,1.821111,2.1469216,2.3732746,2.5961976,3.1792276,4.0229063,4.8322887,5.06893,4.8117113,4.7774153,5.1169443,5.90232,6.694555,7.3290286,7.8949103,8.333898,7.6685576,6.831738,6.279575,5.9743414,6.101236,5.861165,5.593657,5.453044,5.425607,4.9660425,4.897451,5.0140567,5.0346346,4.5990767,4.2766957,3.6765177,2.760818,1.8142518,1.4747226,1.2723769,1.2380811,1.4918705,1.7971039,1.5810398,1.3924125,1.3821237,1.6324836,2.0474637,2.369845,2.5207467,2.4452958,2.2086544,1.8759843,1.5055889,1.1420527,1.0220171,0.88826317,0.64476246,0.33952916,0.19891608,0.1371835,0.14404267,0.22292319,0.36696586,0.52815646,0.6310441,0.6824879,0.69963586,0.72021335,0.7682276,0.7956643,0.8025235,0.7888051,0.7442205,0.6824879,0.61389613,0.52815646,0.44584638,0.42869842,0.4389872,0.47328308,0.65848076,0.97057325,1.2449403,1.488441,1.8142518,1.99602,1.9685832,1.845118,1.7730967,1.7525192,1.7456601,1.7353712,1.7319417,1.9582944,2.1469216,2.3629858,2.6476414,3.0489032,3.309552,3.4810312,3.5702004,3.590778,3.542764,3.3678548,3.117495,2.8019729,2.4898806,2.3218307,2.177788,2.085189,1.9994495,1.978872,2.1469216,2.335549,2.4041407,2.644212,2.9974594,3.0386145,2.651071,2.5893385,2.4761622,2.2120838,1.9720128,1.9925903,2.287535,2.6990852,3.0969174,3.3815732,2.8980014,2.8054025,2.9322972,3.175798,3.4844608,3.6868064,4.081209,4.650521,5.219832,5.4667625,5.686256,5.9743414,6.2075534,6.351596,6.444195,6.5950966,6.715132,7.0032177,7.3839016,7.500508,7.5553813,7.840037,8.375052,9.084977,9.81205,10.597425,11.447963,12.456262,13.591455,14.712931,15.560039,16.204802,17.017612,18.156237,19.572655,20.165974,20.244854,20.03565,19.637817,19.058218,20.045938,21.352612,22.806757,24.158014,25.090862,24.552416,23.626429,22.546108,21.27716,19.548649,18.20082,16.993607,16.060759,15.450292,15.148488,15.055889,14.987297,14.791811,14.445422,14.068168,13.841815,12.579727,10.998687,9.619993,8.748878,7.8983397,7.2535777,6.5950966,5.8405876,5.0140567,4.389872,3.8925817,3.4535947,3.1312134,3.1140654,3.4021509,3.525616,3.40901,3.210094,3.3266997,3.3815732,3.6044965,4.0537724,4.602506,4.9420357,4.9180284,4.773986,4.866585,5.127233,5.0620713,4.887162,4.8322887,5.178677,5.7925735,6.138962,6.2075534,6.701414,7.4765005,8.2310095,8.512236,9.115844,9.602845,10.086417,10.741467,11.842365,12.47341,12.47341,12.106443,11.753197,11.910957,12.202472,12.322508,12.339656,12.566009,13.560589,13.474849,12.713481,9.757176,5.7136927,4.32471,4.2183924,4.3007026,4.6916757,5.4016004,6.324159,7.7714453,12.21619,14.846684,14.79867,15.141628,15.707511,15.844694,15.522313,14.637479,13.001566,12.010415,11.05356,10.336777,10.422516,12.21619,16.386568,18.893597,19.027351,17.809847,17.991615,18.03277,17.785841,17.175373,16.37971,15.824117,15.309678,14.671775,13.639469,12.483699,12.020704,11.856084,11.235329,10.072699,8.831187,8.543102,9.253027,9.431366,9.201583,8.663138,7.870903,6.759717,6.3961806,6.6396813,7.0718093,7.006647,6.3035817,6.1766872,6.385892,6.464772,5.7102633,5.0174866,4.8117113,5.15467,5.813151,6.252138,6.8214493,7.682276,8.872343,10.131001,10.912948,11.036412,11.417097,11.838936,12.034423,11.688034,11.30735,10.782623,10.14129,9.424506,8.683716,7.9257765,7.250148,6.5813785,5.9434752,5.456474,5.535354,6.0052075,6.835168,7.98065,9.366203,9.39021,8.621983,7.610255,7.051232,7.7920227,8.834618,7.949784,6.121814,4.3452873,3.6079261,6.142391,9.836057,12.319078,12.579727,10.9541025,8.158989,6.0875177,4.4859004,3.2066643,2.1915064,1.2792361,0.72021335,0.3566771,0.11317638,0.01371835,0.048014224,0.07888051,0.09602845,0.08573969,0.041155048,0.1097468,0.15433143,0.16119061,0.13032432,0.048014224,0.024007112,0.034295876,0.048014224,0.09259886,0.25378948,0.30866286,0.29494452,0.2469303,0.17490897,0.07888051,0.06859175,0.058302987,0.034295876,0.01371835,0.037725464,0.07545093,0.0548734,0.024007112,0.0034295875,0.0,0.01371835,0.09259886,0.18862732,0.22292319,0.072021335,0.037725464,0.072021335,0.116605975,0.12003556,0.024007112,0.024007112,0.01371835,0.0034295875,0.0,0.006859175,0.058302987,0.1097468,0.15776102,0.20920484,0.26750782,0.18862732,0.08573969,0.0274367,0.024007112,0.030866288,0.020577524,0.0274367,0.034295876,0.041155048,0.05144381,0.061732575,0.058302987,0.041155048,0.017147938,0.0,0.0,0.061732575,0.106317215,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.006859175,0.006859175,0.006859175,0.006859175,0.006859175,0.010288762,0.01371835,0.006859175,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.010288762,0.01371835,0.0,0.0,0.0,0.0274367,0.06859175,0.061732575,0.048014224,0.044584636,0.044584636,0.044584636,0.0548734,0.08573969,0.10288762,0.106317215,0.09259886,0.08573969,0.072021335,0.06859175,0.07545093,0.08916927,0.09602845,0.08916927,0.07545093,0.08573969,0.10288762,0.06859175,0.06859175,0.058302987,0.048014224,0.044584636,0.037725464,0.020577524,0.061732575,0.106317215,0.14061308,0.17490897,0.01371835,0.0034295875,0.0034295875,0.006859175,0.01371835,0.020577524,0.010288762,0.024007112,0.07888051,0.14747226,0.13032432,0.08573969,0.061732575,0.058302987,0.058302987,0.05144381,0.037725464,0.0274367,0.041155048,0.06859175,0.07545093,0.058302987,0.030866288,0.017147938,0.024007112,0.048014224,0.072021335,0.058302987,0.037725464,0.030866288,0.037725464,0.044584636,0.037725464,0.030866288,0.0274367,0.034295876,0.0274367,0.0274367,0.024007112,0.020577524,0.037725464,0.020577524,0.017147938,0.020577524,0.0274367,0.0274367,0.041155048,0.0548734,0.06859175,0.08573969,0.11317638,0.10288762,0.09945804,0.09602845,0.09602845,0.09602845,0.08573969,0.06516216,0.041155048,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.017147938,0.017147938,0.01371835,0.01371835,0.0,0.006859175,0.01371835,0.01371835,0.017147938,0.017147938,0.024007112,0.020577524,0.010288762,0.006859175,0.01371835,0.010288762,0.017147938,0.0274367,0.037725464,0.05144381,0.058302987,0.0548734,0.048014224,0.048014224,0.05144381,0.048014224,0.058302987,0.058302987,0.041155048,0.024007112,0.020577524,0.024007112,0.030866288,0.034295876,0.041155048,0.041155048,0.072021335,0.10288762,0.1097468,0.08916927,0.09945804,0.13032432,0.14404267,0.1371835,0.12689474,0.1371835,0.16462019,0.22292319,0.2709374,0.23664154,0.2194936,0.22292319,0.37382504,0.6379033,0.83681935,0.89855194,0.90541106,0.9362774,1.0048691,1.0700313,1.1214751,1.1694894,1.2003556,1.2175035,1.2620882,1.3581166,1.5741806,1.7730967,1.8862731,1.9068506,2.0268862,2.270387,2.5207467,2.6716487,2.620205,2.5996273,2.6407824,2.750529,2.9906003,3.4981792,3.8274195,4.149801,4.1600895,3.974892,4.1635194,5.0414934,6.433906,7.4627824,7.8606143,7.9875093,7.81603,6.7940125,6.029215,5.936616,6.2555676,6.9552035,6.8214493,6.5162163,6.3824625,6.433906,6.334448,6.40304,6.5882373,6.8111606,6.948344,6.2212715,5.2815647,4.1189346,2.9185789,2.07833,1.7010754,1.5810398,1.7559488,1.99602,1.7936742,1.6496316,1.6804979,1.9720128,2.393852,2.603057,2.633923,2.6613598,2.4452958,1.9720128,1.4815818,1.0906088,1.138623,1.1214751,0.8471081,0.42869842,0.2469303,0.24007112,0.31209245,0.38754338,0.432128,0.5761707,0.69963586,0.7956643,0.881404,0.9945804,1.08032,1.1351935,1.1660597,1.1523414,1.08032,0.96371406,0.83338976,0.7305021,0.6824879,0.71678376,0.7888051,0.90541106,1.1866373,1.5913286,1.8965619,2.0989075,2.435007,2.5996273,2.5241764,2.369845,2.369845,2.4727325,2.5653315,2.603057,2.5756202,2.819121,2.976882,3.100347,3.234101,3.40901,3.5564823,3.7142432,3.8857226,3.9268777,3.549623,3.3061223,3.1346428,2.952875,2.719663,2.4384367,2.2566686,2.2498093,2.3286898,2.4384367,2.5584722,2.551613,2.428148,2.5207467,2.7573884,2.6990852,2.153781,1.8416885,1.6427724,1.5021594,1.4472859,1.670209,2.085189,2.5893385,3.1552205,3.806842,3.4227283,3.2066643,3.1860867,3.3438478,3.6147852,3.82399,4.1155047,4.5442033,4.955754,5.0003386,5.31929,5.6656785,5.885172,6.0154963,6.2727156,6.5230756,6.5127864,6.608815,6.852316,6.9380555,6.992929,7.233,7.630832,8.131552,8.676856,9.448513,10.065839,10.762046,11.667457,12.826657,14.177915,15.4914465,16.808409,18.142517,19.459478,20.244854,20.7833,21.133118,21.11597,20.327166,20.591244,21.246294,22.398636,23.773901,24.720467,24.754763,24.068846,23.053686,21.901346,20.567236,19.109661,17.7927,16.846134,16.283682,15.913286,16.005884,16.21509,16.20137,15.741806,14.723219,14.352823,13.114742,11.787492,10.731179,9.89093,8.7145815,7.740579,6.9826403,6.341307,5.586798,4.931747,4.256118,3.6182148,3.1620796,3.1072063,3.3129816,3.4707425,3.508468,3.5118976,3.7348208,4.033195,4.1463714,4.266407,4.4104495,4.4275975,4.15323,4.0229063,4.1360826,4.48933,4.9694724,5.809721,6.1766872,6.2041235,6.1149545,6.2075534,6.392751,7.1678376,8.131552,8.868914,8.97523,9.342196,9.469091,9.410788,9.541112,10.569988,11.526843,12.21962,12.857523,13.574307,14.445422,14.38369,13.306799,12.075578,11.465111,12.168177,14.263655,14.819247,13.474849,10.669447,7.654839,5.2918534,4.496189,4.705394,5.586798,7.0375133,7.4799304,10.837497,14.503725,17.405157,19.994495,20.814167,20.899906,19.716698,17.250826,13.989287,13.419975,14.291091,13.279363,10.80663,11.043272,14.79524,18.252264,19.442331,18.78042,19.061647,18.759844,18.176813,17.477179,16.942162,16.976458,16.990177,16.767254,16.084764,15.049029,14.095605,13.474849,12.576297,11.290202,9.674867,7.963502,8.004657,8.22758,8.347616,8.080108,7.1266828,6.48535,6.6465406,7.023795,7.4044795,7.9292064,7.8983397,7.291303,7.366754,8.093826,8.14527,7.936065,7.48336,7.284444,7.377043,7.3564653,7.3118806,7.3221693,7.939495,9.448513,11.869802,10.676306,10.024684,9.794902,9.736599,9.455373,9.668007,9.685155,9.225591,8.570539,8.567109,9.033533,9.9698105,12.22648,14.822677,14.908417,12.847235,9.187865,6.509357,5.8200097,6.557371,7.407909,8.1487,7.846896,6.708273,6.0532217,5.535354,5.693115,6.0326443,6.475061,7.3427467,8.879202,11.005547,11.773774,10.4533825,7.5210853,5.6485305,4.698535,3.99204,3.1963756,2.3252604,1.4438564,0.939707,0.5658819,0.2503599,0.09602845,0.048014224,0.030866288,0.020577524,0.01371835,0.024007112,0.11317638,0.17490897,0.18862732,0.14404267,0.048014224,0.030866288,0.044584636,0.08916927,0.21263443,0.5144381,0.4081209,0.3018037,0.20920484,0.14061308,0.07888051,0.041155048,0.020577524,0.010288762,0.020577524,0.037725464,0.072021335,0.044584636,0.017147938,0.01371835,0.01371835,0.037725464,0.14404267,0.2709374,0.31895164,0.17147937,0.034295876,0.061732575,0.116605975,0.11317638,0.017147938,0.017147938,0.006859175,0.0,0.0,0.006859175,0.106317215,0.18862732,0.20920484,0.18519773,0.19548649,0.17490897,0.1097468,0.048014224,0.010288762,0.017147938,0.034295876,0.05144381,0.06859175,0.07888051,0.07545093,0.07545093,0.048014224,0.020577524,0.006859175,0.0,0.0,0.061732575,0.1097468,0.09602845,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.0034295875,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0,0.0034295875,0.010288762,0.044584636,0.09259886,0.09259886,0.07545093,0.06859175,0.07545093,0.07888051,0.07888051,0.09259886,0.106317215,0.1097468,0.106317215,0.09602845,0.08573969,0.07888051,0.08573969,0.09259886,0.09259886,0.09602845,0.082310095,0.082310095,0.106317215,0.116605975,0.12003556,0.106317215,0.10288762,0.10288762,0.09259886,0.07545093,0.11317638,0.15433143,0.18176813,0.20577525,0.01371835,0.0034295875,0.010288762,0.020577524,0.024007112,0.024007112,0.0034295875,0.006859175,0.05144381,0.12346515,0.1920569,0.12003556,0.07545093,0.048014224,0.030866288,0.024007112,0.024007112,0.0274367,0.030866288,0.0274367,0.024007112,0.01371835,0.006859175,0.006859175,0.01371835,0.037725464,0.05144381,0.058302987,0.058302987,0.05144381,0.044584636,0.05144381,0.041155048,0.030866288,0.024007112,0.024007112,0.0274367,0.037725464,0.037725464,0.0274367,0.01371835,0.010288762,0.034295876,0.048014224,0.041155048,0.01371835,0.017147938,0.020577524,0.024007112,0.041155048,0.09259886,0.08573969,0.09945804,0.09602845,0.07545093,0.06859175,0.06516216,0.058302987,0.041155048,0.024007112,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0274367,0.034295876,0.030866288,0.01371835,0.0034295875,0.0034295875,0.010288762,0.01371835,0.010288762,0.0034295875,0.010288762,0.01371835,0.01371835,0.020577524,0.034295876,0.010288762,0.01371835,0.034295876,0.06516216,0.09945804,0.106317215,0.09259886,0.061732575,0.030866288,0.0274367,0.041155048,0.06516216,0.06859175,0.048014224,0.0274367,0.037725464,0.048014224,0.0548734,0.061732575,0.06859175,0.08573969,0.14747226,0.19548649,0.1920569,0.1371835,0.106317215,0.13375391,0.17147937,0.19548649,0.1920569,0.23664154,0.29151493,0.35324752,0.36696586,0.23321195,0.19891608,0.22978236,0.3841138,0.65505123,0.99801,1.2037852,1.313532,1.5261664,1.8519772,2.07833,2.0646117,1.8588364,1.6290541,1.4747226,1.4404267,1.7079345,2.2120838,2.6407824,2.8568463,2.8980014,3.275256,3.8377085,4.3178506,4.4859004,4.125794,3.806842,3.642222,3.625074,3.799983,4.273266,4.057202,3.6113555,3.234101,3.1895163,3.707384,5.099797,7.051232,7.949784,7.466212,6.56766,5.675967,5.4907694,5.761707,6.2727156,6.8557453,7.298162,7.1541195,6.927767,6.8557453,6.90033,7.0546613,7.140401,7.3358874,7.7885933,8.618553,7.3598948,6.1904054,5.0929375,3.9851806,2.6853669,2.1880767,1.9891608,2.0097382,2.0886188,1.9925903,1.9994495,2.1126258,2.4247184,2.836269,3.0420442,3.0729103,3.0420442,2.74367,2.201795,1.6839274,1.2963841,1.3238207,1.3032433,1.0494537,0.6790583,0.39440256,0.44927597,0.5761707,0.6001778,0.42869842,0.51100856,0.65505123,0.85396725,1.0906088,1.3409687,1.4747226,1.5604624,1.6016173,1.605047,1.5570327,1.5330256,1.5330256,1.5501735,1.5981878,1.7010754,1.8382589,2.0234566,2.2841053,2.5756202,2.7882545,2.867135,3.0283258,3.1037767,3.0626216,2.9974594,3.0660512,3.2512488,3.4055803,3.4535947,3.3678548,3.4021509,3.391862,3.333559,3.2272418,3.0660512,3.0454736,3.1312134,3.3369887,3.4021509,2.7985435,2.6304936,2.6407824,2.6853669,2.6545007,2.4658735,2.428148,2.585909,2.726522,2.719663,2.5173173,2.2155135,1.9582944,1.821111,1.7833855,1.7422304,1.611906,1.4198492,1.2758065,1.2380811,1.3203912,1.8588364,2.2635276,2.6236343,3.1209247,4.012617,3.7211025,3.4535947,3.3747141,3.5187566,3.782835,3.9131594,4.0366244,4.2115335,4.4584637,4.756838,5.103226,5.4804807,5.8508763,6.228131,6.684266,7.082098,7.0752387,6.8728933,6.6396813,6.48535,6.691125,6.9620624,7.233,7.4799304,7.73029,8.412778,9.019815,9.688584,10.621432,12.061859,13.824667,15.46744,16.890718,18.005335,18.732407,19.603521,20.570665,21.764162,22.745024,22.504953,22.175713,22.02824,22.53239,23.496103,24.075705,24.164873,23.612709,22.86163,22.072824,21.160555,20.063087,19.061647,18.11165,17.240536,16.527182,16.736387,17.29884,17.583494,16.969599,14.846684,13.71492,12.734058,11.928105,11.187314,10.251037,9.067829,8.008087,7.2192817,6.6533995,6.0532217,5.4496145,4.6676683,3.9680326,3.4913201,3.2718265,3.223812,3.2546785,3.5153272,4.0091877,4.5853586,5.0414934,5.1066556,5.0483527,4.931747,4.636802,4.0434837,3.9783216,4.3349986,5.07236,6.200694,7.857185,8.340756,8.018375,7.394191,7.085528,7.010077,7.274155,8.045813,9.057541,9.595985,9.815479,9.945804,9.674867,9.256456,9.5033865,10.192734,11.05699,12.404818,13.985858,14.96329,15.018164,13.985858,12.926115,12.418536,12.562579,16.13278,18.04992,18.732407,17.95389,14.836395,8.772884,5.8988905,4.605936,4.4413157,6.135532,7.205563,9.091836,12.274493,17.072487,23.612709,25.817934,26.579304,25.228045,21.880768,17.449741,15.971589,18.28999,17.326277,12.566009,10.062409,12.000127,14.915276,17.264544,18.492336,19.006773,18.684393,18.37916,18.241976,18.28313,18.36544,18.420315,18.245405,17.916164,17.28512,15.985307,14.627191,13.454271,12.617453,11.828648,10.336777,9.057541,8.176137,7.706283,7.390761,6.708273,6.6431108,7.181556,7.548522,7.6925645,8.272165,8.790032,7.5279446,7.222711,8.471081,9.743458,10.803201,11.38623,11.423956,10.840926,9.582268,8.097256,6.759717,6.4887795,8.203573,12.8197975,11.201033,10.30591,9.839486,9.338767,8.196714,8.210432,8.567109,8.39563,8.1384115,9.571979,10.861504,12.881531,17.494326,23.10856,24.699888,21.476076,14.685493,8.964942,6.1458206,5.2438393,6.2075534,8.258447,9.575408,9.39021,7.970361,6.975781,7.3701835,8.429926,9.716022,11.087856,10.333347,9.016385,7.2638664,5.0243454,2.061182,1.3375391,1.1660597,1.1351935,1.0631721,0.9877212,0.9294182,0.85739684,0.6824879,0.432128,0.25721905,0.12346515,0.06516216,0.044584636,0.044584636,0.058302987,0.06859175,0.09602845,0.11317638,0.09602845,0.0548734,0.0274367,0.030866288,0.106317215,0.274367,0.5453044,0.23664154,0.06516216,0.0034295875,0.0034295875,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.0,0.010288762,0.020577524,0.024007112,0.0274367,0.0274367,0.07545093,0.18862732,0.31209245,0.37382504,0.30523327,0.116605975,0.08573969,0.07545093,0.041155048,0.041155048,0.041155048,0.020577524,0.0034295875,0.010288762,0.034295876,0.18176813,0.2469303,0.26064864,0.2469303,0.19548649,0.15433143,0.12346515,0.06859175,0.0034295875,0.0034295875,0.030866288,0.061732575,0.10288762,0.14061308,0.16119061,0.12346515,0.048014224,0.006859175,0.0034295875,0.0,0.0,0.0,0.0034295875,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.01371835,0.024007112,0.06516216,0.116605975,0.13032432,0.11317638,0.11317638,0.13032432,0.15090185,0.15090185,0.15090185,0.14061308,0.12689474,0.12003556,0.12003556,0.106317215,0.1097468,0.106317215,0.09602845,0.09602845,0.116605975,0.116605975,0.116605975,0.12346515,0.14404267,0.1371835,0.1371835,0.14404267,0.15090185,0.14061308,0.14061308,0.1371835,0.14747226,0.16462019,0.17147937,0.0,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.017147938,0.058302987,0.106317215,0.13032432,0.12689474,0.1097468,0.08573969,0.061732575,0.061732575,0.041155048,0.024007112,0.01371835,0.0,0.0,0.010288762,0.0274367,0.048014224,0.061732575,0.037725464,0.048014224,0.06859175,0.06859175,0.044584636,0.06859175,0.09602845,0.08916927,0.061732575,0.061732575,0.072021335,0.08573969,0.09259886,0.08573969,0.061732575,0.048014224,0.0548734,0.061732575,0.061732575,0.061732575,0.08573969,0.06516216,0.06516216,0.10288762,0.15090185,0.07888051,0.08916927,0.09945804,0.07888051,0.030866288,0.017147938,0.01371835,0.01371835,0.01371835,0.0,0.01371835,0.01371835,0.010288762,0.0034295875,0.01371835,0.0274367,0.048014224,0.048014224,0.0274367,0.01371835,0.01371835,0.01371835,0.010288762,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.020577524,0.044584636,0.020577524,0.024007112,0.030866288,0.041155048,0.07545093,0.11317638,0.10288762,0.072021335,0.05144381,0.07545093,0.08916927,0.09259886,0.09259886,0.08916927,0.07545093,0.07545093,0.07545093,0.06859175,0.06859175,0.106317215,0.17833854,0.19891608,0.216064,0.2469303,0.26064864,0.20920484,0.216064,0.23664154,0.24007112,0.22978236,0.3018037,0.32924038,0.31895164,0.26750782,0.18176813,0.25721905,0.37382504,0.5453044,0.764798,1.0220171,1.0837497,1.2620882,1.9239986,2.9220085,3.6147852,3.4947495,2.6750782,2.037175,1.8691251,1.8931323,2.2086544,2.8945718,3.5153272,3.899441,4.1189346,4.290414,4.5819287,4.8494368,5.0277753,5.127233,4.9934793,4.9488945,4.914599,4.7602673,4.3349986,4.431027,4.3624353,4.0846386,4.1360826,5.662249,7.6376915,9.414218,9.678296,8.447074,7.0786686,6.385892,6.7322803,6.883182,6.574519,6.4990683,6.7700057,6.944915,7.1095347,7.267296,7.3393173,7.143831,7.140401,7.233,7.3358874,7.3839016,6.1766872,5.2506986,4.537344,3.9440255,3.357566,3.1140654,3.0523329,3.1723683,3.2855449,3.0043187,2.9460156,3.0386145,3.1620796,3.2992632,3.5564823,3.6044965,3.175798,2.6579304,2.2463799,1.9514352,1.7696671,1.4678634,1.1626302,0.89855194,0.64133286,0.39783216,0.44584638,0.5693115,0.6241849,0.5658819,0.5761707,0.7613684,1.0734608,1.4267083,1.6942163,1.8759843,1.99602,2.0440342,2.0577524,2.1057668,2.435007,2.976882,3.474172,3.8137012,3.998899,4.0846386,4.1772375,4.3109913,4.4859004,4.6676683,4.8151407,4.8254294,4.695105,4.461893,4.180667,3.9474552,3.8720043,3.8479972,3.8102717,3.724532,3.4913201,3.2032347,2.8945718,2.603057,2.3972816,2.335549,2.301253,2.277246,2.287535,2.3972816,2.2360911,1.8416885,1.5055889,1.4027013,1.587899,1.978872,2.294394,2.1194851,1.529596,1.1146159,1.3581166,1.8759843,2.335549,2.5721905,2.609916,2.3389788,2.0714707,1.8142518,1.6016173,1.4815818,2.5070283,3.1277838,3.3232703,3.316411,3.5873485,3.3541365,3.0111778,2.784825,2.7711067,2.9288676,3.2821152,3.7553983,4.1429415,4.4275975,4.804852,5.2575574,5.7651367,6.1801167,6.4407654,6.560801,6.5127864,6.574519,6.560801,6.4236174,6.2418494,6.5813785,6.824879,6.999788,7.143831,7.2775846,7.377043,7.6651278,8.213862,9.301042,11.413667,13.392539,15.138199,16.420864,17.254255,17.912735,18.656956,19.586374,21.404055,23.835632,25.619019,26.606739,26.891396,26.452408,25.4544,24.247183,23.36578,22.817045,22.323185,21.723007,20.965069,20.402617,19.70641,18.87645,17.933313,16.907866,16.87014,17.106783,17.487467,17.37429,15.638919,13.893259,12.404818,11.622872,11.410237,11.032983,10.432805,9.688584,8.711152,7.6857057,7.06495,6.7974424,5.693115,4.602506,3.882293,3.4192986,3.0900583,2.9151495,3.0489032,3.5599117,4.4241676,5.0483527,5.73427,6.2967224,6.468202,5.90575,5.086078,4.57164,4.530485,5.1512403,6.6533995,7.8503256,8.862054,9.949233,10.981539,11.444533,11.55428,11.526843,11.629731,11.794352,11.612583,11.135871,11.327928,11.321068,10.844356,10.2236,10.113853,10.672876,11.345076,11.763485,11.763485,11.900668,12.785502,13.978998,14.500296,12.816368,13.732068,15.748666,18.921034,22.038528,22.61127,14.850114,9.421077,5.6073756,3.4364467,3.6936657,5.0003386,6.3035817,8.704293,14.2533655,25.968836,30.399864,29.374416,26.006561,22.223726,18.766703,17.864721,18.296848,17.778982,15.05246,9.904649,10.220171,11.207891,12.6586075,14.404267,16.2974,17.857862,19.651537,21.311457,22.271742,21.757303,20.659836,19.123379,18.108221,17.658945,16.877,15.656067,14.363112,13.896688,14.095605,13.718349,11.97269,10.545981,9.314759,8.210432,7.233,7.1095347,7.281014,7.5553813,7.6376915,7.1266828,6.773435,6.8385973,7.486789,8.207003,7.8263187,10.683165,14.016724,15.755525,14.771234,10.864933,7.2021337,5.1066556,4.2869844,4.557922,5.813151,7.6685576,10.789482,12.600305,12.312219,10.8958,8.820899,8.676856,9.884071,12.027563,14.846684,13.077017,11.982979,11.681175,12.322508,14.1299,14.068168,12.617453,10.412228,8.611694,8.879202,11.211322,14.027013,16.475739,17.761833,17.151367,15.745236,14.140189,12.133881,9.866923,7.8263187,5.3741636,3.1415021,1.6804979,1.0597426,0.84024894,0.7888051,0.7510797,0.67219913,0.53844523,0.36696586,0.30523327,0.37382504,0.45270553,0.47671264,0.42869842,0.30523327,0.2469303,0.216064,0.20577525,0.22978236,0.2777966,0.24350071,0.2194936,0.21263443,0.15090185,0.06859175,0.0548734,0.08573969,0.106317215,0.044584636,0.010288762,0.010288762,0.010288762,0.0,0.0,0.01371835,0.006859175,0.006859175,0.01371835,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.0034295875,0.044584636,0.09602845,0.13375391,0.18176813,0.31895164,0.432128,0.37725464,0.20920484,0.19891608,0.19891608,0.09602845,0.024007112,0.034295876,0.106317215,0.216064,0.18862732,0.17147937,0.2194936,0.30523327,0.09602845,0.017147938,0.006859175,0.01371835,0.01371835,0.0034295875,0.017147938,0.048014224,0.08916927,0.1371835,0.08916927,0.048014224,0.030866288,0.024007112,0.0,0.0,0.0,0.01371835,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.01371835,0.01371835,0.024007112,0.048014224,0.082310095,0.106317215,0.12003556,0.14061308,0.15090185,0.15090185,0.15090185,0.15090185,0.16119061,0.16804978,0.16804978,0.16804978,0.15433143,0.15090185,0.13375391,0.106317215,0.106317215,0.16804978,0.15433143,0.12346515,0.106317215,0.106317215,0.12003556,0.13032432,0.15090185,0.16462019,0.15090185,0.15090185,0.14404267,0.14404267,0.15776102,0.18176813,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.010288762,0.01371835,0.020577524,0.037725464,0.044584636,0.061732575,0.09945804,0.18176813,0.2503599,0.14747226,0.06859175,0.037725464,0.020577524,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.037725464,0.048014224,0.034295876,0.08573969,0.11317638,0.08573969,0.020577524,0.0274367,0.05144381,0.07545093,0.08916927,0.09602845,0.1097468,0.11317638,0.10288762,0.072021335,0.037725464,0.034295876,0.034295876,0.048014224,0.06516216,0.072021335,0.08916927,0.09945804,0.09602845,0.082310095,0.09259886,0.06859175,0.08916927,0.09259886,0.058302987,0.030866288,0.017147938,0.01371835,0.020577524,0.030866288,0.037725464,0.030866288,0.0274367,0.030866288,0.044584636,0.07545093,0.058302987,0.044584636,0.034295876,0.0274367,0.01371835,0.01371835,0.006859175,0.0034295875,0.0,0.0034295875,0.010288762,0.0274367,0.0274367,0.017147938,0.020577524,0.017147938,0.048014224,0.072021335,0.082310095,0.09945804,0.116605975,0.15433143,0.1920569,0.2194936,0.23664154,0.18862732,0.15433143,0.1371835,0.12003556,0.08916927,0.06859175,0.058302987,0.0548734,0.06859175,0.09602845,0.17833854,0.2709374,0.30866286,0.29151493,0.28465575,0.29494452,0.36696586,0.4046913,0.3806842,0.33952916,0.37382504,0.36010668,0.31895164,0.25721905,0.17147937,0.23321195,0.26407823,0.3018037,0.38754338,0.5453044,0.6859175,0.8128122,1.0014396,1.4987297,2.7128036,3.74168,4.3178506,4.201245,3.5873485,3.1243541,3.0797696,3.6010668,4.1943855,4.65395,5.0586414,5.4633327,5.6142344,5.6210938,5.5730796,5.552502,5.809721,6.121814,6.2692857,6.0840883,5.4324665,4.846007,4.4687524,4.3007026,4.5030484,5.40503,6.433906,7.2638664,7.507367,7.377043,7.689135,7.864044,7.997798,7.8949103,7.5690994,7.233,6.9346256,6.632822,6.7631464,7.281014,7.658269,7.257007,6.975781,6.9552035,7.2295704,7.7268605,7.239859,6.3653145,5.456474,4.846007,4.846007,4.5613513,4.2286816,3.8685746,3.566771,3.4810312,3.508468,3.6044965,3.74168,3.8308492,3.724532,3.433017,2.9048605,2.486451,2.2566686,2.0508933,1.8691251,1.646202,1.3443983,0.980862,0.6173257,0.42183927,0.47328308,0.58645946,0.64819205,0.6241849,0.922559,1.2723769,1.646202,2.0028791,2.2806756,2.609916,2.9048605,3.1277838,3.309552,3.532475,3.8034124,4.0949273,4.4104495,4.715683,4.938606,5.051782,5.07236,5.0140567,4.911169,4.839148,4.8288593,4.7842746,4.671098,4.48933,4.280125,4.2526884,4.197815,4.0949273,3.9268777,3.6868064,3.5118976,3.292404,3.0146074,2.6990852,2.3835633,2.194936,2.0268862,1.7833855,1.5501735,1.5913286,1.8313997,2.2463799,2.386993,2.177788,1.8931323,1.5398848,1.5536032,1.587899,1.5638919,1.6770682,2.1915064,2.6407824,3.0146074,3.2958336,3.4398763,3.4844608,3.3952916,3.2203827,2.9700227,2.603057,3.1312134,3.6593697,3.998899,4.1360826,4.2218223,3.7039545,2.7745364,2.07833,1.8691251,1.978872,2.3904223,2.9494452,3.532475,4.0846386,4.6608095,5.2575574,5.5319247,5.6039457,5.5833683,5.5490727,5.861165,6.042933,6.0737996,5.936616,5.6176643,6.2247014,6.6396813,6.866034,6.9723516,7.0958166,7.301592,7.699424,8.436785,9.527394,10.840926,12.593445,14.812388,16.441442,17.250826,17.840714,18.488907,19.346302,20.793589,22.755312,24.703318,26.483274,27.405834,27.416122,26.507282,24.723896,23.451519,22.731306,22.326614,21.891056,20.978786,20.416334,19.87789,19.308577,18.526632,17.247395,16.674654,16.698662,17.134218,17.422304,16.616352,15.426285,14.421415,13.488567,12.689473,12.253916,12.133881,11.55771,10.676306,9.685155,8.858624,8.532814,7.5107965,6.307011,5.2026844,4.2595477,3.6765177,3.1689389,2.7813954,2.620205,2.8637056,3.2615378,3.758828,4.290414,4.6916757,4.695105,4.7774153,5.079219,5.4667625,6.036074,7.130112,8.196714,8.995808,9.774324,10.539123,11.05356,11.046701,11.122152,11.605724,12.576297,13.858963,13.937843,13.728639,12.836946,11.454823,10.347065,10.106995,10.189304,10.600855,11.063849,10.995257,11.266195,11.80464,12.682614,13.289652,12.329367,11.537132,12.164746,14.664916,18.21111,20.697561,19.582945,15.107333,10.734609,7.438775,3.6936657,4.1189346,4.839148,6.2487082,9.191295,14.973578,22.61813,24.994833,23.880217,21.20514,19.047928,18.907316,19.390888,19.11652,17.171944,13.125031,10.854645,9.767465,9.901219,11.067279,12.843805,14.891269,17.151367,20.471207,24.291767,26.641035,23.883648,20.845032,18.499195,17.257685,16.973028,16.05733,15.261664,14.819247,14.692352,14.596324,13.077017,11.691463,10.497967,9.551401,8.916927,8.385342,7.7851634,7.239859,7.0272245,7.589677,8.093826,7.857185,7.589677,7.4284863,6.924337,7.1541195,9.647429,12.847235,15.117621,14.747226,9.784613,7.4970784,6.3790326,5.7582774,5.7754254,6.2075534,7.181556,8.038953,8.745448,9.904649,9.530824,8.755736,8.008087,8.309891,11.30735,13.090735,14.016724,14.023583,13.334236,12.445972,10.947243,9.863494,9.256456,9.225591,9.89436,11.746337,13.227919,14.328816,14.898128,14.647768,13.255356,11.108434,8.700864,6.355026,4.2389703,3.0660512,2.1091962,1.4027013,0.9602845,0.77851635,0.7099246,0.7373613,0.94656616,1.2072148,1.1832076,0.94656616,0.66191036,0.59674823,0.71678376,0.70649505,0.42869842,0.31209245,0.274367,0.2777966,0.3018037,0.45956472,0.5041494,0.41498008,0.2503599,0.14061308,0.11317638,0.09259886,0.072021335,0.041155048,0.010288762,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.0034295875,0.01371835,0.01371835,0.020577524,0.030866288,0.041155048,0.041155048,0.037725464,0.037725464,0.037725464,0.037725464,0.037725464,0.09259886,0.18176813,0.28465575,0.35324752,0.31895164,0.23321195,0.21263443,0.25721905,0.30866286,0.26407823,0.17833854,0.08916927,0.07888051,0.17490897,0.32924038,0.2777966,0.28122616,0.39783216,0.548734,0.53844523,0.19548649,0.06859175,0.07545093,0.15433143,0.2709374,0.12346515,0.037725464,0.006859175,0.0034295875,0.0,0.0,0.006859175,0.020577524,0.0548734,0.15090185,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.006859175,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.017147938,0.024007112,0.01371835,0.034295876,0.041155048,0.061732575,0.09602845,0.12003556,0.14061308,0.16462019,0.17833854,0.17490897,0.16462019,0.14404267,0.12003556,0.11317638,0.12003556,0.13032432,0.12003556,0.1371835,0.15433143,0.15776102,0.16804978,0.17147937,0.15090185,0.12346515,0.11317638,0.13032432,0.15433143,0.14747226,0.14061308,0.14404267,0.15090185,0.17147937,0.16804978,0.16462019,0.16804978,0.18176813,0.006859175,0.006859175,0.0034295875,0.0,0.0034295875,0.010288762,0.01371835,0.01371835,0.017147938,0.024007112,0.041155048,0.058302987,0.072021335,0.11317638,0.16119061,0.14061308,0.07888051,0.044584636,0.017147938,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.06516216,0.058302987,0.061732575,0.058302987,0.044584636,0.01371835,0.024007112,0.030866288,0.05144381,0.08916927,0.116605975,0.09259886,0.10288762,0.11317638,0.106317215,0.08573969,0.08573969,0.08573969,0.08916927,0.09945804,0.10288762,0.12346515,0.14061308,0.13032432,0.11317638,0.15090185,0.12346515,0.08916927,0.06516216,0.0548734,0.030866288,0.041155048,0.07545093,0.07888051,0.048014224,0.037725464,0.037725464,0.0274367,0.024007112,0.030866288,0.044584636,0.044584636,0.030866288,0.020577524,0.020577524,0.01371835,0.030866288,0.030866288,0.020577524,0.010288762,0.017147938,0.030866288,0.024007112,0.01371835,0.006859175,0.006859175,0.020577524,0.05144381,0.07545093,0.09945804,0.13375391,0.16119061,0.18519773,0.216064,0.2469303,0.274367,0.1920569,0.15433143,0.14747226,0.15090185,0.12689474,0.09602845,0.08573969,0.08916927,0.1097468,0.16462019,0.21263443,0.274367,0.3018037,0.29494452,0.29151493,0.32238123,0.40126175,0.41840968,0.36010668,0.31209245,0.32924038,0.34981793,0.32924038,0.26750782,0.20577525,0.26407823,0.26064864,0.2469303,0.26407823,0.32581082,0.45613512,0.490431,0.4698535,0.5590228,1.0666018,2.0406046,2.9082901,3.8479972,4.557922,4.266407,3.8308492,3.5530527,3.6696587,4.1943855,4.945465,5.645101,5.802862,5.7754254,5.744559,5.7239814,5.874883,6.2658563,6.447624,6.183546,5.470192,4.712253,4.2286816,3.9954693,3.998899,4.2526884,5.6142344,7.0203657,8.31675,9.22216,9.318189,9.091836,8.556821,7.7097125,6.8728933,6.684266,6.625963,6.3824625,6.1321025,5.950334,5.796003,5.4599032,5.7582774,6.228131,6.636252,6.9963584,6.742569,6.3207297,5.909179,5.686256,5.830299,5.113515,4.4241676,3.8205605,3.4535947,3.5633414,3.6353626,3.7142432,3.8274195,3.8548563,3.5118976,3.000889,2.4007113,1.9102802,1.6084765,1.471293,1.4644338,1.2517995,1.0597426,0.96714365,0.922559,0.7888051,0.77508676,0.8265306,0.91912943,1.0631721,1.5741806,2.1469216,2.7299516,3.2375305,3.5599117,3.9646032,4.2835546,4.4447455,4.57507,5.0346346,5.4736214,5.8474464,6.217842,6.464772,6.2727156,5.7411294,5.442755,5.2438393,5.079219,4.9660425,4.866585,4.7671266,4.633373,4.461893,4.2766957,4.2046742,4.105216,3.9611735,3.7451096,3.4124396,3.0351849,2.6373527,2.2326615,1.8828435,1.6942163,1.6564908,1.6667795,1.5810398,1.4164196,1.3512574,1.5090185,2.0474637,2.2155135,1.8588364,1.4198492,1.1077567,1.0597426,1.2072148,1.5158776,1.978872,2.3972816,2.8808534,3.316411,3.5702004,3.4638834,3.3815732,3.2272418,3.0386145,2.8499873,2.7093742,2.9665933,3.223812,3.357566,3.3301294,3.199805,2.8019729,2.2738166,1.7902447,1.4815818,1.4472859,1.7799559,2.3664153,3.0454736,3.7348208,4.431027,5.096367,5.267846,5.188966,5.0449233,4.9660425,5.346727,5.593657,5.6999745,5.6039457,5.195825,5.56965,5.9983487,6.495639,6.9860697,7.3050213,7.5450926,7.747438,8.203573,9.054111,10.275044,12.089295,14.078457,15.659496,16.70552,17.528622,18.094503,18.828436,19.668684,20.488356,21.088533,21.959648,22.62156,22.961088,22.916504,22.453508,22.227156,22.210009,22.316326,22.354052,22.02481,21.242865,19.922474,18.989626,18.53692,17.799559,17.223389,16.750105,16.849564,17.329706,17.319416,16.47231,15.446862,14.4145565,13.560589,13.070158,12.97413,12.579727,11.948683,11.14273,10.213311,9.541112,8.546532,7.4044795,6.258997,5.2026844,4.307562,3.4433057,2.7299516,2.2841053,2.2258022,2.428148,2.8122618,3.1723683,3.4192986,3.5804894,4.0606318,4.852866,5.6999745,6.550512,7.5690994,8.611694,9.421077,10.103564,10.624862,10.789482,10.666017,10.834066,11.413667,12.380811,13.560589,13.9309845,13.790371,12.833516,11.358793,10.257896,10.0041065,9.818909,9.853205,9.914937,9.493098,8.951223,8.81404,9.571979,10.97468,12.068718,11.749766,10.88894,11.146159,13.433694,17.902447,18.999914,17.857862,16.19794,13.6086035,7.5553813,6.3790326,6.5024977,6.90033,7.706283,10.209882,14.562028,19.185112,21.390337,20.797018,19.301718,17.600643,17.895588,18.303709,17.693241,15.707511,12.686044,10.203023,8.7145815,8.453933,9.414218,11.4033785,14.006435,17.676094,22.237446,26.884537,24.662163,21.45893,18.37916,16.355703,16.173935,15.63206,14.983868,14.483148,14.249936,14.277372,13.690913,12.768354,11.777204,10.930096,10.374502,9.716022,8.8929205,8.176137,7.7611566,7.7714453,7.939495,8.241299,8.498518,8.495089,7.970361,8.357904,9.623423,10.947243,11.88352,12.373952,11.372512,12.151029,13.231348,13.437123,11.893809,9.314759,8.22758,8.556821,9.750318,10.792912,9.335337,8.025234,7.157549,7.4113383,9.863494,12.596875,15.097044,16.938732,17.576635,16.37285,13.615462,11.177026,9.270175,8.179566,8.251588,9.743458,10.930096,11.571428,11.598865,11.111863,9.829198,8.021805,6.0154963,4.1189346,2.6167753,2.1091962,1.5707511,1.138623,0.8745448,0.7613684,0.58645946,0.5624523,0.6859175,0.85739684,0.8848336,0.7579388,0.59331864,0.5521636,0.65505123,0.77851635,0.66533995,0.5658819,0.4629943,0.39440256,0.4389872,0.5796003,0.61389613,0.5453044,0.41840968,0.34638834,0.2469303,0.18176813,0.12689474,0.07888051,0.044584636,0.024007112,0.01371835,0.010288762,0.006859175,0.0,0.006859175,0.017147938,0.020577524,0.020577524,0.024007112,0.024007112,0.034295876,0.044584636,0.06516216,0.09945804,0.14404267,0.10288762,0.0548734,0.030866288,0.017147938,0.07545093,0.21263443,0.38754338,0.50757897,0.4424168,0.35324752,0.29837412,0.2777966,0.274367,0.26064864,0.18519773,0.14747226,0.15090185,0.19891608,0.29151493,0.36696586,0.37382504,0.36696586,0.37725464,0.42526886,0.24007112,0.12689474,0.07888051,0.082310095,0.12346515,0.0548734,0.01371835,0.0034295875,0.010288762,0.010288762,0.0034295875,0.0034295875,0.006859175,0.024007112,0.072021335,0.01371835,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.01371835,0.010288762,0.01371835,0.024007112,0.024007112,0.030866288,0.034295876,0.041155048,0.05144381,0.061732575,0.07888051,0.08916927,0.10288762,0.12003556,0.13032432,0.14061308,0.15090185,0.15090185,0.1371835,0.10288762,0.072021335,0.05144381,0.048014224,0.061732575,0.10288762,0.09945804,0.1097468,0.12689474,0.14061308,0.14747226,0.13375391,0.12003556,0.1097468,0.1097468,0.12689474,0.14404267,0.13032432,0.116605975,0.1097468,0.116605975,0.12689474,0.13032432,0.1371835,0.15433143,0.17490897,0.0,0.0034295875,0.006859175,0.006859175,0.01371835,0.020577524,0.020577524,0.020577524,0.020577524,0.024007112,0.034295876,0.05144381,0.0548734,0.06859175,0.1097468,0.15776102,0.15090185,0.09602845,0.044584636,0.017147938,0.006859175,0.006859175,0.020577524,0.034295876,0.041155048,0.058302987,0.08573969,0.07545093,0.0548734,0.037725464,0.034295876,0.0274367,0.020577524,0.034295876,0.072021335,0.09602845,0.07888051,0.09945804,0.14404267,0.17490897,0.15776102,0.12003556,0.12689474,0.14404267,0.14404267,0.13375391,0.14061308,0.19548649,0.2469303,0.2777966,0.30866286,0.20920484,0.12346515,0.09259886,0.09259886,0.030866288,0.09259886,0.17147937,0.17147937,0.09945804,0.061732575,0.09259886,0.15433143,0.14747226,0.06516216,0.020577524,0.034295876,0.0274367,0.020577524,0.024007112,0.0274367,0.037725464,0.037725464,0.0274367,0.017147938,0.024007112,0.030866288,0.020577524,0.01371835,0.017147938,0.017147938,0.0274367,0.044584636,0.07888051,0.1371835,0.2194936,0.26064864,0.24007112,0.21263443,0.216064,0.23321195,0.17490897,0.15776102,0.16462019,0.17490897,0.17147937,0.16804978,0.17833854,0.19891608,0.24350071,0.34295875,0.31895164,0.31552204,0.32238123,0.32924038,0.31552204,0.32581082,0.3566771,0.32924038,0.25721905,0.24350071,0.26750782,0.30866286,0.31552204,0.28122616,0.26407823,0.32581082,0.29494452,0.26750782,0.28122616,0.31552204,0.3841138,0.34295875,0.25378948,0.17833854,0.15776102,0.6001778,1.0906088,2.0268862,3.069481,3.1312134,2.877424,2.5756202,2.6922262,3.3198407,4.190956,5.079219,5.6348124,5.7377,5.5593615,5.5833683,5.8165803,6.228131,6.416758,6.2075534,5.6828265,5.07236,4.5956473,4.2869844,4.139512,4.1292233,5.994919,7.936065,9.825768,11.125582,10.899229,9.97324,8.783174,7.4627824,6.385892,6.169828,6.3035817,6.4064693,5.926327,5.07236,4.8185706,5.219832,6.101236,6.6739774,6.677407,6.368744,5.9640527,5.7102633,5.6142344,5.6999745,6.001778,5.195825,4.431027,3.7759757,3.3850029,3.4776018,3.6147852,3.673088,3.5804894,3.2615378,2.6647894,2.1057668,1.6496316,1.3238207,1.1866373,1.313532,1.5673214,1.1626302,0.939707,1.155771,1.471293,1.2415106,1.2175035,1.371835,1.6942163,2.1915064,2.9220085,3.6182148,4.2389703,4.746549,5.0826488,5.439326,5.6965446,5.7754254,5.830299,6.2727156,6.64997,6.8969,7.1232533,7.2295704,6.924337,6.3447366,6.138962,5.8508763,5.3570156,4.8734436,4.7534084,4.5510626,4.3041325,4.0434837,3.7931237,3.625074,3.450165,3.2546785,3.0283258,2.7333813,2.2841053,1.8519772,1.5158776,1.2929544,1.1626302,1.1797781,1.2963841,1.4164196,1.4953002,1.5536032,1.6907866,1.9823016,1.9445761,1.5330256,1.1317638,1.1214751,1.1797781,1.4335675,1.937717,2.6647894,2.5138876,2.6545007,2.9460156,3.2581081,3.4638834,3.1277838,2.6956558,2.4212887,2.469303,2.9288676,3.210094,3.1449318,2.9254382,2.6476414,2.3321195,2.0234566,1.786815,1.5501735,1.3684053,1.3924125,1.7388009,2.2120838,2.7882545,3.4707425,4.280125,4.822,4.938606,4.8151407,4.633373,4.5853586,4.9831905,5.329579,5.5319247,5.456474,4.9523244,4.8905916,5.0757895,5.6348124,6.4544835,7.1884155,7.8194594,8.038953,8.371623,9.102125,10.261326,11.780633,13.255356,14.603184,15.79325,16.87014,17.20624,17.785841,18.38259,18.70497,18.413456,18.530062,18.708399,18.725548,18.735836,19.277712,20.093952,21.02337,21.719578,22.12084,22.44665,22.089973,20.467777,19.133669,18.567787,18.187103,18.28656,17.844143,17.665806,17.940172,18.21111,17.144508,15.858413,14.640909,13.677195,13.059869,12.895248,12.71691,12.435684,11.921246,10.995257,10.000677,8.913498,7.915488,7.023795,6.101236,5.103226,4.0503426,3.1346428,2.4624438,2.0920484,2.1674993,2.411,2.603057,2.6887965,2.784825,3.3541365,4.2183924,5.2026844,6.1732574,7.0203657,7.956643,8.961512,10.189304,11.447963,12.188754,12.521424,12.758065,13.087306,13.5503,14.023583,14.167625,13.533153,12.127021,10.360784,9.06097,9.318189,8.882631,8.323608,7.891481,7.517656,7.1712675,6.8214493,6.9723516,7.9257765,9.757176,10.768905,10.415657,9.589127,9.959522,13.989287,15.302819,15.590904,16.527182,16.62321,11.201033,9.259886,9.249598,9.187865,8.745448,9.225591,10.645439,15.422854,18.862732,19.342873,18.338005,15.604623,15.501736,16.438013,17.093063,16.403717,14.356253,12.308789,10.484249,9.112414,8.436785,9.369633,11.571428,15.090185,19.6241,24.504402,24.247183,21.249723,17.844143,15.536031,15.014734,14.726648,14.2190695,13.80409,13.656617,13.824667,13.598314,13.210771,12.867812,12.672326,12.624311,11.749766,10.693454,10.076128,9.81205,9.112414,8.820899,9.3764925,9.962952,10.244178,10.39508,11.64345,12.061859,11.543991,10.590566,10.299051,11.688034,14.342535,17.154797,19.082224,19.167965,15.830976,13.858963,13.258785,13.680624,14.407697,11.825217,9.6645775,8.81061,9.273604,10.179015,11.749766,14.153908,16.486027,17.86815,17.436022,15.313108,12.689473,10.254466,8.573969,8.080108,8.786603,9.534253,9.774324,9.325048,8.381912,7.7131424,6.5539417,5.079219,3.7176728,3.1689389,2.5447538,1.7593783,1.1420527,0.8162418,0.6962063,0.52815646,0.47328308,0.48014224,0.5212973,0.5624523,0.5555932,0.5212973,0.52472687,0.607037,0.7888051,0.8162418,0.75450927,0.6344737,0.52472687,0.53158605,0.69963586,0.72021335,0.6379033,0.53158605,0.52472687,0.4046913,0.31209245,0.24007112,0.17833854,0.1371835,0.106317215,0.08573969,0.07545093,0.072021335,0.0548734,0.061732575,0.07545093,0.08573969,0.08573969,0.08573969,0.06516216,0.058302987,0.058302987,0.06516216,0.09945804,0.19891608,0.16462019,0.09602845,0.061732575,0.09602845,0.1371835,0.25378948,0.42526886,0.5693115,0.5590228,0.53844523,0.50757897,0.39440256,0.24007112,0.18176813,0.16804978,0.24007112,0.30523327,0.31895164,0.3018037,0.28122616,0.26407823,0.20577525,0.1371835,0.16804978,0.14747226,0.09602845,0.044584636,0.01371835,0.0,0.0,0.0,0.0034295875,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.006859175,0.0,0.006859175,0.010288762,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.010288762,0.01371835,0.024007112,0.024007112,0.030866288,0.044584636,0.058302987,0.072021335,0.09259886,0.10288762,0.11317638,0.12346515,0.1371835,0.14404267,0.12346515,0.1097468,0.09259886,0.072021335,0.041155048,0.017147938,0.010288762,0.010288762,0.017147938,0.0548734,0.058302987,0.061732575,0.072021335,0.08573969,0.09259886,0.08573969,0.07545093,0.07545093,0.08573969,0.09602845,0.106317215,0.10288762,0.10288762,0.106317215,0.1097468,0.1097468,0.11317638,0.12003556,0.13375391,0.15090185,0.0034295875,0.01371835,0.01371835,0.020577524,0.0274367,0.0274367,0.0274367,0.0274367,0.0274367,0.024007112,0.01371835,0.024007112,0.048014224,0.09945804,0.16804978,0.22292319,0.24350071,0.16462019,0.08573969,0.048014224,0.037725464,0.037725464,0.058302987,0.082310095,0.08916927,0.05144381,0.09945804,0.12003556,0.106317215,0.07545093,0.06859175,0.034295876,0.0274367,0.044584636,0.072021335,0.09602845,0.11317638,0.14404267,0.19548649,0.2469303,0.22292319,0.1371835,0.15090185,0.1920569,0.21263443,0.19891608,0.17490897,0.26407823,0.39783216,0.50757897,0.5144381,0.33266997,0.2469303,0.22635277,0.20234565,0.07545093,0.15090185,0.22978236,0.22978236,0.16119061,0.11317638,0.16462019,0.30866286,0.3018037,0.14061308,0.041155048,0.044584636,0.037725464,0.030866288,0.034295876,0.041155048,0.034295876,0.024007112,0.024007112,0.030866288,0.0274367,0.0274367,0.034295876,0.041155048,0.05144381,0.058302987,0.05144381,0.0548734,0.09602845,0.18176813,0.3018037,0.34295875,0.29494452,0.23664154,0.21263443,0.216064,0.21263443,0.20920484,0.20920484,0.216064,0.23321195,0.274367,0.31552204,0.35324752,0.4115505,0.52472687,0.45270553,0.41840968,0.42526886,0.44927597,0.45613512,0.38754338,0.32581082,0.2503599,0.19548649,0.22635277,0.274367,0.32581082,0.36010668,0.3806842,0.42183927,0.47328308,0.432128,0.42869842,0.47671264,0.490431,0.42183927,0.33266997,0.26064864,0.22635277,0.2503599,0.23664154,0.2194936,0.216064,0.29494452,0.5590228,0.823101,1.2037852,1.7730967,2.568761,3.5976372,4.5853586,5.6176643,5.90232,5.562791,5.6519604,6.142391,6.540223,6.680836,6.5367937,6.2247014,5.7582774,5.3158607,5.0449233,5.0346346,5.2781353,7.1678376,8.89635,10.398509,11.379372,11.334786,10.244178,8.903209,7.613684,6.660259,6.3035817,6.3378778,6.694555,6.341307,5.5113473,5.7068334,6.8626046,7.7920227,8.032094,7.548522,6.7528577,6.2247014,5.8405876,5.6245236,5.6142344,5.8543057,5.23698,4.5784993,3.9440255,3.4638834,3.3541365,3.433017,3.3815732,2.9871707,2.270387,1.5090185,1.0460242,0.8711152,0.89512235,1.1043272,1.5741806,2.0577524,1.4815818,1.1592005,1.4953002,1.9685832,1.704505,1.8073926,2.201795,2.836269,3.7039545,4.712253,5.360445,5.7136927,5.9126086,6.1904054,6.4544835,6.684266,6.8557453,7.006647,7.222711,7.431916,7.6445503,7.459353,6.9346256,6.5710897,6.4887795,6.6293926,6.307011,5.429037,4.4756117,4.3041325,3.9714622,3.5976372,3.2512488,2.9631636,2.7368107,2.469303,2.177788,1.9102802,1.7525192,1.471293,1.2346514,1.138623,1.1214751,0.9877212,0.96371406,1.0734608,1.2312219,1.4198492,1.6873571,2.0440342,2.0577524,1.8416885,1.5364552,1.2998136,1.4850113,1.646202,1.9308578,2.452155,3.2855449,2.5653315,2.177788,2.153781,2.503599,3.2272418,2.7882545,2.201795,2.020027,2.4590142,3.4055803,3.7794054,3.4776018,2.9631636,2.4761622,2.037175,1.7353712,1.4232788,1.2620882,1.3169615,1.5570327,2.0131679,2.3149714,2.668219,3.216953,4.057202,4.386442,4.4927597,4.4104495,4.2938433,4.434457,4.9214582,5.4016004,5.6176643,5.4324665,4.8425775,4.4241676,4.2835546,4.6848164,5.6073756,6.7357097,7.8023114,8.375052,8.992378,9.853205,10.827208,11.664027,12.603734,13.6086035,14.671775,15.830976,16.03675,16.55119,17.243965,17.7927,17.689812,17.830425,17.772121,17.178804,16.506605,17.003895,18.149376,19.562366,20.591244,21.211998,22.04539,22.974806,21.966507,20.481497,19.325726,18.667244,19.486916,19.576086,19.438902,19.281141,18.986197,17.405157,15.902997,14.417986,13.077017,12.202472,11.945253,11.924676,11.948683,11.766914,11.06042,10.069269,9.002667,8.261876,7.840037,7.3050213,6.3378778,5.1992545,4.0674906,3.0797696,2.3218307,2.2429502,2.270387,2.352697,2.4315774,2.452155,3.0386145,3.841138,4.712253,5.4804807,5.9126086,6.560801,7.8126,9.80862,12.181894,14.071597,15.244516,15.614912,15.656067,15.608052,15.477728,14.932424,13.255356,10.943813,8.597976,6.917478,7.7748747,7.2638664,6.276145,5.528495,5.5730796,6.2898636,6.334448,5.7308407,5.1821065,6.060081,8.001227,9.8429165,10.014396,9.325048,10.971251,12.048141,11.286773,12.662037,15.196502,12.956982,11.406808,11.640019,11.835506,11.465111,11.279913,12.22648,14.688923,16.352274,16.650646,16.760393,14.781522,13.495427,13.824667,15.055889,14.808959,14.661487,14.2362175,13.423406,12.21962,10.7586155,10.9198065,12.120162,14.757515,18.334574,21.4555,22.714157,19.95677,16.530611,14.249936,13.423406,13.210771,12.919256,12.713481,12.7272,13.066729,12.6929035,12.641459,13.107883,14.009865,14.987297,14.490007,12.97413,12.068718,11.924676,11.204462,11.002116,11.633161,12.360233,13.104454,14.455711,16.060759,16.616352,16.516893,15.88242,14.579176,15.223939,17.384579,19.651537,21.644127,24.03112,22.059107,20.296299,18.427174,16.973028,17.302269,15.175924,12.634601,11.592006,11.869802,11.204462,10.823778,11.588576,12.449403,12.953552,13.207341,13.46799,13.128461,13.200482,13.903547,14.658057,14.802099,14.318527,12.672326,10.189304,8.045813,7.8777623,7.5862474,6.6568294,5.4084597,4.976331,3.8308492,2.5447538,1.5021594,0.90541106,0.7510797,0.64819205,0.5761707,0.5555932,0.58302987,0.6241849,0.6241849,0.5590228,0.5521636,0.64476246,0.8162418,0.8676856,0.83338976,0.7442205,0.64476246,0.5693115,0.77165717,0.7888051,0.66876954,0.53501564,0.5590228,0.5007198,0.42869842,0.3566771,0.3018037,0.26407823,0.2503599,0.23321195,0.2194936,0.20920484,0.17833854,0.16804978,0.17490897,0.18519773,0.18862732,0.18862732,0.14061308,0.106317215,0.07888051,0.0548734,0.048014224,0.15090185,0.16119061,0.116605975,0.08573969,0.18176813,0.19891608,0.26750782,0.4115505,0.5727411,0.607037,0.61389613,0.6379033,0.5007198,0.24350071,0.09602845,0.11317638,0.25378948,0.37039545,0.39440256,0.31895164,0.12003556,0.07888051,0.09602845,0.1097468,0.09602845,0.06859175,0.037725464,0.010288762,0.0,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.01371835,0.020577524,0.072021335,0.07888051,0.037725464,0.01371835,0.006859175,0.0034295875,0.0034295875,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.006859175,0.01371835,0.017147938,0.020577524,0.044584636,0.06516216,0.07545093,0.08916927,0.09945804,0.10288762,0.11317638,0.12689474,0.12689474,0.09259886,0.061732575,0.030866288,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.020577524,0.030866288,0.041155048,0.041155048,0.041155048,0.041155048,0.041155048,0.0548734,0.058302987,0.07888051,0.09945804,0.116605975,0.12346515,0.12689474,0.12003556,0.116605975,0.116605975,0.116605975,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.05144381,0.106317215,0.17490897,0.26064864,0.22292319,0.15776102,0.10288762,0.08573969,0.12346515,0.13375391,0.09259886,0.08573969,0.12346515,0.1371835,0.07545093,0.06859175,0.082310095,0.09259886,0.09259886,0.06859175,0.07888051,0.116605975,0.17147937,0.24350071,0.23321195,0.23664154,0.26407823,0.28465575,0.26064864,0.22292319,0.21263443,0.26750782,0.3566771,0.3806842,0.37039545,0.31895164,0.4046913,0.6001778,0.6859175,0.5521636,0.53844523,0.50757897,0.4046913,0.26064864,0.15090185,0.12346515,0.12689474,0.1371835,0.1371835,0.15090185,0.14404267,0.14404267,0.14061308,0.09259886,0.0548734,0.037725464,0.030866288,0.030866288,0.030866288,0.030866288,0.041155048,0.06516216,0.08916927,0.07545093,0.07545093,0.06859175,0.06859175,0.082310095,0.106317215,0.12003556,0.12346515,0.13375391,0.16804978,0.22978236,0.24007112,0.2709374,0.30866286,0.34981793,0.4115505,0.40126175,0.34295875,0.31895164,0.34295875,0.36696586,0.39097297,0.42526886,0.44927597,0.4629943,0.48700142,0.51100856,0.5178677,0.5693115,0.6893471,0.8848336,0.6276145,0.45613512,0.3566771,0.32238123,0.33609957,0.432128,0.548734,0.67219913,0.77508676,0.823101,0.8471081,0.8711152,0.96371406,1.039165,0.8711152,0.4664239,0.34638834,0.34638834,0.37382504,0.39783216,0.3841138,0.33609957,0.29837412,0.31552204,0.4115505,0.45956472,0.6927767,1.1694894,2.2052248,4.3795834,5.552502,6.2555676,6.6293926,6.824879,7.0203657,7.226141,7.407909,7.2775846,6.800872,6.1629686,5.394741,4.9180284,4.8940215,5.363875,6.2555676,7.500508,8.416207,9.050681,9.417647,9.489669,9.465661,8.985519,7.953213,6.9037595,6.989499,7.0135064,6.992929,7.051232,7.208993,7.3530354,7.56224,7.8263187,8.165848,8.536243,8.803751,8.903209,8.752307,8.330468,7.6342616,6.684266,5.645101,4.746549,4.0057583,3.4776018,3.2203827,2.7813954,2.3218307,1.8828435,1.4472859,0.94656616,0.64133286,0.52815646,0.5418748,0.70649505,1.1592005,1.6736387,1.5364552,1.4198492,1.5913286,1.9068506,2.2978237,2.6990852,3.192946,3.8377085,4.6676683,6.036074,6.5059276,6.2864337,5.874883,6.0566516,6.351596,6.7631464,7.380472,8.004657,8.162418,8.820899,10.2236,9.692014,7.2535777,5.6313825,5.2164025,5.0003386,4.722542,4.280125,3.7553983,3.2889743,2.9082901,2.620205,2.452155,2.4247184,2.170929,1.7936742,1.313532,0.8848336,0.823101,0.7888051,0.7613684,0.6790583,0.61046654,0.7339317,0.9534253,1.2072148,1.1489118,0.85739684,0.8711152,1.4815818,1.5398848,1.4678634,1.4575747,1.4953002,1.5913286,1.5707511,1.5776103,1.7730967,2.335549,2.054323,1.8176813,1.7388009,1.7388009,1.5570327,1.4095604,1.3992717,1.9514352,2.8568463,3.2958336,3.309552,3.0283258,2.4795918,1.8142518,1.3272504,1.2895249,1.1626302,1.0906088,1.1523414,1.371835,1.8005334,2.1194851,2.386993,2.726522,3.309552,3.642222,3.8514268,3.9440255,4.1155047,4.7774153,5.446185,6.025785,5.98463,5.3673043,4.804852,4.3795834,4.273266,4.7191124,5.638242,6.636252,7.1369715,8.141841,9.321619,10.460241,11.4754,11.852654,12.30536,12.830087,13.502286,14.466,15.29596,16.016174,16.523752,16.87357,17.288551,17.641798,17.857862,17.652086,17.247395,17.394867,18.187103,18.862732,19.62753,20.652975,22.093403,24.730755,24.69303,23.321196,21.596113,20.155685,20.303158,20.560377,20.834743,20.53637,18.571217,17.069057,15.704081,14.013294,12.154458,10.909517,10.299051,10.1481495,10.22703,10.326488,10.254466,9.887501,9.47595,9.297611,9.417647,9.674867,8.453933,6.992929,5.4633327,4.0674906,3.0660512,2.5653315,2.2841053,2.2806756,2.4624438,2.609916,3.450165,4.7328305,5.73427,6.142391,6.0566516,6.228131,7.5450926,9.266746,10.971251,12.55915,13.985858,14.754086,15.127911,15.234227,15.076467,13.756075,11.550851,8.934075,6.5162163,5.051782,5.2815647,5.4153185,5.0106273,4.3521466,4.4241676,4.791134,5.377593,5.192395,4.461893,4.6093655,5.8543057,8.855195,11.255906,12.349944,13.107883,14.143619,13.022143,11.941824,12.079007,13.581166,12.617453,12.833516,13.766364,15.234227,17.333136,17.62808,15.45715,13.670336,13.978998,16.96617,17.185663,12.758065,9.949233,10.4533825,11.369082,12.576297,12.483699,12.55915,13.581166,15.656067,18.36544,18.86959,18.598652,18.62609,19.637817,18.941612,16.780972,13.601744,10.799771,10.72775,10.494537,10.299051,10.1652975,10.199594,10.590566,10.967821,10.861504,11.454823,13.046151,15.059319,17.305698,15.2033615,12.682614,11.609154,11.780633,12.524854,14.359683,16.695232,19.095943,21.256582,22.354052,24.494114,28.139765,31.548775,30.790836,31.26755,32.639385,31.418451,27.536158,24.336353,21.750444,20.069946,17.521763,14.143619,11.749766,12.140739,11.688034,11.2593355,11.166737,11.153018,10.189304,9.290752,8.330468,7.507367,7.3255987,9.692014,13.828096,20.296299,28.050596,34.422768,36.06897,33.435047,26.18147,16.96617,11.413667,10.045261,11.197603,11.262765,9.102125,6.025785,4.8322887,3.415869,2.1469216,1.3615463,1.371835,1.0563129,0.85739684,0.78537554,0.7956643,0.8093826,0.69963586,0.5796003,0.5178677,0.58302987,0.84024894,1.0117283,0.9877212,0.8676856,0.7305021,0.65505123,0.64476246,0.6036074,0.5555932,0.51100856,0.47328308,0.4355576,0.41840968,0.4046913,0.39783216,0.39783216,0.432128,0.4424168,0.42869842,0.40126175,0.34981793,0.29151493,0.25721905,0.25721905,0.274367,0.274367,0.22635277,0.17833854,0.13375391,0.09602845,0.061732575,0.037725464,0.030866288,0.041155048,0.072021335,0.12346515,0.25721905,0.4629943,0.64819205,0.6927767,0.47328308,0.26407823,0.13032432,0.06859175,0.058302987,0.044584636,0.044584636,0.06516216,0.08916927,0.1097468,0.12346515,0.15776102,0.09602845,0.106317215,0.22978236,0.34981793,0.2777966,0.15776102,0.0548734,0.0,0.0,0.0,0.017147938,0.061732575,0.08573969,0.0,0.0,0.23664154,0.274367,0.07545093,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.010288762,0.006859175,0.030866288,0.041155048,0.044584636,0.05144381,0.06516216,0.07545093,0.07545093,0.08573969,0.08573969,0.06859175,0.030866288,0.0548734,0.05144381,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.017147938,0.030866288,0.0548734,0.06859175,0.07545093,0.07545093,0.07545093,0.08916927,0.09259886,0.09259886,0.09259886,0.09259886,0.01371835,0.01371835,0.01371835,0.010288762,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.017147938,0.0274367,0.037725464,0.048014224,0.07888051,0.13375391,0.20920484,0.13375391,0.08916927,0.06859175,0.06516216,0.061732575,0.12346515,0.1371835,0.11317638,0.09259886,0.11317638,0.09945804,0.09945804,0.10288762,0.09945804,0.07888051,0.07545093,0.07545093,0.11317638,0.17490897,0.2194936,0.18862732,0.21263443,0.23664154,0.22978236,0.18519773,0.22635277,0.36353627,0.5555932,0.65848076,0.42869842,0.31895164,0.26064864,0.29494452,0.40126175,0.5144381,0.8025235,1.1694894,1.1729189,0.8265306,0.61389613,0.4938606,0.3018037,0.18176813,0.17147937,0.20920484,0.29151493,0.25721905,0.20920484,0.19548649,0.21263443,0.12689474,0.082310095,0.058302987,0.041155048,0.041155048,0.05144381,0.07888051,0.10288762,0.11317638,0.09945804,0.13032432,0.16462019,0.19548649,0.216064,0.24007112,0.18519773,0.1920569,0.22978236,0.274367,0.32581082,0.29151493,0.2777966,0.29151493,0.33266997,0.42526886,0.42183927,0.41840968,0.44584638,0.5041494,0.53844523,0.53158605,0.48357183,0.45613512,0.48357183,0.58645946,0.72707254,0.72707254,0.6962063,0.6927767,0.70306545,0.5624523,0.4389872,0.34638834,0.28808534,0.26407823,0.42869842,0.5761707,0.70649505,0.864256,1.1180456,1.2963841,1.3889829,1.3855534,1.2895249,1.138623,0.86082643,0.607037,0.5007198,0.52472687,0.5178677,0.44927597,0.5178677,0.59674823,0.6276145,0.6207553,0.5693115,0.764798,1.1660597,1.845118,2.9631636,4.0880685,4.8905916,5.188966,5.2438393,5.761707,6.1561093,6.3824625,6.5642304,6.6465406,6.385892,5.857735,5.744559,5.7891436,5.9914894,6.5985265,8.292743,9.040393,9.314759,9.39707,9.3936405,9.242738,8.916927,8.433355,7.9737906,7.891481,7.466212,7.0546613,7.058091,7.455923,7.805741,8.158989,8.519095,8.707723,8.793462,9.071259,9.609704,9.438225,8.635701,7.3358874,5.720552,4.887162,4.15323,3.4810312,2.819121,2.1332035,1.6530612,1.2620882,0.939707,0.6927767,0.5418748,0.41498008,0.32924038,0.40126175,0.64819205,1.0117283,1.4095604,1.5947582,1.7936742,2.1332035,2.6167753,3.3884325,3.9268777,4.40702,4.931747,5.535354,6.1904054,6.5539417,6.725421,6.8866115,7.301592,7.654839,8.131552,8.923786,9.544542,8.834618,7.9600725,7.4696417,6.64997,5.4804807,4.629943,4.1943855,3.806842,3.426158,3.0420442,2.6922262,2.551613,2.386993,2.1846473,1.8999915,1.4850113,1.2689474,1.0631721,0.8265306,0.6001778,0.53158605,0.5418748,0.6173257,0.823101,1.08032,1.1351935,1.0734608,1.1694894,1.2655178,1.313532,1.3958421,1.5158776,1.786815,2.0131679,2.1023371,2.020027,1.7971039,1.5913286,1.4472859,1.4232788,1.6153357,1.6153357,1.6359133,1.6942163,1.6976458,1.4472859,1.2723769,1.2758065,1.6633499,2.2326615,2.369845,1.9994495,1.8073926,1.7559488,1.821111,1.9857311,2.020027,2.486451,3.1346428,3.673088,3.765687,3.4707425,3.3198407,3.3952916,3.6765177,4.0674906,4.201245,4.180667,4.2252517,4.4584637,4.9214582,5.4084597,5.7822843,5.830299,5.6073756,5.4153185,5.3913116,5.5730796,5.8680243,6.1766872,6.4064693,6.526505,7.082098,7.98065,9.174147,10.645439,11.05356,11.249047,11.4754,11.982979,13.025573,14.21564,15.333686,16.235666,16.877,17.312557,17.37429,17.333136,17.254255,17.161655,17.051908,16.732958,17.312557,18.451181,20.02193,22.10712,25.896814,26.822803,24.823355,21.386908,19.54522,19.233126,19.79901,20.388897,20.306587,19.03421,17.580065,16.362562,14.925565,13.282792,11.910957,11.046701,10.861504,10.882081,10.861504,10.779194,10.38479,9.846346,9.352485,9.088407,9.246168,8.601405,7.7577267,6.9620624,6.2247014,5.312431,4.479041,3.707384,3.2546785,3.2375305,3.6113555,4.705394,5.4084597,5.6965446,5.8200097,6.2898636,8.31675,9.962952,11.087856,11.63659,11.64345,13.88983,15.354263,15.649208,14.990726,14.198492,12.713481,10.772334,8.519095,6.217842,4.245829,3.1277838,2.8122618,2.503599,2.085189,2.1297739,2.9082901,4.173808,4.8014226,4.4927597,3.789694,4.448175,6.742569,9.527394,12.010415,13.7526455,14.870691,15.313108,14.88098,13.612033,11.773774,11.101575,12.264205,14.592895,17.765263,21.78817,25.44068,22.04539,18.413456,17.079346,16.321407,16.239098,13.231348,10.333347,9.331907,10.792912,10.676306,10.30934,10.172156,10.7586155,12.579727,16.558048,19.95677,20.70099,19.095943,17.844143,16.307688,14.627191,12.30536,9.801761,8.519095,8.635701,8.553391,8.724871,9.379922,10.504827,11.05699,11.369082,11.96926,13.077017,14.586036,16.245956,16.029892,15.440002,15.357693,16.077906,16.098484,15.172495,15.306249,17.336565,20.96164,24.843931,24.85422,25.711617,28.801676,32.18325,36.555973,41.97129,45.373444,44.38572,37.31391,29.443008,23.36578,18.512913,14.496866,11.077567,9.602845,8.049242,7.085528,6.9689217,7.5416627,8.450503,9.054111,8.80718,8.080108,8.128122,10.096705,12.761495,17.010754,22.60441,28.17406,32.66339,32.546783,28.794817,22.583834,15.282242,14.599753,15.841265,17.014183,16.359133,12.325937,9.030104,6.999788,6.2555676,6.3138704,6.217842,5.658819,5.5079174,5.4770513,5.3913116,5.178677,5.079219,5.020916,4.870014,4.6916757,4.7328305,3.525616,2.3492675,1.3855534,0.805953,0.7407909,0.65162164,0.59331864,0.5693115,0.5590228,0.5212973,0.5624523,0.8779744,1.0425946,0.9328478,0.72707254,0.6173257,0.5658819,0.59331864,0.6790583,0.77851635,0.5007198,0.3566771,0.3018037,0.3018037,0.31209245,0.33952916,0.33952916,0.274367,0.16462019,0.1097468,0.09602845,0.08573969,0.09602845,0.12346515,0.13375391,0.18176813,0.24007112,0.2503599,0.19891608,0.15433143,0.15433143,0.106317215,0.06516216,0.044584636,0.034295876,0.034295876,0.037725464,0.037725464,0.037725464,0.061732575,0.06859175,0.034295876,0.020577524,0.044584636,0.06859175,0.09602845,0.08916927,0.048014224,0.0,0.0,0.0,0.0034295875,0.017147938,0.05144381,0.12346515,0.44584638,0.5521636,0.40126175,0.14404267,0.11317638,0.082310095,0.030866288,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.017147938,0.030866288,0.041155048,0.048014224,0.05144381,0.06516216,0.07545093,0.072021335,0.06516216,0.0548734,0.017147938,0.024007112,0.030866288,0.030866288,0.020577524,0.01371835,0.01371835,0.0034295875,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.020577524,0.034295876,0.041155048,0.041155048,0.041155048,0.05144381,0.061732575,0.061732575,0.058302987,0.06859175,0.01371835,0.030866288,0.024007112,0.010288762,0.0,0.006859175,0.01371835,0.020577524,0.020577524,0.020577524,0.041155048,0.044584636,0.034295876,0.037725464,0.058302987,0.08916927,0.061732575,0.058302987,0.061732575,0.06516216,0.072021335,0.116605975,0.12689474,0.11317638,0.09602845,0.09602845,0.09602845,0.08573969,0.07888051,0.07888051,0.07545093,0.082310095,0.09259886,0.12346515,0.18519773,0.2503599,0.24350071,0.26064864,0.31895164,0.38754338,0.39783216,0.39783216,0.33952916,0.39783216,0.53844523,0.5144381,0.3806842,0.33609957,0.36010668,0.44584638,0.6207553,1.0460242,1.3615463,1.3272504,1.097468,1.1866373,0.881404,0.42869842,0.17833854,0.18862732,0.22978236,0.32581082,0.40126175,0.432128,0.4081209,0.33609957,0.15090185,0.10288762,0.09945804,0.09259886,0.09259886,0.06859175,0.06516216,0.07888051,0.09259886,0.08916927,0.16119061,0.22635277,0.24007112,0.21263443,0.22978236,0.23664154,0.2709374,0.31209245,0.3566771,0.39783216,0.39783216,0.3806842,0.36696586,0.37039545,0.3806842,0.3806842,0.44584638,0.5453044,0.64133286,0.66191036,0.6207553,0.5796003,0.607037,0.70649505,0.8196714,0.881404,0.823101,0.7579388,0.7133542,0.64819205,0.5658819,0.5453044,0.548734,0.5590228,0.5727411,0.72707254,0.9534253,1.1934965,1.4335675,1.704505,1.937717,1.9891608,1.821111,1.5090185,1.2517995,0.96371406,0.70649505,0.6379033,0.72021335,0.72364295,0.65848076,0.70306545,0.78194594,0.85739684,0.90884066,0.88826317,1.1660597,1.587899,2.0646117,2.5824795,2.983741,3.3678548,3.6559403,3.9851806,4.722542,5.192395,5.5593615,6.0223556,6.468202,6.4579134,6.125243,5.809721,5.5730796,5.562791,6.0052075,7.4456344,8.745448,9.702303,10.230459,10.340206,9.825768,9.431366,9.119273,8.855195,8.639131,7.5519514,6.790583,6.9826403,7.9463544,8.680285,9.112414,9.304471,9.105555,8.683716,8.519095,8.659708,8.217292,7.0306544,5.223262,3.199805,2.585909,2.2738166,2.061182,1.7799559,1.2929544,0.9945804,0.7956643,0.6962063,0.6310441,0.48700142,0.36696586,0.31209245,0.5212973,0.9774324,1.4815818,1.9274281,2.1126258,2.386993,2.8980014,3.5976372,4.633373,5.363875,6.0154963,6.725421,7.548522,7.414768,7.442205,7.6171136,7.8674736,8.080108,8.086967,8.035523,7.9943686,7.8126,7.1266828,6.40304,5.90232,5.377593,4.7774153,4.2526884,3.8102717,3.2821152,2.8054025,2.4315774,2.1434922,1.728512,1.5913286,1.5947582,1.5844694,1.3786942,1.0700313,0.8162418,0.66191036,0.6173257,0.6790583,0.75450927,0.8265306,0.8745448,0.88826317,0.86082643,0.864256,0.9568549,1.1283343,1.3546871,1.5913286,1.7593783,2.0234566,2.2052248,2.1915064,1.903421,1.8039631,1.6599203,1.4575747,1.2586586,1.1866373,1.1592005,1.1832076,1.4164196,1.6976458,1.546744,1.2998136,1.3581166,1.5707511,1.7559488,1.7147937,1.3478279,1.4644338,1.7525192,2.020027,2.1983654,2.767677,3.3301294,3.8617156,4.383013,4.98662,4.7602673,4.479041,4.307562,4.314421,4.4859004,4.5510626,4.4584637,4.5510626,4.9008803,5.3158607,5.7274113,6.0669403,6.2898636,6.420188,6.557371,6.725421,6.835168,6.8557453,6.7459984,6.468202,6.3961806,6.708273,7.459353,8.615124,10.024684,10.587136,10.738038,10.882081,11.334786,12.315649,13.745787,15.038741,15.985307,16.53747,16.815268,16.955881,17.165085,17.29198,17.093063,16.235666,15.87213,16.21166,17.137648,18.893597,22.089973,25.553856,26.894825,24.4461,19.651537,17.058767,16.427725,17.532051,18.684393,19.054789,18.684393,17.741257,16.955881,16.023033,14.850114,13.560589,12.298501,11.7257595,11.537132,11.502836,11.46854,11.379372,10.995257,10.14129,9.218731,9.211872,9.1810055,9.105555,9.0369625,8.803751,8.018375,6.8214493,6.245279,5.7411294,5.147811,4.7019644,5.627953,5.778855,5.435896,5.15467,5.7719955,8.680285,10.899229,12.195613,13.011855,14.452282,17.20624,19.233126,19.744135,18.694681,16.798119,14.092175,11.588576,9.287323,7.1678376,5.1683884,3.0489032,2.2052248,1.8039631,1.471293,1.2826657,1.9274281,2.7402403,3.2443898,3.2409601,2.8088322,3.649081,5.7754254,8.940934,12.315649,14.466,15.357693,15.388559,14.723219,13.317088,10.926665,9.678296,10.618003,12.47341,14.939283,18.674105,24.19231,24.377508,22.350622,20.526081,20.61868,19.346302,16.050468,12.188754,9.386781,9.441654,8.999237,8.81404,9.218731,10.093276,10.88551,12.034423,15.683503,18.509483,19.500635,19.967058,18.156237,16.19794,13.924125,11.495977,9.403929,8.920357,8.515666,8.457363,8.98209,10.281903,11.465111,12.63803,13.512574,14.116182,14.778092,15.885849,17.326277,18.718689,19.833303,20.584383,19.473198,18.04306,17.161655,17.189093,17.988186,19.548649,20.090523,21.959648,25.471546,28.914852,32.91375,34.41248,33.129814,29.75167,25.920822,21.098822,16.94902,13.80066,11.585147,9.829198,9.132992,7.5382333,6.001778,5.1855364,5.429037,6.8969,7.970361,8.405919,8.364764,8.433355,10.086417,12.034423,14.105893,16.019604,17.384579,19.017063,19.764713,20.028791,19.716698,18.255693,19.164536,20.875898,21.939072,21.177702,17.682953,11.766914,8.886061,7.970361,7.966932,7.81603,6.7391396,6.1321025,6.0875177,6.3721733,6.427047,6.1321025,5.5902276,4.996909,4.48933,4.1429415,3.175798,2.0406046,1.2106444,0.83681935,0.75450927,0.6379033,0.5658819,0.52815646,0.5178677,0.52472687,0.5555932,0.7990939,1.0082988,1.0254467,0.7990939,0.6962063,0.6207553,0.59331864,0.607037,0.6379033,0.490431,0.39783216,0.34638834,0.33266997,0.32924038,0.34981793,0.36010668,0.32238123,0.2503599,0.19548649,0.16804978,0.14061308,0.13032432,0.13375391,0.12003556,0.106317215,0.09945804,0.07545093,0.044584636,0.058302987,0.12003556,0.12346515,0.09602845,0.06859175,0.048014224,0.06516216,0.05144381,0.0274367,0.01371835,0.037725464,0.06516216,0.058302987,0.037725464,0.0274367,0.0274367,0.048014224,0.037725464,0.017147938,0.0034295875,0.010288762,0.017147938,0.017147938,0.020577524,0.034295876,0.07888051,0.2777966,0.36010668,0.274367,0.10288762,0.0548734,0.041155048,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.041155048,0.072021335,0.09945804,0.10288762,0.082310095,0.044584636,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.020577524,0.037725464,0.05144381,0.06516216,0.061732575,0.072021335,0.06859175,0.061732575,0.058302987,0.05144381,0.037725464,0.037725464,0.034295876,0.0274367,0.01371835,0.024007112,0.020577524,0.017147938,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.006859175,0.006859175,0.006859175,0.010288762,0.01371835,0.01371835,0.010288762,0.01371835,0.020577524,0.020577524,0.020577524,0.020577524,0.034295876,0.041155048,0.041155048,0.037725464,0.041155048,0.01371835,0.030866288,0.020577524,0.006859175,0.0,0.006859175,0.01371835,0.020577524,0.020577524,0.017147938,0.0274367,0.030866288,0.024007112,0.01371835,0.017147938,0.020577524,0.037725464,0.06516216,0.08573969,0.106317215,0.15776102,0.17833854,0.14061308,0.116605975,0.116605975,0.1097468,0.106317215,0.082310095,0.06859175,0.07545093,0.082310095,0.08916927,0.106317215,0.14061308,0.1920569,0.25721905,0.3018037,0.32924038,0.36696586,0.44584638,0.58645946,0.58302987,0.4081209,0.4046913,0.59674823,0.66876954,0.5178677,0.61389613,0.7133542,0.72707254,0.70649505,0.805953,1.1763484,1.3924125,1.3581166,1.3169615,0.9911508,0.5658819,0.31209245,0.28465575,0.3018037,0.36696586,0.4629943,0.5007198,0.44927597,0.34638834,0.18519773,0.15776102,0.17147937,0.18176813,0.18176813,0.09945804,0.06516216,0.061732575,0.06516216,0.05144381,0.16462019,0.2469303,0.26407823,0.23664154,0.2469303,0.29494452,0.34295875,0.37725464,0.4046913,0.44584638,0.48700142,0.48014224,0.4629943,0.44584638,0.4115505,0.40126175,0.490431,0.607037,0.6962063,0.7305021,0.7133542,0.72364295,0.8025235,0.91227025,0.9431366,0.9259886,0.823101,0.7407909,0.72021335,0.7339317,0.7990939,0.9431366,1.1008976,1.2209331,1.2620882,1.2655178,1.5227368,1.8313997,2.1023371,2.3492675,2.760818,2.8156912,2.5550427,2.1023371,1.6907866,1.3306799,1.0288762,0.8471081,0.7956643,0.8265306,0.7990939,0.75450927,0.7956643,0.9362774,1.1111864,1.2586586,1.5638919,1.8519772,2.0474637,2.1469216,2.2258022,2.3767042,2.6613598,3.1620796,3.99204,4.588788,5.137522,5.751418,6.324159,6.543653,6.358455,5.8543057,5.48734,5.4770513,5.809721,6.6225333,7.486789,8.272165,8.865483,9.191295,9.153569,9.270175,9.445084,9.568549,9.506817,8.107545,7.226141,7.4010496,8.405919,9.270175,9.321619,8.779744,7.829748,6.8111606,6.210983,5.960623,5.3741636,4.3109913,2.8637056,1.3684053,0.97400284,0.9362774,1.0117283,1.0151579,0.8162418,0.65162164,0.6173257,0.71678376,0.7888051,0.53158605,0.432128,0.490431,0.8779744,1.5158776,2.07833,2.5241764,2.750529,3.0660512,3.590778,4.2869844,5.2506986,5.9434752,6.6636887,7.5931067,8.803751,8.7317295,8.827758,9.012956,8.985519,8.213862,7.613684,7.0615206,6.5162163,6.012067,5.6656785,5.377593,5.099797,4.6848164,4.1292233,3.57363,3.0523329,2.4967396,2.0268862,1.6770682,1.4164196,1.1146159,0.9774324,0.9328478,0.94656616,1.0254467,0.90198153,0.77851635,0.6824879,0.66191036,0.7682276,0.805953,0.7305021,0.61389613,0.5453044,0.59674823,0.78537554,0.90541106,1.097468,1.3958421,1.7559488,2.0165975,2.201795,2.2463799,2.0646117,1.5433143,1.5330256,1.471293,1.3101025,1.0768905,0.90198153,0.8505377,0.9362774,1.2243627,1.5364552,1.4369972,1.1249046,1.1934965,1.3649758,1.5090185,1.6427724,1.8005334,2.194936,2.5790498,2.8259802,2.9220085,3.4810312,3.806842,4.016047,4.32128,5.0174866,5.1066556,5.07236,4.856296,4.588788,4.57164,4.633373,4.5442033,4.695105,5.1580997,5.693115,6.169828,6.5985265,6.9826403,7.3221693,7.6205435,7.9257765,8.014946,7.888051,7.507367,6.783724,6.475061,6.5127864,7.016936,7.888051,8.803751,9.3079,9.5205345,9.822338,10.432805,11.413667,12.867812,14.723219,16.095055,16.46545,15.680074,16.12935,16.602633,16.842705,16.61292,15.697222,15.426285,15.536031,16.47231,18.557497,22.007662,24.789059,25.831654,23.547548,19.003344,15.923574,14.832966,16.225378,17.984756,19.085653,19.579515,18.722118,17.96761,17.171944,16.177364,14.832966,13.454271,12.566009,12.027563,11.705182,11.482259,11.372512,10.991828,10.14129,9.225591,9.256456,9.908078,10.497967,10.827208,10.710602,9.9698105,8.923786,8.522525,8.097256,7.3873315,6.526505,6.852316,6.6122446,5.9331865,5.4633327,6.351596,8.628842,10.189304,11.235329,12.511135,15.306249,19.078794,21.873909,22.796469,21.626978,18.849012,15.512024,12.795791,10.521975,8.488229,6.4819202,4.0606318,2.6819375,1.961724,1.5673214,1.2209331,1.5090185,1.8416885,2.16064,2.469303,2.8088322,4.0194764,6.060081,9.301042,13.179905,16.187653,16.386568,15.512024,14.071597,12.181894,9.547972,8.344186,8.512236,9.211872,10.5597,13.625751,19.157675,23.002243,23.979675,23.328054,24.682741,24.09971,21.345753,17.086205,12.586586,9.716022,8.652849,7.9292064,8.080108,9.1981535,10.923236,9.705732,11.279913,13.965281,16.753534,19.315437,18.914175,18.005335,16.510035,14.531162,12.363663,10.875222,9.80862,9.273604,9.345626,10.072699,11.297061,12.339656,12.830087,12.792361,12.6586075,14.349394,16.928444,19.558937,21.486366,22.011093,20.673553,19.421753,18.485476,17.971039,17.902447,18.430603,19.908754,23.043398,26.798796,28.403843,26.02714,24.130577,21.719578,19.089085,17.844143,13.087306,10.233889,9.067829,8.889491,8.536243,8.347616,7.191845,5.960623,5.1992545,5.1100855,6.1286726,7.291303,8.378482,9.160428,9.39707,10.343636,11.756626,12.538571,12.164746,10.686595,9.829198,10.405369,12.157887,14.582606,16.914726,18.591793,20.45406,21.85333,22.161995,20.76958,16.239098,13.406258,11.89038,11.032983,9.884071,8.083538,6.8385973,6.2830043,6.217842,6.1149545,5.394741,4.3281393,3.3472774,2.6716487,2.3218307,1.978872,1.4404267,1.0666018,0.91912943,0.77165717,0.6173257,0.53158605,0.48014224,0.4664239,0.53158605,0.61046654,0.6962063,0.84367853,0.96714365,0.83681935,0.72021335,0.6276145,0.5624523,0.5144381,0.490431,0.4629943,0.42183927,0.3806842,0.34638834,0.32238123,0.33266997,0.34638834,0.33952916,0.31209245,0.26750782,0.23664154,0.19548649,0.15776102,0.13032432,0.09602845,0.07888051,0.061732575,0.048014224,0.041155048,0.06859175,0.12346515,0.1371835,0.12346515,0.09602845,0.061732575,0.061732575,0.05144381,0.030866288,0.01371835,0.017147938,0.048014224,0.048014224,0.037725464,0.0274367,0.0274367,0.0274367,0.010288762,0.0,0.0034295875,0.010288762,0.017147938,0.017147938,0.017147938,0.017147938,0.017147938,0.0548734,0.1097468,0.10288762,0.041155048,0.006859175,0.0,0.010288762,0.020577524,0.0274367,0.037725464,0.06516216,0.044584636,0.024007112,0.034295876,0.07888051,0.1097468,0.14061308,0.15776102,0.15090185,0.09945804,0.048014224,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.024007112,0.044584636,0.06516216,0.061732575,0.072021335,0.072021335,0.06516216,0.061732575,0.06859175,0.05144381,0.044584636,0.044584636,0.041155048,0.0274367,0.024007112,0.024007112,0.020577524,0.01371835,0.01371835,0.010288762,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.01371835,0.01371835,0.01371835,0.010288762,0.020577524,0.024007112,0.024007112,0.024007112,0.024007112,0.01371835,0.017147938,0.010288762,0.0034295875,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.024007112,0.024007112,0.020577524,0.020577524,0.030866288,0.05144381,0.07888051,0.10288762,0.14061308,0.23321195,0.23664154,0.17490897,0.14404267,0.16462019,0.15776102,0.14061308,0.10288762,0.082310095,0.08573969,0.08573969,0.08916927,0.12689474,0.16462019,0.1920569,0.22292319,0.32581082,0.4115505,0.42526886,0.4355576,0.6344737,0.65505123,0.5453044,0.6036074,0.8196714,0.8505377,0.7510797,1.0117283,1.2483698,1.2175035,0.7956643,0.34981793,0.9568549,1.5124481,1.4918705,0.97400284,0.9294182,0.764798,0.58302987,0.47328308,0.490431,0.5144381,0.5144381,0.44584638,0.34638834,0.33266997,0.3018037,0.2777966,0.2709374,0.26750782,0.26064864,0.15090185,0.09945804,0.07545093,0.058302987,0.041155048,0.19548649,0.274367,0.30866286,0.31895164,0.32238123,0.34981793,0.38754338,0.4046913,0.41840968,0.4629943,0.5041494,0.51100856,0.51100856,0.50757897,0.5007198,0.490431,0.5761707,0.66191036,0.71678376,0.7922347,0.91227025,1.0151579,1.1008976,1.1249046,0.99801,0.9294182,0.8128122,0.7476501,0.8093826,1.039165,1.4267083,1.8416885,2.1332035,2.2566686,2.2841053,2.1400626,2.3252604,2.551613,2.7299516,2.9734523,3.649081,3.7313912,3.433017,2.942586,2.3904223,1.99602,1.6221949,1.2380811,0.922559,0.89855194,0.84024894,0.70306545,0.70649505,0.89512235,1.1489118,1.4987297,1.8005334,1.8725548,1.7216529,1.5364552,1.8485477,2.0474637,2.301253,2.7711067,3.642222,4.341858,4.996909,5.6073756,6.1561093,6.6225333,6.509357,6.029215,5.7582774,5.874883,6.135532,6.3653145,6.090947,6.0223556,6.39961,6.9792104,7.675417,8.423067,9.153569,9.774324,10.179015,9.153569,8.39563,8.1041155,8.241299,8.512236,7.997798,6.8591747,5.3878818,3.9886103,3.1792276,2.7951138,2.2909644,1.7525192,1.2483698,0.8265306,0.64476246,0.66191036,0.72021335,0.72021335,0.6207553,0.48700142,0.51100856,0.6756287,0.8093826,0.5727411,0.59331864,0.7956643,1.2929544,1.9582944,2.4212887,2.7916842,3.1860867,3.6353626,4.1463714,4.695105,5.271276,5.73427,6.351596,7.2947326,8.628842,9.294182,9.801761,10.069269,9.688584,7.936065,6.8591747,6.125243,5.6965446,5.470192,5.267846,4.962613,4.4687524,3.82399,3.100347,2.4075704,1.8279701,1.3924125,1.0425946,0.7579388,0.53844523,0.7579388,0.6859175,0.42183927,0.20234565,0.39097297,0.607037,0.7407909,0.69963586,0.5761707,0.607037,0.5453044,0.31552204,0.25378948,0.4389872,0.70649505,0.9602845,1.0528834,1.1729189,1.3924125,1.6736387,1.879414,1.978872,1.9239986,1.6667795,1.1214751,1.0220171,0.94656616,0.85396725,0.7442205,0.64476246,0.70649505,0.91227025,1.1111864,1.2072148,1.1797781,1.0734608,1.2277923,1.4987297,1.8073926,2.1469216,2.8945718,3.4055803,3.7622573,3.981751,4.0194764,4.0709205,4.1429415,4.187526,4.266407,4.5784993,4.962613,5.40503,5.3981705,4.9831905,4.7671266,4.7431192,4.6848164,4.8734436,5.3878818,6.077229,6.591667,7.0306544,7.390761,7.699424,7.9943686,8.385342,8.577398,8.433355,7.888051,6.931196,6.39961,6.159539,6.307011,6.708273,7.006647,7.233,7.5862474,8.182996,9.033533,10.041832,11.348505,13.622321,15.409137,15.755525,14.205351,14.928994,15.450292,15.745236,15.762384,15.450292,15.062748,15.062748,16.21166,18.512913,21.208569,23.746464,24.000254,22.220297,19.174824,16.167076,15.0250225,16.304258,18.30028,20.018501,21.167414,20.03222,18.828436,17.686382,16.520323,15.042171,13.845244,12.833516,11.979549,11.273054,10.731179,10.22703,9.530824,8.865483,8.477941,8.663138,9.945804,10.995257,11.530273,11.454823,10.844356,10.285333,9.781183,9.448513,9.132992,8.412778,7.9189177,7.56567,6.944915,6.464772,7.349606,8.014946,8.203573,8.7317295,10.2236,13.094165,18.03277,21.602972,23.125708,22.36434,19.493774,16.780972,14.572317,12.30536,9.829198,7.4044795,5.0757895,3.333559,2.270387,1.7456601,1.3958421,1.371835,1.6393428,2.0268862,2.5413244,3.3541365,4.6265135,6.495639,9.510246,13.505715,17.597214,17.278261,15.971589,13.776653,11.029553,8.31675,7.888051,7.1232533,6.8969,7.8434668,10.357354,14.483148,19.353163,22.803328,24.497543,25.94826,26.68562,25.18689,21.644127,16.825556,12.065289,9.911508,7.881192,6.8969,7.81603,11.417097,10.340206,9.246168,9.510246,11.393089,14.05102,15.3302555,16.63007,17.21653,16.96274,16.352274,14.2533655,12.545431,11.38623,10.796341,10.63858,11.094715,11.019264,10.48082,9.757176,9.338767,11.897239,14.500296,17.302269,19.716698,20.402617,19.53836,18.602083,18.217968,18.718689,20.138538,21.702429,23.478956,26.713057,30.036327,29.460155,19.991066,17.357141,18.37916,19.723558,17.905876,10.106995,6.9071894,6.574519,7.301592,7.2158523,6.948344,6.3001523,5.90575,5.90575,5.9469047,6.420188,7.73029,9.373062,10.6488695,10.652299,10.731179,11.653738,12.140739,11.688034,10.542552,9.825768,9.541112,9.853205,10.72089,11.910957,12.79922,14.044161,16.019604,18.307138,19.70641,20.080235,18.962189,17.648657,16.21509,13.519434,11.149589,9.366203,7.829748,6.478491,5.5319247,4.2869844,2.9665933,1.8828435,1.255229,1.196926,1.2175035,1.2860953,1.2826657,1.1489118,0.8779744,0.6962063,0.58302987,0.4972902,0.4629943,0.5658819,0.7407909,0.77508676,0.84024894,0.9328478,0.8711152,0.6790583,0.58988905,0.5453044,0.5212973,0.52472687,0.4972902,0.45956472,0.4046913,0.34638834,0.30523327,0.31895164,0.32924038,0.33609957,0.33266997,0.29494452,0.274367,0.21263443,0.15433143,0.1097468,0.07888051,0.10288762,0.1097468,0.09945804,0.07888051,0.09602845,0.11317638,0.116605975,0.11317638,0.09259886,0.05144381,0.020577524,0.0274367,0.030866288,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.048014224,0.07545093,0.08573969,0.07545093,0.041155048,0.024007112,0.030866288,0.058302987,0.082310095,0.041155048,0.030866288,0.061732575,0.08573969,0.09259886,0.11317638,0.16804978,0.106317215,0.05144381,0.06516216,0.12346515,0.14061308,0.15776102,0.16119061,0.13032432,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.034295876,0.058302987,0.06859175,0.07545093,0.07545093,0.06859175,0.061732575,0.061732575,0.0548734,0.05144381,0.0548734,0.058302987,0.044584636,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.0034295875,0.006859175,0.01371835,0.010288762,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.010288762,0.0,0.010288762,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.0274367,0.020577524,0.010288762,0.0,0.0,0.01371835,0.006859175,0.006859175,0.020577524,0.044584636,0.06859175,0.058302987,0.041155048,0.030866288,0.030866288,0.041155048,0.037725464,0.037725464,0.061732575,0.12346515,0.09602845,0.1371835,0.20920484,0.26750782,0.24350071,0.19548649,0.1371835,0.08916927,0.061732575,0.061732575,0.08573969,0.16462019,0.20920484,0.19891608,0.19891608,0.31895164,0.5418748,0.7133542,0.7442205,0.61046654,0.52472687,0.4664239,0.44927597,0.5590228,0.9602845,1.1454822,1.2895249,1.6324836,1.8828435,1.2346514,0.7099246,1.3203912,1.5776103,1.1317638,0.77851635,1.2415106,1.0666018,0.77165717,0.66191036,0.8093826,0.881404,0.8265306,0.65162164,0.48014224,0.5658819,0.5521636,0.47671264,0.36010668,0.2469303,0.19891608,0.18519773,0.1371835,0.09602845,0.09259886,0.15090185,0.3841138,0.42526886,0.39440256,0.36010668,0.33609957,0.37382504,0.3806842,0.3806842,0.39097297,0.42869842,0.4389872,0.42526886,0.4355576,0.47671264,0.48700142,0.53844523,0.6962063,0.7990939,0.84367853,0.9774324,1.3786942,1.6256244,1.7113642,1.6187652,1.3272504,1.0837497,0.96714365,0.9842916,1.2003556,1.7250825,2.627064,3.5016088,3.782835,3.5530527,3.5393343,3.6147852,3.5942078,3.5050385,3.4467354,3.6319332,4.3761535,4.307562,3.8788633,3.340418,2.7299516,2.4761622,2.2086544,1.9342873,1.6290541,1.2517995,0.9568549,0.7579388,0.72021335,0.84367853,1.0528834,1.3821237,1.9137098,2.054323,1.7662375,1.5707511,1.9137098,1.9514352,2.136633,2.7162333,3.7519686,4.2183924,4.6916757,5.195825,5.778855,6.4990683,6.3310184,5.885172,5.6142344,5.669108,5.888602,6.121814,6.23499,6.924337,8.100685,8.89635,8.371623,8.1487,8.282454,8.81061,9.750318,9.908078,9.335337,8.128122,6.5333643,4.9591837,4.6916757,4.770556,4.2938433,3.2272418,2.411,1.8142518,1.4438564,1.1146159,0.77851635,0.53501564,0.5453044,0.64133286,0.6893471,0.6207553,0.4115505,0.38754338,0.36353627,0.3566771,0.42869842,0.67219913,0.8676856,1.0906088,1.430138,1.8588364,2.2120838,2.603057,3.1140654,3.8514268,4.722542,5.4153185,5.562791,5.9469047,6.447624,6.9963584,7.5690994,8.399059,8.889491,9.030104,8.738589,7.874333,7.140401,6.492209,6.0326443,5.6348124,4.914599,4.0709205,3.2375305,2.4761622,1.821111,1.2963841,0.9911508,0.7682276,0.58645946,0.41498008,0.24350071,0.4629943,0.51100856,0.41840968,0.32924038,0.48700142,0.548734,0.5453044,0.45613512,0.32581082,0.29151493,0.2777966,0.22978236,0.42526886,0.85396725,1.2209331,1.2209331,1.138623,1.0048691,0.82996017,0.61046654,0.72021335,0.72021335,0.6276145,0.53844523,0.61046654,0.45270553,0.22978236,0.11317638,0.16804978,0.34981793,0.5590228,0.65505123,0.7407909,0.9259886,1.3272504,2.1572106,2.7951138,3.1689389,3.223812,2.9288676,3.234101,3.6970954,4.2389703,4.5819287,4.2252517,4.386442,4.6916757,4.7808447,4.7499785,5.127233,5.785714,6.619104,6.893471,6.4990683,5.950334,5.4976287,5.5147767,5.7822843,6.1972647,6.759717,6.941485,6.9620624,6.8626046,6.8111606,7.0786686,7.3598948,7.5039372,7.2124224,6.5779486,6.0875177,5.720552,5.4736214,5.3844523,5.4187484,5.4941993,5.5559316,6.1629686,6.975781,7.798882,8.591117,9.750318,10.618003,11.269625,11.958971,13.107883,13.694343,14.085316,14.623761,15.097044,14.754086,14.280802,14.352823,15.066177,16.448301,18.4649,21.623549,21.208569,19.28457,17.010754,14.616901,15.2033615,16.13621,17.37772,18.811287,20.265432,19.517782,17.923023,16.335125,15.066177,13.869251,12.723769,11.622872,10.834066,10.350495,9.887501,9.1810055,7.949784,6.8557453,6.2830043,6.3310184,7.9086285,9.270175,10.412228,11.159878,11.183885,10.597425,9.911508,9.654288,9.523964,8.378482,7.267296,7.1987042,6.9792104,6.262427,5.5559316,5.223262,5.830299,7.1095347,8.934075,11.276484,16.002455,19.579515,21.980227,22.755312,21.057667,19.898466,18.471758,15.529172,11.345076,7.720001,4.914599,3.2135234,2.2429502,1.7010754,1.3581166,1.2860953,1.6873571,2.1469216,2.4144297,2.4247184,3.0248961,4.7774153,7.579388,11.163307,15.107333,15.913286,15.107333,12.915827,10.525404,10.086417,9.901219,8.182996,7.8777623,9.403929,10.652299,13.152468,15.728088,19.305147,23.067406,24.459818,21.884197,19.576086,17.54234,15.923574,14.983868,12.22648,9.191295,7.5450926,7.8263187,9.47595,10.539123,9.321619,8.076678,7.5931067,7.2021337,6.4716315,8.742019,12.30536,16.21852,20.29287,19.03764,17.339994,15.337115,13.639469,13.337666,12.836946,12.089295,10.837497,9.668007,10.010965,10.9369545,11.537132,13.591455,16.87357,19.11995,17.741257,17.70696,18.0362,18.173384,17.991615,17.806417,19.408035,22.295748,24.442669,22.292318,17.336565,12.3911,10.566559,10.837497,8.042382,5.1855364,4.928317,5.161529,5.1169443,5.3878818,6.728851,6.385892,5.7822843,5.717122,6.3618846,7.6925645,9.482809,11.458252,12.432255,10.285333,10.295622,11.077567,11.640019,12.006986,13.227919,13.742357,11.993267,10.151579,9.006097,7.98065,6.7494283,6.4304767,7.15069,8.999237,12.041282,15.323397,18.012194,19.939621,20.207129,17.182234,15.0456,13.063298,10.587136,7.7920227,5.693115,4.105216,2.901431,2.07833,1.587899,1.3443983,1.4404267,1.6770682,1.786815,1.6221949,1.1592005,1.0734608,0.90541106,0.69963586,0.5521636,0.6241849,0.77165717,0.94656616,1.0494537,1.0082988,0.7613684,0.5178677,0.47671264,0.5007198,0.52472687,0.548734,0.5624523,0.51100856,0.4355576,0.36696586,0.30523327,0.28122616,0.26407823,0.2777966,0.29494452,0.26064864,0.2469303,0.15090185,0.072021335,0.0548734,0.09259886,0.15090185,0.18519773,0.17490897,0.12346515,0.061732575,0.037725464,0.041155048,0.041155048,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.07545093,0.2469303,0.3806842,0.4355576,0.3841138,0.21263443,0.116605975,0.14747226,0.274367,0.3566771,0.1371835,0.1371835,0.20234565,0.2194936,0.18519773,0.19891608,0.18519773,0.09259886,0.017147938,0.0,0.0,0.0,0.12689474,0.2194936,0.18176813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.06516216,0.09602845,0.106317215,0.082310095,0.06859175,0.061732575,0.061732575,0.061732575,0.072021335,0.07545093,0.06859175,0.058302987,0.044584636,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.010288762,0.0034295875,0.0,0.0,0.0034295875,0.0,0.006859175,0.01371835,0.010288762,0.044584636,0.0548734,0.048014224,0.030866288,0.030866288,0.034295876,0.037725464,0.034295876,0.0274367,0.048014224,0.06516216,0.12689474,0.20234565,0.2469303,0.23321195,0.16462019,0.1371835,0.1371835,0.14404267,0.13375391,0.14747226,0.17490897,0.21263443,0.2503599,0.2709374,0.32581082,0.4355576,0.4938606,0.48014224,0.4629943,0.45613512,0.38754338,0.3841138,0.5453044,0.9362774,1.4815818,1.5124481,1.2826657,1.0906088,1.2723769,1.5193073,1.8382589,1.8348293,1.471293,1.0597426,0.94656616,0.91912943,0.864256,0.7922347,0.8196714,1.0220171,1.1866373,1.1934965,0.9877212,0.61389613,0.4629943,0.37725464,0.32924038,0.28465575,0.19891608,0.16804978,0.16462019,0.21263443,0.29151493,0.32238123,0.4081209,0.5727411,0.6790583,0.6790583,0.6173257,0.48700142,0.42526886,0.42869842,0.5041494,0.64819205,0.58988905,0.5453044,0.5212973,0.548734,0.65848076,0.65848076,0.65162164,0.70306545,0.8265306,1.0014396,1.2072148,1.2826657,1.3375391,1.430138,1.546744,1.6942163,1.9891608,2.428148,3.0111778,3.7519686,4.2938433,4.6745276,4.681387,4.417309,4.307562,4.1772375,4.057202,4.383013,5.0757895,5.5250654,5.7994323,5.861165,5.178677,3.8171308,2.4247184,2.7951138,2.620205,2.194936,1.6907866,1.1660597,0.9911508,0.89169276,0.85396725,0.939707,1.2860953,1.5055889,1.6530612,1.8862731,2.2258022,2.5481834,2.8980014,2.7951138,2.901431,3.4638834,4.314421,4.6436615,4.8254294,5.0586414,5.610805,6.8283086,7.490219,7.7131424,7.438775,6.7940125,6.0840883,5.9469047,6.368744,7.0306544,7.840037,8.944365,10.244178,10.786053,10.6317215,9.897789,8.738589,7.31531,6.1458206,5.1821065,4.4241676,3.9337368,3.9680326,3.8960114,3.2375305,2.177788,1.5433143,1.1523414,0.91227025,0.78537554,0.7407909,0.77851635,0.89855194,0.881404,0.78194594,0.6379033,0.44927597,0.5521636,0.8745448,1.3375391,1.7353712,1.7456601,1.9308578,2.1434922,2.2909644,2.6785078,4.0194764,5.07236,4.914599,4.9214582,5.535354,6.258997,6.8557453,7.2432885,7.548522,7.8366075,8.117833,8.858624,9.108984,8.937505,8.694004,9.009526,8.128122,6.783724,5.579939,4.65395,3.6799474,2.750529,1.9823016,1.3924125,0.94999576,0.6001778,0.39440256,0.30523327,0.2777966,0.2709374,0.25721905,0.41840968,0.50757897,0.52815646,0.5041494,0.48700142,0.42183927,0.34981793,0.31895164,0.32238123,0.31552204,0.28122616,0.22292319,0.38754338,0.78537554,1.1592005,1.1317638,1.0323058,0.922559,0.86082643,0.91569984,0.77165717,0.58988905,0.40126175,0.2503599,0.20920484,0.1371835,0.07545093,0.072021335,0.16804978,0.40126175,0.78194594,1.3272504,1.7971039,2.1332035,2.4384367,3.1209247,3.5393343,3.858286,4.2286816,4.7842746,5.284994,5.830299,6.4098988,6.835168,6.7528577,6.4716315,6.090947,5.7411294,5.446185,5.103226,4.7671266,4.996909,5.2815647,5.4153185,5.5113473,5.2438393,5.5250654,6.060081,6.56766,6.807731,6.756287,6.6431108,6.461343,6.3721733,6.691125,6.9689217,7.0923867,6.8728933,6.358455,5.830299,5.3090014,5.0586414,4.996909,5.0620713,5.223262,5.295283,5.6519604,6.186976,6.9037595,7.932636,9.256456,10.467101,11.369082,12.000127,12.63117,13.186764,13.824667,14.359683,14.678635,14.706071,14.514014,14.863832,15.316538,15.758954,16.386568,16.914726,16.606062,16.005884,15.388559,14.764374,15.12448,15.645778,16.077906,16.2974,16.2974,15.971589,15.63206,15.29253,14.956431,14.589465,13.989287,13.330807,12.607163,11.753197,10.645439,9.6645775,8.628842,7.6514096,6.9346256,6.759717,7.6205435,8.652849,9.239308,9.410788,9.853205,10.4705305,10.755186,10.707172,10.254466,9.294182,7.750868,7.48336,7.6445503,7.630832,7.0786686,6.427047,6.40304,7.1849856,9.088407,12.545431,17.144508,21.424633,23.427511,23.204588,22.827333,22.477516,20.96164,17.943602,13.708061,9.184435,5.3330083,3.1826572,2.0749004,1.6016173,1.6016173,1.646202,1.7422304,1.7662375,1.7902447,2.085189,2.819121,4.1943855,6.842027,10.278474,12.922686,13.718349,13.54687,13.245067,13.241637,13.55373,9.541112,7.267296,7.3564653,9.626852,13.080446,15.621771,17.518333,19.181683,21.260014,24.641586,25.649885,24.720467,21.678423,17.682953,15.241087,13.516005,10.4705305,8.217292,7.64798,8.4264965,8.237869,8.100685,8.255017,8.176137,6.5539417,6.574519,7.9257765,9.242738,10.600855,13.557159,14.555169,13.245067,12.449403,13.543441,16.462019,22.19972,21.585823,19.140528,17.655516,18.163095,16.180794,14.534592,13.594885,14.044161,16.88729,17.88873,18.62609,19.579515,20.683842,21.311457,22.347193,25.389236,28.808535,30.475315,27.748793,18.907316,13.186764,9.853205,8.001227,6.5642304,6.324159,6.327589,5.9571934,5.425607,5.751418,5.9331865,5.6519604,5.8337283,6.5059276,6.790583,7.5245147,8.879202,10.408798,11.640019,12.079007,12.9809885,12.751206,12.020704,11.173596,10.374502,11.091286,12.535142,15.282242,16.94902,12.202472,8.872343,7.2535777,6.708273,7.016936,8.378482,10.703742,13.337666,16.026463,18.36887,19.805868,18.684393,16.510035,13.96185,11.581717,9.80519,8.1487,6.4990683,5.3261495,4.5613513,3.5633414,2.9082901,2.6579304,2.5481834,2.4212887,2.2223728,2.095478,1.8108221,1.5227368,1.3615463,1.3958421,1.6084765,1.5947582,1.4644338,1.3821237,1.5673214,1.255229,0.9328478,0.7373613,0.69963586,0.7442205,0.7373613,0.59331864,0.4698535,0.41840968,0.36696586,0.33266997,0.28465575,0.24350071,0.21263443,0.18519773,0.14404267,0.1097468,0.10288762,0.10288762,0.041155048,0.044584636,0.048014224,0.05144381,0.048014224,0.037725464,0.030866288,0.041155048,0.07545093,0.12689474,0.17490897,0.16119061,0.26750782,0.3566771,0.34295875,0.20920484,0.39440256,0.4389872,0.34981793,0.2503599,0.36696586,0.5212973,0.5761707,0.44584638,0.22292319,0.18519773,0.20920484,0.30866286,0.35324752,0.29494452,0.16462019,0.106317215,0.2709374,0.41840968,0.3841138,0.07545093,0.23321195,0.31209245,0.2503599,0.116605975,0.1371835,0.24350071,0.36696586,0.32924038,0.14747226,0.061732575,0.030866288,0.041155048,0.0548734,0.048014224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.0274367,0.020577524,0.0274367,0.024007112,0.030866288,0.037725464,0.037725464,0.037725464,0.0548734,0.061732575,0.058302987,0.044584636,0.030866288,0.024007112,0.020577524,0.010288762,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.010288762,0.010288762,0.010288762,0.010288762,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.020577524,0.037725464,0.041155048,0.041155048,0.048014224,0.048014224,0.048014224,0.041155048,0.058302987,0.15090185,0.18862732,0.24007112,0.28122616,0.28808534,0.23664154,0.16462019,0.12346515,0.1097468,0.11317638,0.116605975,0.15090185,0.15776102,0.16804978,0.20234565,0.26407823,0.34981793,0.4664239,0.53501564,0.50757897,0.3806842,0.3806842,0.39783216,0.5555932,0.83681935,1.0940384,1.2689474,1.2346514,1.155771,1.2106444,1.5913286,1.5501735,1.5913286,1.6599203,1.6530612,1.430138,1.138623,0.939707,0.84024894,0.89512235,1.2175035,1.3615463,1.0940384,0.86082643,0.764798,0.5693115,0.4389872,0.4355576,0.4389872,0.37382504,0.216064,0.17147937,0.22978236,0.37382504,0.53844523,0.6241849,0.65505123,0.72707254,0.75450927,0.71678376,0.65848076,0.58988905,0.5693115,0.5761707,0.607037,0.6756287,0.6241849,0.67219913,0.7339317,0.7579388,0.7373613,0.77165717,0.764798,0.7682276,0.86082643,1.1523414,1.430138,1.6084765,1.6599203,1.6290541,1.6667795,1.8142518,2.4041407,3.0557625,3.6147852,4.173808,4.5167665,4.4413157,4.1189346,3.7451096,3.5221863,3.9680326,4.4859004,5.336438,6.3310184,6.8214493,6.468202,5.4941993,4.3795834,3.40901,2.6716487,3.069481,2.7951138,2.2841053,1.7936742,1.3546871,1.3101025,1.2483698,1.155771,1.0837497,1.1420527,1.313532,1.488441,1.7799559,2.218943,2.7642474,3.2443898,3.415869,3.7451096,4.3624353,5.0586414,5.360445,5.442755,5.504488,5.7274113,6.307011,7.31531,7.795452,7.599966,6.9792104,6.574519,6.262427,6.2075534,6.783724,8.014946,9.578837,11.228469,11.393089,10.511685,8.944365,6.9723516,5.3741636,4.1360826,3.223812,2.6579304,2.5070283,2.5584722,2.4212887,1.8725548,1.1249046,0.83338976,0.84367853,1.0666018,1.1934965,1.1420527,1.0768905,0.9877212,0.922559,0.8745448,0.84024894,0.83338976,1.1214751,1.4644338,1.8485477,2.194936,2.3424082,2.9665933,3.549623,3.7965534,3.899441,4.5339146,5.1100855,5.1821065,5.346727,5.809721,6.3961806,7.1061053,7.7714453,8.364764,8.868914,9.280463,9.31133,9.0644,8.570539,8.032094,7.8366075,6.883182,5.6142344,4.372724,3.3232703,2.4487255,1.7388009,1.1900668,0.77851635,0.47671264,0.25378948,0.18862732,0.17833854,0.19891608,0.2194936,0.21263443,0.30866286,0.3566771,0.3566771,0.33609957,0.37725464,0.35324752,0.31209245,0.31552204,0.36696586,0.40126175,0.42526886,0.47328308,0.5555932,0.64476246,0.6859175,0.6859175,0.67219913,0.65505123,0.65505123,0.6893471,0.5624523,0.4115505,0.26750782,0.15776102,0.09602845,0.09259886,0.17147937,0.36010668,0.71678376,1.3169615,2.301253,2.843128,3.1620796,3.3987212,3.6147852,3.7691166,4.108646,4.6916757,5.470192,6.2727156,6.7665763,7.143831,7.3187394,7.2158523,6.7631464,6.3790326,6.3378778,6.1561093,5.7274113,5.2987127,5.07236,5.127233,5.31929,5.5662203,5.857735,5.874883,6.3035817,7.0135064,7.6033955,7.39762,7.3084507,7.3393173,7.099246,6.691125,6.684266,6.81802,6.914048,6.824879,6.5333643,6.142391,5.610805,5.2644167,5.06893,5.0243454,5.1580997,5.305572,5.56965,5.950334,6.550512,7.5931067,8.937505,10.446524,11.674315,12.583157,13.536582,14.476289,14.730078,14.908417,15.234227,15.553179,15.162207,15.326826,15.765814,16.417435,17.408587,16.53404,15.419425,14.994157,15.271953,15.367981,15.563468,15.659496,15.46744,15.031882,14.644339,14.740367,14.819247,14.96672,15.230798,15.621771,15.913286,15.769243,15.182784,14.205351,12.96727,11.537132,9.993818,8.745448,7.98408,7.699424,7.9600725,8.405919,8.656279,8.755736,9.174147,10.542552,11.989838,12.96727,13.059869,11.976119,10.731179,9.6817255,8.690575,7.953213,7.98408,7.579388,7.3598948,8.1487,10.31277,13.742357,18.12537,21.77102,23.437801,23.27318,22.820475,22.77589,21.369759,18.752985,15.151917,10.844356,7.366754,4.9248877,3.2786856,2.301253,1.9823016,1.8965619,1.9685832,2.0097382,2.0268862,2.2086544,2.7162333,4.091498,6.3310184,8.97866,11.122152,11.444533,11.585147,11.88352,12.288212,12.349944,9.410788,7.3839016,6.835168,8.711152,14.318527,16.496315,18.79071,20.323736,21.321745,23.087982,23.965958,23.640146,21.476076,17.902447,14.407697,13.337666,12.97413,13.282792,12.984418,9.544542,9.030104,10.185875,11.458252,11.770344,10.532263,8.635701,8.004657,8.344186,9.877212,13.327377,14.421415,12.751206,11.629731,13.2862215,18.862732,19.716698,17.29198,15.388559,15.347404,16.064188,17.03819,19.558937,19.905325,18.135658,18.094503,18.571217,19.010202,19.70641,20.61182,21.314886,22.343761,23.959099,25.389236,26.047716,25.553856,19.325726,14.040731,10.082987,7.675417,6.8557453,6.975781,7.349606,7.442205,7.208993,7.099246,6.183546,5.7994323,6.0154963,6.461343,6.310441,7.1026754,8.865483,11.369082,14.027013,15.896138,16.79126,16.321407,15.858413,15.13134,12.212761,9.949233,10.299051,12.977559,15.6697855,14.030442,10.419086,8.512236,7.414768,7.016936,7.963502,9.678296,11.321068,12.4974165,13.152468,13.5503,13.128461,12.229909,11.005547,9.630281,8.268735,6.7871537,5.892031,5.209543,4.6093655,4.201245,5.0586414,5.5147767,5.5593615,5.15467,4.245829,3.5599117,2.9871707,2.4727325,2.095478,2.0646117,2.0234566,1.845118,1.7662375,1.8519772,1.9994495,1.786815,1.5193073,1.255229,1.0151579,0.7922347,0.8265306,0.8711152,0.9328478,0.91569984,0.64819205,0.50757897,0.42869842,0.3806842,0.36353627,0.4046913,0.42183927,0.4629943,0.48014224,0.4355576,0.2777966,0.25721905,0.31895164,0.39783216,0.4389872,0.39783216,0.22978236,0.14747226,0.18176813,0.29151493,0.36010668,0.36353627,0.4115505,0.5555932,0.70306545,0.6344737,0.45613512,0.39440256,0.37382504,0.3566771,0.3566771,0.47328308,0.6173257,0.64133286,0.5624523,0.59674823,0.7339317,0.72707254,0.6207553,0.48014224,0.3806842,0.2503599,0.41840968,0.6790583,0.8779744,0.922559,1.2346514,1.4267083,1.3649758,1.0940384,0.8162418,0.6893471,0.5727411,0.4046913,0.2709374,0.38754338,0.41840968,0.20577525,0.048014224,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.10288762,0.11317638,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.017147938,0.010288762,0.0,0.0,0.0,0.006859175,0.006859175,0.0034295875,0.010288762,0.010288762,0.020577524,0.030866288,0.041155048,0.06516216,0.058302987,0.034295876,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0034295875,0.006859175,0.006859175,0.01371835,0.01371835,0.01371835,0.024007112,0.041155048,0.048014224,0.037725464,0.030866288,0.024007112,0.020577524,0.01371835,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.0274367,0.034295876,0.041155048,0.041155048,0.037725464,0.034295876,0.058302987,0.15090185,0.20920484,0.2469303,0.26064864,0.25378948,0.24350071,0.17490897,0.11317638,0.08916927,0.10288762,0.12689474,0.16804978,0.17833854,0.18862732,0.22292319,0.30523327,0.4081209,0.4698535,0.5007198,0.47328308,0.33266997,0.33952916,0.4389872,0.65162164,0.9774324,1.3752645,1.4369972,1.2963841,1.2209331,1.3272504,1.5673214,1.4335675,1.3992717,1.4850113,1.5981878,1.529596,1.529596,1.4164196,1.2929544,1.2346514,1.2723769,1.1729189,0.72021335,0.45270553,0.47328308,0.45613512,0.42526886,0.5555932,0.59331864,0.47328308,0.29494452,0.2469303,0.37725464,0.6001778,0.85396725,1.0734608,1.2209331,1.2209331,1.08032,0.864256,0.6824879,0.64819205,0.6893471,0.7407909,0.78194594,0.8196714,0.83681935,0.89512235,0.9568549,0.9877212,0.939707,0.91227025,0.85396725,0.7888051,0.805953,1.0563129,1.3272504,1.6667795,2.0474637,2.294394,2.0817597,2.085189,2.6167753,3.2992632,3.841138,4.029765,3.6868064,3.3198407,3.0214665,2.867135,2.9185789,3.7348208,4.623084,5.5147767,6.1801167,6.210983,5.7239814,4.636802,3.758828,3.3644254,3.1826572,3.2958336,2.8705647,2.4041407,2.1126258,1.9342873,1.978872,1.7971039,1.5227368,1.255229,1.0631721,1.2106444,1.4575747,1.7593783,2.1880767,2.9288676,3.6147852,4.1326528,4.6402316,5.2026844,5.8165803,6.293293,6.4098988,6.3653145,6.2830043,6.217842,6.9380555,7.4524937,7.5759587,7.3221693,6.8969,6.495639,6.108095,6.2692857,7.1849856,8.724871,10.065839,9.897789,8.666568,6.852316,4.996909,4.0366244,3.1346428,2.3492675,1.7593783,1.4507155,1.3169615,1.1660597,0.9259886,0.6962063,0.764798,1.0151579,1.3992717,1.5330256,1.3581166,1.1317638,0.89169276,0.90541106,1.0288762,1.1900668,1.3889829,1.7010754,1.8279701,1.9274281,2.194936,2.8568463,3.5873485,4.180667,4.434457,4.3590055,4.170378,4.1600895,4.4516044,4.938606,5.5490727,6.2555676,7.15069,8.086967,8.937505,9.630281,10.158438,9.455373,8.656279,7.7714453,6.8626046,6.060081,5.1821065,4.2526884,3.199805,2.16064,1.4575747,1.0323058,0.7339317,0.5041494,0.31895164,0.19891608,0.26407823,0.2777966,0.26407823,0.22978236,0.17147937,0.1920569,0.21263443,0.24350071,0.274367,0.29151493,0.28465575,0.31209245,0.41498008,0.548734,0.6036074,0.52815646,0.5453044,0.53501564,0.45613512,0.34981793,0.34638834,0.37382504,0.4081209,0.41498008,0.36696586,0.3018037,0.22635277,0.16462019,0.1371835,0.14061308,0.2194936,0.45956472,0.82996017,1.3443983,2.0646117,3.1826572,3.6319332,3.8788633,4.1772375,4.5784993,4.7808447,5.2335505,5.878313,6.543653,6.914048,7.0889573,7.1266828,7.0032177,6.759717,6.5196457,6.5985265,6.701414,6.5059276,6.018926,5.579939,5.5387836,5.5490727,5.6313825,5.8165803,6.135532,6.23156,6.540223,7.1232533,7.630832,7.3255987,7.281014,7.4970784,7.4010496,6.9792104,6.7871537,6.848886,6.8557453,6.7700057,6.5950966,6.368744,6.042933,5.8234396,5.720552,5.7308407,5.830299,5.9571934,6.118384,6.375603,6.8283086,7.6342616,8.752307,10.398509,12.116733,13.738928,15.405707,16.424294,16.462019,16.307688,16.208231,15.854982,15.8138275,16.12249,16.45516,16.942162,18.176813,17.473747,16.173935,15.700651,16.235666,16.736387,17.29541,17.274832,16.828985,16.167076,15.553179,15.395418,15.357693,15.577187,16.03675,16.554619,17.37772,17.782412,17.391438,16.235666,14.754086,12.854094,10.823778,9.22902,8.258447,7.7131424,7.6616983,7.8023114,8.001227,8.220721,8.525954,10.031544,11.876661,13.649758,14.712931,14.191633,13.262215,11.664027,9.856634,8.443645,8.158989,7.6857057,7.332458,8.097256,10.244178,13.296511,17.45317,20.584383,22.419212,23.012531,22.734735,22.336903,20.827885,18.420315,15.409137,12.185325,9.4862385,6.948344,4.911169,3.5153272,2.7402403,2.3801336,2.428148,2.5961976,2.7333813,2.867135,3.199805,4.506478,6.5059276,8.745448,10.621432,10.871792,11.005547,11.211322,11.413667,11.245617,10.209882,8.515666,7.3084507,7.9943686,12.22648,14.459141,17.758404,20.61525,22.415783,23.465237,23.297188,22.556396,20.917053,18.313997,14.939283,14.05102,15.182784,16.026463,14.685493,9.674867,8.553391,9.465661,11.015835,12.418536,13.498857,12.024134,11.592006,12.281353,13.992717,16.45859,16.890718,16.002455,14.496866,14.071597,17.412016,14.867262,11.97269,10.786053,11.485688,12.367092,13.581166,16.79126,18.001905,16.828985,16.520323,17.12393,17.655516,17.840714,17.809847,18.108221,18.667244,18.982767,18.862732,18.756414,19.761284,18.338005,14.332246,10.429376,8.141841,7.7748747,7.8194594,8.179566,8.491658,8.742019,9.290752,7.9772205,7.0272245,7.366754,8.361334,7.7920227,7.281014,8.025234,10.360784,13.629181,16.208231,17.343424,18.193962,19.243416,19.634388,17.154797,13.114742,11.509696,11.773774,12.854094,13.231348,11.382801,10.696883,10.288762,9.911508,9.959522,10.062409,10.106995,9.640571,8.683716,7.740579,7.257007,7.0272245,6.756287,6.2967224,5.645101,4.8734436,4.6882463,4.3761535,3.9783216,4.3178506,6.0703697,7.298162,7.682276,7.1987042,6.108095,5.178677,4.619654,4.245829,4.016047,4.0229063,3.5221863,3.1312134,2.9151495,2.8705647,2.9460156,2.6579304,2.3801336,2.061182,1.6667795,1.1660597,1.0837497,1.2723769,1.4507155,1.4472859,1.1900668,0.97400284,0.7922347,0.6379033,0.548734,0.61389613,0.69963586,0.7682276,0.8711152,0.89512235,0.5761707,0.5418748,0.7579388,0.89169276,0.84024894,0.70649505,0.4698535,0.30866286,0.29837412,0.41498008,0.5418748,0.61389613,0.58302987,0.6379033,0.7442205,0.65162164,0.42526886,0.40126175,0.39440256,0.32238123,0.18519773,0.29151493,0.6001778,0.7510797,0.70306545,0.72707254,1.0357354,0.96371406,0.7613684,0.6001778,0.5761707,0.41840968,0.548734,0.91569984,1.3615463,1.6359133,1.728512,1.7696671,1.704505,1.4918705,1.097468,0.83338976,0.59331864,0.39440256,0.30523327,0.4355576,0.5041494,0.32924038,0.18519773,0.14404267,0.06859175,0.034295876,0.030866288,0.072021335,0.11317638,0.0548734,0.11317638,0.11317638,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.0274367,0.037725464,0.030866288,0.024007112,0.010288762,0.0,0.006859175,0.0548734,0.1097468,0.13375391,0.11317638,0.05144381,0.030866288,0.034295876,0.041155048,0.048014224,0.06516216,0.061732575,0.037725464,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.020577524,0.030866288,0.024007112,0.024007112,0.020577524,0.01371835,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.020577524,0.024007112,0.0274367,0.030866288,0.030866288,0.030866288,0.041155048,0.1097468,0.13032432,0.13032432,0.14404267,0.22292319,0.16462019,0.10288762,0.08573969,0.12346515,0.18176813,0.216064,0.2469303,0.2777966,0.31895164,0.3806842,0.44584638,0.4115505,0.36696586,0.34295875,0.31895164,0.36353627,0.4664239,0.58988905,0.8505377,1.5193073,1.8313997,1.6427724,1.3684053,1.2277923,1.2415106,1.3752645,1.3615463,1.3169615,1.313532,1.3855534,1.9308578,2.1915064,2.1126258,1.670209,0.8745448,0.548734,0.33266997,0.28122616,0.33266997,0.3018037,0.42526886,0.67219913,0.7339317,0.5693115,0.4115505,0.35324752,0.5212973,0.83681935,1.2277923,1.6256244,1.8279701,1.7662375,1.4747226,1.0563129,0.6893471,0.6962063,0.8128122,0.9534253,1.0425946,1.039165,1.0734608,1.0323058,1.0220171,1.0734608,1.1283343,0.9945804,0.83338976,0.71678376,0.6756287,0.7339317,0.8676856,1.2655178,2.0508933,2.8294096,2.668219,2.7299516,3.0454736,3.525616,3.9200184,3.8377085,2.9254382,2.6579304,2.6579304,2.784825,3.1380725,3.8171308,4.4275975,4.846007,4.9660425,4.6779575,4.633373,4.4996185,4.314421,4.064061,3.6765177,3.3678548,2.8808534,2.5790498,2.5619018,2.6990852,2.877424,2.6167753,2.2086544,1.8416885,1.5913286,1.6393428,1.7696671,1.9582944,2.3252604,3.1277838,3.8788633,4.5270553,5.038064,5.552502,6.3790326,7.3530354,7.7097125,7.675417,7.442205,7.160979,7.4353456,8.052671,8.694004,8.879202,7.98065,7.349606,6.728851,5.977771,5.597087,6.728851,7.675417,7.5759587,6.4579134,4.773986,3.3952916,3.1346428,2.644212,2.0680413,1.4987297,0.9568549,0.64133286,0.52472687,0.6001778,0.84024894,1.1797781,1.4541451,1.6633499,1.6187652,1.3512574,1.0871792,0.8848336,1.0220171,1.2963841,1.587899,1.8691251,1.9342873,1.8108221,1.7353712,2.0303159,3.100347,3.6079261,3.8479972,3.8308492,3.6010668,3.2546785,3.2272418,3.6868064,4.465323,5.4324665,6.495639,7.675417,8.618553,9.294182,9.685155,9.791472,8.673427,7.500508,6.293293,5.1580997,4.3007026,3.5942078,2.952875,2.1503513,1.2963841,0.823101,0.65162164,0.5521636,0.45613512,0.34981793,0.2777966,0.41498008,0.432128,0.38754338,0.31209245,0.22292319,0.21263443,0.2503599,0.34638834,0.42183927,0.3018037,0.24007112,0.31209245,0.4938606,0.6962063,0.77508676,0.67219913,0.5761707,0.490431,0.41498008,0.36010668,0.31209245,0.30523327,0.29494452,0.26750782,0.22292319,0.17833854,0.12346515,0.1097468,0.16119061,0.23664154,0.3841138,0.7922347,1.2998136,1.845118,2.4555845,3.4124396,3.9714622,4.40702,4.8905916,5.4667625,6.0669403,6.5779486,6.989499,7.1712675,6.8763227,6.615674,6.3378778,6.1458206,6.166398,6.5642304,7.3084507,7.2432885,6.8763227,6.4407654,5.888602,5.7068334,5.6176643,5.5902276,5.6176643,5.7377,5.669108,5.7136927,5.970912,6.3173003,6.3824625,6.5779486,7.06495,7.3598948,7.332458,7.2124224,7.2124224,7.0443726,6.8111606,6.619104,6.5779486,6.619104,6.7494283,6.9552035,7.160979,7.2432885,7.267296,7.31531,7.4799304,7.81603,8.333898,9.194724,10.89237,13.059869,15.357693,17.480608,18.331144,18.591793,18.36544,17.62465,16.21852,16.852993,17.672665,17.892159,17.741257,18.485476,18.756414,18.053349,17.645227,17.988186,18.725548,20.059656,20.35803,20.090523,19.44919,18.358582,17.267973,16.657507,16.70552,17.20624,17.559488,18.427174,19.075365,18.722118,17.305698,15.46401,13.327377,11.163307,9.349055,8.035523,7.14726,7.0203657,7.1541195,7.431916,7.73372,7.9257765,8.98209,10.333347,12.236768,14.171056,14.839825,14.246507,12.5145645,10.635151,9.078118,7.8091707,6.893471,6.3618846,6.783724,8.351046,10.878652,14.668345,17.86815,20.296299,21.733295,21.942501,20.814167,19.253704,17.12393,14.757515,12.936404,10.950673,8.711152,6.7219915,5.137522,3.7519686,3.1312134,3.0386145,3.1860867,3.426158,3.7485392,4.280125,5.545643,7.73029,10.31277,12.041282,12.428825,12.082437,11.698323,11.523414,11.345076,12.171606,11.327928,10.082987,9.335337,9.589127,11.763485,15.357693,19.19197,22.43979,24.641586,24.69303,23.485815,21.664703,19.552078,17.165085,16.249386,16.839275,15.971589,12.9809885,9.506817,7.373613,6.684266,7.654839,9.993818,12.895248,13.869251,15.494876,17.689812,19.740705,20.316875,19.349733,20.351171,19.678972,16.894148,14.781522,13.954991,12.325937,11.05699,10.710602,11.262765,9.571979,9.277034,9.469091,10.052121,11.739478,13.29994,14.531162,15.011304,15.13134,16.091625,17.03819,16.191082,14.339106,13.080446,14.808959,16.808409,14.428274,10.882081,8.457363,8.536243,8.913498,8.796892,8.64256,9.012956,10.593996,9.822338,8.663138,9.499957,11.698323,11.595435,8.820899,7.1369715,7.3598948,9.283894,11.694893,13.677195,16.856422,19.768143,21.486366,21.626978,18.921034,17.12736,15.388559,13.594885,12.415107,12.891819,13.728639,14.29452,14.099034,12.785502,10.80663,9.253027,7.881192,6.691125,5.936616,5.086078,4.6745276,4.461893,4.3178506,4.214963,4.2389703,4.386442,4.280125,4.1120753,4.6402316,6.029215,7.4936485,8.186425,7.9429245,7.2878733,6.6122446,6.39961,6.478491,6.6533995,6.701414,5.8988905,5.4839106,5.0174866,4.482471,4.2698364,3.782835,3.3781435,3.000889,2.551613,1.879414,1.5398848,1.6770682,1.9068506,2.0028791,1.8554068,1.5055889,1.2998136,1.097468,0.90884066,0.8505377,0.8471081,0.8779744,1.0768905,1.255229,0.91227025,0.84024894,1.0871792,1.1317638,0.8848336,0.7133542,0.6001778,0.4664239,0.4629943,0.6036074,0.77508676,0.823101,0.7373613,0.64133286,0.5521636,0.36353627,0.42526886,0.51100856,0.42869842,0.19548649,0.044584636,0.17490897,0.5521636,0.6790583,0.5178677,0.47671264,0.8505377,0.8711152,0.7682276,0.69963586,0.7510797,0.61046654,0.6790583,1.039165,1.5604624,1.9102802,1.6153357,1.3443983,1.2758065,1.2758065,0.90198153,0.6241849,0.47328308,0.36010668,0.2503599,0.17833854,0.2194936,0.26750782,0.29494452,0.26407823,0.13375391,0.06516216,0.06516216,0.14747226,0.22635277,0.1097468,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.041155048,0.082310095,0.09602845,0.044584636,0.01371835,0.0,0.0034295875,0.01371835,0.1097468,0.20920484,0.25721905,0.22292319,0.08573969,0.048014224,0.030866288,0.020577524,0.010288762,0.0,0.010288762,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.020577524,0.037725464,0.061732575,0.072021335,0.08573969,0.08573969,0.07888051,0.09259886,0.12689474,0.082310095,0.058302987,0.08916927,0.1371835,0.08916927,0.058302987,0.05144381,0.082310095,0.16804978,0.25378948,0.3018037,0.30866286,0.29494452,0.31895164,0.3566771,0.40126175,0.41498008,0.39440256,0.3806842,0.4424168,0.44927597,0.51100856,0.70306545,1.0666018,1.214074,1.3066728,1.371835,1.3992717,1.3272504,1.155771,0.89512235,0.7407909,0.8745448,1.4335675,2.253239,2.6853669,2.4830213,1.670209,0.53501564,0.4115505,0.29151493,0.18176813,0.12003556,0.16804978,0.48357183,0.77508676,0.83681935,0.66876954,0.47328308,0.37382504,0.45270553,0.90884066,1.6256244,2.1503513,1.8348293,1.4610043,1.1008976,0.77508676,0.45613512,0.83681935,1.1420527,1.3443983,1.3341095,0.9294182,0.7099246,0.65505123,0.70649505,0.7888051,0.823101,0.7888051,0.7339317,0.67219913,0.6241849,0.61046654,0.70649505,0.9602845,1.3752645,1.9720128,2.7779658,3.5839188,4.149801,4.029765,3.5050385,3.6147852,4.091498,4.6402316,4.6676683,4.1635194,3.724532,4.149801,4.064061,4.016047,4.4104495,5.5079174,5.970912,6.060081,5.744559,5.007198,3.8617156,3.0900583,2.760818,2.6819375,2.784825,3.1140654,3.7108135,3.8788633,3.82399,3.6525106,3.3712845,3.0797696,2.8225505,2.620205,2.5653315,2.8225505,3.1037767,3.4295874,3.8925817,4.7671266,6.4990683,8.440215,9.465661,9.661148,9.349055,9.078118,9.81205,11.019264,12.144169,12.668896,12.130451,10.786053,9.043822,6.8283086,5.2026844,6.3618846,7.143831,7.0375133,5.8645945,4.0880685,2.8088322,2.393852,1.8416885,1.3169615,0.90541106,0.6241849,0.48014224,0.45956472,0.5761707,0.84024894,1.2655178,1.6084765,1.8759843,1.8897027,1.6839274,1.5261664,1.4404267,1.5193073,1.6907866,1.8691251,1.9685832,1.5055889,1.4267083,1.5844694,1.8931323,2.318401,3.0523329,3.3266997,2.7711067,1.8862731,2.0440342,2.8877127,4.297273,5.675967,6.835168,7.9943686,9.2153015,9.678296,9.462232,8.618553,7.140401,6.0532217,4.9420357,3.799983,2.760818,2.0920484,1.4918705,0.94999576,0.607037,0.4938606,0.5178677,0.64133286,0.64476246,0.5453044,0.38754338,0.22978236,0.32581082,0.41498008,0.48357183,0.5144381,0.5041494,0.6001778,0.6790583,0.65162164,0.5212973,0.4115505,0.34981793,0.33609957,0.32924038,0.37382504,0.5796003,1.1900668,1.2860953,1.1420527,0.89855194,0.5796003,0.5418748,0.4698535,0.34638834,0.26064864,0.3806842,0.3566771,0.23321195,0.20234565,0.28808534,0.33609957,0.432128,0.91569984,1.5570327,2.2841053,3.1895163,4.897451,6.001778,6.64997,6.917478,6.8214493,6.7459984,6.7391396,6.9380555,7.181556,6.9723516,6.6431108,6.385892,6.0806584,5.7822843,5.720552,6.368744,6.8145905,6.9792104,6.8043017,6.2555676,5.830299,5.5113473,5.2918534,5.003768,4.3349986,4.040054,4.0503426,4.2766957,4.695105,5.3570156,6.3447366,7.4970784,8.351046,8.711152,8.652849,8.261876,7.8434668,7.459353,7.274155,7.5690994,7.9600725,8.340756,8.652849,8.844906,8.879202,8.8929205,8.995808,9.2153015,9.592556,10.179015,11.30049,13.22106,15.313108,17.189093,18.677534,19.898466,20.594673,20.639257,20.111101,19.318867,19.476627,20.440342,21.064526,21.109112,21.256582,21.45207,20.896477,20.412905,20.385468,20.752434,22.53239,23.547548,23.815056,23.218307,21.482935,19.44576,17.682953,17.29198,18.241976,19.377169,20.244854,20.207129,19.325726,17.830425,16.098484,14.30481,12.336226,10.491108,9.026674,8.1487,7.8537555,7.798882,7.9463544,8.1212635,8.011517,8.268735,8.934075,10.487679,12.55915,13.96185,14.4145565,12.538571,10.288762,8.601405,7.431916,6.5162163,5.90232,5.6142344,5.936616,7.4010496,10.329918,13.680624,16.513464,18.012194,17.487467,15.999025,15.340545,14.784951,13.999576,13.046151,11.8115,10.618003,9.170717,7.2158523,4.530485,3.8720043,3.542764,3.40901,3.5290456,4.149801,5.4941993,7.349606,10.278474,13.666906,15.717799,15.217079,13.598314,11.900668,10.696883,10.086417,15.055889,17.154797,16.777542,15.107333,14.1299,14.263655,15.230798,16.45173,18.015623,20.676983,23.753323,24.219748,23.046827,21.133118,19.301718,18.77699,18.965618,18.900457,17.501184,13.594885,10.995257,9.438225,9.482809,10.206452,9.23245,9.074688,10.683165,15.155347,20.731855,22.78275,18.28999,20.351171,22.817045,22.559826,19.469769,20.11796,18.996485,16.407146,13.54687,12.4974165,12.483699,12.939834,12.017275,9.9698105,9.139851,9.273604,10.765475,13.845244,18.410025,24.000254,28.054026,23.20802,15.22051,10.377932,15.518884,16.715809,15.704081,12.250486,8.436785,8.683716,9.695444,8.968371,8.090397,7.7371492,7.675417,8.213862,9.153569,10.587136,12.6586075,15.563468,12.377381,9.163857,6.3138704,4.616225,5.2506986,8.275595,12.895248,16.540901,18.526632,20.066517,21.225718,22.823904,22.714157,20.395756,17.027903,17.223389,16.935303,16.348843,15.470869,14.1299,11.993267,9.719451,7.7920227,6.495639,5.936616,5.7891436,5.8988905,5.593657,4.787704,3.981751,3.7142432,4.3624353,5.171818,5.65539,5.56965,6.948344,8.035523,8.738589,8.81404,7.874333,7.48336,7.531374,7.7268605,7.8126,7.5690994,7.2158523,7.517656,7.3427467,6.307011,4.804852,4.4275975,4.1120753,3.765687,3.2718265,2.503599,1.978872,1.920569,2.4247184,2.952875,2.318401,1.5021594,1.6804979,1.978872,1.937717,1.5090185,0.99801,0.91569984,1.0323058,1.2175035,1.4507155,1.2792361,0.99801,0.6241849,0.31209245,0.33609957,0.44584638,0.53844523,0.8128122,1.1660597,1.1900668,0.7990939,0.64819205,0.61046654,0.607037,0.59674823,0.47328308,0.31552204,0.16119061,0.06859175,0.106317215,0.06859175,0.061732575,0.06859175,0.1097468,0.24350071,0.41498008,0.823101,1.1351935,1.2277923,1.1900668,0.97057325,0.89855194,1.0082988,1.3855534,2.1674993,2.1057668,1.9171394,1.9651536,2.0131679,1.2209331,0.64819205,0.40126175,0.274367,0.16462019,0.09259886,0.0548734,0.0274367,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.116605975,0.14404267,0.106317215,0.044584636,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.006859175,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.034295876,0.05144381,0.05144381,0.037725464,0.048014224,0.048014224,0.06516216,0.09259886,0.06859175,0.06516216,0.05144381,0.061732575,0.09259886,0.09945804,0.082310095,0.058302987,0.058302987,0.07888051,0.106317215,0.14404267,0.216064,0.30523327,0.4115505,0.5521636,0.47328308,0.4081209,0.36696586,0.34295875,0.31895164,0.37039545,0.47671264,0.70649505,1.0425946,1.3992717,1.7010754,1.7079345,1.611906,1.529596,1.4850113,1.8245405,1.6736387,1.1214751,0.6756287,1.2758065,2.4658735,3.6799474,3.3987212,1.8176813,0.84024894,0.65848076,0.41840968,0.2469303,0.19548649,0.25378948,0.5212973,0.7407909,0.85739684,0.8471081,0.7305021,0.61046654,0.59674823,0.82996017,1.2449403,1.5536032,1.6256244,1.5776103,1.3375391,0.96371406,0.66533995,0.90541106,0.9568549,0.90198153,0.7888051,0.65162164,0.5555932,0.548734,0.64133286,0.7476501,0.6790583,0.64133286,0.70306545,0.66533995,0.5727411,0.70649505,1.255229,1.2689474,1.2655178,1.5158776,2.0680413,2.6304936,2.9117198,2.8088322,2.5001693,2.4452958,2.6956558,3.1517909,3.8034124,4.2869844,3.9063,3.1895163,3.858286,4.5270553,4.6265135,4.396731,3.875434,3.8479972,4.0057583,3.9131594,3.0317552,3.0146074,3.2306714,3.2889743,3.175798,3.2718265,3.5564823,3.799983,3.9508848,3.9954693,3.957744,3.8034124,3.4535947,3.117495,2.9631636,3.1517909,3.2375305,3.4707425,3.9954693,4.8494368,5.9880595,7.840037,10.285333,11.698323,11.845795,11.897239,12.298501,11.958971,11.598865,11.543991,11.729189,11.2250395,10.086417,8.31332,6.4373355,5.4976287,4.822,4.1600895,3.2306714,2.1640697,1.5398848,1.4164196,1.3546871,1.214074,0.96371406,0.66191036,0.53501564,0.6379033,0.91227025,1.2483698,1.5090185,1.9514352,2.3321195,2.3972816,2.1812177,2.0131679,1.9274281,1.9720128,2.2635276,2.6716487,2.7985435,1.7010754,1.8862731,2.551613,3.1140654,3.210094,2.9940298,3.0557625,3.525616,4.870014,7.8777623,9.688584,9.873782,9.530824,9.187865,8.81404,8.375052,7.5416627,6.5024977,5.3501563,4.0880685,3.1415021,2.294394,1.5536032,0.9774324,0.6859175,0.4698535,0.30866286,0.25378948,0.28808534,0.31209245,0.33609957,0.34295875,0.34295875,0.34638834,0.36353627,0.432128,0.4972902,0.5658819,0.61389613,0.6001778,0.5521636,0.50757897,0.51100856,0.5212973,0.4115505,0.29151493,0.26407823,0.35324752,0.5555932,0.8128122,1.0906088,0.9945804,0.77165717,0.58645946,0.5418748,0.6927767,0.72364295,0.5624523,0.31895164,0.29494452,0.26064864,0.1920569,0.17833854,0.33609957,0.823101,1.8485477,2.4898806,3.1792276,4.149801,5.422178,6.0395036,6.385892,6.495639,6.433906,6.307011,6.186976,6.077229,6.0086374,5.9812007,5.960623,5.9812007,5.9228973,5.720552,5.425607,5.195825,5.754848,6.3035817,6.776865,7.0272245,6.8283086,6.783724,6.6053853,6.029215,5.137522,4.3590055,4.0366244,4.3521466,4.887162,5.4667625,6.1732574,7.143831,8.131552,8.903209,9.297611,9.239308,9.325048,9.349055,9.256456,9.146709,9.263316,9.568549,10.000677,10.371073,10.583707,10.63858,10.542552,10.868362,11.619442,12.80265,14.424845,15.488017,16.595774,17.655516,18.917604,20.982216,22.312897,23.074265,23.156574,23.02968,23.760181,25.26577,25.821363,25.958548,26.02028,26.136887,26.35295,26.082012,25.574434,25.02227,24.548986,26.126596,27.827673,29.082901,29.59734,29.35727,28.60619,27.364677,27.632187,29.51846,31.219534,30.67766,28.60276,25.797358,22.796469,19.881319,18.008764,16.256245,14.606613,12.864383,10.63858,9.448513,9.283894,9.146709,8.687145,8.207003,8.004657,7.9772205,8.327039,9.050681,9.945804,10.155008,9.73317,9.108984,8.457363,7.723431,6.9552035,6.262427,6.169828,6.8797526,8.268735,10.14129,11.660598,12.682614,13.118172,12.932974,12.079007,12.027563,12.3533745,12.679185,12.703192,12.614022,12.2093315,10.957532,8.927217,6.776865,5.346727,4.650521,4.40359,4.5030484,5.0174866,6.3310184,7.8777623,9.774324,11.849225,13.666906,13.056439,12.0138445,10.909517,9.9801,9.328478,10.587136,11.849225,12.79922,13.461131,14.201921,15.577187,16.523752,18.20082,21.314886,26.143745,26.555296,24.552416,21.016512,17.638369,16.921585,16.084764,15.162207,13.954991,13.567448,16.438013,21.407484,17.693241,12.737488,9.788043,7.9120584,7.9120584,9.318189,11.797781,14.517444,16.12935,16.647217,17.545769,17.003895,14.932424,12.977559,12.325937,12.0138445,11.790922,11.893809,13.070158,17.130789,17.45317,16.71238,17.267973,21.174273,15.402277,10.652299,8.7283,10.847785,17.679523,19.672113,14.997586,10.172156,9.057541,12.867812,18.910746,19.20569,16.667795,13.594885,11.660598,10.515115,9.22902,8.1384115,7.2638664,6.2830043,5.7377,5.439326,5.6176643,6.2727156,7.1678376,6.392751,5.3844523,4.479041,3.9268777,3.9200184,4.671098,6.948344,9.441654,11.129011,11.290202,11.375941,11.97269,13.162757,14.575747,15.405707,16.167076,15.820687,15.12448,14.452282,13.810948,13.581166,11.876661,10.007536,8.868914,8.961512,8.913498,8.988949,9.105555,8.841476,7.449064,6.8763227,7.332458,8.032094,8.587687,9.012956,9.863494,11.317638,12.576297,13.173045,12.97413,10.456812,8.587687,7.2604365,6.3893213,5.919468,5.528495,5.206114,4.5819287,3.8479972,3.7931237,4.431027,4.2389703,3.7211025,3.1483612,2.5756202,2.4624438,3.0111778,3.957744,4.7191124,4.40702,3.899441,3.7794054,4.012617,4.40702,4.5853586,4.297273,3.093488,2.369845,2.5001693,2.8396983,2.603057,2.4590142,2.3458378,2.2292318,2.1160555,1.6221949,1.2826657,1.255229,1.4164196,1.371835,1.2380811,1.2003556,1.1146159,0.9431366,0.75450927,0.58302987,0.5590228,0.5144381,0.3566771,0.082310095,0.07545093,0.09602845,0.1371835,0.21263443,0.36696586,0.5555932,0.7510797,0.91227025,1.0117283,1.0425946,0.980862,0.94656616,1.1592005,1.7010754,2.5207467,2.7539587,2.417859,1.9274281,1.4815818,1.0494537,1.0425946,1.1008976,0.9328478,0.5521636,0.274367,0.1097468,0.06516216,0.0548734,0.034295876,0.01371835,0.01371835,0.0034295875,0.116605975,0.4698535,1.1832076,0.9877212,0.6824879,0.34638834,0.1371835,0.29151493,0.34295875,0.22292319,0.09945804,0.037725464,0.0,0.0,0.017147938,0.041155048,0.05144381,0.044584636,0.01371835,0.010288762,0.017147938,0.024007112,0.024007112,0.024007112,0.024007112,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.006859175,0.0034295875,0.006859175,0.01371835,0.01371835,0.037725464,0.058302987,0.058302987,0.037725464,0.020577524,0.0274367,0.041155048,0.06859175,0.09602845,0.08916927,0.09259886,0.09259886,0.08916927,0.08573969,0.09259886,0.1097468,0.1097468,0.10288762,0.10288762,0.12689474,0.17490897,0.2194936,0.32581082,0.48014224,0.59331864,0.3566771,0.28465575,0.30866286,0.39783216,0.5418748,0.48357183,0.5212973,0.7476501,1.0837497,1.2620882,1.6084765,2.085189,2.07833,1.6256244,1.3992717,1.8382589,1.6530612,1.2003556,0.9602845,1.5193073,2.318401,2.9254382,2.6956558,1.7696671,1.08032,0.7305021,0.45613512,0.28122616,0.2194936,0.26407823,0.4698535,0.6379033,0.7373613,0.7373613,0.61046654,0.61389613,0.7133542,0.9534253,1.2003556,1.1489118,1.1283343,1.097468,0.9602845,0.7442205,0.58988905,0.65162164,0.64476246,0.6036074,0.5590228,0.5418748,0.5624523,0.5624523,0.5796003,0.59331864,0.53158605,0.5761707,0.65505123,0.61046654,0.5041494,0.58645946,0.91569984,0.96371406,1.0837497,1.3958421,1.7730967,2.0303159,2.194936,2.1743584,1.9994495,1.821111,2.170929,2.5893385,3.018037,3.350707,3.4295874,3.2786856,3.8479972,4.2526884,4.2389703,4.184097,4.4687524,4.6127954,4.5167665,3.9474552,2.5310357,2.6716487,2.8877127,2.9254382,2.8054025,2.7985435,3.216953,3.974892,4.3795834,4.3281393,4.280125,4.2218223,4.0606318,3.923448,3.8925817,4.012617,4.297273,4.5167665,4.722542,5.0140567,5.521636,7.051232,9.496528,12.281353,14.685493,15.854982,15.964729,15.604623,15.059319,14.455711,13.759505,11.519984,9.719451,8.097256,6.543653,5.113515,3.9440255,2.942586,2.1057668,1.5193073,1.3478279,1.4164196,1.4027013,1.2517995,0.9842916,0.70649505,0.77508676,0.96371406,1.2380811,1.5501735,1.8382589,2.2566686,2.5996273,2.6785078,2.5138876,2.318401,2.1229146,1.9720128,2.0234566,2.2429502,2.3835633,2.0646117,2.1846473,2.5138876,2.8808534,3.1483612,2.784825,2.976882,3.9783216,5.874883,8.577398,10.065839,10.124143,9.342196,8.196714,7.06838,5.9880595,5.0655007,4.1463714,3.1449318,2.054323,1.4369972,0.939707,0.5624523,0.32924038,0.2709374,0.2503599,0.26064864,0.34295875,0.44927597,0.41498008,0.26750782,0.22292319,0.22635277,0.24350071,0.26064864,0.2777966,0.34981793,0.4424168,0.490431,0.4046913,0.34295875,0.29837412,0.30523327,0.32924038,0.28465575,0.24350071,0.26750782,0.44584638,0.7510797,1.0254467,0.86082643,0.65505123,0.4698535,0.36353627,0.38754338,0.4424168,0.4355576,0.33266997,0.1920569,0.14747226,0.14747226,0.20920484,0.4629943,0.94656616,1.6324836,2.4658735,3.1277838,3.8137012,4.57164,5.295283,5.909179,6.293293,6.3378778,6.138962,5.9983487,6.0154963,6.1629686,6.3961806,6.7391396,7.2638664,7.9292064,8.086967,7.922347,7.5519514,7.0443726,7.222711,7.2775846,7.1884155,7.0032177,6.8283086,6.8900414,6.9380555,6.56766,5.857735,5.3432975,5.1821065,5.161529,5.2918534,5.6039457,6.138962,7.2432885,8.30646,9.256456,10.021255,10.545981,10.782623,10.792912,10.707172,10.690024,10.9541025,11.55428,12.566009,13.423406,13.872682,13.972139,13.666906,14.006435,14.860402,16.108772,17.658945,18.509483,19.20912,19.929333,20.978786,22.806757,24.374079,25.708187,26.702768,27.567024,28.84626,30.286688,31.099499,31.58993,31.830002,31.651663,32.59137,33.462486,34.192986,34.7623,35.22872,35.921497,36.09641,35.97637,35.798035,35.82204,36.720592,35.969513,35.25959,35.050385,34.56338,32.224403,29.34698,26.34266,23.482386,20.910194,19.137098,17.741257,16.300829,14.579176,12.5145645,11.019264,10.786053,10.628291,10.038403,9.2153015,8.340756,7.658269,7.2124224,7.0752387,7.3290286,7.548522,7.7920227,8.110974,8.4093485,8.436785,8.344186,7.4970784,6.7185616,6.392751,6.478491,7.7611566,8.999237,10.106995,10.864933,10.899229,10.5597,10.477389,10.497967,10.597425,10.878652,11.2421875,11.050131,10.275044,9.084977,7.8331776,6.694555,5.9469047,5.504488,5.429037,5.9469047,6.8454566,7.932636,9.287323,10.779194,12.082437,12.247057,12.010415,11.441104,10.676306,9.935514,9.527394,11.540562,14.147048,16.098484,16.756964,21.11597,23.1943,22.717587,21.517231,23.520111,23.821915,23.341772,20.687271,16.588915,13.910407,11.845795,12.874671,14.527733,16.101913,18.653526,22.18943,22.43979,22.823904,21.94936,13.615462,8.680285,6.7940125,7.016936,8.351046,9.705732,11.423956,12.46998,12.867812,12.912396,13.173045,15.426285,17.079346,17.69667,17.000465,14.843254,15.899568,15.789821,16.029892,17.29198,19.387459,15.021593,11.506266,10.6317215,12.823228,17.151367,17.03819,13.275933,9.383351,7.623973,8.992378,12.4802685,13.46799,13.5503,13.083877,11.204462,9.8429165,10.079557,9.822338,8.416207,6.6225333,5.751418,5.453044,5.5387836,5.768566,5.844017,5.5559316,5.271276,5.209543,5.3090014,5.188966,5.2815647,6.23499,7.0615206,7.226141,6.632822,6.697984,7.2947326,8.371623,9.657719,10.652299,11.050131,10.940384,10.861504,11.070708,11.543991,11.869802,11.077567,9.997248,9.541112,10.700313,12.075578,12.041282,11.794352,11.729189,11.427385,12.202472,12.833516,13.011855,12.871242,12.96727,13.004995,13.413116,14.270514,14.928994,14.023583,11.2421875,9.407358,7.953213,6.691125,5.830299,5.909179,5.394741,4.5510626,3.882293,4.1429415,4.2595477,3.8925817,3.4433057,3.0729103,2.6853669,2.7230926,3.350707,4.232111,5.0140567,5.3330083,5.07236,5.3878818,6.4990683,8.110974,9.431366,9.218731,8.018375,6.975781,6.5230756,6.3824625,6.186976,6.327589,6.5162163,6.5333643,6.23499,5.161529,3.9303071,2.9220085,2.270387,1.8588364,1.5947582,1.3615463,1.2758065,1.2620882,1.0666018,1.0597426,1.4610043,1.5913286,1.2517995,0.69963586,0.4115505,0.37039545,0.4698535,0.64476246,0.864256,1.0425946,1.1592005,1.2312219,1.2517995,1.2003556,1.2037852,1.2586586,1.3203912,1.4095604,1.611906,1.6393428,1.3889829,1.0563129,0.7682276,0.59674823,0.67219913,0.84367853,0.9328478,0.805953,0.4115505,0.24007112,0.17833854,0.2503599,0.39783216,0.490431,0.5212973,0.5178677,0.5624523,0.6756287,0.8196714,0.6790583,0.51100856,0.36010668,0.31209245,0.4938606,0.52472687,0.41840968,0.3841138,0.40126175,0.22978236,0.061732575,0.010288762,0.006859175,0.017147938,0.041155048,0.16119061,0.18519773,0.1371835,0.07545093,0.06859175,0.05144381,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.006859175,0.0034295875,0.017147938,0.044584636,0.06859175,0.08573969,0.08916927,0.07888051,0.061732575,0.034295876,0.024007112,0.041155048,0.061732575,0.07545093,0.07545093,0.07888051,0.08573969,0.08573969,0.07888051,0.09259886,0.09259886,0.106317215,0.11317638,0.11317638,0.14747226,0.21263443,0.24007112,0.29151493,0.36353627,0.40126175,0.21263443,0.17490897,0.22978236,0.33609957,0.4938606,0.41498008,0.45270553,0.66876954,0.96371406,1.1008976,1.2758065,1.7422304,1.8142518,1.4164196,1.0871792,1.2998136,1.2175035,1.1146159,1.1626302,1.4575747,1.6359133,1.6256244,1.4747226,1.2209331,0.86082643,0.5796003,0.40126175,0.28122616,0.22635277,0.2777966,0.40126175,0.48700142,0.5453044,0.5658819,0.51100856,0.65162164,0.9568549,1.2723769,1.4335675,1.2449403,1.0288762,0.91569984,0.8025235,0.6756287,0.59674823,0.53501564,0.51100856,0.51100856,0.5212973,0.53844523,0.5727411,0.5418748,0.48700142,0.42869842,0.37725464,0.432128,0.47671264,0.45270553,0.39440256,0.432128,0.548734,0.67219913,0.8745448,1.1214751,1.3032433,1.371835,1.5090185,1.5981878,1.5947582,1.5227368,1.9102802,2.2978237,2.5721905,2.9254382,3.8445675,4.273266,4.32471,4.2389703,4.2046742,4.3178506,4.8905916,4.99005,4.547633,3.549623,2.0234566,2.1400626,2.3252604,2.4624438,2.5173173,2.5070283,2.9117198,3.6696587,4.173808,4.297273,4.389872,4.5613513,4.9008803,5.099797,5.0586414,4.911169,5.1752477,5.4016004,5.504488,5.5147767,5.579939,6.684266,8.450503,11.22161,14.651197,17.720678,19.473198,20.083664,19.401176,17.652086,15.450292,12.524854,10.069269,8.045813,6.416758,5.120374,3.765687,2.5619018,1.7559488,1.4129901,1.4232788,1.4644338,1.2689474,1.0048691,0.78194594,0.64819205,0.8848336,1.1180456,1.3615463,1.646202,1.99602,2.4418662,2.767677,2.8808534,2.7882545,2.6064866,2.3664153,2.1229146,2.0063086,2.061182,2.2360911,2.644212,2.5824795,2.4007113,2.301253,2.3561265,2.5378947,3.2409601,4.6093655,6.3481665,7.7371492,8.285883,8.052671,7.1678376,5.9228973,4.7499785,3.7211025,2.9940298,2.335549,1.6187652,0.84024894,0.5521636,0.33609957,0.20234565,0.16119061,0.216064,0.29494452,0.3841138,0.4664239,0.490431,0.4081209,0.23664154,0.18862732,0.18519773,0.18862732,0.17833854,0.16462019,0.23321195,0.34638834,0.42526886,0.37039545,0.28122616,0.18862732,0.15776102,0.18862732,0.22292319,0.2777966,0.30866286,0.42869842,0.6379033,0.8128122,0.53501564,0.3806842,0.29837412,0.26064864,0.23664154,0.19891608,0.15776102,0.116605975,0.09259886,0.10288762,0.1920569,0.40126175,0.90884066,1.6770682,2.4795918,2.8019729,3.350707,3.9714622,4.4996185,4.756838,5.394741,5.830299,5.8988905,5.7891436,6.0566516,6.550512,6.8454566,7.14726,7.606825,8.296172,9.304471,9.945804,10.251037,10.096705,9.184435,8.831187,8.405919,7.9292064,7.466212,7.1198235,7.140401,7.6376915,7.6685576,7.099246,6.601956,6.3035817,5.9331865,5.7377,5.861165,6.355026,7.599966,8.8929205,10.244178,11.519984,12.415107,12.737488,12.686044,12.562579,12.624311,13.087306,14.119612,15.422854,16.427725,16.88729,16.856422,16.53747,16.88729,17.820137,19.095943,20.306587,21.047379,21.599543,22.306036,23.35206,24.76505,26.298077,27.947708,29.559614,31.078922,32.550213,33.469345,34.299305,34.99208,35.50309,35.808323,37.72203,40.15361,42.365692,43.799263,44.083916,42.588615,40.438267,38.74062,38.123295,38.74062,40.139893,39.433395,37.547123,35.32475,33.52765,30.804554,28.246082,25.968836,23.986534,22.20315,20.95135,20.12139,19.12681,17.785841,16.304258,14.627191,13.982429,13.570878,12.833516,11.430815,9.873782,8.639131,7.781734,7.267296,6.975781,6.9209075,7.0032177,7.349606,7.891481,8.364764,8.827758,8.512236,7.939495,7.257007,6.228131,6.279575,6.6876955,7.599966,8.718011,9.266746,9.609704,9.585697,9.318189,9.040393,9.108984,9.427936,9.263316,8.879202,8.450503,8.052671,7.4113383,6.835168,6.433906,6.368744,6.831738,7.4696417,8.347616,9.489669,10.645439,11.30049,11.153018,11.399949,11.633161,11.602294,11.218181,10.30591,11.838936,14.555169,17.353712,19.318867,24.230036,26.047716,24.209457,20.539799,19.267422,19.140528,20.138538,19.312008,16.088194,12.250486,10.14472,11.543991,14.109323,16.328266,17.54234,18.962189,22.182571,26.8571,29.127487,21.606401,15.954441,10.436234,6.64997,5.192395,5.6348124,7.1781263,8.584257,10.182446,12.044711,14.009865,17.401728,19.764713,20.742146,19.850452,16.492886,15.306249,14.71636,15.021593,15.827546,16.03675,14.263655,13.419975,14.153908,15.5085945,14.894698,12.891819,10.268185,7.750868,6.1561093,6.3618846,7.006647,7.7268605,8.89635,9.9869585,9.541112,8.261876,9.136421,9.654288,8.738589,6.7459984,6.245279,6.4716315,6.8728933,7.4181976,8.594546,8.995808,9.102125,9.818909,11.396519,13.426835,14.472859,13.111313,10.374502,7.4524937,5.703404,5.9160385,7.191845,7.723431,7.1987042,6.7802944,6.608815,6.5367937,6.708273,7.208993,8.083538,8.776315,8.844906,8.745448,9.067829,10.521975,12.699762,13.3033695,13.13532,12.857523,13.008426,14.102464,15.22051,15.690363,15.323397,14.4145565,13.323947,13.035862,13.581166,14.099034,12.833516,10.871792,9.499957,8.203573,6.883182,5.857735,6.0703697,5.6656785,5.0243454,4.5339146,4.5956473,4.3349986,3.9165888,3.5050385,3.1826572,2.9734523,3.0214665,3.3678548,3.9303071,4.5853586,5.195825,5.2815647,6.0154963,7.7131424,10.034973,12.000127,12.415107,11.729189,10.710602,9.921797,9.6988735,9.421077,9.489669,9.657719,9.685155,9.349055,8.244728,6.711703,5.0757895,3.6319332,2.6647894,2.0577524,1.5947582,1.4198492,1.4541451,1.3855534,1.5638919,1.8519772,1.786815,1.3478279,0.9602845,0.8505377,0.9877212,1.2312219,1.4918705,1.7182233,1.8554068,1.8931323,1.8931323,1.8691251,1.7902447,1.7319417,1.7422304,1.6256244,1.3958421,1.2620882,1.1934965,1.097468,0.939707,0.7407909,0.5761707,0.548734,0.64476246,0.89512235,1.1111864,0.864256,0.5144381,0.42869842,0.5727411,0.85739684,1.1489118,1.6736387,1.9274281,1.6736387,1.0563129,0.59674823,0.47328308,0.37039545,0.33952916,0.39783216,0.548734,0.607037,0.5693115,0.5796003,0.61046654,0.490431,0.26407823,0.14404267,0.082310095,0.044584636,0.034295876,0.20920484,0.32238123,0.29494452,0.17833854,0.15090185,0.17147937,0.17833854,0.14404267,0.07888051,0.048014224,0.034295876,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.010288762,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.030866288,0.07888051,0.13032432,0.13032432,0.11317638,0.106317215,0.09945804,0.0548734,0.034295876,0.037725464,0.048014224,0.048014224,0.041155048,0.024007112,0.037725464,0.058302987,0.07888051,0.08916927,0.058302987,0.072021335,0.10288762,0.1371835,0.15090185,0.19548649,0.2194936,0.19891608,0.14747226,0.12346515,0.12346515,0.13375391,0.15776102,0.19548649,0.2194936,0.22978236,0.33266997,0.51100856,0.7339317,0.9431366,0.85739684,0.8676856,0.9568549,0.9945804,0.71678376,0.64819205,0.78194594,0.9602845,1.0597426,0.9877212,0.7407909,0.6173257,0.5418748,0.4629943,0.37382504,0.34638834,0.31552204,0.274367,0.2469303,0.29837412,0.33952916,0.33952916,0.36696586,0.44584638,0.5418748,0.7339317,1.1043272,1.4095604,1.5364552,1.488441,1.2072148,1.0906088,1.0048691,0.89169276,0.764798,0.66191036,0.59331864,0.5590228,0.5590228,0.5624523,0.5418748,0.4698535,0.40126175,0.34981793,0.29151493,0.26407823,0.28122616,0.31209245,0.33952916,0.37382504,0.48700142,0.6173257,0.6790583,0.6756287,0.6927767,0.7305021,0.85396725,0.9945804,1.1317638,1.2895249,1.5981878,1.903421,2.2635276,2.9665933,4.513337,5.2472687,5.1752477,5.0174866,4.9180284,4.4447455,4.149801,3.981751,3.4638834,2.5413244,1.5604624,1.6016173,1.8348293,2.1434922,2.4007113,2.4555845,2.6236343,2.9220085,3.433017,4.029765,4.400161,4.852866,5.689686,6.1492505,6.012067,5.6313825,5.658819,6.029215,6.433906,6.6396813,6.492209,7.3564653,8.484799,10.034973,12.476839,16.585485,20.495214,22.412354,21.78474,19.11995,16.009314,13.783512,11.283342,8.786603,6.608815,5.1066556,3.642222,2.417859,1.6770682,1.3992717,1.2998136,1.155771,0.8196714,0.5555932,0.47671264,0.5212973,0.7922347,1.0185875,1.2860953,1.6599203,2.177788,2.620205,2.9048605,2.9906003,2.9082901,2.7573884,2.5207467,2.253239,2.0989075,2.1194851,2.2909644,2.760818,2.627064,2.277246,1.920569,1.5913286,2.5619018,3.782835,5.2506986,6.5333643,6.773435,6.4098988,5.576509,4.629943,3.7451096,2.9322972,2.218943,1.5981878,1.0597426,0.607037,0.2469303,0.16462019,0.10288762,0.07545093,0.09945804,0.18519773,0.3018037,0.432128,0.4355576,0.31895164,0.23664154,0.20234565,0.28122616,0.33952916,0.31209245,0.20234565,0.17147937,0.216064,0.31209245,0.42526886,0.5041494,0.38754338,0.20577525,0.12689474,0.17833854,0.2503599,0.35324752,0.34638834,0.32238123,0.32238123,0.32924038,0.24350071,0.216064,0.22978236,0.23664154,0.16462019,0.12689474,0.10288762,0.08916927,0.11317638,0.216064,0.41498008,0.7682276,1.3546871,2.1160555,2.8396983,2.8911421,3.3061223,3.8548563,4.3521466,4.6265135,5.0243454,5.305572,5.346727,5.411889,6.166398,7.1129646,7.5450926,7.8331776,8.193284,8.690575,9.369633,10.329918,11.194174,11.430815,10.367643,9.640571,9.023245,8.584257,8.2481575,7.7885933,7.7440085,8.532814,8.820899,8.31332,7.723431,7.0203657,6.615674,6.526505,6.759717,7.3255987,8.64256,10.220171,12.082437,13.838386,14.678635,14.925565,14.79867,14.723219,14.977009,15.71094,16.95931,17.988186,18.62609,18.818146,18.6158,18.62266,19.157675,20.344313,21.801888,22.662714,23.19087,23.69845,24.473536,25.553856,26.740494,28.17406,29.75853,31.33271,32.797146,34.141544,34.64912,35.14984,35.763737,36.706875,38.270767,41.007576,44.529762,47.424335,48.652126,47.53065,43.675797,40.167328,38.133583,38.06156,39.790073,40.462273,39.436825,36.92294,33.91519,32.18325,30.25925,28.633625,27.337242,26.256922,25.125158,24.500973,24.243753,23.85964,23.091412,21.911634,20.093952,18.735836,17.604073,16.283682,14.181344,12.151029,10.55284,9.496528,8.844906,8.196714,7.599966,7.023795,6.7185616,6.824879,7.346176,8.06296,8.707723,9.122703,8.961512,7.706283,6.420188,5.5730796,5.5593615,6.2692857,7.085528,8.169277,8.522525,8.450503,8.182996,7.9017696,7.970361,7.870903,7.7371492,7.6788464,7.805741,7.500508,7.140401,6.9826403,7.116394,7.466212,8.025234,8.858624,9.829198,10.624862,10.755186,9.513676,9.688584,10.63858,11.694893,12.168177,11.5645685,11.190743,12.373952,15.374841,19.387459,22.408924,23.098272,22.007662,19.665255,16.588915,15.611482,16.6335,17.171944,16.074476,13.533153,12.9981365,12.987847,13.588025,14.63062,15.690363,16.554619,18.924463,22.559826,25.845371,25.780209,24.411804,18.015623,10.858074,5.8988905,4.7979927,5.672538,7.0375133,8.875772,11.231899,14.198492,16.400288,17.339994,17.61436,17.353712,16.21852,15.96816,15.436573,15.151917,15.241087,15.412566,14.757515,15.086755,15.560039,14.664916,10.220171,7.610255,6.0052075,5.40503,5.689686,6.5950966,6.351596,6.012067,6.293293,7.4627824,9.328478,8.81747,9.050681,9.071259,8.237869,6.2212715,6.4716315,7.1712675,7.8263187,8.903209,11.828648,13.834956,15.011304,17.247395,21.393766,27.289227,29.806545,25.619019,18.588364,11.89038,8.025234,7.689135,9.277034,9.448513,7.6925645,6.3310184,5.3844523,4.7945633,4.506478,4.5201964,4.870014,5.7994323,6.3961806,7.0272245,7.829748,8.7145815,10.463672,11.893809,12.325937,11.934964,11.732618,11.924676,13.334236,14.565458,14.620332,12.871242,11.159878,11.005547,11.571428,11.910957,10.967821,9.870353,8.862054,7.805741,6.742569,5.895461,5.693115,5.470192,5.3227196,5.195825,4.866585,4.7191124,4.4756117,4.091498,3.7313912,3.7691166,3.99204,3.957744,4.0606318,4.396731,4.770556,5.2301207,6.1561093,7.8126,9.97324,11.914387,13.015285,12.6929035,11.71547,10.830637,10.7586155,10.357354,10.120712,10.038403,9.9801,9.6817255,9.0369625,7.949784,6.4133286,4.7088237,3.4055803,2.5378947,1.9823016,1.6427724,1.5090185,1.6804979,2.2463799,1.8897027,1.2895249,0.939707,1.1351935,1.6221949,2.0886188,2.469303,2.7470996,2.9494452,3.1860867,3.223812,3.0900583,2.9082901,2.8945718,2.9117198,2.74367,2.469303,2.2155135,2.1743584,2.1194851,2.1229146,2.061182,1.8416885,1.4164196,1.2517995,1.2037852,1.3752645,1.6427724,1.6290541,1.0151579,0.85739684,0.9431366,1.1660597,1.5090185,2.4898806,3.0111778,2.568761,1.5055889,1.0014396,0.805953,0.58988905,0.4698535,0.4698535,0.52472687,0.58988905,0.6036074,0.5693115,0.5453044,0.6241849,0.52815646,0.39097297,0.26750782,0.17147937,0.09602845,0.16462019,0.32924038,0.39097297,0.32924038,0.31895164,0.4046913,0.45270553,0.3841138,0.24007112,0.16462019,0.1097468,0.061732575,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.041155048,0.034295876,0.020577524,0.044584636,0.09602845,0.09602845,0.07888051,0.0548734,0.030866288,0.017147938,0.024007112,0.048014224,0.07545093,0.07545093,0.05144381,0.0548734,0.06859175,0.07545093,0.07545093,0.11317638,0.15776102,0.20234565,0.22635277,0.21263443,0.12689474,0.116605975,0.13375391,0.1371835,0.07545093,0.07545093,0.11317638,0.1920569,0.29151493,0.36696586,0.41498008,0.3806842,0.34981793,0.3566771,0.3806842,0.34638834,0.52815646,0.7339317,0.8025235,0.59674823,0.6927767,0.77165717,0.8093826,0.7682276,0.61046654,0.4389872,0.39783216,0.40126175,0.4115505,0.4115505,0.36353627,0.34981793,0.33952916,0.31209245,0.274367,0.274367,0.26407823,0.29151493,0.37039545,0.5041494,0.6001778,0.5796003,0.6241849,0.7579388,0.85396725,0.70649505,0.84367853,1.0288762,1.0837497,0.89855194,0.77851635,0.66533995,0.5796003,0.53844523,0.548734,0.548734,0.47671264,0.42869842,0.42526886,0.4115505,0.32581082,0.39783216,0.4938606,0.53158605,0.45613512,0.5418748,0.6001778,0.5693115,0.51100856,0.59674823,0.6927767,0.72707254,0.72021335,0.7305021,0.84024894,1.2037852,1.2963841,1.4267083,1.8142518,2.609916,4.4756117,5.895461,6.591667,6.228131,4.4104495,3.1277838,2.952875,2.7402403,2.1332035,1.5707511,1.3409687,1.4095604,1.5947582,1.786815,1.9685832,2.1160555,2.527606,3.2889743,4.1429415,4.4859004,4.938606,5.6005163,6.0326443,6.1561093,6.2418494,6.4236174,7.3839016,8.31332,8.711152,8.405919,9.712592,10.9369545,11.976119,12.874671,13.838386,15.707511,18.499195,19.672113,18.608942,16.6335,13.505715,11.537132,9.674867,7.3255987,4.3487167,3.0317552,2.1160555,1.6084765,1.3238207,0.8848336,0.6036074,0.4972902,0.48014224,0.4972902,0.53501564,0.66876954,0.82996017,1.214074,1.9342873,3.0214665,3.1312134,3.0660512,2.8396983,2.5481834,2.3664153,1.9754424,1.4095604,1.0323058,0.9259886,0.90198153,0.99801,1.1214751,1.3478279,1.704505,2.1674993,3.350707,4.32471,5.0929375,5.442755,4.928317,4.280125,3.525616,2.8911421,2.3835633,1.786815,1.0906088,0.65162164,0.36353627,0.17490897,0.07545093,0.05144381,0.0274367,0.01371835,0.041155048,0.1371835,0.22292319,0.31895164,0.31209245,0.22635277,0.21263443,0.28808534,0.69963586,0.9431366,0.77508676,0.21263443,0.16462019,0.15090185,0.17147937,0.23664154,0.3806842,0.3806842,0.29151493,0.20920484,0.18862732,0.21263443,0.33609957,0.34638834,0.32924038,0.31895164,0.30523327,0.2194936,0.17147937,0.15776102,0.17833854,0.21263443,0.17833854,0.12346515,0.13375391,0.24007112,0.4115505,0.66876954,1.1900668,1.6427724,1.8725548,1.9239986,2.287535,2.7642474,3.3747141,4.040054,4.5784993,4.955754,5.2335505,5.312431,5.302142,5.5079174,6.0326443,7.2638664,8.556821,9.582268,10.316199,9.849775,9.846346,10.131001,10.39165,10.1481495,9.6817255,9.119273,8.611694,8.2653055,8.117833,8.141841,8.1487,8.258447,8.457363,8.591117,7.7611566,7.654839,8.032094,8.597976,8.988949,10.2921915,12.092726,14.352823,16.448301,17.182234,16.70552,16.156786,16.21166,17.065628,18.434032,19.263992,19.716698,19.881319,19.884748,19.898466,20.567236,21.650986,23.201159,24.665592,24.871368,24.43238,24.816494,25.61559,26.630747,27.861969,29.950588,31.634514,32.927467,33.798584,34.16555,34.556522,35.057243,36.06211,37.807774,40.359386,43.398,46.21712,47.928486,48.165127,47.105385,43.600346,41.827248,41.429417,42.283382,44.47832,44.516045,43.41858,40.884113,37.468243,34.577103,32.330723,31.34643,30.749681,30.09463,29.374416,28.59247,28.441568,28.479294,28.112328,26.610168,24.987974,23.11542,20.779871,18.135658,15.731518,13.694343,12.003556,10.659158,9.613133,8.759167,7.9292064,6.8866115,5.977771,5.610805,6.2727156,7.222711,7.9909387,8.158989,7.716572,7.0958166,6.5230756,6.358455,5.9743414,5.2438393,4.547633,5.950334,6.7219915,7.06495,7.0718093,6.728851,6.728851,6.8111606,7.0375133,7.3290286,7.4765005,7.466212,7.140401,7.006647,7.208993,7.5382333,7.7097125,8.100685,8.532814,8.862054,8.971801,8.436785,8.090397,8.632272,10.017825,11.458252,12.154458,10.882081,10.569988,12.123591,14.421415,17.264544,19.558937,20.598103,19.54179,15.443433,15.820687,16.657507,17.559488,18.331144,18.965618,20.344313,21.37662,21.273731,20.53637,20.965069,18.986197,18.20082,18.28656,18.70154,18.677534,18.811287,17.727537,14.112752,9.2153015,6.835168,5.895461,6.660259,9.043822,12.747777,17.226818,20.755863,18.752985,15.097044,12.346515,11.749766,12.603734,13.577737,14.308239,14.483148,13.824667,13.629181,13.810948,12.758065,10.624862,9.294182,9.23245,8.327039,7.706283,8.217292,10.4533825,8.656279,7.174697,6.90033,8.755736,13.687484,17.04505,17.514904,14.445422,9.39707,6.1492505,6.9552035,7.596536,8.261876,9.325048,11.351934,15.1862135,18.972477,24.061985,31.034336,39.700905,42.033024,37.471672,29.144634,20.049368,13.029003,10.6145735,10.39508,10.63858,10.566559,10.360784,7.723431,5.8371577,4.8185706,4.417309,4.029765,4.029765,4.650521,5.4153185,6.042933,6.468202,7.301592,7.781734,8.31332,8.988949,9.599416,9.962952,10.487679,11.067279,11.286773,10.405369,10.237319,10.247607,10.590566,10.786053,9.736599,8.244728,7.9737906,7.9429245,7.6651278,7.140401,6.420188,6.111525,6.307011,6.5162163,5.662249,5.1100855,5.038064,5.0277753,5.0757895,5.6005163,6.6739774,6.48535,5.967482,5.610805,5.4770513,6.0635104,7.298162,8.824328,10.511685,12.452832,12.634601,11.818358,10.401938,8.889491,7.888051,7.6925645,7.689135,7.6959944,7.534804,7.034084,6.680836,6.0326443,5.06893,4.0023284,3.2958336,2.6716487,2.253239,1.8142518,1.546744,2.061182,3.7691166,3.0523329,2.1057668,2.0131679,2.7470996,3.4295874,3.8479972,4.1155047,4.341858,4.623084,5.453044,5.8543057,5.4084597,4.5442033,4.530485,5.336438,5.055212,4.5099077,4.125794,3.9063,3.391862,3.3472774,3.7691166,4.1017866,3.234101,2.9048605,2.9220085,2.843128,2.568761,2.3492675,1.8245405,1.4747226,1.2483698,1.08032,0.8848336,0.86082643,0.9568549,1.1694894,1.3786942,1.3443983,1.1489118,0.9259886,0.83338976,0.8162418,0.61046654,0.4389872,0.38754338,0.40126175,0.4389872,0.48700142,0.59674823,0.5796003,0.51100856,0.45270553,0.42869842,0.31895164,0.22635277,0.28808534,0.48014224,0.6241849,0.7099246,0.6790583,0.58645946,0.4698535,0.33609957,0.21263443,0.12003556,0.05144381,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.006859175,0.020577524,0.06859175,0.09602845,0.08573969,0.06859175,0.09259886,0.1097468,0.072021335,0.08916927,0.17833854,0.2469303,0.14404267,0.106317215,0.1097468,0.14061308,0.19891608,0.16804978,0.1371835,0.15090185,0.20234565,0.2503599,0.26407823,0.26064864,0.22978236,0.17147937,0.09945804,0.09945804,0.28465575,0.48014224,0.5178677,0.2194936,0.36696586,0.490431,0.44927597,0.30523327,0.31895164,0.3806842,0.5007198,0.6310441,0.72364295,0.7407909,0.65505123,0.61389613,0.58302987,0.52472687,0.41498008,0.4389872,0.47328308,0.4424168,0.3566771,0.32581082,0.29837412,0.33266997,0.34638834,0.31209245,0.28808534,0.33609957,0.37382504,0.41840968,0.45613512,0.45613512,0.4629943,0.44927597,0.45270553,0.4938606,0.5624523,0.5796003,0.607037,0.6241849,0.6173257,0.5693115,0.4972902,0.50757897,0.5521636,0.5658819,0.45270553,0.40126175,0.37725464,0.34638834,0.33266997,0.38754338,0.4664239,0.5521636,0.5590228,0.48357183,0.37382504,0.50757897,0.5418748,0.5041494,0.45956472,0.4972902,0.64476246,0.77165717,0.6893471,0.5144381,0.64476246,0.980862,1.1523414,1.3169615,1.5536032,1.8759843,2.3286898,4.016047,6.0806584,6.842027,3.8102717,2.510458,2.1126258,1.9068506,1.6187652,1.3889829,1.3238207,1.5433143,1.7079345,1.6839274,1.5638919,1.7902447,2.3252604,3.0866287,3.8548563,4.266407,4.3658648,4.4516044,4.8494368,5.504488,5.960623,6.4064693,7.98408,9.72631,11.14273,12.202472,12.9638405,14.438563,16.345413,17.923023,17.940172,18.608942,19.658396,20.141968,19.524641,17.693241,14.579176,11.327928,8.31332,5.6828265,3.3609958,2.1983654,1.430138,1.0082988,0.7888051,0.5418748,0.41840968,0.3806842,0.48357183,0.67219913,0.77851635,0.84367853,1.097468,1.4781522,1.9480057,2.4967396,2.7128036,2.6853669,2.428148,1.99602,1.4610043,1.0631721,0.7579388,0.77851635,1.0940384,1.4129901,1.704505,1.4472859,1.3272504,1.670209,2.4487255,3.083199,3.6079261,4.0057583,4.0949273,3.5118976,2.9048605,2.2738166,1.704505,1.214074,0.77165717,0.4081209,0.2194936,0.12003556,0.058302987,0.041155048,0.024007112,0.017147938,0.01371835,0.041155048,0.1371835,0.24350071,0.3566771,0.3841138,0.32924038,0.29837412,0.28465575,0.4972902,0.70306545,0.7922347,0.7888051,0.4664239,0.26064864,0.17490897,0.23321195,0.4664239,0.50757897,0.34295875,0.2194936,0.20577525,0.20234565,0.23664154,0.2777966,0.31209245,0.33609957,0.34295875,0.22635277,0.14061308,0.08916927,0.08916927,0.16462019,0.19548649,0.17490897,0.216064,0.37382504,0.6310441,1.0631721,1.4987297,1.978872,2.5481834,3.2409601,4.8082814,5.802862,6.0497923,5.645101,4.979761,4.695105,4.8494368,4.9694724,5.079219,5.717122,7.4113383,8.255017,8.742019,9.174147,9.644,10.1652975,10.868362,11.72233,12.4974165,12.771784,12.277924,11.019264,10.278474,10.264755,10.106995,9.280463,8.879202,8.683716,8.567109,8.457363,7.829748,7.5279446,7.613684,8.203573,9.462232,11.423956,13.972139,16.510035,18.530062,19.634388,19.082224,18.437462,18.28313,19.03764,20.971928,21.44178,21.740154,22.059107,22.467228,22.889067,23.413794,23.955667,24.391226,24.60729,24.480396,24.168303,24.936531,26.366669,28.27352,30.718815,33.078373,34.817173,35.602547,35.42078,34.556522,33.82259,33.565372,34.41248,36.429077,39.128162,42.626343,44.64294,45.568928,45.610085,44.821278,43.847275,43.56262,44.09078,44.97218,45.188244,44.197094,42.221653,39.258488,35.705437,32.34444,29.988314,28.283808,26.918833,25.76992,24.891945,24.326063,24.068846,24.096281,24.127148,23.633287,22.799898,21.53781,20.073376,18.588364,17.20967,16.029892,15.086755,14.160767,12.9707,11.187314,9.791472,8.639131,7.953213,7.6342616,7.2604365,7.0203657,7.205563,7.3530354,7.3427467,7.4113383,8.244728,7.689135,6.3790326,5.0312047,4.413879,4.5682106,4.756838,5.086078,5.597087,6.2418494,6.776865,6.6122446,6.4544835,6.540223,6.660259,6.4133286,6.0875177,5.8337283,5.7651367,5.9880595,6.355026,6.8728933,7.5862474,8.440215,9.301042,9.897789,10.082987,10.683165,11.869802,13.193623,13.574307,12.665466,11.561139,11.170166,12.185325,13.38911,14.599753,15.927004,16.582056,14.891269,13.025573,11.4033785,10.275044,9.860064,10.350495,15.175924,17.113642,17.165085,17.04162,19.157675,17.267973,14.562028,12.6757555,12.466551,14.013294,16.324837,15.46401,14.057879,13.481709,13.855534,11.156448,10.388221,11.146159,13.029003,15.666355,17.072487,16.643787,14.30481,11.609154,11.7257595,13.584596,12.596875,10.854645,9.373062,8.086967,8.069819,9.22902,10.878652,12.188754,12.185325,10.14129,7.0443726,5.2438393,5.8234396,8.584257,11.653738,10.618003,8.460793,6.824879,5.98463,7.1541195,7.9737906,8.272165,8.255017,8.491658,9.249598,10.069269,13.1593275,19.092514,26.781649,35.643703,36.871494,37.59171,40.962994,46.172535,38.994408,34.4845,32.622234,31.490473,27.261791,22.676432,17.844143,14.661487,12.874671,10.079557,5.7822843,3.6936657,2.7916842,2.4830213,2.5996273,2.726522,3.3952916,4.4516044,5.363875,5.223262,5.878313,6.9620624,8.567109,10.377932,11.660598,12.308789,14.668345,16.63007,17.096493,15.971589,17.782412,17.991615,16.6335,14.092175,11.091286,9.493098,9.239308,9.554831,9.770895,9.314759,7.949784,7.164408,6.725421,6.40304,5.977771,5.576509,5.5833683,5.936616,6.5196457,7.160979,7.953213,8.512236,8.488229,8.001227,7.6514096,7.795452,8.2481575,8.580828,8.553391,8.131552,7.9909387,7.6171136,7.0546613,6.5882373,6.728851,7.0135064,7.291303,7.2604365,6.81802,6.046363,4.9008803,4.3933015,4.057202,3.690236,3.333559,3.6765177,3.6936657,3.2032347,2.4727325,2.2429502,3.0454736,4.1292233,5.15467,6.0154963,6.835168,7.2947326,7.64798,8.220721,9.239308,10.847785,9.901219,8.64942,7.164408,5.6965446,4.6779575,4.2252517,3.9611735,3.5770597,3.0317552,2.5893385,2.301253,2.4212887,2.7093742,2.8945718,2.6750782,3.0077481,3.1346428,2.8054025,2.2360911,2.1057668,1.8725548,1.5536032,1.4027013,1.4164196,1.2998136,0.83681935,0.7613684,0.8196714,0.805953,0.5727411,0.64133286,0.6893471,0.6962063,0.64819205,0.53844523,0.5041494,0.5727411,0.75450927,0.9534253,0.96371406,0.4115505,0.18862732,0.13032432,0.14404267,0.20920484,0.33266997,0.45956472,0.61046654,0.7510797,0.8093826,0.7956643,0.71678376,0.58988905,0.44584638,0.31209245,0.18862732,0.116605975,0.06516216,0.020577524,0.0,0.010288762,0.020577524,0.037725464,0.0548734,0.037725464,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.010288762,0.010288762,0.006859175,0.0034295875,0.010288762,0.010288762,0.010288762,0.01371835,0.020577524,0.024007112,0.044584636,0.116605975,0.16462019,0.15090185,0.07888051,0.08916927,0.06516216,0.07545093,0.13375391,0.18862732,0.14747226,0.1097468,0.09602845,0.12689474,0.20234565,0.21263443,0.17147937,0.14404267,0.16119061,0.22292319,0.20920484,0.19548649,0.216064,0.25378948,0.25378948,0.26750782,0.36010668,0.4355576,0.42526886,0.274367,0.41498008,0.45613512,0.36353627,0.22635277,0.23321195,0.26750782,0.30866286,0.36696586,0.42869842,0.45613512,0.39097297,0.3806842,0.37382504,0.34981793,0.3018037,0.39097297,0.42183927,0.39097297,0.34295875,0.38754338,0.4424168,0.51100856,0.44927597,0.30523327,0.31895164,0.4355576,0.39783216,0.33952916,0.30866286,0.28808534,0.4355576,0.47328308,0.432128,0.39783216,0.52472687,0.5555932,0.50757897,0.490431,0.5418748,0.6173257,0.67219913,0.59331864,0.53844523,0.5453044,0.53844523,0.5212973,0.4938606,0.4424168,0.4081209,0.48357183,0.48700142,0.44584638,0.39783216,0.36696586,0.34295875,0.4081209,0.4081209,0.37382504,0.32581082,0.29837412,0.4355576,0.5624523,0.58302987,0.53501564,0.6036074,0.82996017,1.0906088,1.1763484,1.1351935,1.2620882,1.6530612,2.620205,4.033195,5.223262,4.99005,3.7142432,2.7642474,2.0097382,1.5501735,1.728512,1.99602,2.2909644,2.4315774,2.4315774,2.5001693,3.0214665,3.3884325,3.8308492,4.4516044,5.209543,4.98662,4.698535,4.681387,5.0929375,5.8988905,6.852316,8.416207,10.048691,11.533703,12.9981365,14.661487,16.077906,17.343424,18.156237,17.851004,18.756414,19.665255,19.850452,18.752985,15.999025,12.55915,10.1481495,7.956643,5.689686,3.542764,2.0817597,1.2483698,0.84024894,0.6824879,0.6036074,0.5624523,0.58645946,0.77165717,1.0185875,1.0323058,0.96371406,1.2449403,1.6496316,2.0440342,2.4007113,2.2498093,2.1126258,1.9480057,1.6221949,0.9259886,0.58645946,0.4424168,0.53158605,0.78537554,1.0288762,1.2380811,1.1866373,1.313532,1.8108221,2.627064,3.07634,3.2855449,3.2958336,3.0797696,2.5619018,1.978872,1.3649758,0.8676856,0.52472687,0.26407823,0.11317638,0.058302987,0.037725464,0.020577524,0.01371835,0.01371835,0.048014224,0.1097468,0.18862732,0.26407823,0.274367,0.23321195,0.22978236,0.28122616,0.34638834,0.4424168,0.53501564,0.6036074,0.6379033,0.65505123,0.4355576,0.2777966,0.17833854,0.15433143,0.2503599,0.2709374,0.20920484,0.16462019,0.17147937,0.18862732,0.20920484,0.23664154,0.26064864,0.2777966,0.30523327,0.2709374,0.22978236,0.1920569,0.16804978,0.17833854,0.19891608,0.24350071,0.36010668,0.58645946,0.9328478,1.5501735,2.1332035,2.7402403,3.4055803,4.15666,4.756838,4.979761,4.897451,4.5784993,4.0846386,4.1155047,5.0655007,6.183546,7.226141,8.440215,10.151579,10.624862,10.535692,10.456812,10.858074,11.489118,12.144169,12.932974,13.718349,14.140189,13.728639,11.543991,9.897789,9.534253,9.626852,9.040393,8.724871,8.601405,8.673427,9.043822,9.102125,9.290752,9.702303,10.439664,11.622872,13.272504,15.659496,17.902447,19.555508,20.594673,20.7833,21.04052,21.578964,22.710728,24.837072,25.420103,25.413242,24.957108,24.250612,23.554407,22.906214,22.913074,23.180582,23.568125,24.171732,25.138876,26.486704,28.030018,29.51503,30.626217,31.84029,32.91032,33.061222,32.32043,31.521338,31.181808,31.277838,32.1078,33.695698,35.804893,38.627445,40.596027,41.9953,43.055042,43.939873,44.704674,45.349434,46.011345,46.45719,46.086796,44.756115,42.420567,39.16589,35.08125,30.255821,26.966846,24.555847,23.146286,22.470657,21.877338,21.572105,21.623549,22.093403,22.727877,22.961088,22.36434,21.712719,21.009653,20.189981,19.133669,18.434032,17.799559,17.034761,16.009314,14.661487,13.399398,12.0138445,10.950673,10.240748,9.513676,8.98209,8.663138,8.3922,8.179566,8.186425,8.652849,8.114404,6.9209075,5.5662203,4.681387,4.07435,4.0777793,4.5099077,5.2026844,5.9914894,6.5950966,6.475061,6.138962,5.9228973,5.9880595,5.9400454,5.909179,6.0326443,6.310441,6.615674,7.010077,7.500508,7.9429245,8.31332,8.724871,10.213311,11.341646,12.524854,13.773223,14.71636,14.860402,14.311668,13.066729,11.646879,11.094715,10.878652,10.978109,11.80121,13.066729,13.810948,12.950122,11.660598,10.155008,9.273604,10.463672,13.011855,13.516005,13.149038,13.166186,14.908417,15.837835,14.428274,12.319078,10.484249,9.23245,11.149589,12.000127,13.279363,14.96329,15.4914465,13.841815,13.351384,13.375391,13.704632,14.586036,15.385129,14.188204,11.852654,9.856634,10.281903,10.81006,10.131001,9.414218,9.084977,8.831187,8.745448,8.98209,9.613133,10.288762,10.244178,8.841476,7.764586,7.133542,6.8900414,6.773435,8.179566,7.5553813,6.4887795,5.6965446,5.0483527,5.1512403,5.3673043,6.029215,7.0615206,7.98065,8.498518,9.201583,11.393089,15.46401,20.879328,26.167753,27.60818,28.19121,28.966295,29.041746,23.218307,20.745575,20.186552,19.94305,18.252264,18.310568,17.312557,16.777542,16.571766,14.88098,11.252477,8.388771,5.6005163,3.2032347,2.5173173,2.603057,3.275256,4.355576,5.5387836,6.4236174,7.846896,10.419086,13.749216,16.149927,14.668345,12.88839,12.517994,13.245067,13.999576,12.932974,12.758065,12.823228,12.397959,11.4205265,10.477389,9.997248,9.9869585,10.196163,10.377932,10.295622,9.640571,9.098696,8.683716,8.333898,7.9086285,7.3050213,6.9826403,7.1095347,7.682276,8.515666,8.779744,8.800322,8.416207,7.8263187,7.5725293,7.490219,7.613684,7.689135,7.500508,6.8763227,6.444195,6.0875177,5.7754254,5.597087,5.761707,6.0703697,6.2247014,6.0395036,5.518206,4.835718,4.0366244,3.8308492,3.858286,3.9063,3.9097297,4.046913,4.2183924,4.2218223,4.1120753,4.2115335,4.9523244,6.0806584,7.2295704,8.275595,9.321619,10.576848,12.308789,13.059869,12.569438,11.763485,10.285333,8.872343,7.798882,7.205563,7.0752387,6.5710897,6.5470824,7.0135064,7.7542973,8.299602,8.639131,8.169277,7.675417,7.4627824,7.366754,6.914048,6.341307,5.7274113,5.2301207,5.0757895,4.7534084,4.40702,4.417309,4.7842746,5.1100855,4.787704,3.7485392,2.9700227,2.7299516,2.633923,1.7490896,1.1489118,0.7956643,0.61046654,0.47328308,0.42869842,0.48014224,0.65505123,0.84367853,0.7990939,0.33609957,0.13375391,0.09945804,0.16462019,0.2709374,0.52815646,0.70649505,0.805953,0.84024894,0.85396725,0.8471081,0.85739684,0.7682276,0.6036074,0.50757897,0.4938606,0.4664239,0.47328308,0.5624523,0.77851635,0.61389613,0.48357183,0.36696586,0.25378948,0.15433143,0.10288762,0.06516216,0.034295876,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.010288762,0.01371835,0.010288762,0.010288762,0.020577524,0.017147938,0.010288762,0.01371835,0.024007112,0.017147938,0.037725464,0.15090185,0.2709374,0.31209245,0.19548649,0.10288762,0.061732575,0.061732575,0.082310095,0.1097468,0.11317638,0.08573969,0.07545093,0.10288762,0.16462019,0.23664154,0.274367,0.26064864,0.22635277,0.22292319,0.16804978,0.18519773,0.26407823,0.33609957,0.29494452,0.3018037,0.29494452,0.26750782,0.23664154,0.23664154,0.32581082,0.29837412,0.2194936,0.16119061,0.16462019,0.17490897,0.17490897,0.17833854,0.1920569,0.19548649,0.1920569,0.22635277,0.26407823,0.274367,0.25378948,0.28122616,0.2777966,0.26407823,0.26750782,0.33266997,0.4081209,0.45270553,0.37039545,0.24007112,0.31209245,0.45613512,0.4424168,0.36010668,0.2777966,0.25721905,0.41840968,0.4698535,0.4424168,0.42526886,0.5555932,0.5624523,0.5178677,0.53158605,0.6241849,0.7373613,0.8196714,0.6790583,0.5761707,0.59674823,0.64819205,0.5727411,0.5453044,0.5178677,0.4938606,0.51100856,0.4698535,0.39783216,0.36010668,0.3566771,0.34638834,0.30523327,0.28122616,0.25378948,0.2194936,0.17833854,0.26407823,0.37039545,0.4629943,0.5178677,0.48700142,0.65162164,0.9294182,1.0117283,0.91912943,1.0014396,1.4027013,1.6599203,2.2086544,3.2478194,4.7534084,4.2595477,3.6285036,2.9494452,2.4555845,2.5138876,2.6956558,2.8465576,2.8465576,2.8499873,3.275256,4.2081037,4.40702,4.5647807,5.07236,6.0154963,5.7308407,5.4976287,5.456474,5.73427,6.4407654,7.3118806,8.299602,9.482809,10.837497,12.247057,14.140189,15.004445,15.29939,15.237658,14.805529,15.645778,16.715809,17.528622,17.192522,14.417986,11.393089,9.595985,8.042382,6.2727156,4.3624353,2.5653315,1.6187652,1.196926,1.0906088,1.2072148,1.2792361,1.3341095,1.371835,1.371835,1.2758065,1.2998136,1.8416885,2.287535,2.428148,2.4624438,2.2806756,1.9857311,1.6324836,1.2072148,0.58988905,0.38754338,0.36010668,0.44927597,0.59674823,0.7305021,0.86082643,1.0460242,1.3924125,1.9171394,2.5619018,2.7128036,2.6064866,2.301253,1.9274281,1.6770682,1.2380811,0.70306545,0.33266997,0.17490897,0.061732575,0.024007112,0.024007112,0.030866288,0.034295876,0.030866288,0.034295876,0.07888051,0.17490897,0.29494452,0.34638834,0.28465575,0.13032432,0.1097468,0.2469303,0.36696586,0.51100856,0.5555932,0.5555932,0.52815646,0.47328308,0.39783216,0.36353627,0.25721905,0.11317638,0.09602845,0.09259886,0.116605975,0.1371835,0.15090185,0.18176813,0.45270553,0.36010668,0.2469303,0.24350071,0.2503599,0.2503599,0.23321195,0.216064,0.20920484,0.216064,0.25721905,0.3566771,0.5796003,0.9534253,1.4541451,2.1812177,2.8294096,3.4021509,3.899441,4.314421,4.396731,4.417309,4.341858,4.2183924,4.166949,4.6265135,6.3893213,8.416207,10.168727,11.64345,12.205902,12.157887,11.910957,11.7257595,11.712041,11.880091,12.085866,12.367092,12.730629,13.173045,13.38568,11.893809,10.48082,9.839486,9.595985,9.054111,8.673427,8.584257,8.800322,9.2153015,9.410788,9.654288,10.618003,12.295071,14.009865,15.525743,17.521763,19.394318,20.879328,22.041958,22.741594,23.76704,25.324074,27.227495,28.907993,29.01431,27.865398,25.985985,23.907654,22.148275,21.506943,21.60983,22.144846,22.971376,24.123718,26.00999,27.663052,28.637054,28.709076,27.868828,27.248072,27.292658,27.162333,26.747353,26.68219,27.01829,27.546446,28.386696,29.703657,31.692818,34.127827,36.49424,38.675457,40.620033,42.341686,43.446014,44.64294,45.71297,46.49835,46.88246,44.824707,41.840965,38.116436,33.75743,28.784527,25.210897,22.563255,21.215427,20.86218,20.52951,20.382038,20.807306,21.644127,22.566685,23.053686,22.429502,21.915064,21.414345,20.697561,19.390888,18.245405,17.051908,16.095055,15.350834,14.466,13.231348,11.928105,10.861504,10.151579,9.719451,9.469091,9.129561,8.611694,8.035523,7.716572,7.6685576,7.4970784,6.8385973,5.754848,4.7431192,3.9646032,3.875434,4.2218223,4.8185706,5.545643,6.2041235,6.4887795,6.4579134,6.245279,6.0497923,5.888602,6.1492505,6.5642304,6.914048,7.051232,7.1884155,7.613684,8.1041155,8.512236,8.742019,10.419086,12.010415,13.371962,14.38369,14.935853,14.946142,14.476289,13.3033695,11.633161,10.076128,8.762596,8.179566,8.64599,10.048691,11.859513,12.253916,12.003556,11.122152,10.412228,11.47197,11.97269,11.897239,11.509696,11.1393,11.173596,13.368532,13.433694,12.13731,10.0041065,7.346176,7.8434668,8.971801,10.710602,12.432255,12.915827,13.090735,13.402828,13.409687,13.035862,12.593445,13.989287,13.783512,12.703192,11.784062,12.349944,12.538571,12.38424,12.147599,12.291641,13.4645605,14.369971,13.965281,12.932974,12.394529,13.886399,12.243628,10.432805,10.131001,10.55284,8.47451,6.461343,6.077229,6.3138704,6.464772,6.1286726,5.6313825,5.5387836,6.0326443,6.975781,7.9257765,8.032094,8.107545,8.992378,10.909517,13.481709,14.500296,15.268523,15.501736,14.733508,12.30536,9.949233,9.235879,9.253027,9.623423,10.508256,13.841815,16.160215,16.897577,16.249386,15.169065,13.5503,11.266195,8.182996,5.0346346,3.391862,3.1346428,3.3952916,4.139512,5.254128,6.5539417,8.868914,12.250486,15.251375,16.187653,13.128461,10.830637,8.848335,8.049242,8.038953,7.2021337,6.1149545,6.2384195,6.5127864,6.677407,7.274155,7.7577267,8.124693,8.4093485,8.656279,8.916927,9.136421,9.167287,9.126132,9.057541,8.937505,8.553391,8.244728,8.169277,8.412778,9.002667,9.033533,8.429926,7.671987,7.116394,6.992929,6.6568294,6.540223,6.5162163,6.416758,6.0223556,5.638242,5.4187484,5.3261495,5.295283,5.223262,5.3570156,5.305572,5.0277753,4.5853586,4.1463714,3.799983,3.7485392,3.8891523,4.125794,4.372724,4.4687524,4.6436615,4.9831905,5.576509,6.5230756,7.720001,8.604835,9.373062,10.1481495,10.964391,12.027563,13.677195,14.270514,13.279363,11.314209,10.024684,9.119273,8.81747,9.040393,9.427936,9.290752,9.544542,10.545981,11.910957,12.517994,12.915827,12.915827,12.415107,11.495977,10.412228,9.482809,8.687145,8.2310095,8.06639,7.8949103,7.208993,6.742569,6.543653,6.543653,6.5539417,5.960623,4.7979927,4.0503426,3.9543142,3.9886103,2.7779658,1.7971039,1.1077567,0.6927767,0.45613512,0.3566771,0.32924038,0.3841138,0.45613512,0.40126175,0.23321195,0.216064,0.29494452,0.40126175,0.44927597,0.7888051,0.9945804,1.0940384,1.1489118,1.2758065,1.7113642,2.0817597,1.9548649,1.4267083,1.1283343,1.1420527,1.138623,1.1694894,1.255229,1.371835,1.0220171,0.78537554,0.58988905,0.4081209,0.26407823,0.18519773,0.11317638,0.0548734,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.006859175,0.006859175,0.01371835,0.017147938,0.0274367,0.017147938,0.006859175,0.006859175,0.01371835,0.0034295875,0.048014224,0.16119061,0.3018037,0.40126175,0.34638834,0.16119061,0.08916927,0.072021335,0.07888051,0.08573969,0.07545093,0.07545093,0.08573969,0.106317215,0.14061308,0.23321195,0.34638834,0.3841138,0.33266997,0.26407823,0.2194936,0.28122616,0.35324752,0.35324752,0.20920484,0.18519773,0.16119061,0.13032432,0.10288762,0.09259886,0.12346515,0.12003556,0.12003556,0.13375391,0.14404267,0.16119061,0.15090185,0.12346515,0.10288762,0.116605975,0.14404267,0.18862732,0.2469303,0.2777966,0.22978236,0.16462019,0.13032432,0.13032432,0.14747226,0.15776102,0.17147937,0.16462019,0.15090185,0.17490897,0.30866286,0.3806842,0.44927597,0.4389872,0.36696586,0.33266997,0.37039545,0.432128,0.48014224,0.51100856,0.5521636,0.53844523,0.5453044,0.58988905,0.65162164,0.6859175,0.7099246,0.64819205,0.61389613,0.6344737,0.65162164,0.5144381,0.490431,0.5007198,0.490431,0.4389872,0.432128,0.4389872,0.42869842,0.39440256,0.34638834,0.2469303,0.20920484,0.1920569,0.18176813,0.17490897,0.20234565,0.29494452,0.38754338,0.4115505,0.31552204,0.48014224,0.6893471,0.82996017,0.8848336,0.9568549,1.0837497,1.1249046,1.3992717,2.0303159,2.942586,3.5702004,3.9851806,4.081209,3.841138,3.3266997,3.07634,2.9460156,2.7230926,2.644212,3.391862,4.619654,4.863155,4.972902,5.3981705,6.1904054,6.3001523,6.3961806,6.5950966,6.917478,7.281014,7.671987,8.028665,8.7145815,9.791472,11.022695,12.308789,12.325937,11.8869505,11.393089,10.847785,10.995257,11.945253,13.711491,15.073037,13.605173,11.8115,9.952662,8.443645,7.233,5.813151,3.9131594,2.6750782,1.9411465,1.6496316,1.845118,2.037175,2.1057668,1.9308578,1.6324836,1.5810398,1.8348293,2.551613,2.8637056,2.5824795,2.2120838,2.4418662,2.0440342,1.3512574,0.6824879,0.32581082,0.30866286,0.39783216,0.5590228,0.7407909,0.8711152,0.99801,1.2209331,1.5158776,1.845118,2.1469216,1.845118,1.471293,1.0425946,0.71678376,0.7579388,0.5624523,0.2503599,0.058302987,0.030866288,0.01371835,0.01371835,0.024007112,0.041155048,0.061732575,0.07545093,0.072021335,0.09602845,0.18176813,0.28808534,0.29837412,0.24007112,0.09945804,0.09945804,0.2469303,0.32581082,0.38754338,0.4355576,0.4698535,0.48014224,0.44584638,0.432128,0.5041494,0.38754338,0.1371835,0.12346515,0.12003556,0.15433143,0.17147937,0.16804978,0.18519773,0.6962063,0.4938606,0.25378948,0.22292319,0.19891608,0.17490897,0.15433143,0.18176813,0.25378948,0.31552204,0.3841138,0.50757897,0.85396725,1.4575747,2.2292318,3.3198407,4.0503426,4.448175,4.523626,4.2766957,4.588788,5.0106273,5.2987127,5.5833683,6.355026,7.798882,9.695444,11.46854,12.823228,13.72178,12.926115,12.380811,12.154458,12.017275,11.434244,11.146159,11.029553,10.782623,10.508256,10.734609,11.701753,12.195613,12.236768,11.790922,10.789482,9.716022,8.8929205,8.621983,8.827758,9.040393,9.112414,8.958082,10.30591,13.241637,16.20137,18.019053,19.764713,21.393766,22.8582,24.11,24.723896,25.807646,27.84482,30.108349,30.653652,29.401854,26.815945,23.883648,21.314886,19.53836,20.04251,20.680412,21.465788,22.432932,23.616138,25.399525,26.747353,26.69591,25.19718,23.142857,21.242865,20.60839,20.646116,20.999365,21.53781,22.017952,22.552967,23.393215,24.843931,27.248072,29.854559,32.611946,35.129265,37.114994,38.38394,38.98412,40.441696,42.21479,43.98103,45.62723,42.88699,39.31679,35.372765,31.466465,27.961426,25.138876,22.77589,21.37319,20.86904,20.639257,20.724997,21.400625,22.306036,23.125708,23.598991,22.998814,22.131128,21.139977,19.905325,18.04306,15.87213,13.519434,11.938394,11.180455,10.398509,9.160428,8.31675,7.7371492,7.4284863,7.531374,7.73029,7.857185,7.5553813,6.90033,6.4133286,6.258997,6.341307,6.042933,5.2815647,4.5167665,3.9851806,3.7691166,3.8342788,4.190956,4.8905916,5.658819,6.392751,6.8797526,6.9654922,6.540223,6.018926,6.368744,6.8145905,6.9517736,6.7494283,6.48535,6.708273,7.490219,8.556821,9.273604,10.63858,12.103014,13.214201,13.855534,14.249936,14.105893,13.450842,12.315649,10.741467,8.755736,6.8043017,6.0052075,6.4373355,7.747438,9.163857,9.897789,10.576848,10.8958,10.88894,10.943813,11.47197,12.089295,12.127021,11.252477,9.455373,10.052121,10.203023,9.832627,8.98209,7.8023114,7.2638664,7.1884155,7.438775,8.018375,9.043822,10.456812,11.348505,11.622872,11.317638,10.593996,12.689473,14.3974085,15.340545,15.88242,17.130789,18.094503,17.768692,16.45516,15.415996,16.863281,18.728977,18.488907,16.78783,15.762384,19.03421,16.997036,12.8197975,11.907528,13.896688,12.655178,8.913498,8.440215,8.906639,8.64942,6.677407,5.5147767,5.456474,6.0395036,6.9826403,8.186425,8.354475,8.172707,8.769455,10.2236,11.5645685,11.2421875,10.604284,9.932085,9.06097,7.363324,6.385892,6.451054,7.8194594,10.281903,13.169616,15.484588,17.147938,16.37628,13.557159,11.228469,10.772334,9.901219,8.999237,7.9875093,6.3035817,4.5956473,3.7519686,3.7622573,4.3109913,4.8014226,7.226141,10.096705,11.204462,10.182446,8.519095,7.98408,6.5950966,5.0620713,3.8925817,3.391862,3.3129816,3.5633414,3.4398763,3.0866287,3.474172,4.3692946,5.0655007,5.593657,6.025785,6.5024977,7.0306544,7.4970784,7.8846216,8.251588,8.745448,9.115844,9.331907,9.338767,9.160428,8.906639,8.834618,8.083538,7.3564653,6.975781,6.883182,6.3035817,5.9571934,5.7377,5.521636,5.178677,5.137522,5.1992545,5.3330083,5.40503,5.1752477,5.086078,4.9077396,4.6779575,4.437886,4.245829,4.0777793,3.9440255,3.9268777,4.0537724,4.2766957,4.7602673,4.99005,5.3913116,6.2830043,7.9086285,9.4862385,10.360784,10.916377,11.30735,11.489118,11.273054,11.334786,11.547421,11.571428,10.834066,10.113853,9.80862,9.97324,10.336777,10.302481,10.419086,10.871792,11.749766,12.562579,12.229909,12.017275,12.860953,12.812939,11.334786,9.31133,8.927217,8.762596,8.844906,8.964942,8.659708,7.7371492,7.2021337,6.5950966,5.7308407,4.695105,3.5770597,3.1895163,3.234101,3.4398763,3.566771,3.100347,2.2978237,1.5330256,1.0117283,0.7579388,0.7613684,0.7613684,0.67219913,0.51100856,0.4046913,0.4629943,0.72707254,0.9945804,1.1180456,1.0357354,1.3066728,1.5090185,1.6221949,1.7079345,1.9445761,2.9288676,3.542764,3.2855449,2.4041407,1.9068506,1.8245405,1.7765263,1.7456601,1.6633499,1.3924125,0.9842916,0.7442205,0.5761707,0.42869842,0.29837412,0.2194936,0.14747226,0.07545093,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.006859175,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.05144381,0.07888051,0.10288762,0.12689474,0.15090185,0.15090185,0.12346515,0.09602845,0.072021335,0.061732575,0.061732575,0.106317215,0.15433143,0.17833854,0.15090185,0.17833854,0.20234565,0.21263443,0.22978236,0.29151493,0.3018037,0.30523327,0.28122616,0.23664154,0.19891608,0.17490897,0.14061308,0.116605975,0.10288762,0.09259886,0.10288762,0.116605975,0.14061308,0.16804978,0.16804978,0.15433143,0.116605975,0.08573969,0.07888051,0.09259886,0.12689474,0.1920569,0.25378948,0.26407823,0.16804978,0.13032432,0.12346515,0.12346515,0.12346515,0.12346515,0.08573969,0.10288762,0.15776102,0.26064864,0.4424168,0.31895164,0.20920484,0.18176813,0.22292319,0.19891608,0.29494452,0.53158605,0.64819205,0.58988905,0.5041494,0.42869842,0.4389872,0.4629943,0.42869842,0.26064864,0.3806842,0.5041494,0.48014224,0.37039545,0.4424168,0.6001778,0.5418748,0.4355576,0.37725464,0.36696586,0.32924038,0.28465575,0.23664154,0.20920484,0.26064864,0.26064864,0.22292319,0.1920569,0.18519773,0.19891608,0.18519773,0.29151493,0.3841138,0.40126175,0.34981793,0.4972902,0.607037,0.66191036,0.66533995,0.64133286,0.77508676,1.0460242,1.4438564,1.9274281,2.4418662,2.952875,3.7039545,4.2355404,4.2046742,3.3884325,3.1072063,2.8534167,2.5001693,2.393852,3.357566,4.40702,5.007198,5.360445,5.6519604,6.042933,7.1884155,7.3290286,7.006647,6.81802,7.414768,8.1487,8.779744,8.913498,8.934075,10.010965,11.646879,11.129011,10.127572,9.407358,8.820899,8.783174,9.462232,10.738038,11.96926,11.993267,11.334786,10.151579,9.462232,9.242738,8.436785,6.800872,4.6265135,2.7093742,1.5536032,1.3581166,1.529596,1.646202,1.6942163,1.7765263,2.1057668,2.253239,2.1160555,1.7353712,1.2723769,0.9911508,1.4541451,1.1592005,0.58645946,0.12003556,0.044584636,0.20577525,0.44584638,0.7613684,1.0666018,1.1763484,1.2346514,1.3992717,1.5090185,1.488441,1.3443983,0.805953,0.45270553,0.22635277,0.08573969,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.017147938,0.037725464,0.05144381,0.07545093,0.09945804,0.12346515,0.18519773,0.23664154,0.15090185,0.10288762,0.082310095,0.106317215,0.15433143,0.16804978,0.13032432,0.17833854,0.2503599,0.31209245,0.33609957,0.37382504,0.52815646,0.4355576,0.15776102,0.18176813,0.2194936,0.25721905,0.24350071,0.19891608,0.19891608,0.20920484,0.20577525,0.16119061,0.11317638,0.1371835,0.16119061,0.21263443,0.37725464,0.58302987,0.59674823,0.5453044,0.67219913,1.1351935,1.99602,3.2032347,5.6348124,6.992929,7.346176,6.800872,5.5079174,4.7774153,4.4104495,5.171818,7.3221693,10.604284,15.37827,16.187653,15.515453,14.610043,13.488567,13.087306,12.562579,11.842365,11.094715,10.72775,10.847785,11.245617,11.074138,10.295622,9.674867,10.247607,11.482259,12.562579,12.840376,11.842365,10.179015,8.748878,8.107545,8.491658,9.794902,11.091286,11.166737,12.339656,15.237658,18.814716,20.731855,22.419212,23.845922,24.840502,25.084003,25.330933,25.711617,26.572443,27.261791,26.140316,23.149715,20.587814,18.694681,17.573206,17.182234,17.70696,18.303709,18.945042,19.761284,21.04052,21.846472,22.131128,21.20514,19.298288,17.562918,16.70895,16.760393,17.12736,17.422304,17.470318,17.192522,17.322845,18.163095,19.802439,22.11055,24.538698,27.080023,28.945719,30.032898,30.900583,31.850578,33.287575,35.029808,36.898933,38.74405,37.24189,34.67656,31.953466,29.521889,27.374968,25.61559,23.739605,22.340332,21.664703,21.592682,22.456938,23.280039,24.0174,24.723896,25.526419,25.306927,24.044838,22.041958,19.665255,17.333136,14.781522,11.646879,8.940934,7.2604365,6.759717,6.492209,6.159539,5.7754254,5.4804807,5.5559316,5.909179,6.574519,6.9654922,6.9380555,6.8043017,6.464772,5.809721,5.127233,4.6265135,4.4550343,4.149801,3.8274195,3.6868064,3.865145,4.4241676,5.0586414,5.5662203,5.950334,6.1972647,6.2727156,6.001778,6.1458206,6.6225333,7.1061053,7.0203657,6.5779486,6.138962,6.4133286,7.455923,8.652849,10.055551,11.513125,12.8197975,13.845244,14.5414505,13.9309845,13.155897,11.958971,10.124143,7.4627824,5.521636,4.5784993,4.698535,5.5387836,6.3310184,7.174697,9.088407,10.991828,12.089295,11.869802,12.22648,12.459691,12.4802685,11.845795,9.794902,7.610255,6.341307,5.909179,6.0840883,6.48535,6.5710897,6.6293926,6.7459984,7.2124224,8.529384,9.884071,10.947243,11.0981455,10.851214,11.842365,12.782072,11.540562,11.742908,14.4317045,18.080786,17.87501,16.88729,14.942713,12.641459,11.382801,10.700313,10.281903,9.078118,7.438775,7.0958166,9.465661,10.494537,11.05699,11.924676,13.780083,12.116733,11.080997,10.868362,10.206452,6.3481665,4.0537724,3.2135234,3.2512488,3.8891523,5.1580997,7.133542,9.030104,10.323058,10.539123,9.23245,9.829198,11.032983,12.655178,13.834956,13.015285,11.684605,12.394529,14.445422,17.185663,20.018501,19.336014,18.434032,18.04649,17.20967,13.227919,9.688584,8.117833,10.034973,13.639469,13.824667,8.06296,5.24041,4.1120753,3.6525106,3.0660512,3.8102717,5.1512403,6.464772,7.6788464,9.277034,8.947794,6.7974424,5.2026844,4.866585,4.804852,4.3178506,3.9303071,3.474172,3.1792276,3.6936657,5.0003386,5.754848,6.012067,6.1492505,6.883182,6.883182,7.0923867,7.6788464,8.515666,9.184435,10.357354,11.190743,11.465111,10.9541025,9.431366,8.539673,8.021805,7.7542973,7.6033955,7.431916,6.931196,6.56766,6.3173003,6.1904054,6.2418494,6.4236174,6.4236174,6.2898636,6.0052075,5.4941993,5.188966,4.955754,4.9008803,4.9660425,4.928317,4.928317,4.6093655,4.1120753,3.6285036,3.3712845,3.8857226,4.4996185,5.1512403,5.970912,7.2638664,8.299602,8.961512,9.458802,9.757176,9.599416,8.803751,8.56025,8.659708,8.8929205,9.0644,9.126132,9.167287,9.283894,9.3764925,9.156999,9.095266,9.592556,10.062409,10.192734,9.949233,9.2153015,8.107545,6.8866115,5.977771,5.967482,6.831738,7.6171136,8.014946,7.8194594,6.927767,6.608815,6.358455,5.936616,5.0757895,3.4638834,2.8534167,2.6373527,2.4418662,2.3218307,2.760818,3.1517909,2.5001693,1.9068506,1.7936742,1.8931323,2.452155,2.8396983,2.6819375,2.0920484,1.6633499,1.8965619,2.4487255,2.867135,2.9631636,2.7916842,2.585909,2.5961976,2.469303,2.1880767,2.0920484,2.7128036,2.5584722,2.2155135,2.0303159,2.0920484,1.920569,1.704505,1.4815818,1.2689474,1.039165,0.805953,0.61046654,0.45270553,0.32238123,0.21263443,0.26407823,0.26407823,0.17490897,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.0,0.006859175,0.020577524,0.041155048,0.058302987,0.072021335,0.06516216,0.048014224,0.0274367,0.024007112,0.05144381,0.08573969,0.116605975,0.14061308,0.15090185,0.16119061,0.18519773,0.19891608,0.14747226,0.14747226,0.22292319,0.2469303,0.19548649,0.15090185,0.16804978,0.17490897,0.17833854,0.19548649,0.26407823,0.2777966,0.274367,0.25378948,0.22635277,0.19891608,0.16462019,0.12003556,0.08573969,0.06859175,0.06859175,0.06859175,0.09259886,0.14404267,0.18862732,0.17833854,0.14747226,0.09602845,0.06516216,0.07545093,0.12689474,0.17490897,0.21263443,0.2194936,0.18176813,0.09602845,0.12689474,0.14747226,0.14747226,0.14061308,0.17147937,0.22292319,0.29837412,0.29494452,0.21263443,0.16119061,0.19548649,0.18862732,0.19891608,0.26064864,0.39440256,0.5590228,0.7099246,0.72707254,0.61389613,0.48014224,0.38754338,0.32581082,0.3018037,0.3018037,0.29494452,0.37039545,0.4115505,0.4115505,0.3806842,0.3566771,0.4081209,0.4389872,0.432128,0.39097297,0.32924038,0.23321195,0.20234565,0.18862732,0.17490897,0.17490897,0.18519773,0.17833854,0.16462019,0.16804978,0.2469303,0.29494452,0.29837412,0.29151493,0.29151493,0.29151493,0.38754338,0.4698535,0.53158605,0.5590228,0.5418748,0.6962063,0.89169276,1.0597426,1.2517995,1.6496316,2.16064,2.551613,2.8945718,3.175798,3.3129816,2.7882545,2.4898806,2.3664153,2.5996273,3.6147852,4.6916757,5.754848,6.7322803,7.455923,7.641121,7.1095347,6.9826403,7.040943,7.239859,7.720001,8.443645,9.445084,10.878652,12.298501,12.672326,12.21619,10.31277,8.903209,8.64599,8.930646,9.644,8.700864,7.0375133,5.6039457,5.3673043,5.778855,6.5162163,8.018375,9.414218,8.512236,5.909179,6.111525,5.9983487,4.2046742,1.138623,1.5055889,1.8142518,2.0680413,2.2738166,2.4487255,2.2223728,1.6324836,1.1832076,1.0014396,0.85739684,0.83338976,0.64819205,0.39440256,0.18176813,0.16804978,0.4355576,0.7373613,0.9774324,1.1317638,1.2586586,1.1934965,1.1180456,0.9568549,0.70306545,0.4389872,0.22635277,0.16462019,0.18176813,0.20577525,0.15776102,0.09945804,0.034295876,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.010288762,0.01371835,0.116605975,0.15433143,0.1371835,0.09945804,0.09259886,0.10288762,0.09602845,0.21263443,0.432128,0.5693115,0.39783216,0.29151493,0.22292319,0.18176813,0.17833854,0.19548649,0.2503599,0.216064,0.1097468,0.08573969,0.09259886,0.14404267,0.19548649,0.24007112,0.30866286,0.28122616,0.26407823,0.2503599,0.23664154,0.20920484,0.24350071,0.31209245,0.4389872,0.59331864,0.6927767,0.7613684,0.980862,1.8073926,3.4913201,6.0978065,6.701414,6.7459984,6.210983,5.521636,5.545643,5.826869,6.2727156,6.711703,7.2124224,8.06639,9.72288,11.732618,13.423406,13.937843,12.21962,11.876661,11.859513,11.986408,12.157887,12.339656,12.46998,12.38424,12.147599,11.825217,11.506266,10.768905,9.911508,8.903209,8.097256,8.22758,8.327039,8.498518,9.218731,10.340206,11.091286,11.132441,13.46799,16.564907,19.483486,21.877338,22.477516,22.882208,23.166862,23.595562,24.621008,25.450968,25.780209,25.368658,24.147726,22.244305,19.692692,18.005335,17.04162,16.828985,17.573206,17.141079,16.503176,16.280252,16.756964,17.892159,18.855871,17.909306,16.088194,14.078457,12.229909,12.507706,12.768354,12.929544,13.025573,13.210771,13.478279,13.934414,14.767803,15.9750185,17.37429,18.903887,20.971928,23.105131,25.132017,27.138325,28.990303,30.711956,32.17296,33.32873,34.227283,33.476204,31.291555,29.285248,28.043737,27.10403,26.10945,25.039417,24.085993,23.34863,22.837624,23.293758,24.120289,25.512701,27.491573,29.909431,32.015198,31.274408,28.650774,24.792488,20.018501,15.923574,12.857523,10.912948,9.626852,7.956643,6.9071894,6.327589,6.025785,5.892031,5.909179,5.9880595,6.183546,6.3035817,6.262427,6.060081,5.5730796,5.1683884,5.0174866,4.9694724,4.554492,4.064061,3.7451096,3.5221863,3.415869,3.5599117,4.496189,5.144381,5.5250654,5.5730796,5.147811,5.2026844,5.593657,6.210983,6.8043017,6.9826403,6.8454566,7.0958166,7.829748,9.016385,10.508256,11.286773,12.411677,13.742357,14.867262,15.114192,15.453721,16.071047,15.107333,12.260776,8.779744,5.1409516,3.7005248,3.4364467,3.6799474,4.1120753,5.813151,7.881192,9.884071,11.38966,11.96926,12.127021,11.941824,11.818358,11.640019,10.762046,7.442205,5.456474,4.4447455,4.2423997,4.897451,5.411889,5.8645945,6.15268,6.420188,7.06495,7.874333,8.968371,9.73317,10.0041065,10.034973,9.002667,8.193284,8.467651,10.028113,12.418536,13.910407,14.939283,14.79867,13.718349,12.871242,13.155897,14.267084,15.549749,16.87357,18.629519,16.311117,13.564018,11.736049,11.934964,15.011304,17.151367,15.522313,13.656617,12.950122,12.706621,12.130451,10.110424,7.6274023,5.4804807,4.290414,4.9420357,6.3481665,7.301592,7.6685576,8.412778,10.360784,11.509696,12.373952,12.994707,12.977559,14.198492,15.920145,18.310568,21.187992,24.010542,23.533829,19.853882,19.071936,21.829325,23.300617,19.78872,15.289101,11.979549,11.660598,15.741806,12.048141,8.200144,6.2967224,6.3310184,6.1561093,5.8543057,4.8322887,3.8925817,3.4810312,3.6627994,4.437886,5.2266912,6.416758,7.7371492,8.272165,7.891481,7.085528,6.9826403,7.6205435,7.9292064,7.915488,7.7440085,7.1781263,6.2384195,5.171818,7.291303,9.122703,10.271614,10.566559,10.076128,9.784613,9.72288,9.119273,7.949784,6.9517736,7.7714453,8.580828,9.383351,10.1481495,10.837497,10.179015,9.235879,8.423067,7.9737906,7.9257765,8.128122,7.963502,7.7028537,7.442205,7.1026754,6.6225333,6.1732574,5.7754254,5.442755,5.161529,4.955754,4.722542,4.4241676,4.173808,4.2526884,4.8117113,5.422178,5.960623,6.368744,6.677407,7.1987042,7.56224,7.8263187,8.032094,8.193284,8.1041155,7.888051,7.7714453,7.798882,7.8434668,7.6616983,7.795452,8.086967,8.31332,8.189855,7.689135,7.346176,7.414768,8.011517,9.095266,10.1481495,9.071259,7.8503256,7.4765005,7.9429245,8.351046,8.508806,8.3922,7.956643,7.133542,6.759717,6.5127864,6.1492505,5.5833683,4.880303,4.417309,3.7142432,3.2958336,3.5393343,4.7019644,5.5319247,5.744559,5.346727,4.98662,5.9434752,6.468202,5.0277753,3.683377,3.3266997,3.690236,5.0929375,5.6005163,5.3673043,4.4550343,2.8294096,2.1812177,1.9891608,2.0474637,2.1812177,2.2498093,2.3252604,2.0680413,1.8142518,1.7182233,1.7490896,1.6667795,1.5227368,1.3375391,1.1420527,0.9877212,0.83338976,0.67219913,0.6276145,0.66191036,0.5796003,0.30523327,0.17833854,0.09259886,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.017147938,0.01371835,0.01371835,0.030866288,0.0548734,0.072021335,0.07888051,0.06516216,0.037725464,0.020577524,0.030866288,0.0548734,0.06516216,0.06516216,0.072021335,0.09259886,0.1097468,0.14061308,0.17147937,0.16804978,0.22635277,0.29494452,0.29494452,0.22635277,0.17147937,0.16119061,0.14747226,0.14747226,0.17147937,0.22292319,0.2194936,0.20920484,0.19548649,0.18176813,0.17147937,0.14747226,0.12346515,0.10288762,0.09259886,0.116605975,0.1371835,0.15433143,0.18519773,0.2194936,0.22978236,0.21263443,0.17490897,0.13032432,0.12346515,0.2194936,0.25378948,0.24350071,0.2194936,0.19548649,0.17833854,0.2709374,0.26064864,0.22292319,0.21263443,0.3018037,0.31552204,0.32238123,0.26064864,0.14747226,0.082310095,0.12003556,0.15090185,0.16462019,0.17490897,0.22292319,0.31895164,0.45270553,0.5658819,0.5796003,0.39097297,0.3018037,0.25721905,0.22292319,0.19891608,0.21263443,0.274367,0.30866286,0.32581082,0.32238123,0.28122616,0.25378948,0.2503599,0.26064864,0.26750782,0.23664154,0.20920484,0.2469303,0.25721905,0.2194936,0.16119061,0.15776102,0.20234565,0.25721905,0.29494452,0.30523327,0.32924038,0.33609957,0.3566771,0.39097297,0.4115505,0.44584638,0.5041494,0.58645946,0.6859175,0.78537554,0.7956643,0.89855194,1.0597426,1.2449403,1.4232788,1.728512,2.0646117,2.5413244,3.1243541,3.5976372,3.2992632,3.1895163,3.2786856,3.673088,4.5647807,5.1821065,5.7994323,6.5230756,7.233,7.5553813,7.349606,7.630832,8.152129,8.790032,9.527394,10.912948,11.80121,12.370522,12.4802685,11.688034,10.587136,9.091836,8.086967,7.747438,7.5279446,7.2158523,6.0840883,4.605936,3.3438478,2.9665933,3.3712845,4.0674906,5.15467,6.433906,7.394191,7.2021337,6.615674,5.3673043,3.433017,1.0185875,1.4575747,1.9823016,2.5241764,2.8534167,2.5790498,2.0989075,1.4610043,1.039165,0.89512235,0.77851635,0.6893471,0.490431,0.29837412,0.20234565,0.26407823,0.67219913,1.0220171,1.2175035,1.2277923,1.097468,0.8676856,0.66876954,0.4355576,0.20234565,0.08573969,0.33266997,0.40126175,0.37725464,0.31209245,0.216064,0.13032432,0.041155048,0.0,0.0,0.0,0.0,0.044584636,0.07545093,0.07888051,0.06516216,0.12689474,0.16462019,0.16804978,0.12689474,0.030866288,0.041155048,0.12689474,0.274367,0.4389872,0.5418748,0.44584638,0.34638834,0.25721905,0.18862732,0.15433143,0.13032432,0.09602845,0.082310095,0.08573969,0.06859175,0.06859175,0.10288762,0.14747226,0.19891608,0.26407823,0.26407823,0.26407823,0.26407823,0.2777966,0.31895164,0.38754338,0.45613512,0.4972902,0.53844523,0.65162164,0.86082643,1.3581166,2.3389788,3.957744,6.3173003,6.0737996,5.6176643,5.24041,5.178677,5.6005163,6.2692857,7.3393173,8.128122,8.491658,8.820899,9.897789,10.933525,11.506266,11.30049,10.096705,10.662587,11.962401,12.744347,12.682614,12.38424,11.770344,12.466551,13.296511,13.591455,13.207341,12.614022,11.80121,10.768905,9.880642,9.832627,9.856634,9.911508,10.916377,12.754636,14.287662,14.195063,15.810398,17.947031,19.949911,21.69214,22.494663,23.180582,23.808197,24.411804,25.008553,25.032558,23.832203,21.928782,19.69955,17.388008,15.498305,14.208781,13.426835,13.070158,13.056439,12.55229,12.171606,12.247057,12.792361,13.478279,13.749216,12.9638405,11.808069,10.64201,9.5033865,9.523964,9.499957,9.458802,9.534253,9.966381,10.635151,11.30049,11.9040985,12.435684,12.950122,14.695783,16.828985,19.161106,21.654415,24.43238,27.285797,30.152933,32.231262,33.153824,33.01321,30.92116,28.976585,27.639046,27.049156,27.038868,25.968836,24.895376,24.027689,23.410364,22.919933,23.022821,23.626429,24.994833,27.158903,29.899143,33.57909,34.75201,33.990643,30.962317,24.398085,19.140528,15.038741,12.490558,11.111863,9.746887,9.074688,7.970361,7.034084,6.5642304,6.5642304,6.759717,6.8969,6.869464,6.625963,6.186976,5.6176643,5.1340923,4.9591837,4.98662,4.7602673,4.0709205,3.5942078,3.2546785,3.069481,3.1483612,4.170378,5.1512403,5.686256,5.669108,5.2781353,5.099797,5.188966,5.579939,6.1972647,6.8728933,7.164408,7.6685576,8.375052,9.246168,10.237319,11.338216,13.056439,14.627191,15.6869335,16.283682,17.017612,17.470318,16.616352,14.140189,10.456812,6.608815,4.139512,3.0043187,2.8499873,2.9871707,4.0263357,5.6348124,7.606825,9.650859,11.406808,11.362224,11.283342,11.321068,11.410237,11.293632,9.434795,7.675417,6.217842,5.2644167,5.003768,5.086078,5.302142,5.669108,6.3173003,7.5039372,7.2535777,7.438775,8.327039,9.304471,8.868914,7.582818,6.9963584,7.377043,8.694004,10.618003,12.754636,14.027013,14.273943,13.649758,12.641459,12.212761,11.893809,12.531713,13.786942,14.13676,11.22161,10.038403,10.182446,11.626302,14.71636,15.343974,14.400838,14.1299,14.856973,14.96672,13.924125,13.155897,11.327928,8.471081,5.960623,6.1972647,6.701414,7.051232,7.4936485,8.934075,9.897789,10.398509,12.13731,14.71636,15.614912,15.7795315,16.736387,19.239986,23.389786,28.626766,23.238884,18.001905,16.29054,18.560926,22.330044,21.815605,18.735836,15.354263,13.495427,14.534592,12.343085,9.465661,7.4113383,6.5470824,6.094377,6.310441,5.970912,4.8837323,3.4878905,2.8705647,3.0351849,3.6044965,4.461893,5.346727,5.861165,6.4819202,6.608815,6.869464,7.3290286,7.514226,7.6342616,7.689135,6.9380555,5.5662203,4.6916757,6.495639,7.73372,8.179566,7.764586,6.5642304,6.0086374,5.7377,5.346727,4.8837323,4.8597255,6.060081,7.658269,9.112414,10.192734,11.002116,10.6488695,10.069269,9.510246,9.108984,8.89635,8.7283,8.378482,7.9737906,7.56567,7.1061053,6.5127864,6.2418494,5.9812007,5.552502,4.9248877,4.705394,4.537344,4.413879,4.413879,4.681387,5.1238036,5.552502,6.0395036,6.5470824,6.914048,7.2707253,7.5382333,7.7097125,7.798882,7.8606143,7.9017696,7.805741,7.7542973,7.7097125,7.390761,6.715132,6.701414,6.852316,6.866034,6.6225333,6.3618846,6.3447366,6.756287,7.473071,8.083538,8.793462,8.529384,8.467651,9.026674,9.884071,10.213311,9.510246,8.501947,7.8263187,8.011517,7.6342616,7.099246,6.601956,6.2041235,5.802862,5.5730796,5.73427,5.8680243,5.871454,5.9400454,6.0806584,6.0395036,5.6485305,5.1580997,5.2472687,5.1066556,3.981751,3.0043187,2.6750782,2.877424,3.724532,3.8720043,3.542764,2.8705647,1.9137098,1.5673214,1.4850113,1.605047,1.786815,1.821111,1.7319417,1.6153357,1.5398848,1.529596,1.5536032,1.4987297,1.4815818,1.4610043,1.3341095,0.922559,0.7133542,0.61389613,0.64133286,0.7099246,0.64476246,0.37725464,0.39783216,0.41840968,0.29494452,0.0274367,0.01371835,0.010288762,0.010288762,0.006859175,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0274367,0.030866288,0.020577524,0.020577524,0.034295876,0.048014224,0.0548734,0.06516216,0.058302987,0.030866288,0.01371835,0.034295876,0.0548734,0.05144381,0.037725464,0.041155048,0.06859175,0.082310095,0.11317638,0.15776102,0.19891608,0.2777966,0.31552204,0.29837412,0.24007112,0.18862732,0.16462019,0.14404267,0.14404267,0.16804978,0.19891608,0.1920569,0.17833854,0.16119061,0.1371835,0.12689474,0.15090185,0.16804978,0.17490897,0.17833854,0.19548649,0.20234565,0.1920569,0.1920569,0.20920484,0.22978236,0.24350071,0.2469303,0.216064,0.18176813,0.22635277,0.24007112,0.216064,0.19548649,0.20234565,0.22635277,0.32238123,0.33266997,0.29494452,0.26407823,0.31552204,0.274367,0.22978236,0.17147937,0.106317215,0.06859175,0.082310095,0.12003556,0.12346515,0.09259886,0.07545093,0.12689474,0.2503599,0.4046913,0.48700142,0.34295875,0.28465575,0.26407823,0.23321195,0.1920569,0.17147937,0.1920569,0.22635277,0.2469303,0.2503599,0.23664154,0.21263443,0.1920569,0.19548649,0.21263443,0.20234565,0.21263443,0.2503599,0.26407823,0.24007112,0.19891608,0.18519773,0.21263443,0.26750782,0.32581082,0.32924038,0.34981793,0.38754338,0.45613512,0.5212973,0.5212973,0.51100856,0.5590228,0.6859175,0.8711152,1.0460242,0.9431366,0.980862,1.1489118,1.3649758,1.5090185,1.7696671,2.1983654,2.8328393,3.525616,3.9508848,3.9097297,4.091498,4.4104495,4.8734436,5.5730796,5.8680243,6.118384,6.5024977,7.0135064,7.466212,7.905199,8.597976,9.352485,10.072699,10.762046,11.698323,12.130451,11.993267,11.252477,9.918367,9.246168,8.683716,7.6651278,6.334448,5.545643,5.188966,4.355576,3.542764,3.0523329,2.9665933,2.9460156,3.100347,3.4192986,4.0023284,5.038064,5.874883,5.219832,3.8720043,2.4075704,1.1900668,1.5776103,2.095478,2.6545007,3.018037,2.784825,2.1743584,1.4747226,1.0117283,0.823101,0.66191036,0.548734,0.34981793,0.22635277,0.26407823,0.4629943,1.0151579,1.3478279,1.3992717,1.138623,0.58645946,0.39440256,0.2777966,0.14061308,0.0,0.0,0.4081209,0.48357183,0.37382504,0.2194936,0.1371835,0.07888051,0.024007112,0.0,0.0,0.0,0.0,0.061732575,0.1097468,0.116605975,0.11317638,0.16804978,0.20920484,0.22635277,0.19548649,0.072021335,0.07888051,0.19891608,0.31209245,0.36353627,0.39783216,0.3806842,0.33609957,0.2777966,0.216064,0.14404267,0.07888051,0.024007112,0.017147938,0.044584636,0.044584636,0.044584636,0.08916927,0.13375391,0.16804978,0.20234565,0.22635277,0.2469303,0.26750782,0.32924038,0.51100856,0.5761707,0.4972902,0.41840968,0.432128,0.5796003,0.922559,1.786815,2.942586,4.3178506,5.9983487,5.5833683,4.996909,4.8185706,5.188966,5.813151,6.711703,7.6857057,8.556821,9.328478,10.182446,10.556271,10.326488,9.657719,9.132992,9.743458,10.7757635,11.447963,11.712041,11.784062,12.109874,12.915827,14.459141,15.601193,15.54632,13.831526,13.162757,12.699762,12.236768,11.746337,11.375941,11.087856,11.365653,12.703192,14.956431,17.339994,17.53548,17.984756,18.495766,19.202261,20.53294,21.78474,23.019392,23.69159,23.623,23.002243,21.733295,19.757853,17.607502,15.488017,13.262215,11.948683,10.909517,10.055551,9.301042,8.570539,8.1212635,8.114404,8.460793,8.97866,9.379922,9.266746,8.886061,8.351046,7.7577267,7.208993,6.941485,6.7974424,6.7322803,6.807731,7.1952744,7.829748,8.505377,9.033533,9.362774,9.585697,11.38623,13.454271,15.820687,18.533491,21.674994,25.132017,28.918282,31.932888,33.644253,34.07638,31.017189,28.76738,27.042297,25.893385,25.69104,24.548986,23.454948,22.717587,22.343761,22.065966,21.891056,22.237446,23.406935,25.588152,28.859978,33.17097,36.113556,37.307053,35.66428,29.35384,23.35549,18.578075,15.371411,13.526293,12.243628,11.38966,9.97324,8.700864,7.956643,7.822889,7.7440085,7.442205,7.0443726,6.5985265,6.0703697,5.5902276,5.130663,4.839148,4.7019644,4.5339146,3.9303071,3.4535947,3.1140654,2.9494452,3.0454736,3.7553983,4.712253,5.346727,5.501058,5.4496145,4.996909,4.839148,5.038064,5.672538,6.842027,7.4799304,8.06296,8.80718,9.6817255,10.39165,11.207891,12.929544,14.599753,15.8138275,16.746675,17.082775,16.890718,16.026463,14.30481,11.485688,8.666568,6.495639,5.164959,4.4413157,3.666229,3.6044965,4.3521466,5.7719955,7.6616983,9.760606,9.983529,10.089847,10.319629,10.751757,11.30735,11.605724,10.566559,8.985519,7.490219,6.5230756,5.90575,5.4770513,5.442755,6.0052075,7.3393173,7.1369715,6.9552035,7.2947326,7.6959944,6.7459984,6.6225333,6.800872,7.4456344,8.47451,9.578837,11.441104,12.878101,13.855534,14.38026,14.490007,14.959861,13.173045,11.173596,9.794902,8.680285,7.1541195,7.548522,8.680285,10.024684,11.712041,11.324498,11.72233,13.214201,15.268523,16.516893,14.695783,13.114742,10.755186,7.949784,6.3618846,7.64798,8.477941,8.344186,8.018375,9.561689,11.770344,13.845244,16.396858,18.152807,15.9578705,14.987297,15.556609,18.663815,24.051697,30.207806,25.214327,20.004784,17.20967,17.847572,21.335464,20.718138,19.058218,17.809847,16.952452,14.973578,12.343085,9.280463,6.9860697,5.895461,5.686256,6.5024977,7.4044795,7.274155,5.8680243,3.799983,3.0146074,2.9220085,3.5359046,4.57164,5.422178,6.293293,6.7357097,7.1849856,7.7611566,8.268735,8.004657,7.764586,7.0032177,6.0532217,6.1492505,6.7219915,6.3893213,5.6485305,4.756838,3.7313912,3.6696587,3.6696587,3.6765177,3.724532,3.9200184,4.791134,6.193835,7.517656,8.447074,8.958082,8.841476,8.844906,8.786603,8.573969,8.200144,7.9600725,7.682276,7.349606,6.9552035,6.495639,6.293293,6.3961806,6.293293,5.8234396,5.1752477,4.8597255,4.7979927,4.866585,5.038064,5.3844523,5.65539,5.844017,6.1629686,6.680836,7.3187394,7.8194594,8.107545,8.217292,8.196714,8.080108,8.052671,8.080108,8.172707,8.152129,7.623973,6.8728933,6.7459984,6.677407,6.4407654,6.1286726,5.9331865,5.9571934,6.2555676,6.6636887,6.790583,7.130112,7.4936485,7.9772205,8.570539,9.184435,9.39021,8.344186,7.31531,7.1061053,8.049242,7.582818,6.8797526,6.262427,5.888602,5.7411294,5.672538,6.0052075,6.4304767,6.6568294,6.427047,5.6999745,5.411889,5.3913116,5.353586,4.911169,4.3521466,3.7553983,3.2649672,2.9185789,2.6579304,2.411,2.1091962,1.8142518,1.5604624,1.3443983,1.2175035,1.1694894,1.1729189,1.1934965,1.1866373,1.1489118,1.1934965,1.2758065,1.3615463,1.4198492,1.3786942,1.3512574,1.3272504,1.2483698,0.9774324,0.89169276,0.9362774,0.99801,1.0048691,0.9294182,0.6207553,0.64133286,0.66533995,0.5212973,0.17833854,0.082310095,0.0274367,0.010288762,0.006859175,0.0,0.0,0.006859175,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.010288762,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.0274367,0.017147938,0.017147938,0.0274367,0.0274367,0.030866288,0.05144381,0.0548734,0.037725464,0.01371835,0.024007112,0.034295876,0.044584636,0.048014224,0.058302987,0.07888051,0.09259886,0.12346515,0.17490897,0.22635277,0.274367,0.2777966,0.25378948,0.216064,0.18176813,0.15776102,0.14747226,0.15433143,0.17147937,0.19548649,0.19891608,0.1920569,0.16804978,0.13375391,0.12346515,0.18862732,0.24007112,0.26750782,0.26750782,0.25721905,0.216064,0.17833854,0.16119061,0.16462019,0.18176813,0.21263443,0.2469303,0.2469303,0.21263443,0.15090185,0.15090185,0.15433143,0.15776102,0.16804978,0.17833854,0.23321195,0.29837412,0.3018037,0.2469303,0.1920569,0.1371835,0.106317215,0.09602845,0.09259886,0.06859175,0.07888051,0.106317215,0.10288762,0.07888051,0.09602845,0.16462019,0.2503599,0.32924038,0.36696586,0.32581082,0.3018037,0.28808534,0.26750782,0.24007112,0.20234565,0.16804978,0.18176813,0.19548649,0.20234565,0.22978236,0.26064864,0.28122616,0.28465575,0.26407823,0.2194936,0.20920484,0.1920569,0.19548649,0.2194936,0.25378948,0.25721905,0.23321195,0.22635277,0.25378948,0.31895164,0.37382504,0.4389872,0.52815646,0.6036074,0.5693115,0.5521636,0.607037,0.8025235,1.0734608,1.2243627,1.0494537,1.1420527,1.3238207,1.5090185,1.6942163,2.095478,2.651071,3.3815732,4.1189346,4.4996185,4.6676683,5.096367,5.586798,6.046363,6.5024977,6.660259,6.842027,7.0752387,7.414768,7.9429245,8.484799,9.091836,9.822338,10.583707,11.118723,10.926665,10.813489,10.659158,10.233889,9.194724,8.844906,8.546532,7.143831,5.0449233,4.2252517,4.73969,4.0846386,3.350707,3.093488,3.3541365,3.0248961,2.9151495,3.0489032,3.1586502,2.6853669,2.428148,2.7711067,2.7162333,2.0714707,1.4438564,1.728512,2.0577524,2.4041407,2.7333813,3.0146074,2.3801336,1.5536032,0.9842916,0.7476501,0.5555932,0.33609957,0.19891608,0.23664154,0.47328308,0.8848336,1.4232788,1.6084765,1.4061309,0.86082643,0.12346515,0.106317215,0.15776102,0.116605975,0.0,0.0,0.216064,0.28122616,0.22292319,0.13375391,0.15433143,0.10288762,0.034295876,0.0,0.0034295875,0.010288762,0.0034295875,0.037725464,0.06516216,0.08573969,0.13032432,0.24007112,0.29494452,0.29151493,0.2469303,0.20577525,0.2194936,0.29494452,0.34981793,0.35324752,0.34638834,0.30523327,0.2709374,0.23664154,0.18176813,0.08573969,0.017147938,0.010288762,0.010288762,0.0,0.0,0.010288762,0.08916927,0.15776102,0.1920569,0.2194936,0.25378948,0.30866286,0.38754338,0.5178677,0.7442205,0.7339317,0.4424168,0.26750782,0.3566771,0.59674823,1.1077567,2.2566686,3.5873485,4.856296,6.0326443,5.90575,5.518206,5.3981705,5.744559,6.4098988,7.164408,7.407909,7.8674736,8.875772,10.364213,9.928656,9.5205345,9.132992,9.434795,11.770344,12.487128,11.0981455,10.124143,10.593996,12.05157,15.309678,16.901007,17.240536,16.204802,13.128461,12.151029,11.907528,11.739478,11.38966,11.008976,11.14273,12.247057,13.937843,16.029892,18.550638,19.065077,19.154245,18.855871,18.660385,19.521212,20.574095,21.630407,21.544668,20.19341,18.4649,16.427725,14.87755,13.509145,12.044711,10.22703,9.194724,8.357904,7.466212,6.526505,5.7994323,5.3844523,5.353586,5.5147767,5.7925735,6.193835,6.252138,6.0497923,5.5902276,5.038064,4.698535,4.5956473,4.602506,4.633373,4.6745276,4.7774153,5.0655007,5.597087,6.228131,6.842027,7.346176,8.676856,10.340206,12.569438,15.371411,18.533491,22.038528,25.907104,29.501312,32.454185,34.68342,32.1078,29.408712,26.634176,24.243753,23.10856,22.261452,21.397196,20.827885,20.570665,20.340883,20.045938,20.320305,21.434921,23.719027,27.567024,31.490473,35.022945,36.905792,36.13756,31.956896,26.154034,21.726437,18.475187,16.173935,14.555169,13.046151,11.787492,10.827208,10.206452,9.935514,9.39707,8.381912,7.425057,6.7219915,6.1321025,5.6519604,5.23698,4.8425775,4.4584637,4.1017866,3.7759757,3.4810312,3.234101,3.0797696,3.0969174,3.2786856,3.865145,4.4996185,4.99005,5.305572,4.8425775,4.6402316,4.8014226,5.4599032,6.7974424,7.6376915,8.440215,9.510246,10.72775,11.550851,11.8115,12.926115,14.328816,15.608052,16.489456,16.160215,15.388559,14.249936,12.847235,11.317638,10.419086,9.911508,9.1981535,7.9257765,5.9743414,4.9488945,4.6127954,5.0106273,6.0497923,7.4936485,8.30646,8.405919,8.601405,9.283894,10.422516,12.079007,11.982979,10.916377,9.578837,8.580828,7.5245147,6.5882373,5.967482,5.8405876,6.358455,6.8145905,6.7871537,6.276145,5.3570156,4.1635194,5.353586,6.475061,7.449064,8.1487,8.4093485,9.407358,11.153018,13.066729,14.750656,16.002455,18.056778,16.208231,12.312219,8.515666,7.250148,7.143831,7.3873315,7.4456344,7.226141,7.058091,7.610255,9.071259,11.008976,13.416546,16.684942,14.791811,10.827208,6.9620624,4.7602673,5.178677,7.716572,9.22216,8.673427,7.3358874,8.776315,14.2362175,19.507494,22.6147,21.589252,14.466,12.181894,12.730629,16.194511,21.335464,25.591581,25.985985,23.043398,21.157125,21.747015,23.259462,19.754423,17.981327,18.564358,19.87446,18.04306,14.287662,10.511685,7.8674736,6.574519,5.926327,6.9792104,8.676856,9.513676,8.471081,5.007198,3.5050385,3.5016088,4.9831905,7.2432885,8.903209,8.940934,8.742019,9.191295,10.47396,12.055,11.495977,10.127572,8.89635,8.429926,9.040393,8.906639,7.613684,6.1046658,4.979761,4.4584637,4.8905916,5.206114,5.267846,5.0277753,4.5167665,4.5270553,4.9180284,5.4667625,5.926327,6.0326443,5.844017,6.0566516,6.2727156,6.279575,6.029215,6.252138,6.444195,6.451054,6.258997,6.012067,6.392751,6.711703,6.6225333,6.1732574,5.826869,5.435896,5.4976287,5.675967,5.8988905,6.341307,6.7700057,6.869464,6.927767,7.174697,7.795452,8.378482,8.618553,8.639131,8.543102,8.4093485,8.447074,8.591117,8.759167,8.766026,8.31675,8.038953,8.008087,7.8331776,7.421627,6.975781,6.3893213,5.871454,5.5730796,5.552502,5.761707,6.2075534,6.5950966,6.6705475,6.478491,6.385892,6.4373355,5.8234396,5.597087,6.108095,6.9826403,6.5539417,6.042933,5.4633327,5.020916,5.15467,5.518206,5.3501563,5.4839106,6.0223556,6.3378778,5.394741,5.209543,5.6176643,6.1321025,5.9297566,5.411889,4.9077396,4.5647807,4.314421,3.8720043,3.0900583,2.4761622,2.0131679,1.6942163,1.5330256,1.3478279,1.2106444,1.039165,0.86082643,0.8025235,0.8265306,0.90541106,1.0528834,1.2209331,1.3272504,1.3101025,1.1489118,0.9534253,0.85396725,1.0048691,1.1420527,1.3306799,1.4267083,1.4129901,1.3992717,0.99801,0.823101,0.6962063,0.53158605,0.34638834,0.16804978,0.06516216,0.024007112,0.017147938,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.041155048,0.0548734,0.048014224,0.0274367,0.01371835,0.0034295875,0.017147938,0.037725464,0.044584636,0.044584636,0.058302987,0.061732575,0.06859175,0.09259886,0.15090185,0.20234565,0.20577525,0.18176813,0.14404267,0.106317215,0.09602845,0.1097468,0.13375391,0.15776102,0.18176813,0.19548649,0.19891608,0.19891608,0.20920484,0.24350071,0.28122616,0.28122616,0.26750782,0.25721905,0.24350071,0.18176813,0.15090185,0.1371835,0.14404267,0.16804978,0.18176813,0.16462019,0.15090185,0.15090185,0.15090185,0.15090185,0.16119061,0.16119061,0.14061308,0.09259886,0.12689474,0.17490897,0.17490897,0.13032432,0.106317215,0.06859175,0.05144381,0.05144381,0.06859175,0.106317215,0.106317215,0.116605975,0.12689474,0.14404267,0.16804978,0.216064,0.2469303,0.2709374,0.2777966,0.22978236,0.15433143,0.16462019,0.19548649,0.21263443,0.21263443,0.18862732,0.1920569,0.1920569,0.1920569,0.22978236,0.29151493,0.33266997,0.34638834,0.30523327,0.18176813,0.17147937,0.17833854,0.18862732,0.216064,0.29151493,0.34981793,0.39440256,0.3806842,0.32924038,0.30523327,0.39097297,0.48357183,0.58988905,0.66876954,0.65505123,0.65505123,0.7373613,1.039165,1.4061309,1.4198492,1.0906088,1.4541451,1.8759843,2.0097382,1.8142518,2.218943,2.8328393,3.7725463,4.887162,5.768566,6.3653145,6.883182,7.301592,7.6033955,7.7371492,7.394191,7.2535777,7.301592,7.6376915,8.467651,8.529384,8.196714,8.930646,10.714031,12.068718,12.7272,12.343085,11.598865,10.89237,10.329918,8.182996,6.3721733,5.5593615,5.518206,5.127233,4.540774,3.690236,2.9151495,2.352697,1.937717,1.8039631,1.8245405,1.9582944,2.2566686,2.867135,2.6613598,1.8588364,1.2655178,1.138623,1.1763484,1.430138,1.7250825,2.061182,2.4418662,2.867135,2.2841053,1.587899,1.0323058,0.72707254,0.64133286,0.37382504,0.30523327,0.51100856,0.9842916,1.6187652,1.7147937,1.529596,1.0700313,0.6001778,0.6241849,0.53844523,0.5007198,0.29151493,0.0,0.0,0.0,0.20234565,0.45613512,0.66876954,0.77851635,0.51100856,0.17833854,0.0,0.010288762,0.044584636,0.010288762,0.0,0.0,0.034295876,0.16804978,0.32581082,0.39440256,0.37382504,0.31552204,0.29151493,0.31552204,0.3566771,0.42526886,0.490431,0.5041494,0.30866286,0.17833854,0.09602845,0.048014224,0.0,0.0,0.0548734,0.0548734,0.0,0.0,0.048014224,0.116605975,0.19548649,0.28122616,0.36696586,0.4389872,0.5761707,0.8025235,1.0014396,0.91569984,0.72021335,0.432128,0.31895164,0.47328308,0.84024894,1.646202,2.74367,4.0023284,5.2026844,6.0566516,6.5950966,7.06838,7.5245147,7.8366075,7.689135,7.0203657,6.6225333,6.6533995,7.239859,8.484799,9.825768,11.187314,12.524854,13.759505,14.784951,14.994157,13.910407,12.823228,12.271064,12.037852,13.588025,13.903547,13.478279,12.641459,11.5645685,11.650309,12.459691,12.082437,10.64201,10.299051,11.958971,12.960411,13.810948,14.915276,16.585485,17.343424,17.854433,18.28656,18.61923,18.629519,18.324286,17.782412,16.897577,15.707511,14.390549,13.227919,11.941824,10.4705305,8.872343,7.3084507,6.1492505,5.3570156,4.5613513,3.7348208,3.1723683,3.2581081,3.117495,2.9803114,3.069481,3.5702004,3.6696587,3.5839188,3.2889743,2.942586,2.867135,2.9803114,2.952875,2.9220085,2.9460156,3.0077481,3.1895163,3.5839188,4.170378,4.880303,5.6005163,6.492209,7.658269,9.647429,12.442543,15.45715,18.61923,21.644127,24.645016,27.615038,30.410152,29.446438,27.357819,24.641586,22.10712,20.875898,20.594673,19.936192,19.167965,18.410025,17.655516,17.545769,18.159666,19.507494,21.548098,24.185452,26.76107,29.172071,30.149504,29.367558,27.450418,23.787619,20.61182,17.909306,15.848124,14.784951,14.030442,13.426835,13.128461,13.097594,13.121602,13.111313,12.109874,10.789482,9.513676,8.31675,7.143831,6.1732574,5.446185,4.9180284,4.4550343,4.1017866,3.8925817,3.6559403,3.3644254,3.1586502,3.1346428,3.5599117,4.249259,4.9488945,5.3398676,5.2301207,4.8837323,4.972902,5.6245236,6.392751,7.3701835,8.934075,10.477389,11.646879,12.343085,13.992717,15.319967,16.016174,16.269962,16.770683,16.842705,15.570327,13.557159,11.427385,9.825768,11.351934,12.061859,11.917816,10.871792,8.879202,7.0752387,5.5593615,4.962613,5.2987127,5.9812007,6.910619,6.7391396,6.427047,6.6876955,7.98065,9.091836,10.072699,10.628291,10.545981,9.705732,8.9100685,8.501947,8.06296,7.4181976,6.636252,5.7582774,4.852866,4.108646,3.6868064,3.724532,4.1635194,4.914599,5.994919,7.2638664,8.423067,8.471081,9.455373,10.449953,10.487679,8.546532,7.7268605,7.174697,6.4716315,5.5662203,4.7602673,4.32128,4.496189,4.5990767,4.386442,4.0434837,4.605936,5.56965,6.7974424,8.39563,10.72775,9.6645775,7.2124224,5.6313825,5.470192,5.56965,6.48535,5.6245236,4.2698364,3.6147852,4.7602673,10.47396,16.53404,21.28402,22.422644,17.027903,9.5205345,8.258447,9.630281,11.286773,12.116733,11.835506,14.318527,19.270851,23.907654,22.978235,20.488356,18.348293,18.37916,20.141968,20.934202,19.260563,18.643238,16.20137,11.396519,6.012067,7.514226,10.038403,10.645439,8.865483,6.728851,4.482471,4.9934793,7.2638664,10.151579,12.360233,11.46854,10.971251,11.369082,13.1421795,16.753534,19.181683,16.907866,13.944703,12.236768,11.626302,12.7272,12.953552,12.13731,10.645439,9.414218,9.280463,9.301042,8.903209,7.932636,6.6533995,4.9934793,4.3658648,4.1292233,3.957744,3.8617156,3.3472774,2.9082901,2.7813954,3.0626216,3.724532,4.7362604,5.785714,6.2727156,6.193835,6.135532,6.23156,6.1286726,6.018926,5.936616,5.751418,5.813151,5.874883,5.8680243,6.012067,6.8043017,8.354475,8.824328,8.769455,8.64942,8.820899,8.711152,8.573969,8.433355,8.361334,8.484799,9.009526,9.331907,9.424506,9.318189,9.108984,9.438225,9.788043,9.764035,9.174147,8.025234,6.9037595,6.108095,5.8405876,6.0052075,6.2247014,6.15268,6.0978065,5.909179,5.5662203,5.188966,5.504488,5.8508763,5.9228973,5.7754254,5.7994323,6.090947,6.210983,5.9126086,5.422178,5.446185,7.363324,8.080108,7.7748747,6.8763227,6.0566516,6.276145,6.094377,5.8200097,5.552502,5.171818,4.7328305,4.5030484,4.4721823,4.5922174,4.7774153,5.020916,4.448175,3.3438478,2.253239,1.9823016,1.8965619,1.8588364,1.7353712,1.4987297,1.2037852,1.0357354,0.9568549,1.0460242,1.2415106,1.3272504,1.3409687,1.1420527,0.89855194,0.69963586,0.5658819,0.5761707,0.6790583,0.864256,1.1180456,1.4335675,1.2895249,1.0597426,0.71678376,0.3566771,0.19891608,0.1371835,0.13032432,0.12346515,0.09259886,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.030866288,0.0034295875,0.0034295875,0.07545093,0.06859175,0.037725464,0.017147938,0.01371835,0.024007112,0.0274367,0.037725464,0.048014224,0.058302987,0.06859175,0.06516216,0.09259886,0.16462019,0.274367,0.20577525,0.15776102,0.13375391,0.13032432,0.14404267,0.16119061,0.19891608,0.23321195,0.25378948,0.26750782,0.2503599,0.2469303,0.23664154,0.21263443,0.17147937,0.17833854,0.1920569,0.20577525,0.20577525,0.18176813,0.14061308,0.13375391,0.15090185,0.18862732,0.24007112,0.23321195,0.2194936,0.19548649,0.15776102,0.12689474,0.12003556,0.1097468,0.1097468,0.12003556,0.12689474,0.12689474,0.12346515,0.116605975,0.09259886,0.058302987,0.041155048,0.034295876,0.044584636,0.06859175,0.09602845,0.12346515,0.12689474,0.12689474,0.14404267,0.16804978,0.18862732,0.20920484,0.2194936,0.21263443,0.20577525,0.20920484,0.20234565,0.20920484,0.23664154,0.274367,0.24007112,0.21263443,0.17833854,0.17147937,0.26407823,0.32581082,0.31895164,0.28122616,0.23321195,0.17147937,0.15776102,0.17147937,0.19548649,0.22635277,0.29151493,0.39097297,0.50757897,0.53158605,0.45613512,0.40126175,0.40126175,0.4424168,0.50757897,0.5761707,0.6310441,0.8848336,1.2209331,1.6633499,1.99602,1.7730967,1.4815818,1.7490896,2.1023371,2.318401,2.4247184,2.4075704,2.860276,3.707384,4.6779575,5.305572,5.9297566,6.584808,7.164408,7.5588107,7.6616983,7.2124224,6.8283086,6.6396813,6.807731,7.4799304,8.224151,8.855195,9.55826,10.326488,10.957532,11.218181,10.463672,9.506817,8.759167,8.207003,8.361334,7.723431,6.324159,4.695105,3.8445675,3.1895163,2.6064866,2.2429502,2.061182,1.8519772,1.3958421,1.2277923,1.2277923,1.3512574,1.611906,1.5398848,1.2929544,1.08032,1.0323058,1.1866373,1.5981878,1.7113642,1.7833855,1.9685832,2.318401,2.0646117,1.7388009,1.4232788,1.1626302,0.97057325,0.7613684,0.5555932,0.61046654,0.94999576,1.3615463,1.2723769,1.1934965,1.1180456,1.0425946,0.980862,0.922559,0.89855194,0.53501564,0.0,0.0,0.14747226,0.39783216,0.66191036,0.8471081,0.88826317,0.5521636,0.18519773,0.034295876,0.082310095,0.06859175,0.01371835,0.0,0.0548734,0.17147937,0.32581082,0.29151493,0.25721905,0.23321195,0.2469303,0.34981793,0.4629943,0.5727411,0.58645946,0.4938606,0.37039545,0.25378948,0.18519773,0.14404267,0.11317638,0.072021335,0.06516216,0.072021335,0.048014224,0.0,0.0,0.07888051,0.18176813,0.28122616,0.36010668,0.41498008,0.6927767,0.96371406,1.1832076,1.2929544,1.2072148,1.0048691,0.66191036,0.607037,0.9911508,1.7182233,3.1860867,4.8494368,6.619104,8.203573,9.098696,9.829198,10.415657,10.113853,8.98209,7.8983397,7.3427467,7.3873315,7.689135,8.028665,8.275595,8.868914,9.47595,9.849775,10.333347,11.856084,14.30138,15.752095,15.594335,13.612033,10.000677,10.350495,10.576848,10.816919,11.269625,12.188754,12.771784,12.6586075,12.05157,11.348505,11.14273,12.089295,13.059869,14.126471,15.415996,17.086205,17.610931,17.590355,17.350283,17.027903,16.592344,16.071047,15.498305,14.836395,14.068168,13.179905,11.561139,9.853205,8.131552,6.5539417,5.3432975,4.3487167,3.333559,2.452155,1.7936742,1.3684053,1.2860953,1.2792361,1.3786942,1.5501735,1.6770682,1.7079345,1.6942163,1.5844694,1.4369972,1.4027013,1.5433143,1.670209,1.7902447,1.903421,2.0063086,2.1091962,2.3081124,2.7916842,3.5393343,4.3178506,5.1992545,6.392751,8.035523,10.134431,12.566009,15.073037,17.521763,19.915615,22.240875,24.490685,25.34122,24.885086,23.70188,22.254593,20.886189,19.288,17.79613,16.503176,15.577187,15.251375,15.62863,16.420864,17.274832,18.001905,18.605513,18.965618,19.761284,20.27915,20.183123,19.517782,17.837284,16.167076,14.5414505,13.155897,12.356804,11.88352,11.492548,11.05699,10.563129,10.106995,10.329918,10.295622,10.189304,9.983529,9.451943,8.632272,7.630832,7.085528,6.9209075,6.358455,4.8940215,4.1635194,3.7794054,3.5016088,3.2443898,3.2306714,3.450165,3.9543142,4.6127954,5.120374,5.3707337,5.0620713,4.931747,5.305572,6.111525,6.9826403,8.128122,9.47938,10.943813,12.428825,14.263655,16.11906,17.21996,17.394867,17.075916,15.662926,13.954991,12.178465,10.772334,10.374502,11.080997,11.7257595,12.092726,11.989838,11.2593355,9.825768,8.820899,8.032094,7.3598948,6.8111606,6.8591747,6.5196457,5.717122,4.9488945,5.295283,6.1321025,7.2604365,8.361334,9.263316,9.925226,9.921797,9.609704,9.016385,8.186425,7.15069,5.892031,4.6848164,3.8617156,3.4947495,3.3952916,3.649081,4.262977,5.2815647,6.800872,8.985519,9.5205345,9.719451,9.379922,8.80718,8.800322,9.2153015,7.6514096,5.785714,4.513337,3.9303071,3.7553983,3.7691166,3.7794054,3.673088,3.40901,3.649081,4.540774,5.1512403,5.329579,5.6965446,5.9331865,5.6142344,5.2781353,4.979761,4.2869844,4.4413157,4.6436615,4.605936,4.506478,4.979761,6.944915,9.9869585,12.744347,14.212211,13.756075,15.076467,15.79325,13.498857,9.455373,8.577398,10.179015,12.915827,14.637479,14.339106,12.154458,10.765475,10.6488695,11.780633,13.011855,12.099585,11.900668,12.79922,12.075578,9.421077,6.9380555,6.4887795,7.997798,9.757176,10.683165,10.343636,9.102125,8.450503,9.445084,11.314209,11.444533,9.331907,9.417647,11.80121,16.098484,21.428062,23.077694,21.990515,18.54035,15.014734,15.594335,17.082775,17.343424,15.782962,12.758065,9.571979,9.702303,10.508256,11.64345,12.63117,12.854094,11.845795,10.439664,9.249598,8.344186,7.2295704,5.809721,4.616225,3.7211025,3.210094,3.1860867,3.292404,3.433017,3.4913201,3.525616,3.765687,4.2252517,4.7842746,5.1992545,5.3878818,5.411889,5.7925735,6.252138,6.831738,7.8126,9.6988735,11.540562,12.569438,12.572867,11.739478,10.6488695,9.427936,8.594546,8.008087,7.6376915,7.5450926,7.7577267,7.9429245,8.011517,8.114404,8.669997,9.56512,9.56512,9.266746,9.016385,8.906639,8.220721,7.6171136,6.9723516,6.341307,5.9571934,5.970912,6.701414,7.407909,7.6342616,7.1781263,5.8337283,5.411889,5.5250654,5.8508763,6.1286726,5.796003,5.195825,5.302142,6.258997,7.3873315,8.776315,8.4093485,7.4353456,6.5162163,5.826869,5.761707,5.5833683,5.1855364,4.629943,4.1360826,3.9508848,4.1155047,3.99204,3.4295874,2.7745364,2.8637056,2.6545007,2.352697,2.16064,2.311542,2.2086544,1.99602,1.8965619,1.8931323,1.7182233,1.3306799,1.1043272,1.0014396,0.9945804,1.0700313,0.9259886,0.75450927,0.7407909,0.83681935,0.7613684,0.6241849,0.6859175,0.8093826,0.9328478,1.0425946,0.6824879,0.42183927,0.23664154,0.13032432,0.1371835,0.14404267,0.11317638,0.116605975,0.16804978,0.21263443,0.1920569,0.15433143,0.12346515,0.09259886,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.006859175,0.017147938,0.024007112,0.024007112,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044584636,0.044584636,0.061732575,0.061732575,0.037725464,0.0,0.034295876,0.05144381,0.034295876,0.006859175,0.006859175,0.041155048,0.048014224,0.048014224,0.044584636,0.041155048,0.061732575,0.07545093,0.11317638,0.18176813,0.26064864,0.19891608,0.17833854,0.18176813,0.18519773,0.18862732,0.22978236,0.25378948,0.2503599,0.22978236,0.22635277,0.20920484,0.20577525,0.19891608,0.18519773,0.16119061,0.16804978,0.16804978,0.16119061,0.14747226,0.13032432,0.1097468,0.10288762,0.12346515,0.16804978,0.21263443,0.216064,0.1920569,0.15090185,0.106317215,0.08573969,0.07888051,0.082310095,0.09259886,0.106317215,0.1097468,0.08916927,0.082310095,0.07888051,0.07888051,0.06516216,0.05144381,0.044584636,0.048014224,0.06516216,0.082310095,0.09602845,0.09602845,0.11317638,0.14747226,0.18519773,0.20577525,0.20234565,0.17490897,0.14404267,0.14404267,0.16119061,0.16804978,0.16462019,0.15776102,0.16119061,0.15433143,0.1371835,0.12003556,0.12689474,0.1920569,0.26064864,0.28465575,0.26407823,0.2194936,0.17833854,0.1371835,0.14404267,0.17833854,0.23321195,0.30866286,0.35324752,0.4115505,0.4389872,0.44584638,0.5007198,0.53501564,0.5178677,0.5144381,0.5590228,0.66191036,1.0906088,1.4507155,1.7765263,2.0234566,2.0817597,2.0920484,2.287535,2.386993,2.3561265,2.386993,2.469303,3.0077481,3.724532,4.3178506,4.4447455,4.8768735,5.411889,5.994919,6.5779486,7.1129646,7.449064,7.6376915,7.747438,7.8434668,8.011517,8.889491,9.431366,9.496528,9.458802,10.206452,10.912948,11.115293,10.659158,9.647429,8.4264965,7.5039372,6.6739774,5.7068334,4.5922174,3.5702004,2.9151495,2.4727325,2.201795,2.095478,2.177788,2.5070283,2.0714707,1.471293,1.1043272,1.196926,1.1008976,0.99801,0.9602845,1.0254467,1.2072148,1.5364552,1.9068506,2.0440342,1.862266,1.4575747,1.4404267,1.4369972,1.4644338,1.4095604,1.0425946,0.7373613,0.59674823,0.66876954,0.90541106,1.1420527,0.96371406,0.8505377,0.8093826,0.88826317,1.1763484,1.0940384,0.78194594,0.45956472,0.25378948,0.20920484,0.15776102,0.25721905,0.38754338,0.47671264,0.4938606,0.29494452,0.09602845,0.017147938,0.041155048,0.030866288,0.006859175,0.020577524,0.11317638,0.28808534,0.51100856,0.36696586,0.25721905,0.1920569,0.20234565,0.32924038,0.4698535,0.6036074,0.59331864,0.432128,0.24350071,0.17490897,0.13032432,0.10288762,0.09259886,0.09259886,0.07888051,0.048014224,0.041155048,0.061732575,0.082310095,0.12346515,0.17490897,0.24350071,0.33952916,0.48357183,0.7099246,0.94656616,1.1626302,1.2758065,1.1523414,0.9328478,0.7922347,1.1489118,2.1469216,3.6593697,5.6965446,7.2467184,8.203573,9.108984,11.1393,12.000127,10.88551,8.951223,7.0306544,5.6245236,6.0154963,6.2418494,6.358455,6.684266,7.8126,8.851766,9.794902,12.055,15.275383,17.350283,17.29198,17.562918,17.010754,14.953001,11.183885,11.80464,12.908967,14.081886,14.839825,14.651197,13.570878,12.7272,12.1921835,12.020704,12.229909,12.325937,12.679185,13.293081,14.246507,15.693792,16.45516,16.63007,16.427725,16.064188,15.734947,15.923574,15.371411,14.29795,12.80608,10.882081,9.266746,7.997798,6.5950966,5.086078,4.0023284,3.3781435,2.5481834,1.728512,1.0494537,0.548734,0.41840968,0.42183927,0.53158605,0.66876954,0.6824879,0.65848076,0.65162164,0.66533995,0.6927767,0.72707254,0.8128122,0.90884066,1.0151579,1.138623,1.2689474,1.4198492,1.605047,2.0063086,2.651071,3.3850029,4.2698364,5.295283,6.5162163,8.080108,10.237319,12.38424,14.476289,16.259674,17.851004,19.740705,21.78817,22.52896,22.474087,21.860191,20.632399,18.416885,16.29054,14.514014,13.327377,12.946692,13.241637,14.05102,14.675205,14.812388,14.565458,14.935853,15.388559,15.690363,15.851553,16.149927,15.916716,15.350834,14.733508,14.157337,13.533153,12.034423,10.81006,9.719451,8.796892,8.237869,7.9909387,7.7097125,7.610255,7.675417,7.64798,7.6033955,7.3221693,7.1369715,7.010077,6.5333643,5.703404,5.188966,4.7362604,4.2115335,3.6216443,3.199805,3.316411,3.7211025,4.2218223,4.698535,5.0277753,5.0414934,5.0483527,5.2506986,5.7754254,6.451054,7.380472,9.06097,11.413667,13.786942,15.405707,17.425734,19.143957,19.771572,18.440891,16.527182,14.575747,12.881531,11.629731,10.926665,10.563129,11.094715,11.931535,12.723769,13.392539,12.607163,11.756626,10.683165,9.421077,8.200144,7.421627,7.2021337,6.6739774,5.7102633,4.9351764,5.0140567,5.5387836,6.3893213,7.4353456,8.522525,9.355915,10.072699,10.055551,9.246168,8.1384115,6.893471,5.970912,5.3398676,4.7671266,3.7965534,3.5359046,3.7382503,4.482471,5.6656785,6.999788,7.380472,8.05953,8.570539,8.89635,9.451943,9.417647,8.176137,6.557371,5.127233,4.2081037,3.6868064,3.7279615,3.9611735,4.170378,4.2938433,3.8960114,3.865145,3.758828,3.5702004,3.724532,4.2595477,4.73969,4.9180284,4.698535,4.149801,3.858286,4.413879,5.2506986,6.0326443,6.684266,7.1884155,8.083538,9.925226,11.931535,11.996697,11.050131,11.050131,10.041832,8.330468,8.460793,11.231899,13.450842,13.004995,10.237319,7.963502,6.8454566,6.8866115,7.73029,8.721441,8.906639,9.328478,10.14129,10.264755,9.589127,8.964942,8.604835,9.050681,9.993818,10.981539,11.427385,11.451392,11.297061,11.701753,12.46312,12.46998,10.587136,9.5033865,11.06042,14.843254,18.193962,18.921034,18.241976,16.311117,14.287662,14.315098,16.101913,16.70552,14.959861,11.677745,9.657719,10.117283,11.832077,13.927555,15.8138275,17.189093,17.487467,16.55119,14.819247,12.812939,11.1393,9.417647,7.8537555,6.5950966,5.7239814,5.2575574,5.2747054,5.127233,4.880303,4.6265135,4.482471,4.870014,5.521636,6.279575,6.975781,7.431916,7.857185,8.309891,8.838047,9.568549,10.696883,12.421966,13.567448,13.618892,12.689473,11.519984,10.405369,9.863494,9.571979,9.3764925,9.294182,9.472521,9.619993,9.692014,9.853205,10.47396,10.501397,9.345626,8.361334,8.052671,8.090397,8.117833,8.090397,7.922347,7.613684,7.2432885,7.082098,7.239859,7.1369715,6.6739774,6.217842,5.641671,5.439326,5.4941993,5.669108,5.7994323,5.442755,5.15467,5.638242,6.691125,7.222711,7.6171136,7.6959944,7.486789,7.0546613,6.5196457,5.892031,5.453044,5.096367,4.629943,3.7759757,3.3747141,3.4124396,3.2958336,2.843128,2.2909644,1.99602,1.7662375,1.6359133,1.6736387,1.9754424,1.9239986,1.7216529,1.5673214,1.488441,1.3341095,1.0700313,0.90198153,0.8025235,0.7476501,0.7339317,0.67219913,0.64476246,0.72364295,0.86082643,0.881404,0.8265306,0.8025235,0.85396725,0.97400284,1.1008976,0.58302987,0.25721905,0.09602845,0.061732575,0.10288762,0.1371835,0.13032432,0.13032432,0.14061308,0.15090185,0.116605975,0.08573969,0.061732575,0.048014224,0.01371835,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.024007112,0.020577524,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07545093,0.082310095,0.07888051,0.07545093,0.061732575,0.030866288,0.024007112,0.048014224,0.048014224,0.030866288,0.024007112,0.058302987,0.072021335,0.06859175,0.06859175,0.07888051,0.08573969,0.09602845,0.12346515,0.16804978,0.22292319,0.22978236,0.26407823,0.29837412,0.30866286,0.29151493,0.28808534,0.28808534,0.26064864,0.216064,0.18176813,0.16462019,0.15776102,0.16119061,0.16462019,0.15433143,0.15433143,0.14061308,0.12346515,0.09945804,0.08916927,0.09602845,0.09259886,0.106317215,0.1371835,0.15090185,0.15433143,0.13375391,0.10288762,0.07545093,0.06859175,0.06859175,0.07545093,0.09259886,0.106317215,0.10288762,0.08573969,0.072021335,0.06859175,0.06859175,0.06859175,0.061732575,0.058302987,0.06516216,0.082310095,0.09945804,0.116605975,0.12346515,0.13375391,0.14747226,0.16804978,0.18862732,0.1920569,0.17147937,0.14061308,0.12346515,0.12689474,0.14061308,0.12689474,0.09602845,0.09602845,0.11317638,0.09945804,0.08573969,0.09259886,0.12003556,0.18862732,0.24350071,0.26407823,0.24350071,0.20234565,0.14404267,0.13032432,0.15776102,0.20920484,0.2709374,0.26750782,0.29494452,0.34638834,0.42526886,0.548734,0.607037,0.58988905,0.6173257,0.75450927,1.0357354,1.646202,1.9925903,2.177788,2.2978237,2.4247184,2.5481834,2.6236343,2.503599,2.270387,2.2155135,2.411,2.8808534,3.4124396,3.82399,3.9508848,4.273266,4.73969,5.360445,6.012067,6.4716315,7.15069,8.018375,8.752307,9.211872,9.445084,10.007536,9.908078,9.22216,8.656279,9.571979,10.120712,10.251037,10.100135,9.668007,8.803751,7.4353456,6.3378778,5.4496145,4.588788,3.4192986,2.8294096,2.4658735,2.1846473,2.0097382,2.1126258,2.6476414,2.2155135,1.5227368,1.039165,1.0117283,0.83338976,0.69963586,0.6927767,0.823101,1.0185875,1.2277923,1.6221949,1.7388009,1.4095604,0.7579388,0.83681935,0.94656616,1.0768905,1.1146159,0.8128122,0.58302987,0.5727411,0.70649505,0.89855194,1.0323058,0.8093826,0.6824879,0.61389613,0.7305021,1.3066728,1.3101025,0.96714365,0.64476246,0.47328308,0.34638834,0.36696586,0.47328308,0.5521636,0.5212973,0.35324752,0.18176813,0.0548734,0.0,0.0,0.0,0.044584636,0.06516216,0.14061308,0.3018037,0.53158605,0.35324752,0.23321195,0.18519773,0.2194936,0.33609957,0.4389872,0.4972902,0.44927597,0.29151493,0.1097468,0.07888051,0.058302987,0.041155048,0.041155048,0.0548734,0.048014224,0.034295876,0.05144381,0.09602845,0.12003556,0.09602845,0.116605975,0.18176813,0.31895164,0.58645946,0.8025235,1.0494537,1.3169615,1.4918705,1.3478279,1.0288762,1.1934965,1.9823016,3.4433057,5.5250654,7.130112,8.210432,8.81061,9.4862385,11.303921,11.619442,9.403929,7.2192817,6.183546,5.977771,6.0566516,5.874883,5.6656785,6.0840883,8.22758,9.911508,11.190743,14.020154,17.916164,19.980776,18.632948,17.655516,16.585485,15.271953,13.876111,15.271953,17.065628,17.473747,16.177364,14.315098,12.830087,12.22648,12.116733,12.274493,12.634601,12.229909,12.027563,12.168177,12.792361,14.027013,15.165636,15.693792,15.741806,15.488017,15.148488,15.121051,14.246507,12.7272,10.779194,8.625413,7.267296,6.3618846,5.3261495,4.1017866,3.1517909,2.760818,2.0920484,1.3101025,0.61389613,0.274367,0.18862732,0.17490897,0.22292319,0.28808534,0.29837412,0.28122616,0.20920484,0.20234565,0.274367,0.34295875,0.39097297,0.44584638,0.5144381,0.61046654,0.77508676,0.9842916,1.1489118,1.430138,1.8897027,2.49331,3.3369887,4.197815,5.103226,6.2555676,8.021805,9.822338,11.616013,13.011855,14.099034,15.45715,17.717249,19.20569,20.176264,20.519222,19.754423,17.885298,15.697222,13.708061,12.243628,11.430815,11.430815,11.934964,12.397959,12.6929035,13.118172,13.893259,14.260224,14.363112,14.490007,15.069608,15.697222,15.916716,15.940722,15.71094,14.88441,12.902108,11.149589,9.578837,8.31332,7.6616983,7.1369715,6.358455,5.751418,5.456474,5.3330083,5.5730796,5.7239814,5.7925735,5.826869,5.9160385,6.029215,5.844017,5.4324665,4.870014,4.2252517,3.7519686,3.6970954,3.7862647,3.9646032,4.3933015,4.8254294,5.2918534,5.5079174,5.552502,5.861165,6.81802,7.8949103,9.568549,11.729189,13.677195,15.285671,17.357141,19.239986,20.141968,19.12681,17.813278,15.707511,13.7526455,12.394529,11.578287,10.854645,11.074138,11.763485,12.710052,13.9481325,13.954991,13.320518,12.05843,10.343636,8.522525,7.1541195,6.8728933,6.931196,6.7700057,6.025785,5.672538,5.360445,5.5490727,6.307011,7.298162,8.64599,9.918367,10.4533825,10.079557,9.122703,8.296172,7.864044,7.613684,7.2021337,6.1629686,5.425607,4.770556,4.5270553,4.715683,5.0655007,5.456474,6.557371,7.905199,9.030104,9.445084,8.937505,8.56368,7.829748,6.660259,5.40503,4.2355404,3.882293,4.0777793,4.557922,5.0757895,4.715683,3.858286,3.1723683,3.000889,3.3541365,3.8171308,4.32471,4.5819287,4.5682106,4.557922,4.437886,4.8254294,5.545643,6.3618846,6.9826403,7.1369715,7.14726,8.141841,9.613133,9.407358,6.9517736,6.23499,6.560801,7.442205,8.587687,10.803201,12.164746,11.345076,8.862054,7.0958166,6.108095,5.672538,5.6793966,6.0737996,6.8283086,7.3255987,7.9292064,8.529384,9.084977,9.599416,9.469091,9.647429,10.429376,11.516555,12.034423,12.343085,12.435684,12.363663,12.199042,12.048141,10.683165,9.259886,9.551401,11.533703,13.368532,14.099034,13.728639,12.607163,11.293632,10.556271,11.934964,13.087306,12.614022,10.744898,9.342196,9.849775,11.8115,14.400838,16.849564,18.434032,18.670673,18.04649,16.527182,14.534592,12.950122,12.044711,10.672876,8.985519,7.48336,6.992929,7.2432885,7.449064,7.5725293,7.610255,7.582818,7.5519514,7.671987,7.936065,8.255017,8.48137,8.543102,8.618553,8.848335,9.239308,9.6645775,10.624862,11.358793,11.499407,11.159878,10.940384,10.9198065,11.279913,11.592006,11.742908,11.900668,12.281353,12.394529,12.308789,12.116733,11.921246,11.375941,10.251037,9.256456,8.7283,8.615124,8.98209,8.875772,8.748878,8.759167,8.752307,8.752307,8.745448,8.354475,7.606825,6.9620624,6.8626046,6.7219915,6.5813785,6.420188,6.169828,5.8817425,5.8337283,6.200694,6.667118,6.385892,6.307011,6.948344,7.5690994,7.7680154,7.514226,6.2384195,5.425607,4.99005,4.6779575,4.0674906,3.707384,3.5976372,3.3987212,3.0146074,2.5893385,2.1297739,1.7765263,1.5330256,1.4267083,1.5227368,1.4232788,1.2449403,1.0631721,0.91569984,0.7888051,0.6927767,0.6276145,0.58302987,0.5555932,0.52472687,0.59674823,0.70649505,0.85739684,1.0425946,1.2415106,1.2860953,1.1043272,0.96714365,0.9602845,0.9842916,0.5796003,0.33266997,0.22635277,0.22978236,0.28122616,0.31209245,0.31552204,0.29494452,0.25721905,0.20577525,0.15776102,0.116605975,0.08573969,0.061732575,0.037725464,0.020577524,0.010288762,0.0034295875,0.0034295875,0.010288762,0.024007112,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.061732575,0.072021335,0.072021335,0.072021335,0.07545093,0.09259886,0.07888051,0.07545093,0.082310095,0.08573969,0.07545093,0.08573969,0.09259886,0.09602845,0.1097468,0.16119061,0.13375391,0.13375391,0.14404267,0.16119061,0.2194936,0.28465575,0.34981793,0.40126175,0.42526886,0.40126175,0.32924038,0.30523327,0.28122616,0.23664154,0.17833854,0.15090185,0.14061308,0.14747226,0.15776102,0.13032432,0.1097468,0.09945804,0.08916927,0.072021335,0.06516216,0.09602845,0.106317215,0.11317638,0.116605975,0.09945804,0.09259886,0.08916927,0.08573969,0.07888051,0.07888051,0.07545093,0.082310095,0.09259886,0.09945804,0.11317638,0.09945804,0.08573969,0.06859175,0.061732575,0.061732575,0.061732575,0.072021335,0.08916927,0.1097468,0.13375391,0.17490897,0.20234565,0.20234565,0.17490897,0.1371835,0.15433143,0.20920484,0.23664154,0.2194936,0.17833854,0.16804978,0.15433143,0.12003556,0.08573969,0.12003556,0.1371835,0.116605975,0.09259886,0.082310095,0.09259886,0.1371835,0.19548649,0.2469303,0.26750782,0.23321195,0.18862732,0.15090185,0.15090185,0.18519773,0.2194936,0.22635277,0.28808534,0.37725464,0.47328308,0.58645946,0.6344737,0.6756287,0.7956643,1.0700313,1.546744,2.2635276,2.668219,2.8568463,2.8980014,2.8156912,2.8739944,2.8294096,2.603057,2.311542,2.277246,2.3972816,2.5927682,2.9151495,3.357566,3.8685746,4.245829,4.773986,5.4599032,6.0532217,6.0532217,6.427047,7.514226,8.711152,9.695444,10.4533825,10.563129,10.2236,9.499957,8.851766,9.126132,8.923786,8.217292,8.158989,8.762596,8.906639,8.251588,7.0923867,5.7239814,4.3590055,3.1380725,2.603057,2.218943,1.9514352,1.7730967,1.6873571,1.6667795,1.5776103,1.3889829,1.1214751,0.84367853,0.6173257,0.44584638,0.4046913,0.51100856,0.70649505,0.8676856,0.99801,0.99801,0.8505377,0.6241849,0.5796003,0.5727411,0.5761707,0.5590228,0.490431,0.5178677,0.64819205,0.85396725,1.0666018,1.155771,0.89169276,0.8196714,0.7990939,0.88826317,1.3375391,1.5090185,1.4850113,1.1077567,0.5555932,0.34638834,0.7133542,0.864256,0.89855194,0.8025235,0.45270553,0.22635277,0.06859175,0.0,0.0,0.0,0.12346515,0.12346515,0.14061308,0.22978236,0.3806842,0.24350071,0.18519773,0.216064,0.30866286,0.42869842,0.4629943,0.37725464,0.26064864,0.14404267,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.030866288,0.06516216,0.09259886,0.09602845,0.048014224,0.08916927,0.20234565,0.4081209,0.77165717,1.0906088,1.4129901,1.7250825,1.9102802,1.7730967,1.3443983,1.7730967,2.8328393,4.448175,6.725421,7.191845,7.6205435,8.31332,9.115844,9.414218,8.968371,7.0375133,5.98463,6.632822,8.255017,7.3530354,6.8214493,6.708273,7.3598948,9.441654,11.05356,12.096155,13.533153,15.498305,17.326277,17.480608,16.846134,15.981877,15.608052,16.61292,17.936743,19.092514,17.508043,13.708061,11.293632,11.135871,11.413667,11.760056,11.993267,12.120162,11.777204,11.499407,11.574858,12.130451,13.145609,14.2533655,14.675205,14.664916,14.3974085,13.982429,12.898679,11.513125,9.846346,8.1384115,6.835168,5.778855,4.931747,4.1429415,3.3678548,2.6613598,2.1812177,1.5227368,0.78537554,0.22292319,0.2194936,0.216064,0.20234565,0.20234565,0.2194936,0.24350071,0.2503599,0.11317638,0.020577524,0.030866288,0.08916927,0.1371835,0.17833854,0.21263443,0.28808534,0.4698535,0.65162164,0.7476501,0.90198153,1.1900668,1.6324836,2.3664153,3.1415021,3.9063,4.770556,5.9983487,7.425057,8.81061,9.925226,10.751757,11.499407,13.183334,14.887839,16.602633,17.895588,17.902447,17.134218,15.549749,13.814379,12.298501,11.070708,10.744898,10.710602,10.9541025,11.646879,13.169616,13.958421,14.366542,14.5414505,14.685493,15.028452,15.741806,16.153357,16.167076,15.666355,14.5414505,13.145609,11.595435,10.045261,8.718011,7.936065,7.5210853,6.550512,5.504488,4.647091,4.0229063,3.940596,3.9886103,4.0674906,4.2698364,4.880303,5.3878818,5.3981705,5.1992545,4.945465,4.6573796,4.5682106,4.372724,4.105216,3.9611735,4.297273,4.8014226,5.562791,5.960623,5.994919,6.279575,7.548522,8.820899,10.172156,11.413667,12.092726,13.810948,15.988737,17.717249,18.62609,18.897026,18.526632,16.520323,14.311668,12.826657,12.507706,12.229909,12.199042,12.30536,12.583157,13.200482,13.639469,13.3033695,12.21619,10.4705305,8.2310095,6.56766,5.8817425,6.334448,7.3839016,7.7714453,7.31531,6.3481665,5.844017,6.0978065,6.7391396,8.165848,9.304471,10.113853,10.408798,9.866923,9.527394,9.465661,9.55826,9.637141,9.5033865,8.669997,7.301592,5.8817425,4.8597255,4.650521,5.1409516,6.025785,7.2021337,8.220721,8.285883,7.9086285,8.244728,8.433355,8.025234,6.9792104,5.518206,4.3624353,3.9680326,4.297273,4.8494368,5.0757895,4.1120753,3.2889743,3.1620796,3.4981792,3.8377085,4.1017866,4.266407,4.431027,4.822,5.188966,5.267846,5.3090014,5.4599032,5.7582774,5.9469047,6.029215,6.1972647,6.461343,6.6636887,6.5196457,6.042933,6.111525,6.869464,7.716572,8.416207,9.187865,9.403929,8.820899,7.5862474,6.5230756,5.73427,5.1409516,4.7774153,4.7774153,5.0003386,5.5387836,6.169828,6.8626046,7.7714453,7.874333,8.899779,10.576848,12.079007,12.044711,11.763485,11.519984,11.166737,10.72089,10.377932,9.582268,8.89635,8.399059,8.505377,9.962952,11.396519,11.516555,10.30934,8.457363,7.3564653,7.8091707,9.321619,10.72089,11.036412,9.513676,9.914937,11.249047,13.519434,15.954441,16.986746,15.844694,14.802099,13.906977,13.070158,12.05157,12.116733,11.2593355,9.489669,7.671987,7.5245147,8.025234,8.707723,9.438225,10.106995,10.635151,10.220171,9.712592,9.084977,8.412778,7.864044,7.4010496,6.992929,6.9037595,7.140401,7.438775,7.438775,7.5759587,7.81603,8.2653055,9.177576,10.432805,11.7086115,12.672326,13.251926,13.677195,14.205351,14.30481,14.040731,13.399398,12.295071,11.8869505,11.80464,11.417097,10.748327,10.48082,10.583707,9.829198,9.218731,9.163857,9.462232,9.8429165,10.230459,10.398509,10.2236,9.674867,9.270175,8.937505,8.632272,8.268735,7.7131424,7.3427467,7.0546613,6.9209075,6.7974424,6.3447366,6.557371,7.2878733,7.98065,8.296172,8.141841,6.7528577,6.0052075,5.6245236,5.4667625,5.5250654,5.3707337,5.0106273,4.4516044,3.789694,3.1826572,2.7779658,2.3629858,1.9891608,1.6839274,1.4335675,1.2209331,1.0425946,0.90198153,0.7956643,0.72021335,0.6893471,0.67219913,0.66876954,0.6927767,0.75450927,0.8745448,1.0117283,1.1866373,1.4129901,1.7010754,1.7182233,1.3958421,1.0563129,0.8265306,0.65162164,0.5453044,0.5007198,0.5178677,0.5727411,0.65162164,0.66876954,0.64476246,0.59331864,0.53158605,0.45270553,0.37382504,0.30523327,0.24007112,0.17147937,0.09259886,0.05144381,0.024007112,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.07888051,0.116605975,0.15090185,0.14061308,0.1371835,0.1371835,0.1371835,0.1371835,0.1371835,0.12689474,0.12346515,0.1371835,0.19891608,0.15090185,0.18176813,0.20234565,0.19548649,0.24350071,0.28122616,0.30866286,0.34638834,0.37725464,0.36696586,0.34295875,0.30866286,0.26407823,0.21263443,0.15090185,0.116605975,0.12346515,0.14404267,0.14404267,0.106317215,0.09602845,0.072021335,0.061732575,0.06516216,0.07545093,0.08916927,0.09945804,0.11317638,0.11317638,0.07545093,0.07545093,0.07545093,0.082310095,0.09259886,0.09259886,0.07888051,0.07545093,0.06859175,0.06516216,0.07545093,0.06516216,0.06859175,0.06859175,0.061732575,0.061732575,0.061732575,0.07888051,0.09259886,0.09602845,0.12346515,0.18176813,0.24350071,0.28808534,0.28465575,0.19891608,0.23664154,0.34638834,0.38754338,0.33952916,0.29151493,0.2777966,0.22978236,0.15433143,0.09602845,0.106317215,0.106317215,0.08916927,0.082310095,0.09259886,0.09259886,0.07888051,0.12346515,0.18176813,0.23321195,0.24350071,0.2194936,0.19548649,0.19548649,0.23321195,0.30523327,0.39097297,0.45613512,0.52472687,0.61046654,0.7339317,0.82996017,0.91912943,1.0151579,1.1797781,1.5090185,1.961724,2.5413244,2.9803114,3.1826572,3.2203827,3.5016088,3.5050385,3.2272418,2.8499873,2.7779658,2.7539587,2.7642474,2.9220085,3.223812,3.5393343,3.9543142,4.5167665,5.137522,5.7136927,6.1046658,6.444195,6.8969,7.599966,8.4264965,8.988949,9.06097,10.278474,11.4205265,11.396519,9.263316,9.177576,9.760606,10.467101,10.748327,10.041832,8.282454,6.608815,5.1100855,3.9063,3.1140654,2.4418662,1.8348293,1.6324836,1.7730967,1.786815,1.7353712,2.1469216,2.2498093,1.7593783,0.85396725,0.70649505,0.607037,0.5521636,0.5624523,0.67219913,0.82996017,0.99801,1.1934965,1.3684053,1.4027013,0.90198153,0.6790583,0.64133286,0.66191036,0.5658819,0.69963586,1.0151579,1.371835,1.6324836,1.6942163,1.3409687,1.3341095,1.430138,1.4232788,1.1283343,1.313532,1.5673214,1.2860953,0.6036074,0.39783216,0.7613684,0.34295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17147937,0.17833854,0.15776102,0.18519773,0.26064864,0.2469303,0.28122616,0.35324752,0.4629943,0.61046654,0.6344737,0.4389872,0.24350071,0.1371835,0.07545093,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.09602845,0.12346515,0.15776102,0.26750782,0.44584638,0.7099246,1.1146159,1.4815818,1.8108221,1.9685832,1.9308578,1.786815,1.4438564,1.9994495,3.1346428,4.7979927,7.2021337,7.3358874,6.9963584,6.427047,5.960623,5.9983487,6.108095,4.979761,4.2183924,4.5682106,5.936616,6.6431108,7.4627824,8.669997,9.904649,10.161868,10.161868,10.326488,11.273054,13.190193,15.837835,17.473747,18.451181,19.013634,19.068506,18.187103,16.846134,14.918706,12.9809885,11.427385,10.4533825,10.878652,11.2250395,11.38966,11.348505,11.153018,11.348505,11.681175,12.298501,13.059869,13.533153,13.461131,12.627741,11.718901,11.2250395,11.444533,10.467101,9.115844,7.6685576,6.334448,5.2506986,4.307562,3.6799474,3.2032347,2.784825,2.3801336,1.5021594,0.84367853,0.432128,0.24350071,0.18176813,0.2194936,0.20234565,0.19548649,0.2194936,0.24350071,0.17147937,0.12346515,0.09602845,0.08916927,0.1371835,0.18519773,0.116605975,0.07888051,0.14061308,0.274367,0.2503599,0.32581082,0.48014224,0.71678376,1.0837497,1.6804979,2.3972816,3.1243541,3.875434,4.791134,6.012067,6.701414,7.191845,7.689135,8.299602,9.352485,10.600855,12.151029,13.738928,14.740367,15.141628,14.63062,13.7697935,12.854094,11.900668,11.2421875,10.7757635,10.690024,10.984968,11.458252,12.144169,13.505715,14.754086,15.518884,15.824117,15.518884,14.901558,13.937843,12.867812,12.22305,11.63659,10.545981,9.496528,8.690575,7.9943686,7.5931067,6.8866115,5.977771,5.0346346,4.3041325,3.9851806,3.9611735,3.8205605,3.4878905,3.2203827,3.316411,3.525616,3.7759757,4.0091877,4.180667,4.314421,4.3761535,4.3349986,4.249259,4.273266,4.40702,4.897451,5.521636,6.0737996,6.3790326,6.5230756,7.267296,8.889491,10.847785,11.763485,12.922686,15.374841,17.54234,18.71183,19.044498,18.310568,17.103354,15.470869,14.033872,13.96185,14.167625,14.640909,14.640909,13.982429,13.032433,12.6757555,12.30536,12.092726,11.612583,9.8429165,8.1212635,6.8111606,6.9346256,8.285883,9.445084,8.419638,7.3221693,6.4544835,6.0052075,6.042933,7.2158523,8.505377,9.547972,10.172156,10.39165,9.914937,9.80519,9.846346,10.041832,10.590566,10.381361,9.764035,8.546532,7.0546613,6.1046658,5.8234396,6.0086374,6.2041235,6.1972647,6.025785,5.9914894,6.276145,6.975781,7.798882,8.042382,7.6616983,5.9400454,4.3933015,3.6525106,3.433017,3.542764,3.5153272,3.3644254,3.2409601,3.450165,3.5942078,3.7862647,3.9200184,4.0023284,4.149801,4.417309,4.650521,4.835718,5.086078,5.662249,6.0154963,6.1321025,6.3824625,6.8728933,7.4456344,7.7028537,7.64798,7.500508,7.2295704,6.5470824,7.301592,8.536243,9.6817255,10.052121,8.820899,6.632822,5.9126086,5.6828265,5.439326,5.1580997,4.791134,4.479041,4.029765,3.6216443,3.8308492,5.796003,8.594546,10.405369,10.494537,9.201583,8.858624,8.985519,9.266746,9.829198,11.245617,11.756626,10.834066,9.448513,8.279024,7.706283,8.999237,9.6817255,9.846346,9.39707,8.042382,8.004657,9.030104,10.281903,11.358793,12.298501,13.032433,13.224489,13.54687,14.191633,14.863832,13.166186,11.22161,10.336777,10.39165,9.8429165,8.608265,7.9257765,7.6925645,7.795452,8.086967,8.721441,8.934075,9.074688,9.280463,9.47595,9.403929,9.266746,8.8929205,8.268735,7.5210853,7.010077,6.5162163,6.1492505,5.936616,5.813151,5.813151,5.960623,6.210983,6.601956,7.2467184,8.591117,10.014396,11.523414,12.775213,13.090735,13.190193,13.423406,13.419975,13.114742,12.771784,12.295071,11.938394,11.537132,11.067279,10.652299,10.041832,9.321619,8.820899,8.64599,8.683716,8.827758,8.673427,8.687145,9.160428,10.2236,10.456812,10.621432,10.587136,10.340206,10.010965,9.410788,8.738589,8.361334,8.371623,8.591117,9.3593445,9.945804,9.657719,8.604835,7.689135,7.7748747,8.512236,9.091836,9.235879,9.201583,8.515666,7.1369715,5.7479887,4.6608095,3.8308492,3.2683969,2.8705647,2.5721905,2.3252604,2.1057668,1.9582944,1.8485477,1.7833855,1.7319417,1.646202,1.587899,1.5638919,1.5810398,1.6564908,1.8142518,1.8279701,1.7936742,1.786815,1.786815,1.6633499,1.4678634,1.2072148,0.939707,0.72707254,0.64133286,0.64133286,0.70649505,0.8025235,0.90541106,0.9911508,0.9911508,0.94656616,0.8711152,0.78194594,0.67219913,0.52472687,0.432128,0.35324752,0.2503599,0.09259886,0.030866288,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.05144381,0.116605975,0.15090185,0.16119061,0.14061308,0.15776102,0.20920484,0.19891608,0.18862732,0.14747226,0.12346515,0.13375391,0.17490897,0.22292319,0.25721905,0.25721905,0.23664154,0.25721905,0.31209245,0.31552204,0.29494452,0.26750782,0.25721905,0.3018037,0.30523327,0.26407823,0.19891608,0.17833854,0.16804978,0.15776102,0.14061308,0.12003556,0.09602845,0.082310095,0.06859175,0.06516216,0.072021335,0.06516216,0.06516216,0.07545093,0.08916927,0.09602845,0.08916927,0.08916927,0.07545093,0.06859175,0.07545093,0.06859175,0.06516216,0.072021335,0.06859175,0.061732575,0.06516216,0.05144381,0.05144381,0.05144381,0.05144381,0.061732575,0.072021335,0.07545093,0.08916927,0.1097468,0.13375391,0.17490897,0.20920484,0.22292319,0.20920484,0.16119061,0.23664154,0.33609957,0.40126175,0.41498008,0.37382504,0.28465575,0.22978236,0.18176813,0.13032432,0.09602845,0.09602845,0.09259886,0.09602845,0.10288762,0.10288762,0.1097468,0.1371835,0.17833854,0.22292319,0.25721905,0.28122616,0.29837412,0.31895164,0.33609957,0.32924038,0.34638834,0.4115505,0.53158605,0.70306545,0.90198153,1.1660597,1.4575747,1.7525192,1.9823016,2.0474637,2.294394,2.6922262,3.0660512,3.3438478,3.5359046,3.6216443,3.4467354,3.1517909,2.9220085,2.983741,3.2032347,3.474172,3.625074,3.6593697,3.7725463,3.9543142,4.1189346,4.3933015,4.8597255,5.5559316,6.677407,7.720001,8.464222,9.033533,9.877212,10.840926,10.172156,9.304471,8.899779,8.824328,8.423067,8.028665,7.7542973,7.346176,6.169828,4.715683,3.782835,3.199805,2.8808534,2.819121,2.5961976,2.301253,1.9823016,1.762808,1.8348293,1.6770682,1.8108221,1.704505,1.2243627,0.6344737,0.50757897,0.4046913,0.32581082,0.37039545,0.7442205,1.138623,1.6187652,1.821111,1.6599203,1.3546871,0.85396725,0.72364295,0.77508676,0.7888051,0.5144381,0.7956643,1.3478279,1.7525192,1.8965619,1.9857311,1.9754424,1.8931323,1.8039631,1.7662375,1.8245405,1.8519772,1.8142518,1.5433143,1.0768905,0.66533995,0.33952916,0.10288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20920484,0.2709374,0.274367,0.2777966,0.2709374,0.30866286,0.33266997,0.33609957,0.33266997,0.34295875,0.32581082,0.2469303,0.16462019,0.09602845,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.05144381,0.16119061,0.29151493,0.5727411,0.6344737,0.58302987,0.58645946,0.881404,1.2758065,1.7456601,2.0268862,2.0474637,1.9308578,1.5913286,2.4590142,3.9611735,5.689686,7.421627,7.56567,7.298162,7.4799304,8.241299,8.999237,9.537683,8.652849,7.3118806,6.0223556,4.8014226,5.4016004,6.3173003,7.1849856,7.6651278,7.4524937,6.9826403,8.56368,10.573419,12.1921835,13.395968,13.042721,12.627741,12.377381,12.418536,12.782072,12.542002,11.321068,10.093276,9.3079,8.879202,10.545981,11.293632,11.087856,10.388221,10.151579,10.319629,10.820349,11.646879,12.586586,13.21763,12.528283,11.211322,9.541112,8.196714,8.272165,7.870903,7.130112,6.0978065,4.9488945,3.9783216,3.4878905,2.9288676,2.3389788,1.7799559,1.3169615,0.86082643,0.51100856,0.32238123,0.26064864,0.2194936,0.18862732,0.15090185,0.1371835,0.13032432,0.09602845,0.044584636,0.024007112,0.037725464,0.06859175,0.08916927,0.09945804,0.061732575,0.05144381,0.09259886,0.18862732,0.18519773,0.22978236,0.32924038,0.50757897,0.8162418,1.255229,1.9274281,2.6922262,3.4947495,4.3521466,5.329579,5.950334,6.258997,6.4098988,6.677407,7.160979,7.9120584,8.944365,10.1481495,11.286773,12.157887,12.538571,12.662037,12.620882,12.3533745,11.958971,11.430815,11.132441,11.153018,11.338216,11.982979,12.8197975,13.618892,14.153908,14.225929,14.064738,13.903547,13.509145,12.895248,12.308789,11.897239,11.334786,10.847785,10.607714,10.741467,9.764035,8.429926,6.999788,5.7102633,4.804852,4.2526884,3.9714622,3.8171308,3.7313912,3.7451096,3.3644254,3.0626216,2.942586,3.07634,3.5221863,3.998899,4.012617,3.9783216,4.125794,4.4927597,4.4996185,4.695105,5.1340923,5.6965446,6.108095,6.608815,7.531374,8.683716,9.884071,10.995257,12.857523,14.479718,15.680074,16.595774,17.689812,18.235117,18.084215,17.062197,15.549749,14.510585,15.100473,15.683503,15.9613,15.608052,14.277372,13.745787,13.821238,14.105893,13.96871,12.55229,9.578837,7.716572,6.773435,6.543653,6.783724,6.7357097,6.6636887,6.2212715,5.610805,5.579939,6.427047,7.682276,8.803751,9.534253,9.89093,9.668007,9.431366,9.22216,9.280463,10.065839,10.707172,10.525404,9.740028,8.525954,7.006647,6.3447366,6.090947,5.8337283,5.442755,5.086078,5.0620713,5.3981705,6.3961806,7.936065,9.469091,9.187865,8.025234,6.327589,4.7671266,4.32471,4.190956,4.3281393,4.245829,3.8548563,3.4981792,2.959734,2.836269,3.0523329,3.4810312,3.9303071,4.2595477,4.341858,4.3109913,4.262977,4.280125,4.4413157,4.6916757,4.979761,5.3090014,5.7377,6.0532217,6.3653145,6.81802,7.332458,7.596536,7.6788464,8.838047,9.829198,9.952662,9.050681,7.949784,7.034084,6.5813785,6.557371,6.5985265,6.5333643,6.1801167,5.56965,4.8322887,4.2081037,5.2575574,6.0737996,6.2075534,5.645101,4.8185706,4.400161,4.5990767,4.928317,5.329579,6.166398,8.371623,9.523964,10.124143,10.511685,10.854645,11.327928,11.818358,11.8115,11.187314,10.213311,9.873782,9.925226,10.100135,10.364213,10.8958,11.578287,12.140739,13.018714,14.208781,15.241087,15.066177,13.834956,12.116733,10.244178,8.279024,7.6033955,7.8194594,8.158989,8.186425,7.795452,7.7268605,7.442205,7.143831,7.06495,7.473071,7.9772205,8.351046,8.3922,8.093826,7.630832,7.2947326,6.9826403,6.677407,6.3481665,5.970912,5.7754254,5.751418,5.8988905,6.1801167,6.5024977,6.9689217,7.48336,8.241299,9.22902,10.261326,11.413667,12.555719,13.708061,15.066177,17.017612,17.69667,16.849564,15.357693,13.697772,11.945253,10.717461,9.777754,9.218731,8.937505,8.632272,8.241299,7.534804,7.034084,7.0306544,7.5759587,8.255017,8.81404,9.122703,9.088407,8.64256,8.680285,8.772884,8.844906,8.913498,9.102125,8.954653,8.543102,8.090397,7.781734,7.7748747,8.467651,9.156999,9.270175,8.7283,7.932636,6.917478,5.8337283,4.8768735,4.15323,3.683377,3.4913201,3.4227283,3.4844608,3.5770597,3.4844608,3.3781435,3.3198407,3.2203827,3.0214665,2.7230926,2.435007,2.253239,2.1297739,2.0234566,1.8897027,1.7353712,1.6084765,1.5158776,1.4438564,1.371835,1.1454822,0.8848336,0.70649505,0.65162164,0.70306545,0.77851635,0.9362774,1.1317638,1.2895249,1.2963841,1.1489118,0.980862,0.823101,0.69963586,0.59674823,0.5212973,0.41498008,0.29151493,0.16804978,0.07888051,0.048014224,0.030866288,0.024007112,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.030866288,0.020577524,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.044584636,0.06859175,0.09602845,0.12003556,0.13375391,0.14061308,0.12003556,0.12346515,0.16804978,0.21263443,0.20920484,0.16119061,0.15090185,0.18176813,0.20577525,0.2194936,0.25378948,0.2777966,0.29151493,0.30523327,0.30866286,0.28465575,0.25378948,0.23321195,0.22978236,0.274367,0.24350071,0.1920569,0.15776102,0.14747226,0.12346515,0.106317215,0.09602845,0.08916927,0.072021335,0.037725464,0.044584636,0.05144381,0.05144381,0.061732575,0.11317638,0.09602845,0.082310095,0.116605975,0.20920484,0.1097468,0.08573969,0.08573969,0.082310095,0.06859175,0.06859175,0.07545093,0.06859175,0.061732575,0.06859175,0.06516216,0.048014224,0.041155048,0.05144381,0.06859175,0.082310095,0.08573969,0.082310095,0.082310095,0.09259886,0.106317215,0.11317638,0.18176813,0.30523327,0.40126175,0.28122616,0.36696586,0.5693115,0.72364295,0.59674823,0.45270553,0.33952916,0.25721905,0.20577525,0.16462019,0.15090185,0.16462019,0.18519773,0.1920569,0.17147937,0.23321195,0.33952916,0.40126175,0.4081209,0.41498008,0.4355576,0.41840968,0.38754338,0.35324752,0.30866286,0.4046913,0.5693115,0.77508676,1.0151579,1.2929544,1.6633499,1.8313997,1.961724,2.1297739,2.318401,2.6236343,2.9082901,3.0146074,2.9803114,3.059192,3.1620796,3.210094,3.1723683,3.059192,2.9460156,3.0660512,3.234101,3.3609958,3.4844608,3.765687,4.0709205,4.122364,4.2698364,4.6779575,5.3432975,6.0532217,6.807731,7.500508,8.361334,9.935514,11.773774,12.55229,12.346515,11.458252,10.425946,8.841476,7.490219,6.5024977,5.785714,5.020916,4.2183924,3.6765177,3.1895163,2.7093742,2.335549,2.1812177,2.0337453,1.8588364,1.7010754,1.6530612,1.5604624,1.6187652,1.5810398,1.3684053,1.0734608,0.78537554,0.5555932,0.3841138,0.36696586,0.6790583,0.9774324,1.2860953,1.8176813,2.3595562,2.277246,1.1180456,0.7339317,0.70649505,0.7133542,0.5590228,0.8745448,1.3649758,1.8759843,2.2292318,2.2258022,1.8142518,1.8999915,2.0131679,1.8828435,1.4575747,1.3443983,1.2758065,1.2175035,1.0734608,0.70649505,0.17490897,0.017147938,0.0,0.034295876,0.16462019,0.034295876,0.0,0.07888051,0.20920484,0.23664154,0.31895164,0.33952916,0.32581082,0.29151493,0.22978236,0.36696586,0.42526886,0.3841138,0.28122616,0.22978236,0.19548649,0.17147937,0.1371835,0.08573969,0.0,0.0,0.0,0.0034295875,0.006859175,0.0,0.0,0.06516216,0.18176813,0.33266997,0.490431,0.6344737,0.6859175,0.6893471,0.6859175,0.70649505,1.1214751,1.8554068,2.2498093,2.1469216,1.8691251,1.3649758,2.3835633,4.1360826,5.7925735,6.468202,6.8214493,7.1541195,8.1487,9.729739,11.06042,11.9040985,10.539123,8.340756,6.293293,4.9831905,5.4907694,6.4373355,7.4181976,8.025234,7.8194594,6.8454566,7.0752387,7.6857057,8.323608,9.115844,9.023245,8.834618,8.471081,8.158989,8.4264965,8.742019,8.608265,8.210432,7.596536,6.691125,8.344186,9.3079,9.187865,8.536243,8.841476,9.606275,10.347065,10.988399,11.434244,11.5645685,10.597425,9.678296,8.951223,8.440215,8.052671,7.380472,6.509357,5.4016004,4.1463714,2.9665933,2.784825,2.369845,1.7593783,1.1420527,0.84367853,0.58988905,0.34981793,0.216064,0.18519773,0.16462019,0.116605975,0.08573969,0.082310095,0.07888051,0.024007112,0.0034295875,0.0,0.010288762,0.024007112,0.030866288,0.05144381,0.048014224,0.041155048,0.0548734,0.10288762,0.15433143,0.23664154,0.33952916,0.4938606,0.7579388,1.1900668,1.7730967,2.4487255,3.210094,4.105216,4.880303,5.456474,5.7274113,5.768566,5.8508763,6.001778,6.550512,7.31531,8.158989,9.002667,9.609704,10.076128,10.576848,11.070708,11.303921,11.324498,11.204462,11.170166,11.31078,11.543991,12.164746,12.79922,13.371962,13.783512,13.896688,13.906977,13.821238,13.588025,13.231348,12.833516,12.788932,12.6586075,12.504276,12.264205,11.739478,10.439664,8.851766,7.332458,6.077229,5.137522,4.698535,4.448175,4.3487167,4.2595477,3.9474552,3.57363,3.5187566,3.4535947,3.3061223,3.2546785,3.3061223,3.4227283,3.7451096,4.249259,4.729401,4.7431192,4.6093655,4.722542,5.144381,5.6210938,6.3961806,7.4044795,8.519095,9.822338,11.581717,13.018714,13.786942,14.147048,14.562028,15.683503,17.772121,18.667244,18.598652,17.761833,16.304258,16.702091,17.463459,17.899017,17.573206,16.29054,14.726648,14.589465,14.843254,14.760944,13.896688,11.190743,9.054111,7.98065,7.6959944,7.143831,6.334448,6.540223,6.728851,6.5779486,6.468202,6.461343,6.7665763,7.431916,8.309891,9.06097,9.561689,10.100135,10.39508,10.463672,10.611144,11.091286,11.05356,10.545981,9.517105,7.8263187,6.601956,6.1046658,6.1972647,6.715132,7.4627824,6.447624,5.90232,5.967482,6.7048435,8.114404,8.635701,8.687145,7.9292064,6.608815,5.5730796,4.7774153,4.372724,4.081209,3.7691166,3.4364467,2.8019729,2.201795,2.2258022,2.9185789,3.7931237,4.7499785,5.1512403,5.195825,5.0243454,4.705394,4.6402316,4.715683,5.0312047,5.4736214,5.703404,5.470192,5.90575,6.667118,7.4284863,7.8846216,7.6685576,7.864044,8.261876,8.553391,8.351046,8.025234,7.6685576,7.5039372,7.56567,7.671987,7.7131424,7.56567,7.250148,6.8043017,6.2898636,6.3961806,6.464772,6.2898636,5.844017,5.288424,4.9008803,4.7774153,4.6573796,4.5099077,4.530485,5.4496145,6.4098988,7.599966,9.0644,10.700313,11.101575,11.921246,13.094165,14.246507,14.685493,14.490007,13.200482,12.024134,11.530273,11.650309,12.133881,12.96727,14.352823,15.824117,16.249386,16.20137,15.724659,14.46257,12.535142,10.542552,10.034973,9.925226,9.801761,9.458802,8.882631,8.450503,7.8503256,7.414768,7.3084507,7.5210853,7.870903,8.213862,8.440215,8.498518,8.3922,8.378482,8.405919,8.333898,8.107545,7.7680154,7.349606,6.992929,6.7528577,6.6876955,6.8557453,6.8454566,6.8454566,7.143831,7.8366075,8.855195,10.22703,11.533703,12.929544,14.589465,16.698662,17.559488,17.436022,16.726099,15.63206,14.153908,12.614022,11.358793,10.336777,9.489669,8.738589,8.282454,7.764586,7.407909,7.2124224,6.975781,6.8626046,6.944915,7.0272245,7.016936,6.927767,6.989499,7.205563,7.466212,7.73029,8.021805,7.8777623,7.06838,6.3378778,6.018926,6.001778,6.5367937,6.927767,6.9792104,6.6533995,6.077229,5.3501563,4.496189,3.8514268,3.4947495,3.2718265,3.1209247,3.0729103,3.100347,3.1312134,3.0351849,2.8980014,2.7916842,2.750529,2.7333813,2.6064866,2.3149714,2.0680413,1.8725548,1.7490896,1.7250825,1.5947582,1.4335675,1.5124481,1.8005334,1.9651536,1.8348293,1.4472859,1.0494537,0.82996017,0.94656616,1.1317638,1.3512574,1.4438564,1.3821237,1.255229,1.0700313,0.85396725,0.65162164,0.4938606,0.38754338,0.31895164,0.2503599,0.17490897,0.10288762,0.06859175,0.058302987,0.044584636,0.030866288,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.017147938,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072021335,0.08573969,0.1371835,0.14747226,0.116605975,0.12346515,0.13032432,0.12689474,0.13032432,0.15776102,0.2194936,0.20577525,0.17833854,0.18862732,0.23664154,0.2777966,0.26407823,0.26064864,0.28808534,0.33609957,0.34638834,0.2777966,0.2469303,0.24007112,0.24350071,0.22292319,0.22978236,0.18862732,0.15090185,0.14061308,0.12689474,0.08573969,0.05144381,0.041155048,0.044584636,0.037725464,0.006859175,0.017147938,0.034295876,0.048014224,0.06859175,0.09259886,0.082310095,0.07545093,0.1097468,0.20577525,0.106317215,0.08916927,0.09259886,0.09259886,0.12003556,0.08916927,0.07888051,0.06859175,0.061732575,0.058302987,0.058302987,0.044584636,0.041155048,0.0548734,0.06516216,0.072021335,0.072021335,0.06516216,0.058302987,0.06859175,0.061732575,0.05144381,0.116605975,0.25721905,0.3806842,0.24350071,0.32581082,0.53501564,0.71678376,0.6344737,0.5418748,0.44927597,0.37039545,0.30866286,0.26407823,0.23321195,0.22292319,0.2194936,0.20920484,0.18176813,0.28465575,0.42869842,0.52472687,0.5521636,0.5796003,0.6001778,0.53844523,0.47328308,0.4424168,0.42869842,0.548734,0.7579388,1.0288762,1.3272504,1.5981878,1.9068506,1.961724,2.0131679,2.1915064,2.503599,2.750529,2.8705647,2.7573884,2.534465,2.534465,2.668219,2.8945718,2.9906003,2.8808534,2.6407824,2.726522,2.8705647,3.07634,3.309552,3.5153272,3.7759757,3.865145,4.197815,4.856296,5.6073756,5.8371577,6.3138704,6.989499,7.846896,8.899779,10.988399,13.63604,14.057879,11.982979,9.661148,8.597976,7.0752387,5.586798,4.695105,5.0277753,4.6745276,3.9474552,3.1860867,2.551613,2.037175,2.0337453,1.903421,1.7456601,1.6256244,1.5673214,1.5604624,1.6016173,1.5227368,1.3101025,1.1043272,0.84367853,0.59674823,0.42869842,0.4355576,0.764798,1.1317638,1.4369972,1.8588364,2.2395205,2.0920484,0.94999576,0.6036074,0.5796003,0.58988905,0.5418748,0.91227025,1.3889829,1.9857311,2.4590142,2.3218307,1.5913286,1.6633499,1.8485477,1.7388009,1.2277923,1.0014396,0.8779744,0.85739684,0.8265306,0.5693115,0.17147937,0.17833854,0.28465575,0.36696586,0.5007198,0.37725464,0.36010668,0.45270553,0.5693115,0.52472687,0.42526886,0.37382504,0.35324752,0.34981793,0.36353627,0.39097297,0.3806842,0.31552204,0.21263443,0.12003556,0.09602845,0.09259886,0.07888051,0.05144381,0.0,0.0,0.0,0.006859175,0.024007112,0.037725464,0.048014224,0.14404267,0.2709374,0.39440256,0.5041494,0.490431,0.5418748,0.64133286,0.7510797,0.8196714,1.214074,1.862266,2.170929,2.0097382,1.7147937,1.1832076,2.136633,3.8857226,5.422178,5.4153185,6.169828,7.534804,8.872343,9.873782,10.528833,10.748327,9.318189,7.366754,5.936616,6.001778,6.6705475,7.455923,8.008087,8.124693,7.740579,6.883182,6.324159,6.1046658,6.341307,7.2535777,7.4970784,7.349606,6.9071894,6.358455,5.977771,5.579939,5.878313,6.1732574,5.9983487,5.096367,5.9400454,6.6053853,6.852316,7.006647,7.956643,9.331907,10.100135,10.422516,10.388221,10.024684,9.043822,8.354475,8.176137,8.241299,7.81603,7.250148,6.217842,4.9831905,3.7348208,2.5824795,2.4144297,2.0920484,1.5604624,0.9877212,0.72707254,0.5007198,0.32581082,0.22635277,0.17490897,0.1097468,0.08573969,0.06516216,0.06516216,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.041155048,0.0548734,0.061732575,0.06859175,0.072021335,0.13375391,0.21263443,0.31552204,0.4664239,0.6962063,1.2106444,1.7593783,2.386993,3.1380725,4.0846386,4.804852,5.3398676,5.5662203,5.5250654,5.411889,5.4496145,5.871454,6.478491,7.133542,7.750868,8.14527,8.457363,8.906639,9.47938,9.932085,10.329918,10.768905,11.297061,11.828648,12.144169,12.627741,13.070158,13.577737,14.105893,14.466,14.284232,13.893259,13.416546,13.063298,13.138749,13.13189,12.795791,12.538571,12.288212,11.509696,10.199594,8.80718,7.5416627,6.4716315,5.5113473,5.2266912,5.206114,5.127233,4.7945633,4.166949,3.6765177,3.7108135,3.758828,3.590778,3.275256,3.069481,3.1860867,3.5976372,4.139512,4.4927597,4.4687524,4.3590055,4.4584637,4.8734436,5.5113473,6.4133286,7.4353456,8.81404,10.597425,12.63117,13.7526455,13.917266,13.735497,13.780083,14.610043,17.089634,18.650097,19.277712,19.03764,18.056778,18.259123,18.8593,19.150816,18.773561,17.737827,15.920145,15.271953,15.059319,14.874121,14.623761,13.330807,11.427385,10.124143,9.499957,8.491658,7.006647,6.701414,6.8866115,7.15069,7.366754,7.2775846,6.989499,7.164408,7.915488,8.786603,9.465661,10.134431,10.456812,10.456812,10.525404,10.995257,11.22161,11.05699,10.388221,9.139851,7.274155,6.2692857,6.193835,6.8728933,7.8846216,6.917478,6.2658563,5.895461,5.8988905,6.5024977,7.0135064,7.4936485,7.5553813,7.051232,6.0806584,5.2747054,4.7979927,4.4104495,3.981751,3.474172,2.8911421,2.2120838,2.0474637,2.6133456,3.7313912,5.127233,6.169828,6.7494283,6.893471,6.7631464,6.550512,6.3653145,6.392751,6.5539417,6.509357,6.090947,6.341307,6.9209075,7.5245147,7.874333,7.6959944,7.455923,7.48336,7.7577267,7.891481,8.049242,8.299602,8.405919,8.347616,8.337327,8.3922,8.423067,8.405919,8.344186,8.2481575,7.881192,7.5862474,7.3221693,7.006647,6.5470824,6.1149545,5.7754254,5.442755,5.096367,4.804852,4.698535,5.0655007,5.9434752,7.301592,9.040393,9.873782,10.456812,11.619442,13.37882,14.935853,15.5085945,14.767803,13.917266,13.55373,13.684054,13.975569,14.400838,15.29253,16.348843,16.6335,16.640358,16.678083,16.146498,14.925565,13.375391,12.590015,12.795791,12.843805,12.188754,10.902658,10.381361,9.757176,9.273604,8.98209,8.718011,8.495089,8.357904,8.320179,8.347616,8.351046,8.443645,8.656279,8.879202,9.047252,9.126132,8.947794,8.632272,8.23444,7.8777623,7.73029,7.7268605,7.8023114,8.128122,8.7283,9.5033865,10.460241,11.207891,11.876661,12.569438,13.354814,13.7526455,13.992717,14.033872,13.96871,14.013294,13.649758,13.351384,12.679185,11.619442,10.600855,10.1652975,9.757176,9.3764925,8.964942,8.385342,7.9600725,7.9017696,7.534804,6.7974424,6.2384195,6.0566516,6.210983,6.550512,6.869464,6.917478,6.7219915,5.919468,5.353586,5.254128,5.2472687,5.209543,5.3090014,5.4187484,5.363875,4.9180284,4.4996185,3.9714622,3.6799474,3.6799474,3.7485392,3.9200184,3.8342788,3.5976372,3.2615378,2.8396983,2.5927682,2.452155,2.4452958,2.527606,2.5824795,2.510458,2.2635276,1.9925903,1.8245405,1.8416885,1.7456601,1.611906,1.7388009,2.0646117,2.16064,1.9274281,1.5501735,1.1660597,0.939707,1.0563129,1.1146159,1.1592005,1.1008976,0.94656616,0.78537554,0.64476246,0.490431,0.34638834,0.23321195,0.16804978,0.12003556,0.10288762,0.1097468,0.12689474,0.10288762,0.058302987,0.044584636,0.06516216,0.13032432,0.24350071,0.17147937,0.1097468,0.06516216,0.037725464,0.017147938,0.0034295875,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.037725464,0.06516216,0.061732575,0.048014224,0.024007112,0.017147938,0.030866288,0.048014224,0.020577524,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09602845,0.10288762,0.15776102,0.15776102,0.1097468,0.12346515,0.15433143,0.17147937,0.18862732,0.20920484,0.23664154,0.20920484,0.20577525,0.2194936,0.25721905,0.32581082,0.33952916,0.29837412,0.28808534,0.32238123,0.32924038,0.23321195,0.216064,0.23321195,0.24350071,0.20234565,0.16804978,0.16119061,0.15090185,0.13032432,0.1097468,0.072021335,0.024007112,0.0,0.0,0.0,0.0,0.0,0.020577524,0.05144381,0.061732575,0.01371835,0.037725464,0.06516216,0.072021335,0.072021335,0.082310095,0.082310095,0.072021335,0.08573969,0.18176813,0.116605975,0.07545093,0.06516216,0.058302987,0.030866288,0.024007112,0.030866288,0.044584636,0.05144381,0.041155048,0.044584636,0.044584636,0.041155048,0.041155048,0.061732575,0.0548734,0.048014224,0.0548734,0.07888051,0.12003556,0.15090185,0.20920484,0.29151493,0.3806842,0.45270553,0.47328308,0.48014224,0.45613512,0.4081209,0.35324752,0.31895164,0.25721905,0.19891608,0.15090185,0.13375391,0.22635277,0.33609957,0.44584638,0.5453044,0.61046654,0.64819205,0.59331864,0.5555932,0.5761707,0.64133286,0.70649505,0.88826317,1.1866373,1.5124481,1.7216529,1.8348293,1.862266,1.9823016,2.2223728,2.4967396,2.5653315,2.5619018,2.4624438,2.318401,2.2669573,2.3492675,2.5481834,2.5790498,2.4041407,2.2258022,2.4041407,2.668219,2.976882,3.1860867,3.0489032,3.1380725,3.3781435,4.0194764,4.9934793,5.90575,6.135532,6.6431108,7.31531,7.8194594,7.606825,9.287323,12.325937,12.542002,9.640571,7.1952744,7.606825,6.917478,5.703404,4.9008803,5.802862,5.2609873,3.9131594,2.8019729,2.287535,2.0440342,2.270387,2.0508933,1.7182233,1.5158776,1.6016173,1.6942163,1.7456601,1.4815818,0.9774324,0.67219913,0.607037,0.45956472,0.37039545,0.47328308,0.8711152,1.5707511,2.153781,2.0406046,1.3306799,0.7990939,0.4115505,0.40126175,0.48357183,0.5178677,0.4972902,1.0151579,1.6084765,2.1915064,2.534465,2.2841053,1.5913286,1.4678634,1.5227368,1.5536032,1.5398848,1.2277923,0.94999576,0.7442205,0.61046654,0.4972902,0.40126175,0.6036074,0.8128122,0.89512235,0.8711152,0.8676856,0.8848336,0.91227025,0.89512235,0.7099246,0.45956472,0.34981793,0.33952916,0.39783216,0.51100856,0.36010668,0.2469303,0.17833854,0.12346515,0.017147938,0.017147938,0.006859175,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.024007112,0.06516216,0.09602845,0.12003556,0.24007112,0.33609957,0.36010668,0.34981793,0.32581082,0.40126175,0.52472687,0.72364295,1.1214751,1.4507155,1.6736387,1.7730967,1.7799559,1.7799559,1.3992717,2.037175,3.3609958,4.6436615,4.729401,5.909179,8.076678,9.273604,9.047252,8.457363,7.5416627,6.5230756,5.562791,5.3330083,7.010077,8.080108,8.64599,8.433355,7.6445503,6.9620624,6.725421,6.6465406,6.7219915,7.040943,7.805741,7.6651278,7.0375133,6.451054,5.9640527,5.164959,3.7553983,3.875434,4.5956473,5.1580997,4.98662,5.0003386,5.147811,5.8062916,6.989499,8.330468,9.81205,10.230459,10.100135,9.712592,9.129561,8.31675,7.531374,7.0546613,6.8763227,6.6739774,6.416758,5.4016004,4.2046742,3.1792276,2.4487255,2.1640697,1.9137098,1.5501735,1.1008976,0.7442205,0.4664239,0.34638834,0.2777966,0.19548649,0.07888051,0.08916927,0.07888051,0.07545093,0.06859175,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.037725464,0.072021335,0.09259886,0.10288762,0.08573969,0.106317215,0.12689474,0.20920484,0.36010668,0.5693115,1.1729189,1.7799559,2.4590142,3.2683969,4.2252517,5.0312047,5.5079174,5.6485305,5.4976287,5.161529,5.2026844,5.4667625,5.960623,6.601956,7.208993,7.6788464,7.939495,8.207003,8.580828,9.023245,9.626852,10.467101,11.530273,12.548861,13.029003,13.4645605,13.817808,14.332246,14.949572,15.319967,14.7369375,13.978998,13.114742,12.528283,12.919256,12.699762,11.845795,11.228469,11.008976,10.652299,9.678296,8.786603,7.8949103,6.9654922,6.025785,5.7308407,5.9126086,5.8543057,5.353586,4.7499785,3.9200184,3.5942078,3.5461934,3.5770597,3.5118976,3.5530527,3.5804894,3.7176728,3.9131594,3.9474552,3.841138,3.9886103,4.32128,4.8494368,5.65539,6.5127864,7.455923,9.040393,11.166737,13.080446,14.352823,14.448852,14.184773,14.088745,14.424845,15.875561,17.580065,18.526632,18.584934,18.492336,18.71526,19.017063,19.226267,19.150816,18.571217,17.514904,16.410576,15.580616,15.189643,15.237658,15.37827,14.188204,12.710052,11.482259,10.542552,9.129561,7.857185,7.281014,7.473071,8.014946,8.467651,8.203573,8.06296,8.416207,9.129561,9.4862385,9.561689,9.39707,9.3079,9.89436,10.491108,10.960961,11.180455,11.080997,10.6488695,8.721441,7.239859,6.375603,6.090947,6.138962,6.060081,6.111525,6.252138,6.341307,6.111525,5.6793966,5.5387836,5.7136927,5.960623,5.7479887,5.56965,5.4941993,5.127233,4.3761535,3.450165,2.867135,2.4795918,2.270387,2.428148,3.3644254,4.629943,6.118384,7.3084507,8.076678,8.687145,8.790032,8.790032,8.625413,8.323608,8.014946,7.7028537,7.596536,7.7611566,8.134981,8.532814,8.621983,8.621983,8.529384,8.3922,8.30646,8.584257,9.026674,9.170717,8.971801,8.80718,8.824328,8.855195,8.940934,9.102125,9.342196,9.091836,8.611694,8.169277,7.81603,7.394191,6.842027,6.3653145,6.0669403,5.9434752,5.8817425,5.9400454,6.1766872,6.5985265,7.191845,7.9120584,8.766026,8.412778,8.347616,9.249598,11.002116,12.349944,13.454271,14.239647,14.832966,15.553179,15.776102,15.354263,14.973578,15.066177,15.827546,16.496315,16.87357,16.852993,16.307688,15.097044,13.80409,14.531162,15.121051,14.486577,12.641459,12.332796,12.072148,11.760056,11.321068,10.700313,10.038403,9.455373,8.992378,8.632272,8.327039,8.001227,7.9600725,8.237869,8.769455,9.403929,9.781183,9.846346,9.637141,9.23245,8.772884,8.913498,9.290752,9.8429165,10.463672,11.005547,11.321068,11.327928,11.108434,10.672876,9.942374,9.547972,9.489669,9.702303,10.388221,12.0309925,13.474849,14.695783,14.96329,14.287662,13.423406,13.073587,12.607163,12.020704,11.406808,10.950673,10.864933,10.9541025,10.264755,8.766026,7.3393173,6.7391396,6.7871537,7.0478024,7.1026754,6.540223,6.108095,5.576509,5.48734,5.826869,6.0395036,5.4907694,5.3398676,5.394741,5.3570156,4.8322887,4.5510626,4.40702,4.4516044,4.6436615,4.8322887,5.3432975,5.40503,5.0414934,4.3590055,3.5599117,3.316411,3.1140654,2.9494452,2.8739944,2.9734523,3.1792276,2.9391565,2.5721905,2.2738166,2.095478,1.9891608,1.903421,1.920569,1.9514352,1.728512,1.2758065,1.0254467,0.864256,0.77165717,0.823101,0.64476246,0.4355576,0.30866286,0.25721905,0.17147937,0.1097468,0.07888051,0.061732575,0.058302987,0.07545093,0.05144381,0.06516216,0.12689474,0.19548649,0.15433143,0.07545093,0.10288762,0.22292319,0.4081209,0.6310441,0.5624523,0.4629943,0.30866286,0.16119061,0.16462019,0.1920569,0.11317638,0.034295876,0.006859175,0.010288762,0.0034295875,0.0034295875,0.006859175,0.01371835,0.020577524,0.0274367,0.024007112,0.01371835,0.006859175,0.0034295875,0.0034295875,0.0274367,0.09259886,0.15433143,0.1371835,0.09945804,0.05144381,0.037725464,0.06516216,0.1097468,0.05144381,0.020577524,0.006859175,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.106317215,0.09602845,0.09945804,0.106317215,0.1097468,0.12346515,0.18176813,0.216064,0.22292319,0.22292319,0.26064864,0.2709374,0.25721905,0.23664154,0.22978236,0.22978236,0.3018037,0.31209245,0.26407823,0.19548649,0.18176813,0.18176813,0.18176813,0.17833854,0.16462019,0.15090185,0.14061308,0.12689474,0.10288762,0.061732575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.061732575,0.061732575,0.061732575,0.061732575,0.07888051,0.0548734,0.037725464,0.18176813,0.14747226,0.0548734,0.037725464,0.07888051,0.030866288,0.006859175,0.0,0.01371835,0.030866288,0.030866288,0.041155048,0.044584636,0.0274367,0.0,0.0,0.024007112,0.041155048,0.06516216,0.106317215,0.16804978,0.17833854,0.14747226,0.16462019,0.24350071,0.30523327,0.31895164,0.36696586,0.42183927,0.45270553,0.42869842,0.39097297,0.31895164,0.23321195,0.15776102,0.12346515,0.14747226,0.216064,0.30866286,0.37725464,0.36696586,0.40126175,0.4664239,0.5212973,0.5693115,0.64133286,0.72707254,0.9568549,1.2620882,1.5638919,1.7696671,1.7456601,1.6393428,1.6393428,1.7765263,1.9239986,2.0680413,2.3081124,2.5138876,2.5241764,2.1194851,2.0474637,2.1400626,2.1469216,2.0406046,2.0303159,2.1400626,2.3595562,2.5619018,2.620205,2.4247184,2.8156912,3.391862,3.9886103,4.57507,5.2335505,5.892031,6.451054,6.9826403,7.5107965,8.011517,9.132992,10.192734,10.48082,9.856634,8.759167,7.5382333,8.357904,9.373062,9.441654,8.1487,6.464772,4.5510626,3.1723683,2.5207467,2.2292318,2.277246,1.8691251,1.4472859,1.2860953,1.4815818,1.7971039,1.978872,1.704505,1.097468,0.7339317,0.61046654,0.45956472,0.36353627,0.36010668,0.45613512,1.4575747,2.1743584,1.9068506,0.922559,0.45613512,0.37382504,0.38754338,0.45956472,0.5590228,0.65505123,1.4369972,2.0920484,2.4795918,2.527606,2.1983654,1.6736387,1.5604624,1.6393428,1.7971039,2.0303159,1.6393428,1.2380811,0.89855194,0.7305021,0.89855194,1.1077567,1.2243627,1.2175035,1.1146159,0.9911508,0.881404,0.8265306,0.8505377,0.8711152,0.6859175,0.3566771,0.25721905,0.22635277,0.18176813,0.106317215,0.24007112,0.29151493,0.23664154,0.12689474,0.09259886,0.07888051,0.030866288,0.0,0.01371835,0.061732575,0.01371835,0.0,0.06859175,0.15433143,0.106317215,0.14404267,0.42869842,0.5796003,0.48357183,0.29151493,0.36353627,0.52815646,0.6241849,0.7339317,1.1592005,1.4267083,1.3581166,1.4850113,1.961724,2.5481834,2.3046827,2.352697,2.6647894,3.2786856,4.3041325,5.5593615,7.0752387,8.1487,8.567109,8.591117,7.6857057,6.5367937,5.223262,4.7019644,6.790583,8.241299,8.916927,9.019815,8.793462,8.498518,8.488229,8.244728,7.8366075,7.2707253,6.4990683,5.8405876,5.3570156,5.0140567,4.7774153,4.5922174,4.5201964,4.996909,5.830299,6.660259,6.927767,7.1849856,7.4936485,8.337327,9.661148,10.8958,11.5645685,11.194174,10.2236,9.139851,8.467651,7.932636,7.438775,7.0443726,6.6122446,5.844017,4.513337,3.3747141,2.369845,1.6187652,1.4335675,1.3855534,1.3821237,1.2346514,0.939707,0.67219913,0.45270553,0.26064864,0.11317638,0.030866288,0.030866288,0.030866288,0.048014224,0.072021335,0.09259886,0.09259886,0.017147938,0.0,0.0,0.0,0.0,0.0,0.072021335,0.09259886,0.048014224,0.061732575,0.061732575,0.07888051,0.13375391,0.25378948,0.47328308,1.0460242,1.7765263,2.5927682,3.457024,4.3487167,5.288424,5.669108,5.7377,5.576509,5.1100855,5.0757895,5.192395,5.6142344,6.2692857,6.866034,7.414768,7.8263187,8.193284,8.573969,8.988949,9.561689,10.299051,11.4033785,12.758065,13.9309845,14.942713,15.765814,16.252815,16.259674,15.6252,15.100473,14.54831,13.694343,12.710052,12.22305,12.2093315,11.72233,11.067279,10.432805,9.873782,9.578837,9.129561,8.330468,7.3427467,6.684266,6.0978065,6.0978065,6.23156,6.2384195,6.042933,5.079219,4.2423997,3.758828,3.6970954,3.9508848,4.4516044,4.5853586,4.513337,4.3041325,3.9371665,3.8377085,3.8788633,4.105216,4.5442033,5.2026844,5.888602,6.5779486,7.740579,9.5033865,11.688034,13.066729,13.88983,14.167625,13.985858,13.474849,13.351384,14.750656,16.019604,16.46888,16.359133,16.688372,17.336565,18.46147,19.668684,20.03565,19.596663,18.434032,17.315987,16.554619,16.005884,15.738377,15.443433,15.172495,14.949572,14.754086,13.694343,11.677745,10.1652975,9.56512,9.246168,9.270175,8.882631,8.512236,8.546532,9.338767,9.935514,10.103564,10.134431,10.247607,10.590566,10.247607,10.271614,10.63858,11.0981455,11.183885,10.978109,10.100135,8.954653,7.8606143,7.0786686,6.2864337,6.2247014,6.989499,7.870903,7.3701835,6.3310184,5.4599032,5.06893,5.1752477,5.4941993,5.4804807,5.103226,4.4859004,3.7211025,2.8534167,2.218943,1.9239986,1.8005334,1.786815,1.9239986,2.4967396,3.3369887,4.307562,5.4770513,7.1266828,8.663138,10.127572,11.008976,11.149589,10.772334,9.746887,9.472521,9.685155,10.288762,11.351934,11.742908,11.55771,10.9541025,10.199594,9.674867,9.541112,9.541112,9.633711,9.6988735,9.551401,9.441654,9.287323,9.321619,9.585697,9.901219,10.124143,10.069269,9.901219,9.712592,9.506817,8.944365,7.805741,7.099246,7.040943,7.06495,7.1129646,7.548522,8.388771,9.304471,9.595985,8.436785,7.3050213,7.2878733,8.378482,9.47595,10.209882,11.005547,12.055,13.4645605,15.258235,15.601193,14.980438,13.924125,13.227919,13.9481325,15.937293,16.890718,17.147938,16.780972,15.608052,14.071597,12.761495,12.085866,12.017275,12.116733,12.432255,13.015285,13.557159,13.824667,13.639469,13.457702,13.347955,13.073587,12.466551,11.427385,9.89093,8.903209,8.48137,8.64942,9.431366,9.846346,10.069269,10.086417,9.9698105,9.873782,9.493098,9.462232,9.6817255,10.028113,10.347065,10.419086,10.545981,10.967821,11.358793,10.834066,9.650859,9.582268,10.175586,11.163307,12.4802685,13.457702,13.975569,14.13676,14.085316,14.023583,14.119612,14.126471,13.9309845,13.526293,13.001566,12.524854,11.746337,11.183885,10.878652,10.39165,9.047252,8.748878,8.543102,7.9189177,6.8214493,6.711703,6.5813785,6.4716315,6.4407654,6.5779486,6.186976,5.6485305,5.3261495,5.284994,5.3090014,5.212973,5.2609873,5.346727,5.2815647,4.804852,4.537344,5.164959,5.3913116,4.9180284,4.4413157,4.7328305,4.201245,3.4878905,3.0454736,3.1449318,3.350707,3.0351849,2.5721905,2.1332035,1.6942163,1.5947582,1.4987297,1.5638919,1.6907866,1.4953002,1.1900668,0.90198153,0.5624523,0.23664154,0.15433143,0.14061308,0.12003556,0.106317215,0.09602845,0.061732575,0.048014224,0.072021335,0.116605975,0.17490897,0.26064864,0.18519773,0.15090185,0.15090185,0.15433143,0.106317215,0.14404267,0.40126175,0.6756287,0.8162418,0.71678376,1.1077567,1.2243627,0.88826317,0.42183927,0.64133286,0.922559,0.5624523,0.17833854,0.034295876,0.044584636,0.020577524,0.024007112,0.041155048,0.06859175,0.106317215,0.14404267,0.116605975,0.06859175,0.0274367,0.01371835,0.01371835,0.034295876,0.07545093,0.11317638,0.07545093,0.0274367,0.006859175,0.01371835,0.037725464,0.061732575,0.061732575,0.05144381,0.034295876,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.082310095,0.09945804,0.12003556,0.13032432,0.13032432,0.12346515,0.13375391,0.15433143,0.18519773,0.23321195,0.30866286,0.31209245,0.31552204,0.32581082,0.33609957,0.32581082,0.31209245,0.2709374,0.21263443,0.15090185,0.1097468,0.12003556,0.13032432,0.13375391,0.13032432,0.12689474,0.106317215,0.09945804,0.08573969,0.05144381,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030866288,0.048014224,0.037725464,0.0,0.0,0.044584636,0.072021335,0.072021335,0.072021335,0.072021335,0.041155048,0.010288762,0.006859175,0.037725464,0.030866288,0.041155048,0.037725464,0.017147938,0.006859175,0.0,0.0,0.0034295875,0.006859175,0.006859175,0.017147938,0.020577524,0.037725464,0.072021335,0.1097468,0.037725464,0.0274367,0.072021335,0.16462019,0.3018037,0.23664154,0.19891608,0.216064,0.31895164,0.52472687,0.41840968,0.36696586,0.35324752,0.36010668,0.35324752,0.33609957,0.30523327,0.29837412,0.30866286,0.28122616,0.2469303,0.23664154,0.24350071,0.25721905,0.25721905,0.28465575,0.34638834,0.4424168,0.5590228,0.64133286,0.71678376,0.9328478,1.1592005,1.3238207,1.4027013,1.5261664,1.6084765,1.7113642,1.8382589,1.9342873,2.0714707,2.1674993,2.1915064,2.1126258,1.9137098,2.0063086,2.0886188,2.0268862,1.8554068,1.786815,1.7971039,1.9480057,2.0817597,2.1023371,1.9857311,2.8739944,3.7485392,4.4687524,5.1512403,6.1629686,7.0546613,7.085528,7.010077,7.174697,7.4970784,7.606825,7.6857057,7.956643,8.447074,8.97866,9.0369625,8.097256,7.1884155,6.660259,6.2075534,4.8254294,3.6319332,2.867135,2.4418662,1.9342873,1.8759843,1.4781522,1.1249046,1.0220171,1.1866373,1.5536032,1.6804979,1.4095604,0.9259886,0.7442205,0.7579388,0.90884066,0.9945804,0.939707,0.7613684,0.9911508,1.1592005,1.1008976,0.84024894,0.5796003,0.41498008,0.50757897,0.7133542,0.9259886,1.0837497,1.786815,2.311542,2.5447538,2.4418662,2.0131679,1.605047,1.8382589,2.1126258,2.1674993,2.07833,1.7353712,1.3409687,0.922559,0.59331864,0.5590228,0.6379033,0.7682276,0.7990939,0.6927767,0.490431,0.50757897,0.5521636,0.6276145,0.6790583,0.5658819,0.274367,0.21263443,0.20234565,0.16462019,0.12003556,0.116605975,0.12689474,0.12003556,0.08573969,0.017147938,0.017147938,0.006859175,0.0,0.01371835,0.061732575,0.07888051,0.09259886,0.072021335,0.09602845,0.33952916,0.51100856,0.29494452,0.116605975,0.1371835,0.25378948,0.28808534,0.37725464,0.4938606,0.7682276,1.4781522,2.0303159,2.1983654,2.3321195,2.5481834,2.74367,2.6064866,2.6613598,2.9460156,3.7108135,5.4016004,6.893471,7.4044795,8.004657,9.129561,10.580277,9.705732,8.584257,7.164408,5.9812007,6.1561093,6.7185616,7.9909387,9.026674,9.462232,9.499957,7.9257765,7.160979,7.2947326,7.73029,7.1952744,6.7322803,6.451054,6.3035817,6.23499,6.1801167,6.2830043,6.8454566,7.8126,8.790032,9.040393,9.314759,9.746887,10.175586,10.47396,10.55284,10.131001,9.537683,8.882631,8.255017,7.7131424,7.1061053,6.2692857,5.4667625,4.773986,4.07435,3.1037767,2.270387,1.5398848,0.9774324,0.72707254,0.61046654,0.64133286,0.6241849,0.4972902,0.31895164,0.22292319,0.1371835,0.06516216,0.017147938,0.006859175,0.006859175,0.010288762,0.01371835,0.017147938,0.017147938,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.01371835,0.017147938,0.010288762,0.01371835,0.041155048,0.06859175,0.09602845,0.19548649,0.48357183,0.9911508,1.7388009,2.6064866,3.5221863,4.4721823,5.302142,5.7308407,5.809721,5.597087,5.171818,4.9214582,4.8768735,5.147811,5.689686,6.3173003,6.9723516,7.507367,7.966932,8.388771,8.803751,9.386781,10.268185,11.22161,12.106443,12.867812,13.999576,15.148488,16.283682,17.117071,17.12736,16.678083,15.6697855,14.562028,13.605173,12.843805,12.627741,12.0309925,11.180455,10.302481,9.702303,9.465661,9.640571,9.3936405,8.56368,7.658269,7.1129646,7.058091,7.284444,7.390761,6.7871537,5.90232,4.9523244,4.372724,4.3007026,4.5853586,4.9214582,5.0929375,5.1238036,4.99005,4.633373,4.506478,4.4859004,4.629943,4.98662,5.6073756,6.1904054,6.800872,7.56224,8.567109,9.89436,11.050131,12.027563,12.878101,13.581166,14.033872,13.502286,14.102464,15.097044,15.923574,16.173935,16.767254,17.562918,18.307138,18.828436,19.058218,19.222837,18.653526,17.70696,16.578627,15.29939,14.589465,14.534592,14.589465,14.452282,14.071597,12.754636,11.533703,10.652299,10.031544,9.283894,9.1810055,9.619993,9.822338,9.568549,9.1810055,8.9100685,9.095266,9.5205345,9.925226,10.0041065,9.866923,9.853205,10.401938,11.331357,11.856084,11.461681,11.05356,10.535692,9.788043,8.656279,7.891481,7.7783046,8.285883,9.06097,9.421077,8.625413,7.6171136,6.927767,6.725421,6.800872,6.7974424,7.0443726,6.7631464,5.7377,4.2938433,3.1209247,2.4418662,2.1263442,2.0508933,2.1194851,2.2806756,2.5207467,2.9185789,3.5016088,4.2218223,4.8322887,5.967482,7.31531,8.64942,9.832627,10.329918,10.707172,11.180455,11.797781,12.439114,12.723769,13.008426,13.197053,13.049581,12.164746,11.4033785,10.672876,10.302481,10.299051,10.357354,10.316199,10.05898,9.822338,9.80519,10.172156,10.39165,10.460241,10.491108,10.501397,10.408798,10.696883,10.446524,9.760606,8.992378,8.711152,9.366203,10.501397,11.269625,11.303921,10.707172,9.499957,8.64256,8.344186,8.529384,8.827758,9.033533,9.499957,10.203023,11.173596,12.500846,13.224489,13.210771,12.740917,12.30193,12.603734,14.116182,15.587475,16.640358,17.075916,16.890718,15.645778,14.205351,12.902108,11.952112,11.444533,11.712041,12.6929035,13.9138365,14.928994,15.302819,14.572317,14.030442,13.416546,12.555719,11.393089,10.010965,9.040393,8.738589,9.023245,9.441654,9.506817,9.499957,9.445084,9.410788,9.517105,9.695444,9.9801,10.401938,10.796341,10.820349,10.425946,10.731179,11.413667,12.322508,13.457702,13.886399,13.567448,13.190193,13.13532,13.505715,13.605173,13.426835,13.128461,12.823228,12.607163,13.152468,13.834956,14.181344,14.174485,14.246507,14.30481,13.327377,12.168177,11.355364,11.063849,10.72432,10.275044,9.839486,9.318189,8.39563,8.433355,8.309891,7.7851634,6.992929,6.4407654,6.060081,5.857735,5.9228973,6.1286726,6.1149545,5.7925735,5.5593615,5.346727,5.144381,4.99005,4.955754,5.164959,5.329579,5.2747054,4.9660425,4.887162,4.4104495,3.9165888,3.683377,3.8891523,3.9474552,3.7211025,3.7794054,3.9680326,3.391862,2.218943,1.6633499,1.3443983,1.0700313,0.83681935,0.6859175,0.58645946,0.4938606,0.4081209,0.37382504,0.34981793,0.3566771,0.37382504,0.36696586,0.28122616,0.22978236,0.31895164,0.4424168,0.50757897,0.41840968,0.7442205,0.91227025,0.78537554,0.4938606,0.4355576,0.6276145,0.78537554,0.91227025,0.9568549,0.7888051,0.9842916,1.1180456,0.9842916,0.6962063,0.70306545,1.5193073,1.5501735,1.0494537,0.48014224,0.5212973,0.37039545,0.29151493,0.4115505,0.61389613,0.53501564,0.2777966,0.14747226,0.09259886,0.07888051,0.07545093,0.058302987,0.061732575,0.09259886,0.12003556,0.11317638,0.082310095,0.082310095,0.06859175,0.037725464,0.024007112,0.044584636,0.041155048,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14061308,0.12003556,0.12346515,0.1371835,0.14747226,0.15090185,0.14061308,0.14061308,0.15433143,0.18176813,0.22978236,0.30866286,0.34295875,0.33952916,0.31209245,0.28808534,0.24350071,0.18519773,0.14404267,0.12003556,0.09259886,0.10288762,0.106317215,0.09945804,0.09602845,0.09602845,0.08573969,0.082310095,0.058302987,0.020577524,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.048014224,0.020577524,0.0,0.030866288,0.0548734,0.05144381,0.041155048,0.07545093,0.06859175,0.0274367,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.006859175,0.017147938,0.034295876,0.0548734,0.017147938,0.01371835,0.034295876,0.072021335,0.13375391,0.13032432,0.13032432,0.15090185,0.2194936,0.39783216,0.44584638,0.33609957,0.2503599,0.24350071,0.24350071,0.24007112,0.2194936,0.20234565,0.19548649,0.20234565,0.18862732,0.17490897,0.16804978,0.17833854,0.1920569,0.26750782,0.33609957,0.4115505,0.4938606,0.5590228,0.6241849,0.7579388,0.94656616,1.1592005,1.3409687,1.4472859,1.6187652,1.8485477,2.0165975,1.9102802,1.8485477,1.7971039,1.7525192,1.704505,1.6599203,1.7662375,1.8313997,1.8279701,1.7936742,1.8245405,1.9308578,2.170929,2.3561265,2.428148,2.452155,3.093488,3.789694,4.482471,5.3158607,6.64997,7.3530354,6.7459984,6.3207297,6.5882373,7.058091,6.159539,6.0566516,6.852316,7.9463544,8.045813,8.018375,7.4799304,7.160979,7.298162,7.6171136,5.826869,4.386442,3.3438478,2.644212,2.1263442,1.7422304,1.2860953,0.9774324,0.8848336,0.94999576,1.0871792,1.1729189,1.1660597,1.0494537,0.8196714,0.7305021,0.881404,0.9602845,0.84367853,0.6001778,0.6001778,0.58645946,0.5418748,0.47671264,0.4355576,0.4355576,0.5796003,0.8093826,1.0460242,1.2072148,1.6359133,2.0028791,2.3149714,2.4075704,1.9411465,1.5844694,1.8897027,2.2635276,2.4315774,2.4658735,1.937717,1.4198492,0.939707,0.5727411,0.4355576,0.4355576,0.6824879,0.86082643,0.83681935,0.66876954,0.48357183,0.35324752,0.29837412,0.29494452,0.2777966,0.19548649,0.19891608,0.19548649,0.15433143,0.09602845,0.10288762,0.11317638,0.11317638,0.09259886,0.06516216,0.07888051,0.116605975,0.116605975,0.072021335,0.034295876,0.061732575,0.08573969,0.09602845,0.1371835,0.2777966,0.37382504,0.28122616,0.20920484,0.23664154,0.29837412,0.29494452,0.36696586,0.5555932,0.90541106,1.4815818,2.061182,2.5378947,2.901431,3.1380725,3.223812,3.707384,4.064061,4.1635194,4.4584637,5.970912,7.459353,6.8969,6.5813785,7.5759587,9.712592,9.702303,9.578837,9.403929,8.879202,7.3530354,5.751418,7.1849856,8.735159,9.006097,8.1041155,6.7219915,6.0840883,6.526505,7.407909,7.1232533,6.4887795,6.090947,5.8200097,5.627953,5.5147767,6.2384195,7.1232533,7.9943686,8.683716,9.043822,9.369633,9.544542,9.496528,9.191295,8.608265,8.097256,7.6445503,7.298162,7.0203657,6.697984,6.2898636,5.5319247,4.6573796,3.7691166,2.836269,2.1400626,1.5398848,0.99801,0.5521636,0.31209245,0.23664154,0.24007112,0.24007112,0.19548649,0.1097468,0.07888051,0.05144381,0.034295876,0.024007112,0.017147938,0.010288762,0.0034295875,0.0,0.006859175,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.037725464,0.09259886,0.24007112,0.5624523,1.0871792,1.728512,2.4590142,3.2718265,4.2081037,5.1100855,5.768566,5.909179,5.5593615,5.079219,4.5613513,4.4550343,4.65395,5.0929375,5.7582774,6.509357,7.1884155,7.7440085,8.224151,8.786603,9.510246,10.556271,11.588576,12.401388,12.905538,13.786942,14.764374,15.909856,17.027903,17.638369,17.820137,16.914726,15.6526375,14.4145565,13.248496,12.751206,12.250486,11.537132,10.655728,9.904649,9.31133,9.235879,9.105555,8.772884,8.525954,8.282454,8.203573,8.176137,7.9600725,7.191845,6.2247014,5.435896,4.928317,4.8117113,5.219832,5.6176643,5.926327,5.9160385,5.586798,5.137522,4.8185706,4.787704,4.928317,5.1992545,5.641671,6.166398,6.742569,7.39762,8.162418,9.06097,9.962952,10.878652,11.8115,12.590015,12.88496,12.754636,13.210771,14.143619,15.2033615,15.772673,16.407146,16.6335,16.516893,16.341984,16.588915,16.88386,16.901007,16.753534,16.438013,15.806969,14.953001,14.417986,14.099034,14.088745,14.678635,14.171056,13.419975,12.483699,11.46854,10.545981,10.30934,10.401938,10.39508,10.185875,10.000677,9.56512,9.259886,9.338767,9.72288,10.014396,10.412228,10.696883,11.204462,11.955542,12.665466,12.30536,11.780633,11.327928,10.864933,9.97324,8.711152,7.949784,7.6274023,7.7851634,8.543102,8.769455,8.947794,8.889491,8.831187,9.451943,10.350495,10.052121,8.947794,7.4524937,5.9914894,4.8014226,3.9680326,3.309552,2.767677,2.4041407,2.3492675,2.3801336,2.5413244,2.8019729,3.0626216,3.3678548,4.0057583,4.979761,6.1801167,7.3839016,8.255017,9.160428,10.192734,11.269625,12.144169,12.668896,13.179905,13.941273,14.79867,15.175924,15.162207,14.757515,14.191633,13.588025,12.96727,12.415107,11.962401,11.609154,11.38623,11.382801,11.279913,11.153018,11.05699,11.084427,11.358793,11.742908,11.869802,11.8115,11.691463,11.698323,11.681175,12.315649,13.066729,13.368532,12.624311,11.499407,10.47396,9.740028,9.338767,9.1810055,8.841476,8.827758,9.1810055,9.863494,10.7586155,11.077567,10.768905,10.326488,10.069269,10.161868,11.149589,12.4974165,13.903547,15.145059,16.084764,16.04018,15.37827,14.325387,13.13532,12.072148,12.020704,12.782072,14.044161,15.247946,15.614912,15.13134,14.3974085,13.474849,12.411677,11.235329,10.624862,10.271614,10.360784,10.762046,11.008976,10.9198065,10.443094,9.914937,9.56512,9.513676,10.100135,10.477389,10.710602,10.827208,10.786053,10.515115,10.6317215,10.988399,11.588576,12.566009,14.1299,14.417986,13.762935,12.812939,12.535142,12.171606,11.399949,10.930096,11.039842,11.574858,12.250486,12.922686,13.440554,13.732068,13.797231,13.598314,12.723769,11.993267,11.787492,12.061859,12.05157,11.351934,10.381361,9.571979,9.3764925,9.4862385,9.297611,8.779744,8.025234,7.2707253,6.9346256,6.5882373,6.4064693,6.509357,6.931196,6.711703,6.1904054,5.7136927,5.4016004,5.144381,5.1855364,5.223262,5.2026844,5.1169443,5.0243454,5.0277753,4.911169,4.9180284,5.147811,5.5490727,5.4976287,5.446185,5.5113473,5.535354,5.079219,4.420738,3.8205605,3.2409601,2.726522,2.4007113,1.8588364,1.5193073,1.4472859,1.4781522,1.2415106,1.1077567,1.3238207,1.5364552,1.5810398,1.4541451,1.214074,1.1146159,0.9945804,0.89512235,1.0631721,1.4747226,1.4747226,1.3272504,1.2037852,1.1763484,1.0871792,1.0323058,1.1043272,1.2072148,1.0734608,1.2209331,1.4953002,1.4644338,1.1043272,0.7990939,1.7147937,2.037175,1.7902447,1.2415106,0.88826317,0.5521636,0.4629943,0.52815646,0.6036074,0.4938606,0.28122616,0.17147937,0.11317638,0.12003556,0.26407823,0.37382504,0.29494452,0.17833854,0.09945804,0.048014224,0.048014224,0.0548734,0.06516216,0.08573969,0.13375391,0.20920484,0.35324752,0.45956472,0.52472687,0.6241849,0.75450927,0.72707254,0.65505123,0.607037,0.61389613,0.51100856,0.34295875,0.22978236,0.19548649,0.17490897,0.12346515,0.09945804,0.08916927,0.08573969,0.09259886,0.08573969,0.07545093,0.06859175,0.061732575,0.0548734,0.0548734,0.0548734,0.05144381,0.044584636,0.037725464,0.15090185,0.12003556,0.106317215,0.09945804,0.09259886,0.09945804,0.13375391,0.14747226,0.15776102,0.17833854,0.1920569,0.32581082,0.4698535,0.48014224,0.35324752,0.20920484,0.16462019,0.12003556,0.09945804,0.09259886,0.08573969,0.09259886,0.08916927,0.07888051,0.06516216,0.044584636,0.044584636,0.044584636,0.0274367,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.024007112,0.0034295875,0.020577524,0.020577524,0.0034295875,0.024007112,0.0548734,0.06859175,0.058302987,0.044584636,0.07545093,0.044584636,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.01371835,0.05144381,0.08916927,0.1097468,0.12346515,0.17147937,0.31209245,0.28122616,0.1920569,0.12689474,0.116605975,0.116605975,0.1097468,0.10288762,0.12003556,0.18862732,0.18519773,0.16804978,0.15090185,0.14747226,0.15433143,0.22292319,0.29837412,0.36696586,0.41840968,0.44927597,0.5007198,0.59674823,0.83681935,1.1866373,1.4507155,1.488441,1.5981878,1.7559488,1.8485477,1.6667795,1.6016173,1.6153357,1.6667795,1.7422304,1.8416885,2.0131679,1.8588364,1.6324836,1.5364552,1.7319417,2.0097382,2.3732746,2.6373527,2.7985435,3.0454736,3.5873485,4.0606318,4.57164,5.3090014,6.557371,6.910619,6.2041235,5.9983487,6.660259,7.3530354,6.615674,6.4373355,6.8111606,7.1129646,6.0669403,5.895461,6.3961806,7.0443726,7.5725293,7.9600725,6.3001523,4.770556,3.4433057,2.411,1.786815,1.3443983,1.1317638,1.039165,0.9911508,0.96714365,0.78537554,0.7407909,0.8162418,0.89855194,0.7956643,0.72707254,0.8025235,0.805953,0.66191036,0.47328308,0.48700142,0.4355576,0.31895164,0.22635277,0.33266997,0.45956472,0.58988905,0.78537554,1.0494537,1.313532,1.7113642,2.1572106,2.6064866,2.8259802,2.4041407,1.9891608,1.8897027,1.9274281,2.0063086,2.1229146,1.8588364,1.4575747,0.9431366,0.48014224,0.36353627,0.37382504,0.6173257,0.823101,0.8779744,0.8265306,0.52815646,0.30866286,0.18519773,0.14747226,0.17833854,0.20920484,0.21263443,0.18862732,0.15090185,0.09945804,0.07888051,0.07888051,0.07545093,0.06516216,0.06516216,0.12346515,0.17147937,0.16462019,0.10288762,0.010288762,0.05144381,0.09945804,0.17833854,0.26064864,0.26407823,0.24007112,0.2777966,0.30866286,0.30866286,0.29151493,0.274367,0.3806842,0.69963586,1.1934965,1.6907866,2.2498093,2.8808534,3.4604537,3.923448,4.266407,4.6093655,4.8117113,4.9591837,5.329579,6.420188,7.5450926,6.8557453,6.324159,6.941485,8.711152,9.122703,9.493098,10.041832,10.14472,8.351046,5.7377,6.2658563,7.2467184,7.3598948,6.680836,5.919468,5.442755,5.9914894,7.1369715,7.257007,6.601956,5.7994323,4.976331,4.266407,3.782835,4.5956473,5.579939,6.375603,6.8969,7.3564653,7.699424,7.8194594,7.716572,7.3118806,6.4373355,5.9640527,5.5902276,5.439326,5.4187484,5.2472687,4.8151407,4.2081037,3.5050385,2.7333813,1.8897027,1.3684053,0.89512235,0.50757897,0.23664154,0.09259886,0.06859175,0.058302987,0.05144381,0.041155048,0.017147938,0.010288762,0.010288762,0.01371835,0.017147938,0.017147938,0.010288762,0.0034295875,0.0,0.006859175,0.0274367,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.037725464,0.15090185,0.37039545,0.6893471,1.2689474,1.8073926,2.3458378,2.9940298,3.9097297,4.804852,5.535354,5.689686,5.2781353,4.729401,4.1360826,3.9714622,4.091498,4.4584637,5.171818,5.977771,6.7528577,7.431916,8.045813,8.742019,9.469091,10.463672,11.530273,12.445972,12.953552,13.63261,14.4317045,15.426285,16.530611,17.497755,17.905876,17.425734,16.503176,15.354263,13.96871,13.042721,12.562579,12.017275,11.235329,10.381361,9.901219,9.671436,9.499957,9.3079,9.14328,8.834618,8.8929205,8.940934,8.759167,8.279024,7.466212,6.7871537,6.0806584,5.56965,5.8680243,6.351596,6.5196457,6.3378778,5.90232,5.446185,5.1683884,5.1992545,5.453044,5.8200097,6.166398,6.5642304,7.085528,7.6788464,8.303031,8.927217,9.47938,10.100135,10.803201,11.379372,11.365653,11.290202,11.753197,12.5145645,13.214201,13.392539,14.164196,14.555169,14.493437,14.249936,14.421415,14.527733,14.7369375,15.059319,15.440002,15.765814,15.117621,14.335675,13.917266,14.037301,14.55174,13.872682,13.097594,12.21962,11.4376745,11.149589,11.022695,10.813489,10.690024,10.714031,10.861504,10.618003,10.271614,10.213311,10.532263,11.036412,11.629731,12.055,12.38767,12.713481,13.104454,12.734058,12.490558,12.490558,12.521424,12.010415,10.4705305,8.886061,7.500508,6.601956,6.5162163,6.7871537,7.3187394,7.6376915,7.9737906,9.239308,10.408798,9.918367,8.776315,7.596536,6.5882373,5.552502,4.729401,3.9783216,3.2992632,2.8568463,2.8156912,2.9631636,3.069481,3.0557625,3.0043187,3.1483612,3.4398763,3.974892,4.6882463,5.336438,6.077229,7.160979,8.543102,10.034973,11.30049,11.567999,11.852654,12.466551,13.526293,14.939283,15.978448,16.643787,16.832415,16.602633,16.170506,15.395418,14.88441,14.531162,14.249936,13.982429,13.639469,13.251926,12.943263,12.847235,13.111313,13.454271,13.920695,14.651197,15.371411,15.371411,14.678635,14.30138,14.428274,14.754086,14.472859,13.337666,12.271064,11.509696,11.022695,10.491108,9.8429165,9.853205,10.045261,10.124143,9.983529,9.949233,9.517105,9.0369625,8.721441,8.64942,9.050681,9.750318,10.72432,11.88352,13.083877,13.906977,14.222499,14.092175,13.629181,12.9809885,12.912396,13.155897,13.776653,14.520873,14.805529,15.117621,15.001016,14.345964,13.289652,12.181894,11.664027,11.38966,11.447963,11.787492,12.22648,12.175035,11.712041,11.266195,11.029553,10.964391,11.434244,11.461681,11.2593355,11.019264,10.899229,10.72775,10.618003,10.676306,10.9369545,11.365653,12.634601,13.262215,13.063298,12.367092,12.017275,11.547421,10.714031,10.22703,10.374502,11.019264,11.626302,12.116733,12.600305,13.046151,13.282792,12.953552,12.30193,12.034423,12.319078,12.788932,12.874671,12.524854,11.8869505,11.194174,10.779194,10.371073,9.791472,9.366203,9.091836,8.611694,8.14527,7.6959944,7.3839016,7.39762,7.9875093,8.2481575,8.292743,7.915488,7.2192817,6.6225333,6.9209075,6.7631464,6.276145,5.7102633,5.425607,5.686256,6.358455,6.8385973,6.9826403,7.1095347,7.281014,7.239859,6.948344,6.5882373,6.5539417,6.560801,6.2384195,5.802862,5.4016004,5.1409516,4.945465,4.664239,4.4104495,4.07435,3.333559,2.8534167,2.9185789,3.0626216,3.0660512,2.9220085,2.4830213,2.1297739,1.7490896,1.5673214,2.153781,2.5138876,2.037175,1.6153357,1.5604624,1.6290541,1.6427724,1.5193073,1.313532,1.138623,1.1489118,1.2826657,1.3443983,1.2072148,0.91569984,0.6790583,1.1523414,1.3855534,1.3409687,1.0871792,0.8025235,0.6207553,0.6310441,0.65848076,0.6241849,0.52472687,0.34295875,0.2469303,0.2469303,0.34295875,0.53501564,0.66533995,0.5590228,0.39097297,0.2503599,0.13375391,0.29151493,0.39783216,0.39440256,0.36353627,0.50757897,0.7373613,1.0185875,1.2689474,1.4987297,1.7765263,2.0749004,2.1126258,1.8965619,1.5913286,1.5364552,1.5055889,1.2998136,1.1523414,1.1489118,1.2346514,1.0666018,0.91227025,0.84367853,0.85739684,0.85396725,0.8265306,0.77165717,0.69963586,0.6207553,0.52472687,0.45270553,0.37725464,0.30523327,0.23664154,0.17833854,0.09602845,0.09259886,0.08573969,0.05144381,0.010288762,0.017147938,0.1097468,0.15776102,0.1920569,0.22292319,0.22292319,0.32581082,0.5418748,0.58302987,0.38754338,0.14404267,0.12003556,0.11317638,0.106317215,0.09259886,0.07545093,0.06516216,0.061732575,0.0548734,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.020577524,0.061732575,0.020577524,0.0034295875,0.0,0.01371835,0.061732575,0.06516216,0.07545093,0.07888051,0.072021335,0.061732575,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.030866288,0.05144381,0.09259886,0.1097468,0.07888051,0.01371835,0.08916927,0.18176813,0.15433143,0.030866288,0.01371835,0.01371835,0.024007112,0.058302987,0.13375391,0.2469303,0.23664154,0.21263443,0.18176813,0.15090185,0.15090185,0.15433143,0.22635277,0.3018037,0.34295875,0.34295875,0.3841138,0.53844523,0.9259886,1.3992717,1.5810398,1.5330256,1.5124481,1.5021594,1.4747226,1.4095604,1.4747226,1.6290541,1.8073926,1.9857311,2.1812177,2.417859,1.9857311,1.4575747,1.2655178,1.6839274,2.1126258,2.5310357,2.784825,2.959734,3.3815732,4.1120753,4.633373,4.9934793,5.312431,5.7925735,6.0532217,6.0669403,6.701414,7.8434668,8.381912,8.124693,7.781734,7.205563,6.2041235,4.5510626,4.5510626,5.5559316,6.427047,6.6705475,6.4579134,5.3844523,4.173808,2.9322972,1.8073926,1.0117283,0.7990939,0.9534253,1.1489118,1.2209331,1.1694894,0.72021335,0.53158605,0.4938606,0.5555932,0.72021335,0.7888051,0.7956643,0.77508676,0.7407909,0.6790583,0.64476246,0.5418748,0.37725464,0.2503599,0.36696586,0.48014224,0.5555932,0.69963586,0.9602845,1.3169615,1.903421,2.5207467,2.9940298,3.1963756,3.0626216,2.651071,1.961724,1.4404267,1.2586586,1.3066728,1.6599203,1.5673214,1.0460242,0.41840968,0.32924038,0.4115505,0.6173257,0.7476501,0.72364295,0.61046654,0.52815646,0.44584638,0.37382504,0.32924038,0.33266997,0.31209245,0.24007112,0.17147937,0.13032432,0.1097468,0.034295876,0.020577524,0.0274367,0.034295876,0.037725464,0.12689474,0.14747226,0.13032432,0.09259886,0.01371835,0.082310095,0.16462019,0.2709374,0.37039545,0.3566771,0.29494452,0.28465575,0.28465575,0.2709374,0.24007112,0.23321195,0.36353627,0.75450927,1.3821237,2.0680413,2.8705647,3.5393343,4.180667,4.8425775,5.4941993,4.9077396,4.4584637,5.0106273,6.341307,7.140401,7.291303,7.040943,6.917478,7.2604365,8.23444,8.652849,9.026674,9.441654,9.561689,8.652849,6.601956,5.645101,5.2506986,5.2506986,5.8234396,5.5730796,5.295283,5.878313,7.1026754,7.613684,7.1369715,5.844017,4.2766957,2.8945718,2.0646117,2.369845,3.1243541,3.8274195,4.3041325,4.705394,5.0346346,5.3501563,5.535354,5.3981705,4.6676683,4.201245,3.8445675,3.7108135,3.690236,3.4398763,2.877424,2.386993,1.9274281,1.488441,1.0768905,0.6927767,0.31895164,0.09602845,0.030866288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010288762,0.082310095,0.26064864,0.53844523,0.864256,1.4438564,1.9274281,2.3424082,2.8499873,3.7279615,4.540774,5.0826488,5.1580997,4.7774153,4.1600895,3.6970954,3.4878905,3.532475,3.8720043,4.5819287,5.377593,6.169828,6.944915,7.6959944,8.429926,9.050681,9.839486,10.803201,11.790922,12.4974165,13.176475,13.920695,14.7369375,15.673215,16.80155,17.072487,17.106783,16.808409,16.081335,14.812388,13.54687,12.950122,12.46998,11.832077,11.043272,10.984968,10.844356,10.539123,10.041832,9.362774,9.009526,9.414218,9.966381,10.237319,9.993818,9.39707,8.690575,7.7268605,6.831738,6.824879,7.15069,6.9517736,6.5985265,6.258997,5.885172,5.813151,5.919468,6.2727156,6.7631464,7.1026754,7.3187394,7.7097125,8.152129,8.580828,8.971801,9.177576,9.366203,9.695444,10.062409,10.086417,9.678296,9.962952,10.257896,10.189304,9.695444,10.635151,11.893809,12.710052,12.905538,12.874671,12.88839,13.059869,13.323947,13.766364,14.616901,14.616901,14.2533655,14.164196,14.229359,13.6086035,11.910957,10.751757,10.086417,9.97667,10.621432,10.899229,10.871792,10.906088,11.067279,11.122152,11.180455,11.345076,11.55428,11.869802,12.432255,12.97413,13.334236,13.488567,13.416546,13.13532,12.761495,13.162757,14.027013,14.812388,14.771234,13.423406,11.406808,9.304471,7.4044795,5.717122,4.8425775,4.372724,4.2698364,4.6676683,5.8543057,6.351596,6.375603,6.3173003,6.2075534,5.7239814,4.9214582,4.32128,3.8720043,3.5839188,3.532475,3.7862647,4.15666,4.2286816,3.9508848,3.6696587,3.5873485,3.690236,3.9680326,4.3178506,4.5201964,5.055212,5.970912,7.2775846,8.834618,10.347065,10.285333,10.374502,10.484249,10.820349,11.931535,13.347955,14.836395,16.084764,17.014183,17.78927,17.62808,17.442883,17.305698,17.21996,17.099922,16.938732,16.582056,16.21166,15.920145,15.728088,15.951012,16.609491,17.682953,18.602083,18.224829,17.329706,16.252815,15.635489,15.676644,16.146498,15.337115,14.459141,13.831526,13.341095,12.439114,11.746337,12.010415,12.048141,11.355364,10.14129,9.993818,9.908078,9.685155,9.349055,9.119273,8.80718,8.512236,8.484799,8.796892,9.321619,10.131001,10.947243,11.701753,12.343085,12.830087,13.179905,13.193623,13.186764,13.334236,13.687484,14.640909,15.470869,15.604623,15.0078745,14.2190695,13.2862215,12.644889,12.415107,12.665466,13.413116,13.265644,13.114742,13.121602,13.258785,13.313659,13.38225,13.025573,12.524854,12.061859,11.732618,11.204462,10.827208,10.72775,10.858074,11.019264,11.211322,11.688034,12.188754,12.521424,12.576297,12.277924,11.900668,11.574858,11.382801,11.324498,11.677745,12.092726,12.531713,13.008426,13.588025,13.375391,12.864383,12.614022,12.699762,12.713481,12.71691,13.090735,13.485138,13.433694,12.3533745,11.30735,10.374502,10.05898,10.237319,10.179015,9.489669,9.057541,8.865483,8.958082,9.458802,10.2236,11.132441,11.091286,10.13786,9.424506,9.942374,9.578837,8.704293,7.7268605,7.085528,7.507367,8.707723,9.328478,9.0644,8.680285,9.040393,8.793462,8.124693,7.5519514,7.936065,8.158989,8.244728,8.323608,8.416207,8.447074,9.002667,9.1810055,8.985519,8.378482,7.250148,6.385892,5.878313,5.579939,5.3878818,5.2301207,4.6916757,4.2183924,3.8034124,3.666229,4.2355404,4.3178506,3.40901,2.6304936,2.4075704,2.469303,2.651071,2.4315774,1.7971039,1.1351935,1.2106444,1.2517995,0.8711152,0.52815646,0.42869842,0.5041494,0.36696586,0.2709374,0.24007112,0.29837412,0.48014224,0.64133286,0.7442205,0.77851635,0.75450927,0.70306545,0.5624523,0.5212973,0.64133286,0.86082643,0.980862,1.039165,1.1317638,1.1729189,1.1180456,0.94999576,1.2072148,1.3375391,1.2758065,1.2037852,1.5364552,2.0303159,2.2292318,2.4041407,2.6785078,3.0317552,3.3369887,3.4981792,3.2203827,2.6887965,2.5721905,2.8225505,2.7230926,2.5824795,2.5893385,2.7951138,2.5550427,2.2738166,2.1400626,2.1469216,2.0920484,2.0097382,1.862266,1.6770682,1.471293,1.2243627,1.0220171,0.823101,0.64819205,0.5007198,0.37039545,0.061732575,0.08573969,0.09945804,0.082310095,0.0548734,0.09259886,0.16462019,0.18176813,0.18862732,0.19891608,0.19891608,0.17490897,0.14061308,0.116605975,0.106317215,0.106317215,0.13032432,0.17490897,0.18519773,0.15090185,0.07545093,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.061732575,0.061732575,0.061732575,0.024007112,0.0,0.01371835,0.061732575,0.072021335,0.06859175,0.037725464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.030866288,0.041155048,0.037725464,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.01371835,0.0274367,0.05144381,0.07545093,0.11317638,0.13032432,0.14404267,0.16119061,0.19891608,0.22292319,0.25721905,0.26407823,0.24350071,0.24350071,0.30523327,0.61389613,1.1694894,1.6770682,1.5570327,1.371835,1.3924125,1.5021594,1.6290541,1.7388009,1.5330256,1.4335675,1.4472859,1.5364552,1.6324836,1.646202,1.3443983,1.2723769,1.6599203,2.4418662,2.9288676,3.2443898,3.2615378,3.1723683,3.4776018,4.0537724,5.0826488,5.7136927,5.4736214,4.3041325,5.3158607,6.7700057,8.656279,10.127572,9.506817,7.1369715,6.8763227,7.1129646,6.992929,6.392751,6.3447366,6.495639,6.742569,6.7494283,5.9812007,4.5167665,3.40901,2.49331,1.6942163,1.0220171,0.84024894,0.77508676,0.94656616,1.2175035,1.2037852,0.6207553,0.52815646,0.6379033,0.7682276,0.85396725,0.805953,0.6756287,0.8162418,1.1797781,1.3272504,0.8505377,0.6036074,0.50757897,0.47671264,0.42869842,0.45270553,0.548734,0.6173257,0.65848076,0.7922347,1.2826657,1.5947582,1.8039631,2.0989075,2.8088322,2.843128,2.194936,1.6393428,1.488441,1.587899,2.037175,1.978872,1.4644338,0.7922347,0.48700142,0.548734,1.1420527,1.3478279,0.8676856,0.0,0.51100856,0.7339317,0.72021335,0.58988905,0.5041494,0.4046913,0.25378948,0.13032432,0.061732575,0.0,0.061732575,0.09602845,0.13032432,0.17147937,0.18176813,0.19548649,0.17833854,0.15433143,0.12346515,0.07545093,0.12346515,0.1920569,0.2469303,0.28465575,0.31895164,0.4046913,0.41840968,0.4355576,0.4355576,0.29151493,0.3018037,0.34295875,0.48700142,0.94656616,2.0440342,3.7519686,4.619654,5.1512403,5.579939,5.857735,4.7842746,3.8479972,5.0449233,7.7028537,8.484799,6.691125,5.6828265,5.284994,5.5730796,6.866034,8.220721,9.585697,10.213311,9.959522,9.263316,7.798882,6.351596,5.0449233,4.197815,4.3349986,4.7499785,5.336438,6.0875177,6.831738,7.2467184,6.7219915,5.2644167,3.3369887,1.6873571,1.3581166,1.4061309,1.8142518,2.0886188,2.1194851,2.1674993,2.4830213,2.7470996,2.9494452,3.0900583,3.1895163,3.2512488,3.275256,2.9803114,2.352697,1.6324836,1.5090185,1.2620882,0.90198153,0.52815646,0.31895164,0.16119061,0.07545093,0.034295876,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1371835,0.37039545,0.6790583,1.0837497,1.4987297,1.9308578,2.3767042,2.8980014,3.6319332,4.5099077,4.7774153,4.6676683,4.2698364,3.525616,3.2066643,3.0626216,3.1723683,3.532475,4.0434837,4.7499785,5.4770513,6.2041235,6.9037595,7.5382333,8.296172,9.06097,9.877212,10.738038,11.581717,12.397959,12.932974,13.354814,14.003006,15.395418,16.225378,16.616352,16.403717,15.693792,14.860402,13.896688,13.207341,12.713481,12.30193,11.825217,11.286773,10.768905,10.103564,9.400499,9.033533,10.045261,10.978109,11.97269,12.47341,11.214751,10.14129,9.424506,8.988949,8.766026,8.666568,8.251588,7.9189177,7.6925645,7.486789,7.0958166,6.8763227,6.931196,7.0889573,7.2604365,7.431916,7.5416627,7.6685576,7.881192,8.165848,8.423067,8.519095,8.388771,8.333898,8.512236,8.927217,8.889491,8.615124,8.131552,7.6925645,7.7680154,8.464222,9.764035,10.72089,10.984968,10.789482,11.495977,12.103014,12.370522,12.4802685,13.032433,14.239647,14.860402,14.843254,14.339106,13.718349,12.459691,11.002116,9.959522,9.606275,9.887501,10.755186,11.026124,10.971251,10.755186,10.436234,10.741467,11.22161,11.574858,11.859513,12.4802685,13.581166,14.102464,14.222499,13.965281,13.183334,13.173045,13.560589,14.771234,16.407146,17.271402,16.355703,15.011304,13.351384,11.4033785,9.108984,7.239859,5.5387836,4.2766957,3.474172,2.8980014,2.702515,3.1140654,3.9611735,4.6265135,4.029765,3.724532,3.7005248,3.8479972,4.108646,4.4859004,5.353586,5.689686,5.5730796,5.219832,4.99005,4.6608095,4.3933015,4.307562,4.420738,4.65395,5.1409516,5.796003,6.6636887,7.8091707,9.321619,10.569988,11.657167,12.109874,11.787492,10.8958,11.091286,11.495977,12.144169,13.138749,14.664916,16.20137,16.997036,17.518333,18.015623,18.54035,19.246845,19.678972,19.6241,19.147387,18.584934,18.084215,18.115082,18.293419,18.296848,17.881868,16.96617,16.438013,16.571766,17.319416,18.293419,19.236557,18.427174,16.993607,15.587475,14.404267,13.7697935,13.317088,12.641459,11.777204,11.214751,10.72775,10.971251,11.533703,11.938394,11.657167,10.398509,8.988949,8.169277,7.9909387,7.781734,7.829748,8.018375,8.40249,9.033533,9.949233,10.875222,11.794352,12.55915,13.149038,13.687484,13.906977,14.520873,15.302819,15.951012,16.098484,15.87899,15.721229,15.9921665,16.62321,17.134218,16.108772,15.433144,14.949572,14.582606,14.328816,14.5585985,14.856973,14.836395,14.407697,13.749216,12.171606,11.183885,10.679735,10.542552,10.666017,11.238758,11.732618,12.147599,12.538571,13.015285,13.087306,13.197053,13.413116,13.54687,13.169616,12.984418,13.471419,14.0750265,14.527733,14.846684,14.321958,13.649758,12.977559,12.284782,11.382801,10.762046,11.091286,11.718901,12.257345,12.572867,12.229909,11.97269,11.948683,12.034423,11.825217,11.214751,10.576848,10.271614,10.532263,11.458252,12.020704,12.079007,12.024134,12.061859,12.205902,12.109874,11.828648,11.509696,11.235329,11.015835,11.273054,11.207891,11.324498,11.595435,11.4754,10.984968,10.460241,9.918367,9.537683,9.657719,9.89093,10.213311,10.844356,11.646879,12.144169,11.900668,12.425395,13.38911,14.123041,13.612033,12.854094,11.794352,10.89237,10.343636,10.100135,9.709162,9.448513,9.379922,9.239308,8.423067,7.654839,6.992929,6.4990683,6.1321025,5.751418,4.715683,3.7794054,2.983741,2.393852,2.0920484,1.8108221,1.4918705,1.2037852,0.9911508,0.8711152,0.77165717,0.70306545,0.66533995,0.66191036,0.6859175,0.66191036,0.6001778,0.5521636,0.5555932,0.64133286,0.97057325,1.2346514,1.4747226,1.6873571,1.845118,2.0063086,2.7230926,3.3678548,3.6113555,3.4021509,3.1826572,2.8637056,2.7539587,3.059192,3.8891523,4.7088237,4.3349986,3.8102717,3.6079261,3.6319332,3.4981792,3.6285036,3.6765177,3.5976372,3.6456516,4.170378,4.0366244,3.6765177,3.391862,3.357566,3.3198407,3.2375305,3.1346428,3.0077481,2.8396983,2.6167753,2.3629858,2.0817597,1.7730967,1.4198492,1.138623,0.8848336,0.6962063,0.5658819,0.4424168,0.061732575,0.07545093,0.07545093,0.06516216,0.058302987,0.06859175,0.10288762,0.13032432,0.18176813,0.22635277,0.19891608,0.17490897,0.16119061,0.15776102,0.15776102,0.16804978,0.16462019,0.16119061,0.1097468,0.041155048,0.06516216,0.05144381,0.048014224,0.0548734,0.058302987,0.048014224,0.048014224,0.020577524,0.020577524,0.037725464,0.0,0.037725464,0.020577524,0.0034295875,0.01371835,0.01371835,0.01371835,0.0034295875,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.006859175,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.006859175,0.01371835,0.041155048,0.09602845,0.10288762,0.09602845,0.09602845,0.11317638,0.1371835,0.17833854,0.23664154,0.30523327,0.35324752,0.4046913,0.5727411,0.8196714,1.039165,1.0425946,1.0082988,1.0117283,1.1008976,1.2517995,1.3615463,1.3684053,1.4987297,1.6976458,1.8176813,1.6324836,1.4507155,1.2175035,1.1763484,1.3752645,1.6976458,1.9308578,2.4007113,2.9871707,3.415869,3.2718265,3.758828,5.147811,6.012067,5.8680243,5.192395,6.3721733,7.1198235,7.4936485,7.6616983,7.9086285,7.822889,7.4010496,7.010077,6.8214493,6.807731,5.4016004,4.5990767,4.804852,5.4667625,5.079219,4.091498,3.1689389,2.3801336,1.7902447,1.4507155,1.2963841,1.2106444,1.2586586,1.3272504,1.1214751,0.64133286,0.53844523,0.6001778,0.7099246,0.85396725,1.0014396,1.1077567,1.2723769,1.4404267,1.3992717,0.9945804,0.6962063,0.5007198,0.39783216,0.37725464,0.4115505,0.45270553,0.47671264,0.5041494,0.61046654,0.922559,1.2826657,1.6393428,1.9651536,2.2326615,2.1640697,1.8005334,1.8108221,2.2669573,2.6476414,2.1812177,1.6804979,1.1146159,0.6276145,0.53844523,0.51100856,0.6036074,0.607037,0.45613512,0.24350071,0.51100856,0.6790583,0.7579388,0.77165717,0.7339317,0.6173257,0.25721905,0.0274367,0.0274367,0.072021335,0.106317215,0.12346515,0.09259886,0.034295876,0.037725464,0.037725464,0.1371835,0.216064,0.22978236,0.20920484,0.26750782,0.32238123,0.36353627,0.39440256,0.4424168,0.4389872,0.490431,0.5212973,0.5007198,0.4115505,0.5521636,0.6001778,0.70306545,1.1077567,2.1674993,4.012617,5.0895076,5.6245236,5.597087,4.7362604,3.8479972,3.083199,3.6936657,5.284994,5.8234396,4.5167665,4.431027,4.99005,5.7925735,6.5985265,7.2124224,7.641121,7.641121,7.174697,6.4304767,5.3261495,4.3007026,3.350707,2.5481834,2.037175,2.0646117,2.651071,3.8171308,5.3673043,6.9071894,7.610255,7.250148,6.012067,4.513337,3.8102717,3.175798,2.5619018,2.085189,1.7971039,1.6770682,1.4198492,1.2655178,1.2723769,1.4164196,1.6016173,1.7593783,1.845118,1.7593783,1.4850113,1.1077567,0.7990939,0.5178677,0.30866286,0.18176813,0.09945804,0.041155048,0.01371835,0.006859175,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01371835,0.020577524,0.01371835,0.01371835,0.01371835,0.16462019,0.42869842,0.7682276,1.1317638,1.4404267,1.6564908,1.9582944,2.4144297,2.9734523,3.6765177,3.99204,4.0194764,3.7759757,3.2066643,2.8499873,2.7573884,2.8705647,3.1449318,3.532475,4.1600895,4.8322887,5.5490727,6.2864337,6.989499,7.6857057,8.512236,9.386781,10.264755,11.105004,11.660598,12.113303,12.500846,12.922686,13.55373,14.003006,14.164196,14.2190695,14.273943,14.363112,13.992717,13.591455,13.083877,12.504276,12.006986,11.598865,11.067279,10.425946,9.729739,9.071259,8.988949,9.030104,9.297611,9.55826,9.239308,8.711152,8.299602,8.021805,8.025234,8.580828,8.916927,9.132992,9.057541,8.697433,8.217292,7.7920227,7.56224,7.390761,7.222711,7.0889573,7.140401,7.394191,7.81603,8.337327,8.838047,8.906639,8.906639,8.872343,8.848335,8.903209,8.786603,8.354475,8.073249,8.200144,8.793462,8.81404,8.906639,9.139851,9.493098,9.822338,10.326488,11.190743,11.780633,11.8115,11.334786,11.770344,12.295071,12.6929035,12.788932,12.459691,11.838936,10.947243,10.22703,9.942374,10.192734,11.129011,11.605724,11.609154,11.276484,10.899229,10.484249,10.408798,10.751757,11.616013,13.114742,14.606613,15.892709,16.149927,15.501736,15.001016,15.145059,15.398848,15.680074,15.782962,15.367981,14.562028,13.80409,13.341095,12.943263,11.917816,10.566559,9.623423,8.875772,8.011517,6.5985265,5.40503,4.4447455,3.923448,3.7519686,3.5633414,3.6319332,3.5839188,3.590778,3.782835,4.280125,5.360445,6.848886,7.795452,7.963502,7.8091707,7.06838,6.7219915,6.6396813,6.697984,6.8145905,7.0889573,7.205563,7.4010496,7.781734,8.309891,9.22216,10.367643,11.629731,12.600305,12.579727,12.521424,12.264205,12.123591,12.267634,12.710052,13.4474125,14.147048,15.011304,15.995596,16.79469,17.590355,18.492336,19.167965,19.486916,19.500635,18.725548,18.30028,18.430603,18.722118,18.187103,17.652086,16.859852,16.287111,16.448301,17.892159,17.37772,15.728088,14.538021,14.325387,14.538021,13.512574,12.905538,12.775213,12.991278,13.241637,12.898679,12.082437,11.5645685,11.55428,11.694893,10.525404,10.062409,10.155008,10.47396,10.539123,9.983529,9.719451,9.575408,9.39707,9.033533,9.561689,10.38479,11.211322,11.784062,11.893809,12.288212,13.310229,14.435134,15.313108,15.7795315,15.981877,16.009314,16.153357,16.496315,16.938732,16.774113,16.595774,16.324837,15.9578705,15.573756,15.199932,15.073037,15.079896,15.011304,14.565458,13.831526,13.344524,13.193623,13.296511,13.399398,13.035862,12.956982,12.943263,12.912396,12.919256,13.598314,14.033872,14.212211,14.393978,15.110763,15.247946,15.234227,15.254805,15.436573,15.858413,16.067617,15.666355,15.138199,14.826107,14.946142,14.589465,14.345964,14.424845,14.856973,15.525743,14.658057,13.543441,12.761495,12.404818,12.068718,11.4205265,11.125582,10.88894,10.755186,11.105004,11.71547,11.976119,12.154458,12.425395,12.867812,13.255356,13.426835,13.227919,12.826657,12.7272,13.852104,14.634049,14.922135,14.836395,14.781522,14.363112,13.972139,13.622321,13.334236,13.125031,12.88839,12.860953,13.214201,13.828096,14.270514,14.424845,14.7369375,15.196502,15.683503,15.940722,16.112202,16.383139,16.400288,16.071047,15.594335,15.426285,15.484588,15.621771,15.80011,16.074476,14.935853,13.320518,12.048141,11.327928,10.744898,9.451943,8.049242,6.842027,5.895461,5.0312047,4.623084,4.400161,4.1360826,3.7691166,3.3712845,3.2066643,3.0900583,2.9974594,2.9185789,2.836269,2.6922262,2.4555845,2.218943,2.037175,1.9480057,2.0337453,2.1640697,2.3561265,2.5550427,2.627064,2.620205,2.8499873,3.292404,3.8857226,4.537344,4.962613,5.147811,5.2781353,5.4804807,5.830299,6.3378778,6.1046658,5.65539,5.2918534,5.120374,5.055212,4.931747,4.65395,4.3178506,4.2218223,4.619654,4.7808447,4.57164,4.07435,3.5873485,3.2889743,3.117495,3.000889,2.8637056,2.6545007,2.386993,2.1091962,1.8348293,1.5741806,1.3443983,1.1832076,1.039165,0.91912943,0.8162418,0.72364295,0.05144381,0.06516216,0.058302987,0.06859175,0.10288762,0.116605975,0.12003556,0.1371835,0.17490897,0.21263443,0.18862732,0.16462019,0.14747226,0.1371835,0.13375391,0.1371835,0.12346515,0.12003556,0.08916927,0.048014224,0.061732575,0.061732575,0.037725464,0.0274367,0.037725464,0.061732575,0.0548734,0.037725464,0.041155048,0.0548734,0.037725464,0.0548734,0.024007112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.037725464,0.0548734,0.072021335,0.09259886,0.12003556,0.1371835,0.16462019,0.20920484,0.26407823,0.31895164,0.3806842,0.4938606,0.66533995,0.8745448,1.08032,0.939707,0.82996017,0.88826317,1.097468,1.2655178,1.3855534,1.546744,1.6804979,1.6942163,1.4575747,1.3203912,1.2380811,1.3684053,1.646202,1.7662375,1.5501735,2.2360911,3.2615378,3.9783216,3.6868064,4.1429415,5.2747054,5.9434752,5.878313,5.672538,6.6225333,6.728851,6.159539,5.5662203,6.0875177,6.6876955,6.992929,6.944915,6.619104,6.2247014,4.8254294,4.0057583,3.9886103,4.4241676,4.40359,3.8445675,2.7882545,1.8588364,1.3306799,1.1180456,1.1111864,1.1454822,1.2723769,1.3546871,1.097468,0.6756287,0.5796003,0.65162164,0.805953,1.0460242,1.0528834,1.1043272,1.3752645,1.7147937,1.6667795,1.2106444,0.91912943,0.7099246,0.53844523,0.40126175,0.4389872,0.5007198,0.53158605,0.52815646,0.5453044,0.6036074,0.96371406,1.4164196,1.7490896,1.7250825,1.8382589,2.0234566,2.2258022,2.3904223,2.4830213,2.1674993,1.7182233,1.1660597,0.6927767,0.6036074,0.5178677,0.4389872,0.47671264,0.64133286,0.85396725,0.64476246,0.7099246,1.0117283,1.2929544,1.0871792,0.7682276,0.274367,0.0,0.01371835,0.06516216,0.07545093,0.07545093,0.044584636,0.0,0.0,0.10288762,0.16462019,0.19548649,0.2194936,0.23664154,0.26064864,0.28465575,0.33609957,0.432128,0.58302987,0.6310441,0.7407909,0.77508676,0.6824879,0.5144381,0.69963586,0.83338976,1.2072148,1.9548649,3.0489032,4.5784993,4.8288593,4.431027,3.858286,3.4295874,3.0111778,2.5927682,3.0454736,4.15666,4.6265135,3.2306714,3.2546785,4.1600895,5.5079174,6.9620624,7.682276,7.589677,6.8591747,5.7377,4.5510626,3.82399,3.2409601,2.8019729,2.4007113,1.8313997,1.5364552,1.7010754,2.4212887,3.625074,5.0620713,6.0840883,6.427047,6.018926,5.099797,4.2423997,3.3198407,2.6304936,2.0406046,1.4747226,0.90541106,0.607037,0.42869842,0.3806842,0.42869842,0.52815646,0.64476246,0.6790583,0.65505123,0.59674823,0.53844523,0.38754338,0.2469303,0.14404267,0.07545093,0.0274367,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.006859175,0.08916927,0.25378948,0.4938606,0.7956643,1.1008976,1.2929544,1.5330256,1.879414,2.311542,2.8637056,3.2203827,3.292404,3.0969174,2.7711067,2.5138876,2.49331,2.6167753,2.8465576,3.192946,3.7862647,4.4721823,5.23698,6.042933,6.8043017,7.4970784,8.309891,9.163857,9.97667,10.655728,11.077567,11.369082,11.567999,11.736049,11.955542,12.288212,12.517994,12.768354,13.087306,13.440554,13.46799,13.361672,13.077017,12.668896,12.291641,12.089295,11.880091,11.650309,11.372512,10.981539,10.878652,10.902658,10.593996,9.798331,8.687145,8.340756,8.64256,9.541112,10.460241,10.30934,10.021255,9.921797,9.767465,9.510246,9.287323,8.64942,8.049242,7.623973,7.431916,7.442205,7.764586,8.193284,8.711152,9.249598,9.6645775,9.571979,9.3593445,9.112414,8.937505,8.951223,9.122703,8.721441,8.292743,8.182996,8.546532,8.333898,8.056101,8.220721,8.790032,9.1810055,8.752307,9.009526,9.499957,9.918367,10.124143,10.4533825,10.593996,10.933525,11.482259,11.862943,11.993267,11.712041,11.201033,10.820349,11.094715,11.4754,11.345076,10.964391,10.511685,10.093276,9.595985,9.352485,9.688584,10.786053,12.689473,14.606613,15.896138,16.321407,16.012743,15.4742985,15.306249,15.306249,15.71094,16.0539,15.175924,13.231348,11.924676,10.984968,10.131001,9.095266,8.824328,9.078118,9.235879,8.800322,7.4113383,5.627953,4.2183924,3.2306714,2.7368107,2.836269,2.819121,2.6785078,2.867135,3.4604537,4.15323,4.8494368,5.8337283,6.5950966,7.085528,7.7371492,7.699424,7.5519514,7.613684,7.9463544,8.361334,9.263316,9.836057,10.161868,10.251037,10.069269,10.014396,10.456812,11.262765,12.154458,12.706621,12.871242,12.744347,12.586586,12.528283,12.562579,12.71691,13.125031,13.697772,14.318527,14.846684,15.488017,16.283682,17.226818,18.252264,19.215979,19.78872,19.613811,19.11995,18.389448,17.147938,16.832415,16.46888,15.999025,15.597764,15.693792,14.616901,13.858963,13.618892,13.708061,13.536582,13.008426,12.579727,12.699762,13.279363,13.701202,13.684054,13.505715,13.457702,13.598314,13.7526455,12.737488,11.910957,11.670886,11.993267,12.421966,12.260776,12.113303,11.852654,11.423956,10.827208,10.63858,10.947243,11.447963,11.808069,11.646879,11.821788,12.22305,12.627741,13.039291,13.677195,13.975569,13.886399,13.896688,14.201921,14.7026415,14.767803,14.668345,14.311668,13.807519,13.495427,13.344524,13.265644,13.317088,13.540011,13.954991,13.965281,13.786942,13.615462,13.591455,13.828096,14.160767,13.944703,13.660047,13.574307,13.725209,14.411126,14.96329,15.0250225,14.815818,15.138199,15.539461,15.618341,15.604623,15.71094,16.13278,16.62321,17.103354,17.388008,17.53891,17.844143,18.238546,18.427174,18.475187,18.410025,18.20768,17.741257,17.1205,16.510035,16.077906,16.012743,15.6526375,15.2033615,14.819247,14.479718,13.982429,13.478279,13.320518,13.200482,12.977559,12.6929035,13.440554,13.9138365,13.900118,13.687484,14.068168,15.412566,16.362562,17.099922,17.71039,18.21111,17.844143,17.326277,16.527182,15.645778,15.193072,15.13134,14.911846,14.815818,14.953001,15.285671,15.536031,15.844694,16.221949,16.62664,16.983316,17.28169,17.521763,17.511473,17.274832,17.031332,17.024471,17.154797,17.21653,17.189093,17.240536,16.489456,15.391989,14.393978,13.639469,12.9809885,11.88352,10.703742,9.719451,8.988949,8.330468,7.840037,7.4113383,6.9723516,6.5333643,6.186976,5.9812007,5.857735,5.7754254,5.7274113,5.73427,5.7479887,5.675967,5.576509,5.456474,5.284994,5.1340923,5.0003386,4.976331,5.0346346,5.0483527,5.0346346,5.1580997,5.3913116,5.7308407,6.193835,6.4373355,6.550512,6.677407,6.8214493,6.848886,6.893471,6.6533995,6.307011,6.0052075,5.857735,5.744559,5.4941993,5.144381,4.7534084,4.400161,4.3624353,4.32471,4.170378,3.882293,3.5564823,3.2032347,2.983741,2.8294096,2.6887965,2.5001693,2.277246,2.0714707,1.8759843,1.7010754,1.5570327,1.4369972,1.313532,1.1866373,1.0563129,0.90198153,0.0274367,0.058302987,0.061732575,0.07545093,0.11317638,0.14747226,0.14747226,0.15090185,0.16462019,0.17833854,0.17147937,0.13032432,0.12346515,0.116605975,0.106317215,0.09945804,0.09259886,0.09602845,0.09259886,0.07888051,0.061732575,0.041155048,0.01371835,0.0,0.006859175,0.037725464,0.030866288,0.0274367,0.030866288,0.037725464,0.037725464,0.037725464,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0274367,0.05144381,0.082310095,0.11317638,0.13375391,0.15433143,0.17490897,0.20920484,0.29151493,0.37725464,0.44927597,0.607037,0.86082643,1.1351935,0.91912943,0.78537554,0.84024894,1.0494537,1.2415106,1.4678634,1.7902447,1.9239986,1.7593783,1.3478279,1.4369972,1.5330256,1.7319417,1.9411465,1.8759843,1.5090185,2.301253,3.3712845,4.0537724,3.8891523,4.1635194,4.6848164,4.870014,4.7191124,4.787704,5.5147767,5.6245236,5.2747054,4.9591837,5.4907694,6.1458206,6.910619,7.157549,6.7322803,5.9400454,4.5339146,3.899441,3.8479972,4.1326528,4.4756117,4.0434837,2.6956558,1.5741806,1.08032,0.90198153,1.0460242,1.1180456,1.138623,1.0940384,0.9328478,0.6927767,0.6276145,0.805953,1.2312219,1.8416885,1.6016173,1.3786942,1.313532,1.3924125,1.4404267,1.3101025,1.1077567,0.881404,0.65162164,0.39783216,0.39440256,0.42869842,0.4424168,0.42183927,0.42526886,0.42183927,0.72364295,1.1043272,1.3478279,1.2346514,1.471293,1.903421,2.0886188,1.9685832,1.862266,1.8554068,1.5638919,1.1111864,0.7682276,0.939707,1.08032,1.1729189,1.1797781,1.1146159,1.0563129,0.66876954,0.69963586,1.0837497,1.4472859,1.0940384,0.66533995,0.25721905,0.041155048,0.020577524,0.034295876,0.0274367,0.024007112,0.0274367,0.030866288,0.024007112,0.12346515,0.14747226,0.16462019,0.20234565,0.2469303,0.23321195,0.23664154,0.28808534,0.4115505,0.6241849,0.77165717,0.9294182,0.9842916,0.8848336,0.6379033,0.764798,0.9294182,1.6221949,2.8568463,4.1600895,5.5559316,5.360445,4.3933015,3.391862,2.9974594,2.7711067,2.7402403,3.0969174,3.6627994,3.8891523,2.7882545,2.9048605,3.9371665,5.2987127,6.1321025,6.3790326,6.1972647,5.48734,4.3590055,3.1449318,2.7230926,2.5070283,2.5721905,2.6887965,2.318401,1.8656956,1.7010754,1.920569,2.5378947,3.4810312,4.2835546,4.7842746,4.7259717,4.122364,3.2855449,2.352697,1.8416885,1.4267083,0.94999576,0.42869842,0.25721905,0.12689474,0.061732575,0.048014224,0.06516216,0.12346515,0.12003556,0.106317215,0.1097468,0.15776102,0.14747226,0.12346515,0.09259886,0.05144381,0.020577524,0.020577524,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.010288762,0.0034295875,0.020577524,0.09945804,0.2469303,0.4664239,0.7305021,0.922559,1.097468,1.3306799,1.7079345,2.1297739,2.4761622,2.568761,2.4315774,2.270387,2.16064,2.194936,2.311542,2.5241764,2.8980014,3.4810312,4.214963,5.038064,5.895461,6.7322803,7.4181976,8.179566,8.97866,9.743458,10.347065,10.762046,10.933525,10.991828,11.019264,11.06042,11.348505,11.653738,12.010415,12.404818,12.775213,13.004995,13.145609,13.162757,13.077017,12.939834,12.874671,12.830087,12.830087,12.795791,12.545431,12.195613,12.123591,11.705182,10.672876,9.102125,8.457363,8.512236,9.5205345,10.827208,10.864933,10.436234,10.206452,10.014396,9.897789,10.134431,9.815479,9.023245,8.385342,8.169277,8.272165,8.844906,9.441654,10.113853,10.672876,10.696883,10.168727,9.897789,9.6645775,9.373062,9.067829,9.136421,8.81404,8.385342,8.069819,8.008087,7.689135,7.380472,7.442205,7.822889,8.080108,7.4113383,7.1952744,7.514226,8.22758,8.999237,9.472521,9.606275,9.942374,10.600855,11.293632,11.657167,11.657167,11.406808,11.166737,11.331357,10.984968,10.521975,10.220171,10.052121,9.6645775,9.1981535,8.80718,8.97523,9.921797,11.567999,13.574307,14.891269,15.638919,15.844694,15.443433,15.011304,14.706071,14.997586,15.580616,15.361122,13.375391,11.821788,10.199594,8.488229,7.1541195,7.143831,7.3084507,7.257007,6.7665763,5.7822843,4.2526884,2.9734523,2.0886188,1.6804979,1.7662375,1.6667795,1.5604624,1.8108221,2.4727325,3.2992632,3.8891523,4.5339146,5.0346346,5.456474,6.118384,6.3790326,6.591667,7.1232533,7.905199,8.440215,9.767465,11.509696,12.795791,13.279363,13.152468,12.9981365,13.015285,12.96727,12.908967,13.190193,13.37882,13.738928,14.05102,14.184773,14.123041,13.9138365,13.848674,13.773223,13.649758,13.560589,13.642899,14.109323,15.001016,16.328266,18.03963,19.744135,20.584383,20.237995,18.931322,17.436022,16.925014,16.486027,15.854982,14.970149,13.978998,12.922686,12.740917,12.977559,13.183334,12.915827,12.579727,12.46312,12.898679,13.900118,15.141628,15.741806,15.361122,14.977009,14.987297,15.206791,14.565458,13.865822,13.725209,14.119612,14.387119,14.277372,14.171056,14.088745,14.085316,14.246507,13.701202,13.512574,13.533153,13.519434,13.128461,12.88496,12.531713,12.161317,11.924676,12.024134,11.986408,11.736049,11.760056,12.130451,12.517994,12.425395,12.229909,11.838936,11.375941,11.180455,11.146159,11.087856,11.197603,11.598865,12.349944,12.603734,12.531713,12.281353,12.085866,12.264205,12.874671,12.88839,12.744347,12.703192,12.836946,13.4645605,14.081886,14.325387,14.356253,14.874121,15.7795315,15.854982,15.693792,15.662926,15.892709,16.407146,17.29884,18.180243,18.945042,19.771572,21.057667,21.335464,21.11597,20.773012,20.550089,20.86904,21.167414,21.253153,21.208569,21.393766,21.1194,20.248285,19.28457,18.482046,17.864721,17.305698,17.46003,17.487467,17.051908,16.321407,16.39,16.2974,15.899568,15.512024,15.909856,16.835844,17.53548,18.416885,19.54522,20.632399,19.792149,18.996485,18.221397,17.562918,17.237106,17.312557,17.165085,17.093063,17.333136,18.04306,18.053349,17.981327,17.86815,17.778982,17.813278,18.019053,18.091074,18.04649,17.936743,17.86815,18.012194,18.265984,18.36544,18.228258,17.971039,17.501184,16.894148,16.225378,15.584045,15.076467,14.342535,13.55373,12.850664,12.257345,11.694893,11.067279,10.449953,9.873782,9.400499,9.132992,8.879202,8.608265,8.40249,8.299602,8.303031,8.282454,8.296172,8.378482,8.464222,8.354475,8.193284,8.162418,8.196714,8.237869,8.213862,8.162418,8.186425,8.182996,8.128122,8.093826,7.936065,7.7028537,7.5553813,7.5039372,7.4284863,7.1849856,6.831738,6.5950966,6.526505,6.5059276,6.2418494,5.8988905,5.535354,5.1409516,4.6436615,4.3041325,4.046913,3.8514268,3.6799474,3.5016088,3.2135234,3.0043187,2.843128,2.702515,2.5413244,2.369845,2.2120838,2.0577524,1.9068506,1.7525192,1.6084765,1.4472859,1.2792361,1.097468,0.89169276,0.01371835,0.06859175,0.07888051,0.07545093,0.08573969,0.12689474,0.15090185,0.14747226,0.14061308,0.14061308,0.1371835,0.09259886,0.106317215,0.11317638,0.09945804,0.08573969,0.09602845,0.1097468,0.09945804,0.06859175,0.048014224,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.034295876,0.05144381,0.06859175,0.09602845,0.11317638,0.12689474,0.16804978,0.28808534,0.37382504,0.41840968,0.5727411,0.83338976,1.0220171,0.8505377,0.82996017,0.91912943,1.0768905,1.2586586,1.546744,2.0406046,2.253239,2.0131679,1.4644338,1.7250825,1.903421,1.9925903,1.9823016,1.8691251,1.7765263,2.4487255,3.1620796,3.542764,3.5873485,3.5393343,3.6079261,3.6765177,3.7176728,3.7965534,4.214963,4.6265135,5.1100855,5.6965446,6.3447366,7.208993,7.98408,8.038953,7.298162,6.2487082,4.5030484,3.9851806,4.0777793,4.3761535,4.6848164,4.0537724,2.5824795,1.5741806,1.3341095,1.1729189,1.3306799,1.2758065,1.0220171,0.7339317,0.7305021,0.7305021,0.7099246,1.0014396,1.6873571,2.609916,2.1915064,1.7525192,1.2620882,0.8745448,0.9362774,1.2037852,1.0837497,0.84024894,0.61046654,0.36010668,0.29494452,0.25378948,0.21263443,0.18862732,0.23664154,0.33952916,0.61389613,0.90884066,1.1146159,1.1763484,1.2449403,1.3649758,1.4095604,1.3684053,1.3478279,1.3855534,1.1797781,0.8676856,0.7305021,1.1934965,1.646202,2.0680413,1.9823016,1.3786942,0.6962063,0.52815646,0.607037,0.8848336,1.1283343,0.8848336,0.5796003,0.30866286,0.12346515,0.034295876,0.017147938,0.006859175,0.010288762,0.034295876,0.061732575,0.05144381,0.048014224,0.08573969,0.14061308,0.20234565,0.2709374,0.28465575,0.28808534,0.33609957,0.45270553,0.6344737,0.7922347,0.9259886,0.99801,0.9568549,0.7373613,0.7579388,0.864256,1.7902447,3.4913201,5.161529,6.691125,6.783724,6.0086374,4.856296,3.7279615,3.2135234,3.2649672,3.3541365,3.2718265,3.1243541,2.860276,3.2203827,4.125794,4.8837323,4.1772375,3.590778,3.7142432,3.7382503,3.3061223,2.5241764,2.0680413,1.845118,2.0920484,2.551613,2.4624438,2.1194851,1.9548649,1.978872,2.2155135,2.6990852,3.1072063,3.3987212,3.2443898,2.6579304,2.0063086,1.2758065,0.8779744,0.6276145,0.45613512,0.4046913,0.31895164,0.18519773,0.09602845,0.07545093,0.06859175,0.09259886,0.09602845,0.082310095,0.061732575,0.037725464,0.020577524,0.020577524,0.024007112,0.0274367,0.0274367,0.024007112,0.017147938,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0548734,0.17147937,0.32238123,0.490431,0.6241849,0.70649505,0.8265306,1.1660597,1.4953002,1.7730967,1.8931323,1.8554068,1.762808,1.7696671,1.8245405,1.937717,2.153781,2.5619018,3.1209247,3.882293,4.7328305,5.6142344,6.5162163,7.2158523,7.936065,8.700864,9.469091,10.14472,10.63858,10.813489,10.861504,10.875222,10.861504,11.070708,11.362224,11.742908,12.164746,12.521424,12.840376,13.152468,13.416546,13.612033,13.745787,13.762935,13.670336,13.591455,13.4645605,13.046151,12.236768,11.856084,11.674315,11.297061,10.155008,8.985519,8.042382,7.9737906,8.827758,10.062409,10.436234,10.669447,10.497967,10.168727,10.446524,10.703742,10.100135,9.513676,9.349055,9.541112,10.14472,10.618003,11.194174,11.629731,11.2250395,10.295622,10.175586,10.22703,10.055551,9.530824,9.335337,8.954653,8.532814,8.107545,7.623973,7.2192817,6.9209075,6.6636887,6.495639,6.5813785,6.495639,6.375603,6.6465406,7.2878733,7.8263187,8.47451,9.132992,9.740028,10.264755,10.703742,10.683165,10.477389,10.278474,10.158438,10.065839,9.345626,9.129561,9.438225,9.928656,9.904649,9.499957,9.067829,9.071259,9.626852,10.511685,12.003556,13.327377,14.277372,14.733508,14.644339,14.085316,13.474849,13.155897,13.327377,14.054449,13.426835,12.620882,11.290202,9.668007,8.543102,7.81603,6.64997,5.439326,4.4516044,3.8102717,2.9734523,1.978872,1.2655178,0.94999576,0.7922347,0.71678376,0.7373613,0.864256,1.2003556,1.9514352,2.6887965,3.5153272,4.0777793,4.2835546,4.3281393,4.3452873,4.787704,5.6999745,6.756287,7.2638664,8.536243,11.026124,13.029003,13.96871,14.400838,15.014734,15.302819,14.953001,14.198492,13.821238,13.828096,14.54831,15.350834,15.865272,15.995596,15.858413,15.515453,14.970149,14.277372,13.505715,12.80265,12.713481,13.200482,14.287662,16.067617,17.995045,19.912186,20.580954,19.908754,18.972477,18.214539,17.29541,16.235666,15.093615,13.954991,13.183334,12.734058,12.627741,12.785502,13.022143,12.576297,12.641459,13.279363,14.620332,16.856422,17.95389,16.756964,15.542891,15.313108,15.772673,15.738377,15.830976,16.256245,16.777542,16.691803,16.191082,15.830976,15.892709,16.444872,17.339994,16.650646,16.067617,15.560039,15.100473,14.678635,14.263655,13.780083,13.190193,12.452832,11.509696,10.984968,10.645439,10.672876,11.026124,11.430815,11.492548,11.094715,10.566559,10.131001,9.884071,9.753747,9.695444,9.856634,10.196163,10.463672,10.39508,10.511685,10.624862,10.693454,10.840926,10.899229,11.063849,11.132441,11.036412,10.840926,11.324498,11.835506,12.336226,13.042721,14.445422,15.868701,16.05733,15.930434,15.927004,16.019604,16.287111,17.003895,18.193962,19.60695,20.70099,21.839613,21.53781,20.899906,20.6907,21.338894,22.172283,22.995384,23.677872,24.175161,24.535269,24.336353,23.331484,22.000803,21.019941,21.253153,21.733295,22.631847,23.084553,22.865059,22.388348,21.589252,20.580954,19.44919,18.574646,18.650097,18.79414,18.79414,19.325726,20.53294,22.052248,20.574095,19.685833,19.600092,19.9602,19.86417,19.733847,19.733847,19.991066,20.61182,21.69214,21.592682,21.153696,20.45063,19.744135,19.459478,19.634388,19.750994,19.805868,19.775002,19.6241,19.757853,20.045938,20.231136,20.189981,19.925903,19.315437,18.78385,18.310568,17.885298,17.511473,17.034761,16.513464,15.947581,15.3302555,14.634049,13.924125,13.289652,12.703192,12.205902,11.907528,11.595435,11.135871,10.717461,10.419086,10.189304,9.928656,9.818909,9.908078,10.086417,10.069269,10.048691,10.31277,10.569988,10.683165,10.662587,10.521975,10.39165,10.2236,9.97667,9.616563,9.153569,8.615124,8.134981,7.81603,7.7268605,7.425057,6.9723516,6.776865,6.8797526,6.944915,6.615674,6.2658563,5.90232,5.521636,5.103226,4.746549,4.431027,4.139512,3.8617156,3.6079261,3.3987212,3.223812,3.0660512,2.9117198,2.7470996,2.5721905,2.3972816,2.2120838,2.0097382,1.7833855,1.5707511,1.3512574,1.1283343,0.90884066,0.6927767,0.061732575,0.09602845,0.08916927,0.06859175,0.06859175,0.09259886,0.10288762,0.09602845,0.09259886,0.08916927,0.07545093,0.08916927,0.1097468,0.1097468,0.08573969,0.061732575,0.1097468,0.14061308,0.09259886,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.01371835,0.0274367,0.044584636,0.044584636,0.034295876,0.041155048,0.058302987,0.09259886,0.15090185,0.20234565,0.28808534,0.5007198,0.77851635,0.90198153,0.8265306,0.90884066,1.0631721,1.2449403,1.4644338,1.5981878,1.6873571,1.7662375,1.8416885,1.8931323,1.879414,1.8142518,1.7147937,1.7490896,2.2120838,2.5653315,2.8465576,3.0111778,3.0626216,3.0351849,2.7573884,3.2992632,4.763697,6.310441,6.1629686,5.6142344,5.3673043,5.6005163,6.3824625,7.675417,9.458802,10.618003,10.134431,8.251588,6.468202,4.773986,4.4859004,4.5339146,4.232111,3.2821152,2.3149714,1.371835,1.3169615,1.903421,1.7696671,1.6359133,1.3924125,1.097468,0.8745448,0.89855194,0.91227025,0.91569984,1.0940384,1.4267083,1.6942163,1.2655178,1.1763484,1.3855534,1.5947582,1.2655178,0.90198153,0.6241849,0.47328308,0.42183927,0.39783216,0.31209245,0.23664154,0.18176813,0.15090185,0.15090185,0.16462019,0.65162164,1.2758065,1.8588364,2.393852,1.920569,1.2415106,0.99801,1.214074,1.313532,1.2037852,1.0117283,0.77165717,0.5453044,0.4115505,0.6310441,1.1249046,1.1866373,0.72021335,0.24350071,0.34295875,0.47671264,0.6276145,0.83681935,1.1900668,1.2277923,0.6962063,0.20920484,0.017147938,0.030866288,0.017147938,0.01371835,0.01371835,0.01371835,0.01371835,0.041155048,0.06516216,0.09602845,0.15090185,0.26064864,0.48014224,0.48700142,0.5796003,0.78194594,0.85396725,0.7579388,0.7339317,0.7339317,0.72707254,0.70306545,0.70306545,0.70306545,1.7593783,3.8548563,5.90575,7.3564653,7.7680154,7.4353456,6.550512,5.1580997,4.046913,3.3198407,2.8637056,2.5756202,2.3801336,2.8088322,3.1072063,3.199805,3.1277838,3.0660512,3.1517909,3.8788633,4.4413157,4.417309,3.7691166,2.5241764,1.4335675,1.0631721,1.3409687,1.5707511,1.7662375,1.8519772,1.8965619,1.9411465,2.0131679,2.1983654,2.435007,2.4418662,2.1880767,1.9068506,1.5913286,1.2620882,0.939707,0.6756287,0.5658819,0.48014224,0.3566771,0.25378948,0.18862732,0.15090185,0.12689474,0.11317638,0.09945804,0.08573969,0.061732575,0.037725464,0.01371835,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.048014224,0.16462019,0.33609957,0.44584638,0.48357183,0.45613512,0.45613512,0.64133286,0.922559,1.1283343,1.2689474,1.3375391,1.313532,1.3478279,1.4027013,1.5433143,1.7936742,2.136633,2.6373527,3.3369887,4.149801,5.0140567,5.90575,6.7219915,7.4936485,8.289313,9.105555,9.887501,10.460241,10.789482,10.923236,10.933525,10.909517,10.984968,11.238758,11.581717,11.948683,12.312219,12.778643,13.186764,13.509145,13.7697935,14.037301,14.270514,14.291091,14.140189,13.814379,13.289652,13.094165,12.891819,12.72034,12.425395,11.657167,10.340206,9.441654,8.947794,9.122703,10.511685,11.698323,12.734058,12.442543,10.957532,9.750318,9.774324,9.880642,10.089847,10.518545,11.396519,11.763485,11.279913,10.734609,10.405369,10.041832,9.489669,9.345626,9.595985,10.1652975,10.909517,11.495977,10.717461,9.510246,8.354475,7.2947326,6.927767,6.5882373,6.135532,5.6793966,5.56965,5.7651367,6.1629686,6.5470824,6.7665763,6.728851,7.5725293,8.906639,9.9869585,10.508256,10.604284,10.017825,9.194724,8.182996,7.2467184,6.866034,6.7459984,6.8969,7.548522,8.625413,9.736599,9.794902,9.993818,10.281903,10.5597,10.679735,10.875222,11.31078,11.670886,11.80121,11.705182,10.813489,9.959522,9.287323,8.903209,8.865483,9.242738,10.117283,10.947243,11.458252,11.64345,10.31277,8.378482,6.869464,6.0223556,5.2644167,4.3007026,3.199805,2.0886188,1.196926,0.85396725,0.67219913,0.6344737,0.77508676,1.0597426,1.3889829,1.6084765,2.0303159,2.5619018,3.1449318,3.7553983,4.2286816,4.3041325,4.5167665,5.127233,6.1046658,7.3358874,8.176137,8.450503,8.457363,8.958082,9.678296,10.755186,11.694893,12.22305,12.284782,12.562579,12.9638405,13.646329,14.565458,15.45715,16.287111,16.595774,16.54776,16.095055,14.983868,13.7526455,12.528283,12.034423,12.404818,13.200482,14.870691,16.46888,17.881868,18.838724,18.934752,18.862732,18.440891,17.734396,16.811838,15.762384,15.223939,14.640909,13.865822,13.13189,13.046151,13.365103,13.186764,13.173045,13.704632,14.87755,15.388559,15.776102,16.232237,16.832415,17.518333,18.176813,18.259123,18.149376,18.231688,18.890167,18.718689,18.019053,17.652086,17.669235,17.302269,15.704081,14.534592,13.437123,12.603734,12.785502,13.152468,13.756075,13.738928,12.816368,11.290202,10.803201,10.377932,9.962952,10.0041065,11.444533,13.114742,12.308789,10.871792,9.764035,9.016385,9.297611,9.743458,9.945804,9.757176,9.294182,8.597976,9.585697,11.149589,12.562579,13.488567,13.402828,12.833516,12.271064,11.89038,11.537132,11.180455,11.029553,11.029553,11.369082,12.466551,13.673765,15.2033615,16.540901,17.46003,18.019053,17.604073,18.362011,20.340883,22.127699,20.858751,18.845583,17.96761,17.703531,17.785841,18.187103,18.492336,18.752985,19.089085,19.593233,20.323736,21.129688,21.167414,21.208569,21.825895,23.376068,23.828773,23.959099,23.77733,23.485815,23.499533,24.243753,23.760181,22.631847,21.726437,22.19972,21.750444,20.28944,20.155685,21.757303,23.588703,22.552967,22.340332,22.875349,23.489244,22.902784,22.306036,22.062536,21.925352,21.77788,21.668133,22.546108,23.132568,23.18744,22.899355,22.889067,23.084553,22.913074,22.594122,22.251163,21.894485,21.479506,21.112541,20.923914,20.79016,20.340883,19.44919,19.298288,19.469769,19.45262,18.646667,18.022482,17.576635,17.21996,16.88043,16.46545,16.050468,15.560039,15.018164,14.483148,14.068168,13.725209,13.413116,12.991278,12.421966,11.763485,11.482259,11.231899,10.97468,10.72775,10.542552,10.446524,10.374502,10.326488,10.30934,10.347065,10.2236,10.120712,10.113853,10.103564,9.81205,9.163857,8.673427,8.275595,7.922347,7.5690994,7.239859,6.8626046,6.5470824,6.3481665,6.2864337,6.3481665,6.23499,6.001778,5.7479887,5.6142344,5.394741,5.055212,4.6916757,4.338428,3.998899,3.789694,3.5633414,3.333559,3.100347,2.867135,2.6236343,2.3904223,2.1503513,1.903421,1.6496316,1.3684053,1.0871792,0.82996017,0.607037,0.4115505,0.072021335,0.08916927,0.09259886,0.082310095,0.07545093,0.07888051,0.09259886,0.08573969,0.07888051,0.06516216,0.01371835,0.08573969,0.12346515,0.13032432,0.12346515,0.1097468,0.08916927,0.06859175,0.037725464,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.0034295875,0.010288762,0.024007112,0.037725464,0.044584636,0.044584636,0.037725464,0.05144381,0.082310095,0.10288762,0.14404267,0.26407823,0.47671264,0.7339317,0.9259886,0.9877212,0.97400284,0.99801,1.1111864,1.2826657,1.5055889,1.7010754,1.8554068,2.0165975,2.318401,2.6579304,2.5413244,2.3561265,2.3732746,2.750529,2.819121,2.8328393,2.867135,3.069481,3.6593697,4.9214582,5.020916,4.6265135,4.0537724,3.2855449,3.2512488,4.2046742,5.1238036,5.6210938,5.9297566,4.9488945,4.9351764,5.871454,7.0375133,6.9826403,6.351596,5.1066556,3.9200184,3.0866287,2.534465,2.7128036,2.3767042,2.1297739,2.1229146,2.037175,1.8931323,1.786815,1.5124481,1.1592005,1.0940384,1.1866373,1.3752645,1.4369972,1.3169615,1.1454822,0.6790583,0.5007198,0.5453044,0.7305021,0.94999576,0.9534253,0.6927767,0.4355576,0.29837412,0.22635277,0.16804978,0.1371835,0.12003556,0.14404267,0.26407823,0.4389872,0.8471081,1.2620882,1.587899,1.821111,1.4541451,1.0357354,0.96371406,1.2072148,1.3238207,1.3615463,1.2723769,1.1317638,0.9877212,0.864256,0.84024894,0.89855194,1.0048691,1.097468,1.097468,0.7373613,0.70649505,0.9362774,1.1694894,0.94656616,0.6790583,0.36696586,0.14747226,0.05144381,0.006859175,0.0034295875,0.010288762,0.020577524,0.030866288,0.041155048,0.07545093,0.07888051,0.08573969,0.116605975,0.18519773,0.37725464,0.5624523,0.7888051,1.0254467,1.1489118,1.097468,0.9774324,0.83338976,0.7442205,0.7888051,0.7956643,0.7476501,1.3924125,2.9048605,4.866585,8.584257,9.362774,7.606825,4.846007,3.7279615,3.0077481,2.6373527,2.5413244,2.6579304,2.9288676,2.6545007,2.4041407,2.2086544,2.16064,2.4315774,3.0043187,3.3712845,3.5530527,3.5599117,3.4021509,2.585909,1.6770682,1.155771,1.0871792,1.1317638,1.4061309,1.4747226,1.4541451,1.4678634,1.6496316,1.7833855,1.8245405,2.177788,2.8705647,3.5564823,2.4384367,1.5604624,0.9602845,0.6344737,0.5041494,0.41840968,0.37725464,0.32238123,0.22292319,0.07888051,0.07545093,0.072021335,0.07888051,0.08916927,0.072021335,0.058302987,0.058302987,0.058302987,0.048014224,0.041155048,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.048014224,0.0548734,0.08573969,0.15090185,0.274367,0.30523327,0.28122616,0.25378948,0.2777966,0.37382504,0.61389613,0.7956643,0.9328478,1.0185875,1.0323058,1.0666018,1.138623,1.2826657,1.5124481,1.8073926,2.218943,2.7539587,3.40901,4.180667,5.0620713,5.967482,6.8214493,7.6788464,8.549961,9.400499,10.0041065,10.491108,10.779194,10.899229,10.984968,11.084427,11.348505,11.694893,12.079007,12.483699,12.830087,13.049581,13.29994,13.615462,13.903547,13.893259,13.917266,13.989287,14.054449,13.999576,14.006435,13.862392,13.612033,13.289652,12.891819,12.569438,12.418536,12.264205,12.147599,12.308789,12.181894,11.941824,11.640019,11.513125,11.982979,11.958971,11.80464,11.540562,11.211322,10.909517,10.858074,10.662587,10.353925,9.938945,9.417647,9.14328,9.14328,9.445084,9.949233,10.4705305,10.247607,9.506817,8.601405,7.740579,6.999788,6.2830043,5.638242,5.2815647,5.3432975,5.8508763,6.691125,7.2535777,7.531374,7.7028537,8.14527,8.820899,9.033533,9.006097,8.916927,8.89635,8.700864,8.663138,8.309891,7.658269,7.2192817,7.116394,7.0272245,7.006647,7.2467184,8.06296,8.838047,9.455373,10.096705,10.779194,11.341646,11.125582,10.768905,10.2921915,9.873782,9.822338,9.606275,8.752307,7.764586,6.914048,6.252138,6.64997,7.2295704,7.6274023,7.8331776,8.162418,8.453933,8.351046,8.035523,7.3530354,5.813151,4.5853586,3.6147852,2.6373527,1.6873571,1.1111864,1.5227368,1.7971039,1.8691251,1.7799559,1.670209,1.5947582,1.6290541,1.9445761,2.5756202,3.4124396,4.170378,4.396731,4.3109913,4.3658648,5.223262,6.358455,6.9826403,7.473071,8.086967,8.958082,9.091836,9.208443,9.280463,9.318189,9.39021,9.719451,10.13786,10.679735,11.334786,12.037852,12.596875,12.915827,12.984418,12.778643,12.274493,11.609154,10.988399,10.6145735,10.64201,11.173596,12.044711,12.960411,13.762935,14.339106,14.603184,14.812388,14.863832,14.671775,14.167625,13.334236,12.46312,11.732618,11.190743,10.89237,10.875222,10.878652,10.820349,10.813489,10.97468,11.434244,11.965831,12.723769,13.498857,14.212211,14.904987,15.621771,16.386568,17.185663,17.916164,18.389448,18.228258,18.21111,18.28313,18.413456,18.571217,18.732407,18.163095,17.274832,16.37628,15.690363,15.337115,14.843254,14.147048,13.238208,12.171606,12.072148,12.199042,12.22305,12.133881,12.22648,12.315649,12.487128,12.905538,13.413116,13.557159,13.615462,13.680624,13.985858,14.273943,13.821238,13.368532,12.792361,12.240198,11.808069,11.523414,12.277924,13.039291,13.852104,14.7369375,15.662926,16.410576,17.309128,17.823566,17.703531,16.993607,17.031332,17.271402,17.607502,18.005335,18.509483,19.137098,20.045938,21.033659,21.4555,20.234566,18.924463,17.929884,17.1205,16.46888,16.04018,16.462019,16.46545,16.170506,15.834405,15.834405,15.817257,15.817257,16.023033,16.441442,16.907866,17.309128,18.094503,18.612371,18.564358,18.02934,18.255693,18.413456,18.38259,18.293419,18.516342,18.54378,18.156237,18.060207,18.482046,19.171394,19.812727,20.79016,21.568676,21.678423,20.680412,20.35803,20.594673,21.088533,21.716148,22.53239,23.060547,23.129137,22.919933,22.676432,22.69358,22.683292,22.395206,22.052248,21.757303,21.482935,21.143406,20.779871,20.430052,20.052797,19.53493,18.965618,18.574646,18.145947,17.641798,17.20624,16.739817,16.13278,15.656067,15.354263,15.035312,14.4145565,13.780083,13.145609,12.566009,12.140739,11.818358,11.550851,11.2421875,10.871792,10.494537,10.323058,10.189304,10.065839,9.914937,9.712592,9.527394,9.297611,9.057541,8.841476,8.673427,8.543102,8.471081,8.48137,8.508806,8.433355,8.213862,8.021805,7.864044,7.73372,7.6033955,7.596536,7.6925645,7.534804,7.082098,6.591667,6.358455,6.245279,6.1801167,6.0669403,5.785714,5.470192,5.0826488,4.6916757,4.338428,4.033195,3.8274195,3.6593697,3.4433057,3.1312134,2.7333813,2.4007113,2.1091962,1.8279701,1.5398848,1.2449403,0.96371406,0.72021335,0.5178677,0.34981793,0.20577525,0.06859175,0.09259886,0.09602845,0.08573969,0.07545093,0.07545093,0.044584636,0.061732575,0.07545093,0.06859175,0.037725464,0.041155048,0.05144381,0.07888051,0.11317638,0.09602845,0.044584636,0.020577524,0.010288762,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.024007112,0.0274367,0.041155048,0.048014224,0.06859175,0.09602845,0.1097468,0.12346515,0.28465575,0.52472687,0.78194594,1.0048691,1.0425946,0.922559,0.8676856,0.9602845,1.1351935,1.4747226,1.6599203,1.7010754,1.7696671,2.177788,2.585909,2.5138876,2.5001693,2.8088322,3.4433057,3.1415021,2.901431,2.7573884,2.867135,3.532475,4.972902,4.7602673,4.180667,4.3795834,6.355026,6.159539,5.06893,4.506478,4.7191124,4.7774153,3.508468,3.4295874,4.431027,5.562791,5.0414934,4.3761535,3.542764,2.8465576,2.417859,2.2223728,2.1229146,2.0474637,2.352697,2.7745364,2.4452958,1.8005334,1.6736387,1.5981878,1.4781522,1.5741806,1.5536032,1.5055889,1.3238207,1.0494537,0.8779744,0.7990939,0.7133542,0.6824879,0.78537554,1.1249046,1.1077567,0.7476501,0.41840968,0.25721905,0.16462019,0.18176813,0.18176813,0.1920569,0.24350071,0.39097297,0.58988905,0.90198153,1.1900668,1.3889829,1.4953002,1.0597426,0.71678376,0.88826317,1.4335675,1.6667795,1.6153357,1.488441,1.3169615,1.1043272,0.8196714,0.72707254,0.7339317,0.84024894,0.9911508,1.0460242,0.7099246,0.67219913,0.86082643,1.0734608,0.9842916,0.7990939,0.44927597,0.18176813,0.06859175,0.037725464,0.01371835,0.01371835,0.020577524,0.034295876,0.044584636,0.061732575,0.12003556,0.1920569,0.24350071,0.26750782,0.33609957,0.41840968,0.5796003,0.78537554,0.91912943,0.91227025,0.823101,0.69963586,0.6173257,0.67219913,0.72021335,0.77165717,1.2758065,2.3424082,3.7485392,6.142391,7.291303,7.3839016,6.90033,6.6053853,6.142391,4.9831905,3.858286,3.1346428,2.7916842,2.5001693,2.318401,2.1434922,2.037175,2.2360911,2.719663,2.8534167,2.9048605,3.0900583,3.5599117,3.018037,1.9548649,1.2312219,1.0871792,1.1214751,1.546744,1.7319417,1.7490896,1.6667795,1.5638919,1.3958421,1.0940384,1.1832076,1.7696671,2.5584722,1.7388009,1.1077567,0.7373613,0.58302987,0.50757897,0.4424168,0.36696586,0.274367,0.16462019,0.05144381,0.037725464,0.0274367,0.034295876,0.044584636,0.041155048,0.0274367,0.034295876,0.037725464,0.030866288,0.0274367,0.024007112,0.01371835,0.010288762,0.010288762,0.017147938,0.0034295875,0.0,0.006859175,0.01371835,0.010288762,0.0034295875,0.0,0.0034295875,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.017147938,0.024007112,0.0274367,0.037725464,0.06859175,0.14061308,0.16119061,0.14061308,0.13375391,0.16119061,0.21263443,0.40126175,0.5624523,0.70649505,0.823101,0.86082643,0.86082643,0.90198153,1.0048691,1.1900668,1.4781522,1.8691251,2.3321195,2.884283,3.542764,4.3041325,5.2026844,6.111525,7.006647,7.888051,8.783174,9.517105,10.127572,10.580277,10.906088,11.183885,11.434244,11.773774,12.205902,12.655178,12.96727,13.152468,13.176475,13.238208,13.399398,13.560589,13.80066,13.972139,13.924125,13.71492,13.6086035,13.38911,13.265644,13.179905,13.049581,12.758065,12.751206,13.035862,13.272504,13.341095,13.334236,12.874671,12.435684,12.233338,12.411677,13.056439,13.166186,13.059869,12.603734,11.72233,10.38479,9.839486,9.568549,9.3079,8.944365,8.529384,8.381912,8.683716,9.201583,9.757176,10.206452,9.89436,9.187865,8.289313,7.363324,6.543653,5.950334,5.6965446,5.744559,6.0395036,6.5162163,7.1884155,7.589677,7.5725293,7.2295704,6.9071894,7.459353,7.7542973,7.9600725,8.06639,7.9017696,7.7577267,7.8091707,7.7268605,7.5416627,7.64798,7.8949103,8.008087,8.090397,8.207003,8.39563,8.687145,9.582268,10.618003,11.365653,11.413667,10.971251,10.422516,9.839486,9.338767,9.088407,8.783174,8.128122,7.3393173,6.5127864,5.638242,5.394741,5.446185,5.439326,5.3432975,5.442755,5.9434752,6.2727156,6.1801167,5.6005163,4.650521,4.016047,3.292404,2.5619018,1.9651536,1.6873571,1.9857311,2.386993,2.4761622,2.1674993,1.6770682,1.5364552,1.4472859,1.4610043,1.670209,2.2086544,2.7162333,3.0146074,3.3815732,4.0606318,5.2335505,6.1766872,6.776865,7.0306544,7.2021337,7.822889,8.073249,8.30646,8.621983,8.868914,8.656279,8.625413,8.766026,9.205012,9.832627,10.288762,10.415657,10.484249,10.467101,10.353925,10.158438,9.904649,9.702303,9.623423,9.729739,10.062409,10.484249,10.827208,11.039842,11.156448,11.286773,11.413667,11.47197,11.369082,11.05356,10.528833,9.921797,9.414218,9.06097,8.862054,8.783174,8.711152,8.666568,8.628842,8.618553,8.680285,8.8929205,9.256456,9.637141,9.993818,10.350495,10.762046,11.38966,12.157887,12.936404,13.533153,13.937843,14.472859,15.062748,15.704081,16.46545,16.907866,17.171944,17.418875,17.53891,17.141079,16.715809,15.899568,15.001016,14.328816,14.212211,14.263655,13.920695,13.430264,13.008426,12.860953,12.956982,13.564018,14.54831,15.704081,16.736387,17.117071,17.600643,18.173384,18.663815,18.763273,18.567787,18.190533,18.091074,18.094503,17.384579,15.697222,15.083325,15.100473,15.429714,15.868701,16.777542,18.053349,19.133669,19.754423,19.95677,20.502073,20.330595,19.95334,19.62067,19.353163,19.147387,19.21255,19.257133,19.047928,18.434032,18.331144,17.87501,17.274832,16.811838,16.86671,17.024471,17.147938,16.979887,16.45516,15.707511,15.302819,15.199932,15.357693,15.590904,15.580616,15.642348,16.005884,16.245956,16.263103,16.259674,16.722668,17.089634,17.333136,17.480608,17.604073,17.53548,17.518333,17.62122,17.833855,18.073925,18.814716,19.744135,20.19684,20.045938,19.685833,20.70442,22.007662,22.666143,22.53925,22.247734,22.628418,22.803328,22.659285,22.299177,22.03167,21.85333,21.489796,21.009653,20.491785,20.02193,19.792149,19.53493,19.215979,18.818146,18.324286,17.86815,17.53891,17.20281,16.818697,16.424294,15.954441,15.343974,14.7369375,14.188204,13.690913,13.179905,12.730629,12.288212,11.862943,11.537132,11.324498,11.156448,10.933525,10.645439,10.360784,10.244178,10.134431,9.983529,9.794902,9.616563,9.451943,9.256456,9.043822,8.81747,8.584257,8.429926,8.330468,8.292743,8.299602,8.289313,8.2310095,8.162418,8.076678,7.9600725,7.798882,7.716572,7.795452,7.8263187,7.630832,7.0615206,6.48535,6.101236,5.8234396,5.5662203,5.2438393,4.9660425,4.695105,4.4447455,4.2046742,3.9337368,3.6079261,3.333559,3.0557625,2.74367,2.4075704,2.0989075,1.8005334,1.5124481,1.2312219,0.9602845,0.70306545,0.4938606,0.32924038,0.1920569,0.08916927,0.0548734,0.082310095,0.08573969,0.082310095,0.07545093,0.07545093,0.044584636,0.061732575,0.07545093,0.06516216,0.037725464,0.006859175,0.0,0.024007112,0.06516216,0.06516216,0.0274367,0.01371835,0.006859175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.01371835,0.01371835,0.041155048,0.061732575,0.08916927,0.11317638,0.12346515,0.14061308,0.34638834,0.6001778,0.8128122,0.9602845,0.9568549,0.85739684,0.85739684,1.0082988,1.2209331,1.5638919,1.6256244,1.5158776,1.4541451,1.7593783,2.0817597,2.177788,2.2600982,2.469303,2.8808534,2.6819375,2.620205,2.6819375,2.860276,3.1415021,3.9303071,4.245829,4.437886,5.0895076,7.0306544,6.6122446,4.99005,4.1292233,4.331569,4.2423997,3.1860867,3.1620796,3.7005248,4.0263357,3.069481,2.4658735,2.2600982,2.2463799,2.277246,2.2841053,1.8245405,1.7593783,2.194936,2.7779658,2.6887965,1.9480057,1.704505,1.6393428,1.6324836,1.7593783,1.6187652,1.4232788,1.2106444,1.0425946,1.0082988,1.1454822,1.2209331,1.2209331,1.1454822,1.0220171,0.8471081,0.5590228,0.33609957,0.23664154,0.17833854,0.22978236,0.274367,0.31552204,0.3841138,0.5624523,0.7442205,0.94999576,1.1008976,1.1489118,1.1111864,0.7990939,0.66191036,1.0597426,1.7422304,1.8313997,1.4815818,1.5398848,1.6221949,1.4541451,0.85739684,0.64819205,0.61046654,0.66876954,0.7407909,0.7407909,0.5418748,0.53501564,0.66191036,0.8196714,0.8711152,0.8025235,0.5212973,0.2709374,0.15433143,0.12346515,0.08573969,0.06859175,0.0548734,0.044584636,0.05144381,0.061732575,0.16119061,0.2709374,0.32924038,0.31209245,0.35324752,0.41498008,0.48700142,0.5590228,0.6241849,0.6824879,0.72021335,0.75450927,0.7922347,0.8676856,0.91912943,0.9568549,1.1694894,1.6016173,2.1434922,3.532475,5.0414934,6.680836,8.141841,8.81404,9.054111,7.39762,5.3981705,3.865145,2.867135,2.702515,2.7333813,2.5893385,2.2566686,2.095478,2.1160555,2.1263442,2.218943,2.4898806,3.0283258,2.767677,1.9754424,1.4815818,1.5261664,1.7388009,1.9548649,2.0406046,2.0337453,1.9239986,1.646202,1.2929544,0.7956643,0.53158605,0.65162164,1.0734608,0.78194594,0.5624523,0.45613512,0.4355576,0.41498008,0.3841138,0.31209245,0.22292319,0.14061308,0.06516216,0.024007112,0.01371835,0.01371835,0.01371835,0.01371835,0.006859175,0.006859175,0.010288762,0.010288762,0.010288762,0.010288762,0.01371835,0.01371835,0.017147938,0.024007112,0.010288762,0.0034295875,0.0034295875,0.010288762,0.01371835,0.006859175,0.006859175,0.010288762,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006859175,0.037725464,0.072021335,0.07888051,0.08573969,0.106317215,0.12346515,0.23664154,0.36010668,0.5041494,0.64133286,0.72021335,0.6962063,0.69963586,0.7407909,0.86082643,1.1351935,1.5124481,1.9720128,2.5001693,3.0866287,3.7348208,4.5784993,5.4667625,6.3653145,7.2775846,8.23444,9.057541,9.767465,10.38479,10.9198065,11.372512,11.763485,12.168177,12.665466,13.186764,13.509145,13.55373,13.423406,13.275933,13.173045,13.063298,13.155897,13.173045,12.97413,12.651748,12.5145645,12.555719,12.740917,12.874671,12.871242,12.723769,12.79922,13.173045,13.488567,13.564018,13.368532,12.97413,12.734058,12.740917,12.956982,13.207341,13.001566,12.5145645,11.653738,10.39165,8.772884,7.9292064,7.599966,7.4284863,7.2535777,7.1026754,7.332458,7.9189177,8.608265,9.211872,9.599416,9.489669,8.89635,8.052671,7.143831,6.3310184,5.9571934,5.9571934,6.2487082,6.684266,7.034084,7.3255987,7.366754,7.0615206,6.5230756,6.077229,6.509357,6.999788,7.4353456,7.699424,7.675417,8.001227,8.241299,8.354475,8.405919,8.549961,8.539673,8.738589,9.026674,9.163857,8.786603,8.834618,9.678296,10.405369,10.566559,10.175586,9.914937,9.626852,9.379922,9.253027,9.331907,9.235879,8.748878,7.9772205,7.023795,5.970912,5.2335505,4.852866,4.6916757,4.7328305,5.0895076,5.641671,5.442755,4.756838,3.9097297,3.3026927,3.1689389,2.8739944,2.49331,2.1572106,2.054323,2.1023371,2.2155135,2.0989075,1.7833855,1.5913286,1.587899,1.5021594,1.3272504,1.1592005,1.214074,1.3992717,1.670209,2.2978237,3.2992632,4.4413157,5.2164025,5.8337283,6.0497923,5.9812007,6.118384,6.385892,6.773435,7.5107965,8.309891,8.371623,8.309891,8.152129,8.155559,8.357904,8.577398,8.577398,8.604835,8.621983,8.611694,8.577398,8.529384,8.522525,8.597976,8.745448,8.903209,9.057541,9.084977,9.019815,8.923786,8.916927,8.906639,8.868914,8.735159,8.498518,8.196714,7.8777623,7.596536,7.363324,7.1781263,7.051232,6.975781,6.914048,6.842027,6.7494283,6.636252,6.5470824,6.4887795,6.461343,6.4887795,6.5985265,6.7391396,6.989499,7.332458,7.740579,8.186425,8.834618,9.496528,10.237319,11.087856,12.05843,12.535142,12.826657,13.200482,13.629181,13.80409,13.522863,12.737488,12.370522,12.710052,13.38911,12.850664,12.000127,11.218181,10.696883,10.456812,10.621432,11.22161,12.120162,13.227919,14.496866,15.22051,16.002455,16.736387,17.412016,18.104792,18.61923,19.263992,20.179693,20.971928,20.724997,18.70497,17.508043,17.058767,17.058767,16.990177,17.099922,18.03963,19.061647,20.35803,23.070835,25.238335,25.557285,24.84736,23.653864,22.234016,21.891056,21.561817,21.211998,20.86561,20.587814,20.556948,20.61525,20.570665,20.474638,20.632399,20.683842,20.457489,19.895037,19.075365,18.221397,17.693241,17.339994,17.226818,17.247395,17.12736,17.075916,17.034761,16.945591,16.931873,17.309128,17.909306,18.396307,18.934752,19.418324,19.483486,19.078794,18.996485,19.137098,19.380598,19.582945,19.730417,19.980776,19.987637,19.792149,19.833303,21.013083,22.244305,22.751883,22.491234,22.168854,22.271742,21.959648,21.465788,20.923914,20.395756,19.905325,19.329155,18.646667,17.936743,17.36057,17.113642,16.911295,16.695232,16.444872,16.167076,15.848124,15.63206,15.429714,15.172495,14.819247,14.452282,14.037301,13.567448,13.080446,12.6586075,12.377381,12.144169,11.9040985,11.660598,11.454823,11.358793,11.252477,11.05356,10.772334,10.518545,10.398509,10.30934,10.161868,9.949233,9.73317,9.626852,9.499957,9.280463,8.985519,8.707723,8.525954,8.405919,8.333898,8.285883,8.23444,8.186425,8.141841,8.05953,7.9120584,7.682276,7.4627824,7.3564653,7.332458,7.274155,6.941485,6.447624,5.936616,5.453044,5.0312047,4.681387,4.4687524,4.262977,4.0949273,3.9303071,3.6593697,3.216953,2.8396983,2.5241764,2.2635276,2.0303159,1.704505,1.3615463,1.1351935,1.039165,0.9362774,0.6036074,0.36010668,0.1920569,0.08573969,0.034295876,0.044584636,0.0548734,0.06516216,0.07545093,0.07545093,0.06516216,0.072021335,0.06516216,0.0548734,0.037725464,0.0,0.0,0.0,0.0034295875,0.020577524,0.0548734,0.048014224,0.034295876,0.017147938,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.01371835,0.041155048,0.06859175,0.09602845,0.11317638,0.116605975,0.17833854,0.4081209,0.6344737,0.7682276,0.7956643,0.77851635,0.7990939,0.9328478,1.1660597,1.3992717,1.6187652,1.529596,1.3546871,1.2758065,1.4267083,1.6736387,1.9720128,2.020027,1.8108221,1.6427724,1.8485477,2.1297739,2.510458,2.7951138,2.568761,2.5893385,3.7039545,4.6745276,4.866585,4.266407,4.1600895,4.139512,4.214963,4.262977,4.0194764,3.2032347,3.0557625,3.093488,2.9151495,2.2052248,2.0337453,2.1126258,2.2841053,2.428148,2.4761622,2.1743584,2.1263442,2.201795,2.3767042,2.6990852,2.2909644,1.9342873,1.6839274,1.5673214,1.5570327,1.4232788,1.3341095,1.3032433,1.3821237,1.670209,2.0028791,2.0714707,1.9274281,1.5124481,0.67219913,0.4081209,0.34981793,0.31552204,0.2469303,0.21263443,0.26407823,0.40126175,0.5041494,0.5727411,0.7305021,0.89169276,1.0460242,1.0631721,0.90884066,0.64476246,0.72364295,0.90541106,1.3375391,1.8005334,1.7216529,1.3512574,1.6530612,1.9823016,1.8588364,0.9877212,0.64819205,0.52815646,0.53158605,0.5727411,0.5624523,0.41840968,0.42183927,0.52472687,0.66533995,0.77165717,0.78194594,0.6173257,0.44584638,0.34638834,0.29151493,0.24007112,0.19548649,0.1371835,0.07545093,0.06859175,0.08573969,0.18519773,0.28808534,0.32924038,0.2709374,0.36353627,0.50757897,0.5521636,0.5041494,0.5212973,0.71678376,0.90884066,1.0906088,1.2243627,1.2346514,1.214074,1.1592005,1.0254467,0.8093826,0.5521636,2.1743584,3.8548563,5.6210938,7.349606,8.748878,9.873782,9.050681,7.56567,5.9400454,3.9440255,3.391862,3.3472774,3.1689389,2.6887965,2.201795,1.5810398,1.4095604,1.5055889,1.704505,1.8828435,1.937717,1.8279701,1.879414,2.1812177,2.585909,2.2326615,1.961724,1.9137098,1.9823016,1.8142518,1.4781522,1.1180456,0.8196714,0.59331864,0.37382504,0.274367,0.26750782,0.2709374,0.25721905,0.2469303,0.22635277,0.20577525,0.1920569,0.16804978,0.09259886,0.034295876,0.0274367,0.030866288,0.024007112,0.024007112,0.020577524,0.010288762,0.0034295875,0.0034295875,0.0034295875,0.0034295875,0.010288762,0.01371835,0.017147938,0.017147938,0.017147938,0.006859175,0.0,0.006859175,0.01371835,0.01371835,0.01371835,0.01371835,0.010288762,0.0,0.0,0.0034295875,0.0034295875,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.0548734,0.06516216,0.072021335,0.061732575,0.09945804,0.17490897,0.28808534,0.42526886,0.5453044,0.53158605,0.5144381,0.51100856,0.58302987,0.8093826,1.1523414,1.6256244,2.1674993,2.74367,3.3472774,4.1292233,4.9488945,5.8371577,6.7871537,7.7714453,8.608265,9.39707,10.13786,10.799771,11.341646,11.808069,12.21619,12.686044,13.214201,13.649758,13.666906,13.536582,13.327377,13.066729,12.7272,12.264205,11.893809,11.622872,11.458252,11.406808,11.931535,12.3911,12.624311,12.6757555,12.80265,12.915827,13.169616,13.37882,13.365103,12.977559,12.826657,12.63803,12.627741,12.71691,12.542002,11.578287,10.275044,8.923786,7.6959944,6.632822,5.9469047,5.669108,5.5250654,5.453044,5.6142344,6.3035817,7.0032177,7.6925645,8.292743,8.659708,8.738589,8.405919,7.8983397,7.3393173,6.7357097,6.368744,6.2144127,6.375603,6.715132,6.8454566,6.893471,6.7322803,6.39961,6.142391,6.4098988,6.927767,7.466212,7.857185,8.06639,8.213862,8.999237,9.5205345,9.815479,9.873782,9.654288,8.882631,8.796892,9.050681,9.2153015,8.81404,9.249598,9.619993,9.400499,8.7283,8.3922,8.7283,9.160428,9.352485,9.383351,9.740028,10.106995,9.716022,8.848335,7.720001,6.5024977,5.675967,5.2506986,5.2266912,5.5902276,6.307011,6.989499,6.228131,5.003768,3.8925817,3.0489032,2.7916842,2.7230926,2.5378947,2.2395205,2.1469216,2.1057668,1.7730967,1.3958421,1.2586586,1.704505,1.8965619,1.8416885,1.611906,1.3272504,1.1351935,1.214074,1.3478279,1.704505,2.2806756,2.8980014,3.5530527,4.1292233,4.5030484,4.5956473,4.3795834,4.40702,4.647091,5.429037,6.5642304,7.366754,7.682276,7.4524937,6.9517736,6.509357,6.5127864,6.691125,6.8969,7.058091,7.143831,7.1849856,7.1781263,7.205563,7.2467184,7.284444,7.301592,7.291303,7.257007,7.2124224,7.1781263,7.14726,7.099246,7.0375133,6.9209075,6.7494283,6.550512,6.3447366,6.1561093,5.9880595,5.844017,5.7274113,5.65539,5.576509,5.4804807,5.353586,5.195825,4.99005,4.791134,4.633373,4.5647807,4.6402316,4.695105,4.6916757,4.698535,4.770556,4.9351764,5.4804807,5.809721,6.0806584,6.4579134,7.1061053,7.6445503,7.349606,6.914048,6.7974424,7.2192817,7.174697,6.6739774,7.0546613,8.323608,9.187865,8.069819,7.239859,6.7322803,6.4407654,6.1286726,5.9640527,6.1904054,6.7357097,7.517656,8.467651,9.451943,10.240748,10.998687,11.784062,12.555719,13.6086035,14.853543,16.071047,17.089634,17.772121,17.933313,17.69667,17.754974,18.180243,18.413456,17.981327,18.03963,18.115082,19.089085,23.19087,26.291218,27.27208,26.846811,25.591581,23.94538,24.662163,24.888515,24.94339,24.895376,24.53184,23.76361,24.085993,24.555847,24.682741,24.411804,24.127148,22.985096,21.52066,20.334024,20.069946,19.94305,19.493774,19.095943,18.849012,18.591793,18.560926,18.427174,18.276272,18.245405,18.516342,18.989626,19.586374,20.443771,21.28059,21.386908,20.985645,21.033659,21.19828,21.301168,21.318316,21.050808,20.714708,20.313446,19.912186,19.648108,19.696121,19.757853,19.884748,20.19341,20.879328,20.598103,19.507494,18.509483,17.902447,17.343424,16.602633,15.865272,15.13134,14.479718,14.030442,13.708061,13.502286,13.371962,13.3033695,13.306799,13.207341,13.077017,12.88496,12.655178,12.46312,12.325937,12.181894,12.037852,11.9040985,11.80121,11.694893,11.55771,11.413667,11.269625,11.135871,11.105004,10.988399,10.768905,10.487679,10.244178,10.072699,10.024684,9.949233,9.760606,9.448513,9.3764925,9.270175,8.995808,8.601405,8.303031,8.131552,8.032094,7.963502,7.888051,7.7783046,7.689135,7.6033955,7.4936485,7.3358874,7.1061053,6.8797526,6.64997,6.427047,6.3001523,6.468202,6.56766,6.046363,5.360445,4.770556,4.3487167,4.125794,3.8617156,3.6525106,3.4638834,3.1483612,2.6304936,2.2223728,1.920569,1.704505,1.529596,1.2037852,0.8711152,0.75450927,0.84024894,0.8711152,0.5144381,0.26064864,0.09945804,0.024007112,0.017147938,0.044584636,0.044584636,0.044584636,0.06516216,0.07545093,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.0,0.024007112,0.06859175,0.09259886,0.0548734,0.0274367,0.010288762,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0034295875,0.01371835,0.041155048,0.0548734,0.06859175,0.07888051,0.09259886,0.20234565,0.3841138,0.5418748,0.6379033,0.6859175,0.6379033,0.6790583,0.84024894,1.0563129,1.1900668,1.2620882,1.1523414,1.1180456,1.2792361,1.6324836,1.9994495,2.318401,2.428148,2.3492675,2.287535,2.287535,2.16064,1.9651536,1.7388009,1.4953002,1.5433143,1.8313997,2.428148,3.3026927,4.3041325,5.6348124,5.8474464,4.8322887,3.4467354,3.4947495,3.957744,3.882293,3.5290456,3.0111778,2.3046827,2.2669573,2.3321195,2.3561265,2.3286898,2.3664153,2.5721905,3.0077481,3.2546785,3.1140654,2.6236343,2.16064,1.8142518,1.546744,1.371835,1.371835,1.4472859,1.5090185,1.546744,1.8519772,3.0351849,4.40359,3.9474552,2.9048605,1.8931323,0.91569984,0.7682276,0.8162418,0.6927767,0.3841138,0.21263443,0.32238123,0.6344737,0.85396725,0.8745448,0.77851635,0.864256,1.1592005,1.196926,0.8505377,0.34981793,0.84024894,1.1249046,1.1317638,1.1111864,1.6496316,2.4795918,2.4007113,1.961724,1.4027013,0.67219913,0.47671264,0.47328308,0.5453044,0.61046654,0.61046654,0.4389872,0.4424168,0.5590228,0.84367853,1.4815818,1.6736387,1.2483698,0.8162418,0.6344737,0.61046654,0.5007198,0.3806842,0.25378948,0.14061308,0.09259886,0.09259886,0.20234565,0.31209245,0.34638834,0.26064864,0.23664154,0.23664154,0.29151493,0.42526886,0.65505123,1.1454822,1.3958421,1.4747226,1.371835,0.9911508,0.78537554,0.9328478,0.9945804,0.78537554,0.3806842,1.4061309,2.726522,4.5613513,6.636252,8.162418,9.239308,11.245617,12.607163,11.670886,6.715132,4.5030484,3.6765177,3.542764,3.5564823,3.309552,2.0646117,1.3512574,1.0666018,1.1249046,1.4815818,1.8108221,2.0028791,2.1846473,2.4144297,2.6716487,1.8416885,1.2209331,1.3238207,1.9239986,2.0440342,1.6907866,1.903421,2.1674993,1.9720128,0.823101,0.33609957,0.26750782,0.28808534,0.2469303,0.19891608,0.08916927,0.061732575,0.09259886,0.12689474,0.09259886,0.041155048,0.041155048,0.05144381,0.061732575,0.061732575,0.037725464,0.020577524,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.01371835,0.017147938,0.030866288,0.030866288,0.01371835,0.006859175,0.01371835,0.01371835,0.0034295875,0.0,0.0,0.0,0.0,0.0,0.010288762,0.01371835,0.01371835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.037725464,0.09259886,0.16804978,0.29151493,0.31552204,0.31895164,0.33952916,0.4046913,0.5658819,0.8711152,1.3032433,1.8108221,2.369845,3.0043187,3.7382503,4.5990767,5.4907694,6.3653145,7.233,8.100685,8.9100685,9.654288,10.302481,10.803201,11.290202,11.616013,11.921246,12.284782,12.710052,12.943263,13.128461,13.255356,13.279363,13.107883,12.583157,12.175035,11.80464,11.46854,11.2593355,11.039842,10.803201,10.820349,11.14273,11.581717,11.619442,11.838936,12.332796,12.991278,13.502286,13.906977,13.255356,12.329367,11.55428,11.015835,9.517105,7.675417,6.540223,6.2658563,6.118384,6.3001523,6.0086374,5.381023,4.8837323,5.3090014,5.7754254,6.2555676,6.773435,7.3290286,7.905199,8.001227,8.134981,8.378482,8.529384,8.100685,7.298162,6.883182,6.550512,6.077229,5.3570156,5.40503,5.7925735,6.012067,6.042933,6.3481665,7.6171136,8.639131,9.4862385,9.932085,9.445084,9.091836,9.156999,9.39707,9.6817255,10.010965,9.119273,8.457363,8.39563,8.9100685,9.582268,10.388221,9.846346,8.934075,8.30646,8.330468,9.47938,11.249047,11.547421,10.179015,8.851766,8.776315,8.584257,8.309891,7.8091707,6.759717,5.9914894,6.1732574,6.4236174,6.3207297,5.90575,5.9914894,6.0395036,5.960623,5.6348124,4.928317,3.7931237,2.9322972,2.2978237,2.0097382,2.3664153,2.4144297,2.2429502,2.1743584,2.2909644,2.4247184,2.5961976,2.5310357,2.2429502,2.0028791,2.318401,2.6236343,2.4898806,2.318401,2.301253,2.411,2.8980014,3.333559,3.4192986,3.2066643,3.0969174,3.1449318,3.2958336,3.5530527,4.046913,5.0346346,5.535354,5.6519604,5.4941993,5.195825,4.914599,5.1683884,5.3158607,5.353586,5.329579,5.3398676,5.363875,5.4084597,5.439326,5.446185,5.4324665,5.394741,5.360445,5.3398676,5.3398676,5.3398676,5.353586,5.3570156,5.336438,5.2815647,5.171818,5.0620713,4.9351764,4.8254294,4.73969,4.65395,4.5819287,4.48933,4.389872,4.280125,4.1360826,3.974892,3.789694,3.6627994,3.642222,3.7382503,3.7622573,3.7862647,4.0023284,4.4584637,5.0826488,6.0086374,5.7651367,4.897451,4.0674906,4.0434837,3.9954693,3.9200184,3.8445675,3.799983,3.799983,4.262977,4.5442033,4.557922,4.4516044,4.623084,4.9420357,4.791134,4.6127954,4.664239,5.003768,4.722542,4.2698364,4.32471,5.0277753,5.967482,7.455923,8.543102,9.3764925,9.846346,9.551401,9.3079,9.129561,9.410788,10.22703,11.338216,11.619442,11.907528,12.22648,12.79922,14.068168,15.8138275,14.805529,13.203912,12.264205,12.315649,12.583157,12.943263,13.773223,15.059319,16.39,17.778982,19.089085,20.327166,21.136547,20.7833,20.759293,21.338894,21.911634,22.227156,22.384918,20.237995,18.252264,16.671225,15.868701,16.359133,17.87158,18.139088,17.857862,17.309128,16.359133,15.758954,15.306249,15.12448,15.206791,15.426285,16.050468,16.53404,16.914726,17.274832,17.761833,18.530062,19.912186,20.69413,20.392326,19.257133,19.572655,19.589804,18.69811,17.192522,16.266533,15.923574,15.501736,15.055889,14.616901,14.191633,13.814379,13.433694,13.097594,12.80265,12.4974165,12.168177,11.873232,11.612583,11.393089,11.245617,11.111863,10.957532,10.844356,10.792912,10.803201,10.840926,10.875222,10.9198065,10.960961,10.984968,10.97468,10.916377,10.830637,10.72775,10.604284,10.456812,10.319629,10.182446,10.038403,9.904649,9.791472,9.637141,9.441654,9.208443,8.927217,8.694004,8.656279,8.594546,8.399059,8.056101,7.936065,7.829748,7.6651278,7.449064,7.2775846,7.191845,7.143831,7.1198235,7.1061053,7.0958166,6.9860697,6.783724,6.5779486,6.39961,6.2418494,6.1801167,6.0737996,5.919468,6.0052075,6.8969,7.7748747,6.8866115,5.6073756,4.6402316,4.0434837,3.6525106,3.2992632,3.0043187,2.7230926,2.318401,1.7216529,1.3169615,1.0117283,0.77165717,0.6241849,0.5658819,0.6036074,0.53844523,0.30866286,0.01371835,0.08916927,0.12346515,0.11317638,0.06859175,0.030866288;
 } 
